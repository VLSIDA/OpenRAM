VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 107980.0 by 207952.5 ;
END  MacroSite
MACRO sram_1rw_32b_512w_1bank_freepdk45
   CLASS BLOCK ;
   SIZE 107980.0 BY 207952.5 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  17512.5 35.0 17582.5 175.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  20332.5 35.0 20402.5 175.0 ;
      END
   END DATA[1]
   PIN DATA[2]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  23152.5 35.0 23222.5 175.0 ;
      END
   END DATA[2]
   PIN DATA[3]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  25972.5 35.0 26042.5 175.0 ;
      END
   END DATA[3]
   PIN DATA[4]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  28792.5 35.0 28862.5 175.0 ;
      END
   END DATA[4]
   PIN DATA[5]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  31612.5 35.0 31682.5 175.0 ;
      END
   END DATA[5]
   PIN DATA[6]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  34432.5 35.0 34502.5 175.0 ;
      END
   END DATA[6]
   PIN DATA[7]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  37252.5 35.0 37322.5 175.0 ;
      END
   END DATA[7]
   PIN DATA[8]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  40072.5 35.0 40142.5 175.0 ;
      END
   END DATA[8]
   PIN DATA[9]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  42892.5 35.0 42962.5 175.0 ;
      END
   END DATA[9]
   PIN DATA[10]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  45712.5 35.0 45782.5 175.0 ;
      END
   END DATA[10]
   PIN DATA[11]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  48532.5 35.0 48602.5 175.0 ;
      END
   END DATA[11]
   PIN DATA[12]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  51352.5 35.0 51422.5 175.0 ;
      END
   END DATA[12]
   PIN DATA[13]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  54172.5 35.0 54242.5 175.0 ;
      END
   END DATA[13]
   PIN DATA[14]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  56992.5 35.0 57062.5 175.0 ;
      END
   END DATA[14]
   PIN DATA[15]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  59812.5 35.0 59882.5 175.0 ;
      END
   END DATA[15]
   PIN DATA[16]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  62632.5 35.0 62702.5 175.0 ;
      END
   END DATA[16]
   PIN DATA[17]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  65452.5 35.0 65522.5 175.0 ;
      END
   END DATA[17]
   PIN DATA[18]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  68272.5 35.0 68342.5 175.0 ;
      END
   END DATA[18]
   PIN DATA[19]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  71092.5 35.0 71162.5 175.0 ;
      END
   END DATA[19]
   PIN DATA[20]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  73912.5 35.0 73982.5 175.0 ;
      END
   END DATA[20]
   PIN DATA[21]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  76732.5 35.0 76802.5 175.0 ;
      END
   END DATA[21]
   PIN DATA[22]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  79552.5 35.0 79622.5 175.0 ;
      END
   END DATA[22]
   PIN DATA[23]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  82372.5 35.0 82442.5 175.0 ;
      END
   END DATA[23]
   PIN DATA[24]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  85192.5 35.0 85262.5 175.0 ;
      END
   END DATA[24]
   PIN DATA[25]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  88012.5 35.0 88082.5 175.0 ;
      END
   END DATA[25]
   PIN DATA[26]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  90832.5 35.0 90902.5 175.0 ;
      END
   END DATA[26]
   PIN DATA[27]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  93652.5 35.0 93722.5 175.0 ;
      END
   END DATA[27]
   PIN DATA[28]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  96472.5 35.0 96542.5 175.0 ;
      END
   END DATA[28]
   PIN DATA[29]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  99292.5 35.0 99362.5 175.0 ;
      END
   END DATA[29]
   PIN DATA[30]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  102112.5 35.0 102182.5 175.0 ;
      END
   END DATA[30]
   PIN DATA[31]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  104932.5 35.0 105002.5 175.0 ;
      END
   END DATA[31]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 11782.5 4655.0 11852.5 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 11077.5 4655.0 11147.5 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 10372.5 4655.0 10442.5 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 9667.5 4655.0 9737.5 ;
      END
   END ADDR[3]
   PIN ADDR[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 8962.5 4655.0 9032.5 ;
      END
   END ADDR[4]
   PIN ADDR[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 8257.5 4655.0 8327.5 ;
      END
   END ADDR[5]
   PIN ADDR[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 7552.5 4655.0 7622.5 ;
      END
   END ADDR[6]
   PIN ADDR[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6847.5 4655.0 6917.5 ;
      END
   END ADDR[7]
   PIN ADDR[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6142.5 4655.0 6212.5 ;
      END
   END ADDR[8]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1187.5 34240.0 1257.5 34380.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1892.5 34240.0 1962.5 34380.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.5 34240.0 552.5 34380.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  3340.0 34240.0 3475.0 34430.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  107630.0 35.0 107980.0 207987.5 ;
         LAYER metal1 ;
         RECT  4175.0 35.0 4525.0 207987.5 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  15102.5 35.0 15452.5 207987.5 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  4317.5 41945.0 4382.5 42150.0 ;
      RECT  8890.0 34695.0 8955.0 34760.0 ;
      RECT  8890.0 34422.5 8955.0 34487.5 ;
      RECT  8820.0 34695.0 8922.5 34760.0 ;
      RECT  8890.0 34455.0 8955.0 34727.5 ;
      RECT  8922.5 34422.5 9025.0 34487.5 ;
      RECT  14177.5 34695.0 14242.5 34760.0 ;
      RECT  14177.5 34207.5 14242.5 34272.5 ;
      RECT  11315.0 34695.0 14210.0 34760.0 ;
      RECT  14177.5 34240.0 14242.5 34727.5 ;
      RECT  14210.0 34207.5 17105.0 34272.5 ;
      RECT  8890.0 36130.0 8955.0 36195.0 ;
      RECT  8890.0 36402.5 8955.0 36467.5 ;
      RECT  8820.0 36130.0 8922.5 36195.0 ;
      RECT  8890.0 36162.5 8955.0 36435.0 ;
      RECT  8922.5 36402.5 9025.0 36467.5 ;
      RECT  14177.5 36130.0 14242.5 36195.0 ;
      RECT  14177.5 36617.5 14242.5 36682.5 ;
      RECT  11315.0 36130.0 14210.0 36195.0 ;
      RECT  14177.5 36162.5 14242.5 36650.0 ;
      RECT  14210.0 36617.5 17105.0 36682.5 ;
      RECT  8890.0 37385.0 8955.0 37450.0 ;
      RECT  8890.0 37112.5 8955.0 37177.5 ;
      RECT  8820.0 37385.0 8922.5 37450.0 ;
      RECT  8890.0 37145.0 8955.0 37417.5 ;
      RECT  8922.5 37112.5 9025.0 37177.5 ;
      RECT  14177.5 37385.0 14242.5 37450.0 ;
      RECT  14177.5 36897.5 14242.5 36962.5 ;
      RECT  11315.0 37385.0 14210.0 37450.0 ;
      RECT  14177.5 36930.0 14242.5 37417.5 ;
      RECT  14210.0 36897.5 17105.0 36962.5 ;
      RECT  8890.0 38820.0 8955.0 38885.0 ;
      RECT  8890.0 39092.5 8955.0 39157.5 ;
      RECT  8820.0 38820.0 8922.5 38885.0 ;
      RECT  8890.0 38852.5 8955.0 39125.0 ;
      RECT  8922.5 39092.5 9025.0 39157.5 ;
      RECT  14177.5 38820.0 14242.5 38885.0 ;
      RECT  14177.5 39307.5 14242.5 39372.5 ;
      RECT  11315.0 38820.0 14210.0 38885.0 ;
      RECT  14177.5 38852.5 14242.5 39340.0 ;
      RECT  14210.0 39307.5 17105.0 39372.5 ;
      RECT  8890.0 40075.0 8955.0 40140.0 ;
      RECT  8890.0 39802.5 8955.0 39867.5 ;
      RECT  8820.0 40075.0 8922.5 40140.0 ;
      RECT  8890.0 39835.0 8955.0 40107.5 ;
      RECT  8922.5 39802.5 9025.0 39867.5 ;
      RECT  14177.5 40075.0 14242.5 40140.0 ;
      RECT  14177.5 39587.5 14242.5 39652.5 ;
      RECT  11315.0 40075.0 14210.0 40140.0 ;
      RECT  14177.5 39620.0 14242.5 40107.5 ;
      RECT  14210.0 39587.5 17105.0 39652.5 ;
      RECT  8890.0 41510.0 8955.0 41575.0 ;
      RECT  8890.0 41782.5 8955.0 41847.5 ;
      RECT  8820.0 41510.0 8922.5 41575.0 ;
      RECT  8890.0 41542.5 8955.0 41815.0 ;
      RECT  8922.5 41782.5 9025.0 41847.5 ;
      RECT  14177.5 41510.0 14242.5 41575.0 ;
      RECT  14177.5 41997.5 14242.5 42062.5 ;
      RECT  11315.0 41510.0 14210.0 41575.0 ;
      RECT  14177.5 41542.5 14242.5 42030.0 ;
      RECT  14210.0 41997.5 17105.0 42062.5 ;
      RECT  8890.0 42765.0 8955.0 42830.0 ;
      RECT  8890.0 42492.5 8955.0 42557.5 ;
      RECT  8820.0 42765.0 8922.5 42830.0 ;
      RECT  8890.0 42525.0 8955.0 42797.5 ;
      RECT  8922.5 42492.5 9025.0 42557.5 ;
      RECT  14177.5 42765.0 14242.5 42830.0 ;
      RECT  14177.5 42277.5 14242.5 42342.5 ;
      RECT  11315.0 42765.0 14210.0 42830.0 ;
      RECT  14177.5 42310.0 14242.5 42797.5 ;
      RECT  14210.0 42277.5 17105.0 42342.5 ;
      RECT  8890.0 44200.0 8955.0 44265.0 ;
      RECT  8890.0 44472.5 8955.0 44537.5 ;
      RECT  8820.0 44200.0 8922.5 44265.0 ;
      RECT  8890.0 44232.5 8955.0 44505.0 ;
      RECT  8922.5 44472.5 9025.0 44537.5 ;
      RECT  14177.5 44200.0 14242.5 44265.0 ;
      RECT  14177.5 44687.5 14242.5 44752.5 ;
      RECT  11315.0 44200.0 14210.0 44265.0 ;
      RECT  14177.5 44232.5 14242.5 44720.0 ;
      RECT  14210.0 44687.5 17105.0 44752.5 ;
      RECT  8890.0 45455.0 8955.0 45520.0 ;
      RECT  8890.0 45182.5 8955.0 45247.5 ;
      RECT  8820.0 45455.0 8922.5 45520.0 ;
      RECT  8890.0 45215.0 8955.0 45487.5 ;
      RECT  8922.5 45182.5 9025.0 45247.5 ;
      RECT  14177.5 45455.0 14242.5 45520.0 ;
      RECT  14177.5 44967.5 14242.5 45032.5 ;
      RECT  11315.0 45455.0 14210.0 45520.0 ;
      RECT  14177.5 45000.0 14242.5 45487.5 ;
      RECT  14210.0 44967.5 17105.0 45032.5 ;
      RECT  8890.0 46890.0 8955.0 46955.0 ;
      RECT  8890.0 47162.5 8955.0 47227.5 ;
      RECT  8820.0 46890.0 8922.5 46955.0 ;
      RECT  8890.0 46922.5 8955.0 47195.0 ;
      RECT  8922.5 47162.5 9025.0 47227.5 ;
      RECT  14177.5 46890.0 14242.5 46955.0 ;
      RECT  14177.5 47377.5 14242.5 47442.5 ;
      RECT  11315.0 46890.0 14210.0 46955.0 ;
      RECT  14177.5 46922.5 14242.5 47410.0 ;
      RECT  14210.0 47377.5 17105.0 47442.5 ;
      RECT  8890.0 48145.0 8955.0 48210.0 ;
      RECT  8890.0 47872.5 8955.0 47937.5 ;
      RECT  8820.0 48145.0 8922.5 48210.0 ;
      RECT  8890.0 47905.0 8955.0 48177.5 ;
      RECT  8922.5 47872.5 9025.0 47937.5 ;
      RECT  14177.5 48145.0 14242.5 48210.0 ;
      RECT  14177.5 47657.5 14242.5 47722.5 ;
      RECT  11315.0 48145.0 14210.0 48210.0 ;
      RECT  14177.5 47690.0 14242.5 48177.5 ;
      RECT  14210.0 47657.5 17105.0 47722.5 ;
      RECT  8890.0 49580.0 8955.0 49645.0 ;
      RECT  8890.0 49852.5 8955.0 49917.5 ;
      RECT  8820.0 49580.0 8922.5 49645.0 ;
      RECT  8890.0 49612.5 8955.0 49885.0 ;
      RECT  8922.5 49852.5 9025.0 49917.5 ;
      RECT  14177.5 49580.0 14242.5 49645.0 ;
      RECT  14177.5 50067.5 14242.5 50132.5 ;
      RECT  11315.0 49580.0 14210.0 49645.0 ;
      RECT  14177.5 49612.5 14242.5 50100.0 ;
      RECT  14210.0 50067.5 17105.0 50132.5 ;
      RECT  8890.0 50835.0 8955.0 50900.0 ;
      RECT  8890.0 50562.5 8955.0 50627.5 ;
      RECT  8820.0 50835.0 8922.5 50900.0 ;
      RECT  8890.0 50595.0 8955.0 50867.5 ;
      RECT  8922.5 50562.5 9025.0 50627.5 ;
      RECT  14177.5 50835.0 14242.5 50900.0 ;
      RECT  14177.5 50347.5 14242.5 50412.5 ;
      RECT  11315.0 50835.0 14210.0 50900.0 ;
      RECT  14177.5 50380.0 14242.5 50867.5 ;
      RECT  14210.0 50347.5 17105.0 50412.5 ;
      RECT  8890.0 52270.0 8955.0 52335.0 ;
      RECT  8890.0 52542.5 8955.0 52607.5 ;
      RECT  8820.0 52270.0 8922.5 52335.0 ;
      RECT  8890.0 52302.5 8955.0 52575.0 ;
      RECT  8922.5 52542.5 9025.0 52607.5 ;
      RECT  14177.5 52270.0 14242.5 52335.0 ;
      RECT  14177.5 52757.5 14242.5 52822.5 ;
      RECT  11315.0 52270.0 14210.0 52335.0 ;
      RECT  14177.5 52302.5 14242.5 52790.0 ;
      RECT  14210.0 52757.5 17105.0 52822.5 ;
      RECT  8890.0 53525.0 8955.0 53590.0 ;
      RECT  8890.0 53252.5 8955.0 53317.5 ;
      RECT  8820.0 53525.0 8922.5 53590.0 ;
      RECT  8890.0 53285.0 8955.0 53557.5 ;
      RECT  8922.5 53252.5 9025.0 53317.5 ;
      RECT  14177.5 53525.0 14242.5 53590.0 ;
      RECT  14177.5 53037.5 14242.5 53102.5 ;
      RECT  11315.0 53525.0 14210.0 53590.0 ;
      RECT  14177.5 53070.0 14242.5 53557.5 ;
      RECT  14210.0 53037.5 17105.0 53102.5 ;
      RECT  8890.0 54960.0 8955.0 55025.0 ;
      RECT  8890.0 55232.5 8955.0 55297.5 ;
      RECT  8820.0 54960.0 8922.5 55025.0 ;
      RECT  8890.0 54992.5 8955.0 55265.0 ;
      RECT  8922.5 55232.5 9025.0 55297.5 ;
      RECT  14177.5 54960.0 14242.5 55025.0 ;
      RECT  14177.5 55447.5 14242.5 55512.5 ;
      RECT  11315.0 54960.0 14210.0 55025.0 ;
      RECT  14177.5 54992.5 14242.5 55480.0 ;
      RECT  14210.0 55447.5 17105.0 55512.5 ;
      RECT  8890.0 56215.0 8955.0 56280.0 ;
      RECT  8890.0 55942.5 8955.0 56007.5 ;
      RECT  8820.0 56215.0 8922.5 56280.0 ;
      RECT  8890.0 55975.0 8955.0 56247.5 ;
      RECT  8922.5 55942.5 9025.0 56007.5 ;
      RECT  14177.5 56215.0 14242.5 56280.0 ;
      RECT  14177.5 55727.5 14242.5 55792.5 ;
      RECT  11315.0 56215.0 14210.0 56280.0 ;
      RECT  14177.5 55760.0 14242.5 56247.5 ;
      RECT  14210.0 55727.5 17105.0 55792.5 ;
      RECT  8890.0 57650.0 8955.0 57715.0 ;
      RECT  8890.0 57922.5 8955.0 57987.5 ;
      RECT  8820.0 57650.0 8922.5 57715.0 ;
      RECT  8890.0 57682.5 8955.0 57955.0 ;
      RECT  8922.5 57922.5 9025.0 57987.5 ;
      RECT  14177.5 57650.0 14242.5 57715.0 ;
      RECT  14177.5 58137.5 14242.5 58202.5 ;
      RECT  11315.0 57650.0 14210.0 57715.0 ;
      RECT  14177.5 57682.5 14242.5 58170.0 ;
      RECT  14210.0 58137.5 17105.0 58202.5 ;
      RECT  8890.0 58905.0 8955.0 58970.0 ;
      RECT  8890.0 58632.5 8955.0 58697.5 ;
      RECT  8820.0 58905.0 8922.5 58970.0 ;
      RECT  8890.0 58665.0 8955.0 58937.5 ;
      RECT  8922.5 58632.5 9025.0 58697.5 ;
      RECT  14177.5 58905.0 14242.5 58970.0 ;
      RECT  14177.5 58417.5 14242.5 58482.5 ;
      RECT  11315.0 58905.0 14210.0 58970.0 ;
      RECT  14177.5 58450.0 14242.5 58937.5 ;
      RECT  14210.0 58417.5 17105.0 58482.5 ;
      RECT  8890.0 60340.0 8955.0 60405.0 ;
      RECT  8890.0 60612.5 8955.0 60677.5 ;
      RECT  8820.0 60340.0 8922.5 60405.0 ;
      RECT  8890.0 60372.5 8955.0 60645.0 ;
      RECT  8922.5 60612.5 9025.0 60677.5 ;
      RECT  14177.5 60340.0 14242.5 60405.0 ;
      RECT  14177.5 60827.5 14242.5 60892.5 ;
      RECT  11315.0 60340.0 14210.0 60405.0 ;
      RECT  14177.5 60372.5 14242.5 60860.0 ;
      RECT  14210.0 60827.5 17105.0 60892.5 ;
      RECT  8890.0 61595.0 8955.0 61660.0 ;
      RECT  8890.0 61322.5 8955.0 61387.5 ;
      RECT  8820.0 61595.0 8922.5 61660.0 ;
      RECT  8890.0 61355.0 8955.0 61627.5 ;
      RECT  8922.5 61322.5 9025.0 61387.5 ;
      RECT  14177.5 61595.0 14242.5 61660.0 ;
      RECT  14177.5 61107.5 14242.5 61172.5 ;
      RECT  11315.0 61595.0 14210.0 61660.0 ;
      RECT  14177.5 61140.0 14242.5 61627.5 ;
      RECT  14210.0 61107.5 17105.0 61172.5 ;
      RECT  8890.0 63030.0 8955.0 63095.0 ;
      RECT  8890.0 63302.5 8955.0 63367.5 ;
      RECT  8820.0 63030.0 8922.5 63095.0 ;
      RECT  8890.0 63062.5 8955.0 63335.0 ;
      RECT  8922.5 63302.5 9025.0 63367.5 ;
      RECT  14177.5 63030.0 14242.5 63095.0 ;
      RECT  14177.5 63517.5 14242.5 63582.5 ;
      RECT  11315.0 63030.0 14210.0 63095.0 ;
      RECT  14177.5 63062.5 14242.5 63550.0 ;
      RECT  14210.0 63517.5 17105.0 63582.5 ;
      RECT  8890.0 64285.0 8955.0 64350.0 ;
      RECT  8890.0 64012.5 8955.0 64077.5 ;
      RECT  8820.0 64285.0 8922.5 64350.0 ;
      RECT  8890.0 64045.0 8955.0 64317.5 ;
      RECT  8922.5 64012.5 9025.0 64077.5 ;
      RECT  14177.5 64285.0 14242.5 64350.0 ;
      RECT  14177.5 63797.5 14242.5 63862.5 ;
      RECT  11315.0 64285.0 14210.0 64350.0 ;
      RECT  14177.5 63830.0 14242.5 64317.5 ;
      RECT  14210.0 63797.5 17105.0 63862.5 ;
      RECT  8890.0 65720.0 8955.0 65785.0 ;
      RECT  8890.0 65992.5 8955.0 66057.5 ;
      RECT  8820.0 65720.0 8922.5 65785.0 ;
      RECT  8890.0 65752.5 8955.0 66025.0 ;
      RECT  8922.5 65992.5 9025.0 66057.5 ;
      RECT  14177.5 65720.0 14242.5 65785.0 ;
      RECT  14177.5 66207.5 14242.5 66272.5 ;
      RECT  11315.0 65720.0 14210.0 65785.0 ;
      RECT  14177.5 65752.5 14242.5 66240.0 ;
      RECT  14210.0 66207.5 17105.0 66272.5 ;
      RECT  8890.0 66975.0 8955.0 67040.0 ;
      RECT  8890.0 66702.5 8955.0 66767.5 ;
      RECT  8820.0 66975.0 8922.5 67040.0 ;
      RECT  8890.0 66735.0 8955.0 67007.5 ;
      RECT  8922.5 66702.5 9025.0 66767.5 ;
      RECT  14177.5 66975.0 14242.5 67040.0 ;
      RECT  14177.5 66487.5 14242.5 66552.5 ;
      RECT  11315.0 66975.0 14210.0 67040.0 ;
      RECT  14177.5 66520.0 14242.5 67007.5 ;
      RECT  14210.0 66487.5 17105.0 66552.5 ;
      RECT  8890.0 68410.0 8955.0 68475.0 ;
      RECT  8890.0 68682.5 8955.0 68747.5 ;
      RECT  8820.0 68410.0 8922.5 68475.0 ;
      RECT  8890.0 68442.5 8955.0 68715.0 ;
      RECT  8922.5 68682.5 9025.0 68747.5 ;
      RECT  14177.5 68410.0 14242.5 68475.0 ;
      RECT  14177.5 68897.5 14242.5 68962.5 ;
      RECT  11315.0 68410.0 14210.0 68475.0 ;
      RECT  14177.5 68442.5 14242.5 68930.0 ;
      RECT  14210.0 68897.5 17105.0 68962.5 ;
      RECT  8890.0 69665.0 8955.0 69730.0 ;
      RECT  8890.0 69392.5 8955.0 69457.5 ;
      RECT  8820.0 69665.0 8922.5 69730.0 ;
      RECT  8890.0 69425.0 8955.0 69697.5 ;
      RECT  8922.5 69392.5 9025.0 69457.5 ;
      RECT  14177.5 69665.0 14242.5 69730.0 ;
      RECT  14177.5 69177.5 14242.5 69242.5 ;
      RECT  11315.0 69665.0 14210.0 69730.0 ;
      RECT  14177.5 69210.0 14242.5 69697.5 ;
      RECT  14210.0 69177.5 17105.0 69242.5 ;
      RECT  8890.0 71100.0 8955.0 71165.0 ;
      RECT  8890.0 71372.5 8955.0 71437.5 ;
      RECT  8820.0 71100.0 8922.5 71165.0 ;
      RECT  8890.0 71132.5 8955.0 71405.0 ;
      RECT  8922.5 71372.5 9025.0 71437.5 ;
      RECT  14177.5 71100.0 14242.5 71165.0 ;
      RECT  14177.5 71587.5 14242.5 71652.5 ;
      RECT  11315.0 71100.0 14210.0 71165.0 ;
      RECT  14177.5 71132.5 14242.5 71620.0 ;
      RECT  14210.0 71587.5 17105.0 71652.5 ;
      RECT  8890.0 72355.0 8955.0 72420.0 ;
      RECT  8890.0 72082.5 8955.0 72147.5 ;
      RECT  8820.0 72355.0 8922.5 72420.0 ;
      RECT  8890.0 72115.0 8955.0 72387.5 ;
      RECT  8922.5 72082.5 9025.0 72147.5 ;
      RECT  14177.5 72355.0 14242.5 72420.0 ;
      RECT  14177.5 71867.5 14242.5 71932.5 ;
      RECT  11315.0 72355.0 14210.0 72420.0 ;
      RECT  14177.5 71900.0 14242.5 72387.5 ;
      RECT  14210.0 71867.5 17105.0 71932.5 ;
      RECT  8890.0 73790.0 8955.0 73855.0 ;
      RECT  8890.0 74062.5 8955.0 74127.5 ;
      RECT  8820.0 73790.0 8922.5 73855.0 ;
      RECT  8890.0 73822.5 8955.0 74095.0 ;
      RECT  8922.5 74062.5 9025.0 74127.5 ;
      RECT  14177.5 73790.0 14242.5 73855.0 ;
      RECT  14177.5 74277.5 14242.5 74342.5 ;
      RECT  11315.0 73790.0 14210.0 73855.0 ;
      RECT  14177.5 73822.5 14242.5 74310.0 ;
      RECT  14210.0 74277.5 17105.0 74342.5 ;
      RECT  8890.0 75045.0 8955.0 75110.0 ;
      RECT  8890.0 74772.5 8955.0 74837.5 ;
      RECT  8820.0 75045.0 8922.5 75110.0 ;
      RECT  8890.0 74805.0 8955.0 75077.5 ;
      RECT  8922.5 74772.5 9025.0 74837.5 ;
      RECT  14177.5 75045.0 14242.5 75110.0 ;
      RECT  14177.5 74557.5 14242.5 74622.5 ;
      RECT  11315.0 75045.0 14210.0 75110.0 ;
      RECT  14177.5 74590.0 14242.5 75077.5 ;
      RECT  14210.0 74557.5 17105.0 74622.5 ;
      RECT  8890.0 76480.0 8955.0 76545.0 ;
      RECT  8890.0 76752.5 8955.0 76817.5 ;
      RECT  8820.0 76480.0 8922.5 76545.0 ;
      RECT  8890.0 76512.5 8955.0 76785.0 ;
      RECT  8922.5 76752.5 9025.0 76817.5 ;
      RECT  14177.5 76480.0 14242.5 76545.0 ;
      RECT  14177.5 76967.5 14242.5 77032.5 ;
      RECT  11315.0 76480.0 14210.0 76545.0 ;
      RECT  14177.5 76512.5 14242.5 77000.0 ;
      RECT  14210.0 76967.5 17105.0 77032.5 ;
      RECT  8890.0 77735.0 8955.0 77800.0 ;
      RECT  8890.0 77462.5 8955.0 77527.5 ;
      RECT  8820.0 77735.0 8922.5 77800.0 ;
      RECT  8890.0 77495.0 8955.0 77767.5 ;
      RECT  8922.5 77462.5 9025.0 77527.5 ;
      RECT  14177.5 77735.0 14242.5 77800.0 ;
      RECT  14177.5 77247.5 14242.5 77312.5 ;
      RECT  11315.0 77735.0 14210.0 77800.0 ;
      RECT  14177.5 77280.0 14242.5 77767.5 ;
      RECT  14210.0 77247.5 17105.0 77312.5 ;
      RECT  8890.0 79170.0 8955.0 79235.0 ;
      RECT  8890.0 79442.5 8955.0 79507.5 ;
      RECT  8820.0 79170.0 8922.5 79235.0 ;
      RECT  8890.0 79202.5 8955.0 79475.0 ;
      RECT  8922.5 79442.5 9025.0 79507.5 ;
      RECT  14177.5 79170.0 14242.5 79235.0 ;
      RECT  14177.5 79657.5 14242.5 79722.5 ;
      RECT  11315.0 79170.0 14210.0 79235.0 ;
      RECT  14177.5 79202.5 14242.5 79690.0 ;
      RECT  14210.0 79657.5 17105.0 79722.5 ;
      RECT  8890.0 80425.0 8955.0 80490.0 ;
      RECT  8890.0 80152.5 8955.0 80217.5 ;
      RECT  8820.0 80425.0 8922.5 80490.0 ;
      RECT  8890.0 80185.0 8955.0 80457.5 ;
      RECT  8922.5 80152.5 9025.0 80217.5 ;
      RECT  14177.5 80425.0 14242.5 80490.0 ;
      RECT  14177.5 79937.5 14242.5 80002.5 ;
      RECT  11315.0 80425.0 14210.0 80490.0 ;
      RECT  14177.5 79970.0 14242.5 80457.5 ;
      RECT  14210.0 79937.5 17105.0 80002.5 ;
      RECT  8890.0 81860.0 8955.0 81925.0 ;
      RECT  8890.0 82132.5 8955.0 82197.5 ;
      RECT  8820.0 81860.0 8922.5 81925.0 ;
      RECT  8890.0 81892.5 8955.0 82165.0 ;
      RECT  8922.5 82132.5 9025.0 82197.5 ;
      RECT  14177.5 81860.0 14242.5 81925.0 ;
      RECT  14177.5 82347.5 14242.5 82412.5 ;
      RECT  11315.0 81860.0 14210.0 81925.0 ;
      RECT  14177.5 81892.5 14242.5 82380.0 ;
      RECT  14210.0 82347.5 17105.0 82412.5 ;
      RECT  8890.0 83115.0 8955.0 83180.0 ;
      RECT  8890.0 82842.5 8955.0 82907.5 ;
      RECT  8820.0 83115.0 8922.5 83180.0 ;
      RECT  8890.0 82875.0 8955.0 83147.5 ;
      RECT  8922.5 82842.5 9025.0 82907.5 ;
      RECT  14177.5 83115.0 14242.5 83180.0 ;
      RECT  14177.5 82627.5 14242.5 82692.5 ;
      RECT  11315.0 83115.0 14210.0 83180.0 ;
      RECT  14177.5 82660.0 14242.5 83147.5 ;
      RECT  14210.0 82627.5 17105.0 82692.5 ;
      RECT  8890.0 84550.0 8955.0 84615.0 ;
      RECT  8890.0 84822.5 8955.0 84887.5 ;
      RECT  8820.0 84550.0 8922.5 84615.0 ;
      RECT  8890.0 84582.5 8955.0 84855.0 ;
      RECT  8922.5 84822.5 9025.0 84887.5 ;
      RECT  14177.5 84550.0 14242.5 84615.0 ;
      RECT  14177.5 85037.5 14242.5 85102.5 ;
      RECT  11315.0 84550.0 14210.0 84615.0 ;
      RECT  14177.5 84582.5 14242.5 85070.0 ;
      RECT  14210.0 85037.5 17105.0 85102.5 ;
      RECT  8890.0 85805.0 8955.0 85870.0 ;
      RECT  8890.0 85532.5 8955.0 85597.5 ;
      RECT  8820.0 85805.0 8922.5 85870.0 ;
      RECT  8890.0 85565.0 8955.0 85837.5 ;
      RECT  8922.5 85532.5 9025.0 85597.5 ;
      RECT  14177.5 85805.0 14242.5 85870.0 ;
      RECT  14177.5 85317.5 14242.5 85382.5 ;
      RECT  11315.0 85805.0 14210.0 85870.0 ;
      RECT  14177.5 85350.0 14242.5 85837.5 ;
      RECT  14210.0 85317.5 17105.0 85382.5 ;
      RECT  8890.0 87240.0 8955.0 87305.0 ;
      RECT  8890.0 87512.5 8955.0 87577.5 ;
      RECT  8820.0 87240.0 8922.5 87305.0 ;
      RECT  8890.0 87272.5 8955.0 87545.0 ;
      RECT  8922.5 87512.5 9025.0 87577.5 ;
      RECT  14177.5 87240.0 14242.5 87305.0 ;
      RECT  14177.5 87727.5 14242.5 87792.5 ;
      RECT  11315.0 87240.0 14210.0 87305.0 ;
      RECT  14177.5 87272.5 14242.5 87760.0 ;
      RECT  14210.0 87727.5 17105.0 87792.5 ;
      RECT  8890.0 88495.0 8955.0 88560.0 ;
      RECT  8890.0 88222.5 8955.0 88287.5 ;
      RECT  8820.0 88495.0 8922.5 88560.0 ;
      RECT  8890.0 88255.0 8955.0 88527.5 ;
      RECT  8922.5 88222.5 9025.0 88287.5 ;
      RECT  14177.5 88495.0 14242.5 88560.0 ;
      RECT  14177.5 88007.5 14242.5 88072.5 ;
      RECT  11315.0 88495.0 14210.0 88560.0 ;
      RECT  14177.5 88040.0 14242.5 88527.5 ;
      RECT  14210.0 88007.5 17105.0 88072.5 ;
      RECT  8890.0 89930.0 8955.0 89995.0 ;
      RECT  8890.0 90202.5 8955.0 90267.5 ;
      RECT  8820.0 89930.0 8922.5 89995.0 ;
      RECT  8890.0 89962.5 8955.0 90235.0 ;
      RECT  8922.5 90202.5 9025.0 90267.5 ;
      RECT  14177.5 89930.0 14242.5 89995.0 ;
      RECT  14177.5 90417.5 14242.5 90482.5 ;
      RECT  11315.0 89930.0 14210.0 89995.0 ;
      RECT  14177.5 89962.5 14242.5 90450.0 ;
      RECT  14210.0 90417.5 17105.0 90482.5 ;
      RECT  8890.0 91185.0 8955.0 91250.0 ;
      RECT  8890.0 90912.5 8955.0 90977.5 ;
      RECT  8820.0 91185.0 8922.5 91250.0 ;
      RECT  8890.0 90945.0 8955.0 91217.5 ;
      RECT  8922.5 90912.5 9025.0 90977.5 ;
      RECT  14177.5 91185.0 14242.5 91250.0 ;
      RECT  14177.5 90697.5 14242.5 90762.5 ;
      RECT  11315.0 91185.0 14210.0 91250.0 ;
      RECT  14177.5 90730.0 14242.5 91217.5 ;
      RECT  14210.0 90697.5 17105.0 90762.5 ;
      RECT  8890.0 92620.0 8955.0 92685.0 ;
      RECT  8890.0 92892.5 8955.0 92957.5 ;
      RECT  8820.0 92620.0 8922.5 92685.0 ;
      RECT  8890.0 92652.5 8955.0 92925.0 ;
      RECT  8922.5 92892.5 9025.0 92957.5 ;
      RECT  14177.5 92620.0 14242.5 92685.0 ;
      RECT  14177.5 93107.5 14242.5 93172.5 ;
      RECT  11315.0 92620.0 14210.0 92685.0 ;
      RECT  14177.5 92652.5 14242.5 93140.0 ;
      RECT  14210.0 93107.5 17105.0 93172.5 ;
      RECT  8890.0 93875.0 8955.0 93940.0 ;
      RECT  8890.0 93602.5 8955.0 93667.5 ;
      RECT  8820.0 93875.0 8922.5 93940.0 ;
      RECT  8890.0 93635.0 8955.0 93907.5 ;
      RECT  8922.5 93602.5 9025.0 93667.5 ;
      RECT  14177.5 93875.0 14242.5 93940.0 ;
      RECT  14177.5 93387.5 14242.5 93452.5 ;
      RECT  11315.0 93875.0 14210.0 93940.0 ;
      RECT  14177.5 93420.0 14242.5 93907.5 ;
      RECT  14210.0 93387.5 17105.0 93452.5 ;
      RECT  8890.0 95310.0 8955.0 95375.0 ;
      RECT  8890.0 95582.5 8955.0 95647.5 ;
      RECT  8820.0 95310.0 8922.5 95375.0 ;
      RECT  8890.0 95342.5 8955.0 95615.0 ;
      RECT  8922.5 95582.5 9025.0 95647.5 ;
      RECT  14177.5 95310.0 14242.5 95375.0 ;
      RECT  14177.5 95797.5 14242.5 95862.5 ;
      RECT  11315.0 95310.0 14210.0 95375.0 ;
      RECT  14177.5 95342.5 14242.5 95830.0 ;
      RECT  14210.0 95797.5 17105.0 95862.5 ;
      RECT  8890.0 96565.0 8955.0 96630.0 ;
      RECT  8890.0 96292.5 8955.0 96357.5 ;
      RECT  8820.0 96565.0 8922.5 96630.0 ;
      RECT  8890.0 96325.0 8955.0 96597.5 ;
      RECT  8922.5 96292.5 9025.0 96357.5 ;
      RECT  14177.5 96565.0 14242.5 96630.0 ;
      RECT  14177.5 96077.5 14242.5 96142.5 ;
      RECT  11315.0 96565.0 14210.0 96630.0 ;
      RECT  14177.5 96110.0 14242.5 96597.5 ;
      RECT  14210.0 96077.5 17105.0 96142.5 ;
      RECT  8890.0 98000.0 8955.0 98065.0 ;
      RECT  8890.0 98272.5 8955.0 98337.5 ;
      RECT  8820.0 98000.0 8922.5 98065.0 ;
      RECT  8890.0 98032.5 8955.0 98305.0 ;
      RECT  8922.5 98272.5 9025.0 98337.5 ;
      RECT  14177.5 98000.0 14242.5 98065.0 ;
      RECT  14177.5 98487.5 14242.5 98552.5 ;
      RECT  11315.0 98000.0 14210.0 98065.0 ;
      RECT  14177.5 98032.5 14242.5 98520.0 ;
      RECT  14210.0 98487.5 17105.0 98552.5 ;
      RECT  8890.0 99255.0 8955.0 99320.0 ;
      RECT  8890.0 98982.5 8955.0 99047.5 ;
      RECT  8820.0 99255.0 8922.5 99320.0 ;
      RECT  8890.0 99015.0 8955.0 99287.5 ;
      RECT  8922.5 98982.5 9025.0 99047.5 ;
      RECT  14177.5 99255.0 14242.5 99320.0 ;
      RECT  14177.5 98767.5 14242.5 98832.5 ;
      RECT  11315.0 99255.0 14210.0 99320.0 ;
      RECT  14177.5 98800.0 14242.5 99287.5 ;
      RECT  14210.0 98767.5 17105.0 98832.5 ;
      RECT  8890.0 100690.0 8955.0 100755.0 ;
      RECT  8890.0 100962.5 8955.0 101027.5 ;
      RECT  8820.0 100690.0 8922.5 100755.0 ;
      RECT  8890.0 100722.5 8955.0 100995.0 ;
      RECT  8922.5 100962.5 9025.0 101027.5 ;
      RECT  14177.5 100690.0 14242.5 100755.0 ;
      RECT  14177.5 101177.5 14242.5 101242.5 ;
      RECT  11315.0 100690.0 14210.0 100755.0 ;
      RECT  14177.5 100722.5 14242.5 101210.0 ;
      RECT  14210.0 101177.5 17105.0 101242.5 ;
      RECT  8890.0 101945.0 8955.0 102010.0 ;
      RECT  8890.0 101672.5 8955.0 101737.5 ;
      RECT  8820.0 101945.0 8922.5 102010.0 ;
      RECT  8890.0 101705.0 8955.0 101977.5 ;
      RECT  8922.5 101672.5 9025.0 101737.5 ;
      RECT  14177.5 101945.0 14242.5 102010.0 ;
      RECT  14177.5 101457.5 14242.5 101522.5 ;
      RECT  11315.0 101945.0 14210.0 102010.0 ;
      RECT  14177.5 101490.0 14242.5 101977.5 ;
      RECT  14210.0 101457.5 17105.0 101522.5 ;
      RECT  8890.0 103380.0 8955.0 103445.0 ;
      RECT  8890.0 103652.5 8955.0 103717.5 ;
      RECT  8820.0 103380.0 8922.5 103445.0 ;
      RECT  8890.0 103412.5 8955.0 103685.0 ;
      RECT  8922.5 103652.5 9025.0 103717.5 ;
      RECT  14177.5 103380.0 14242.5 103445.0 ;
      RECT  14177.5 103867.5 14242.5 103932.5 ;
      RECT  11315.0 103380.0 14210.0 103445.0 ;
      RECT  14177.5 103412.5 14242.5 103900.0 ;
      RECT  14210.0 103867.5 17105.0 103932.5 ;
      RECT  8890.0 104635.0 8955.0 104700.0 ;
      RECT  8890.0 104362.5 8955.0 104427.5 ;
      RECT  8820.0 104635.0 8922.5 104700.0 ;
      RECT  8890.0 104395.0 8955.0 104667.5 ;
      RECT  8922.5 104362.5 9025.0 104427.5 ;
      RECT  14177.5 104635.0 14242.5 104700.0 ;
      RECT  14177.5 104147.5 14242.5 104212.5 ;
      RECT  11315.0 104635.0 14210.0 104700.0 ;
      RECT  14177.5 104180.0 14242.5 104667.5 ;
      RECT  14210.0 104147.5 17105.0 104212.5 ;
      RECT  8890.0 106070.0 8955.0 106135.0 ;
      RECT  8890.0 106342.5 8955.0 106407.5 ;
      RECT  8820.0 106070.0 8922.5 106135.0 ;
      RECT  8890.0 106102.5 8955.0 106375.0 ;
      RECT  8922.5 106342.5 9025.0 106407.5 ;
      RECT  14177.5 106070.0 14242.5 106135.0 ;
      RECT  14177.5 106557.5 14242.5 106622.5 ;
      RECT  11315.0 106070.0 14210.0 106135.0 ;
      RECT  14177.5 106102.5 14242.5 106590.0 ;
      RECT  14210.0 106557.5 17105.0 106622.5 ;
      RECT  8890.0 107325.0 8955.0 107390.0 ;
      RECT  8890.0 107052.5 8955.0 107117.5 ;
      RECT  8820.0 107325.0 8922.5 107390.0 ;
      RECT  8890.0 107085.0 8955.0 107357.5 ;
      RECT  8922.5 107052.5 9025.0 107117.5 ;
      RECT  14177.5 107325.0 14242.5 107390.0 ;
      RECT  14177.5 106837.5 14242.5 106902.5 ;
      RECT  11315.0 107325.0 14210.0 107390.0 ;
      RECT  14177.5 106870.0 14242.5 107357.5 ;
      RECT  14210.0 106837.5 17105.0 106902.5 ;
      RECT  8890.0 108760.0 8955.0 108825.0 ;
      RECT  8890.0 109032.5 8955.0 109097.5 ;
      RECT  8820.0 108760.0 8922.5 108825.0 ;
      RECT  8890.0 108792.5 8955.0 109065.0 ;
      RECT  8922.5 109032.5 9025.0 109097.5 ;
      RECT  14177.5 108760.0 14242.5 108825.0 ;
      RECT  14177.5 109247.5 14242.5 109312.5 ;
      RECT  11315.0 108760.0 14210.0 108825.0 ;
      RECT  14177.5 108792.5 14242.5 109280.0 ;
      RECT  14210.0 109247.5 17105.0 109312.5 ;
      RECT  8890.0 110015.0 8955.0 110080.0 ;
      RECT  8890.0 109742.5 8955.0 109807.5 ;
      RECT  8820.0 110015.0 8922.5 110080.0 ;
      RECT  8890.0 109775.0 8955.0 110047.5 ;
      RECT  8922.5 109742.5 9025.0 109807.5 ;
      RECT  14177.5 110015.0 14242.5 110080.0 ;
      RECT  14177.5 109527.5 14242.5 109592.5 ;
      RECT  11315.0 110015.0 14210.0 110080.0 ;
      RECT  14177.5 109560.0 14242.5 110047.5 ;
      RECT  14210.0 109527.5 17105.0 109592.5 ;
      RECT  8890.0 111450.0 8955.0 111515.0 ;
      RECT  8890.0 111722.5 8955.0 111787.5 ;
      RECT  8820.0 111450.0 8922.5 111515.0 ;
      RECT  8890.0 111482.5 8955.0 111755.0 ;
      RECT  8922.5 111722.5 9025.0 111787.5 ;
      RECT  14177.5 111450.0 14242.5 111515.0 ;
      RECT  14177.5 111937.5 14242.5 112002.5 ;
      RECT  11315.0 111450.0 14210.0 111515.0 ;
      RECT  14177.5 111482.5 14242.5 111970.0 ;
      RECT  14210.0 111937.5 17105.0 112002.5 ;
      RECT  8890.0 112705.0 8955.0 112770.0 ;
      RECT  8890.0 112432.5 8955.0 112497.5 ;
      RECT  8820.0 112705.0 8922.5 112770.0 ;
      RECT  8890.0 112465.0 8955.0 112737.5 ;
      RECT  8922.5 112432.5 9025.0 112497.5 ;
      RECT  14177.5 112705.0 14242.5 112770.0 ;
      RECT  14177.5 112217.5 14242.5 112282.5 ;
      RECT  11315.0 112705.0 14210.0 112770.0 ;
      RECT  14177.5 112250.0 14242.5 112737.5 ;
      RECT  14210.0 112217.5 17105.0 112282.5 ;
      RECT  8890.0 114140.0 8955.0 114205.0 ;
      RECT  8890.0 114412.5 8955.0 114477.5 ;
      RECT  8820.0 114140.0 8922.5 114205.0 ;
      RECT  8890.0 114172.5 8955.0 114445.0 ;
      RECT  8922.5 114412.5 9025.0 114477.5 ;
      RECT  14177.5 114140.0 14242.5 114205.0 ;
      RECT  14177.5 114627.5 14242.5 114692.5 ;
      RECT  11315.0 114140.0 14210.0 114205.0 ;
      RECT  14177.5 114172.5 14242.5 114660.0 ;
      RECT  14210.0 114627.5 17105.0 114692.5 ;
      RECT  8890.0 115395.0 8955.0 115460.0 ;
      RECT  8890.0 115122.5 8955.0 115187.5 ;
      RECT  8820.0 115395.0 8922.5 115460.0 ;
      RECT  8890.0 115155.0 8955.0 115427.5 ;
      RECT  8922.5 115122.5 9025.0 115187.5 ;
      RECT  14177.5 115395.0 14242.5 115460.0 ;
      RECT  14177.5 114907.5 14242.5 114972.5 ;
      RECT  11315.0 115395.0 14210.0 115460.0 ;
      RECT  14177.5 114940.0 14242.5 115427.5 ;
      RECT  14210.0 114907.5 17105.0 114972.5 ;
      RECT  8890.0 116830.0 8955.0 116895.0 ;
      RECT  8890.0 117102.5 8955.0 117167.5 ;
      RECT  8820.0 116830.0 8922.5 116895.0 ;
      RECT  8890.0 116862.5 8955.0 117135.0 ;
      RECT  8922.5 117102.5 9025.0 117167.5 ;
      RECT  14177.5 116830.0 14242.5 116895.0 ;
      RECT  14177.5 117317.5 14242.5 117382.5 ;
      RECT  11315.0 116830.0 14210.0 116895.0 ;
      RECT  14177.5 116862.5 14242.5 117350.0 ;
      RECT  14210.0 117317.5 17105.0 117382.5 ;
      RECT  8890.0 118085.0 8955.0 118150.0 ;
      RECT  8890.0 117812.5 8955.0 117877.5 ;
      RECT  8820.0 118085.0 8922.5 118150.0 ;
      RECT  8890.0 117845.0 8955.0 118117.5 ;
      RECT  8922.5 117812.5 9025.0 117877.5 ;
      RECT  14177.5 118085.0 14242.5 118150.0 ;
      RECT  14177.5 117597.5 14242.5 117662.5 ;
      RECT  11315.0 118085.0 14210.0 118150.0 ;
      RECT  14177.5 117630.0 14242.5 118117.5 ;
      RECT  14210.0 117597.5 17105.0 117662.5 ;
      RECT  8890.0 119520.0 8955.0 119585.0 ;
      RECT  8890.0 119792.5 8955.0 119857.5 ;
      RECT  8820.0 119520.0 8922.5 119585.0 ;
      RECT  8890.0 119552.5 8955.0 119825.0 ;
      RECT  8922.5 119792.5 9025.0 119857.5 ;
      RECT  14177.5 119520.0 14242.5 119585.0 ;
      RECT  14177.5 120007.5 14242.5 120072.5 ;
      RECT  11315.0 119520.0 14210.0 119585.0 ;
      RECT  14177.5 119552.5 14242.5 120040.0 ;
      RECT  14210.0 120007.5 17105.0 120072.5 ;
      RECT  8890.0 120775.0 8955.0 120840.0 ;
      RECT  8890.0 120502.5 8955.0 120567.5 ;
      RECT  8820.0 120775.0 8922.5 120840.0 ;
      RECT  8890.0 120535.0 8955.0 120807.5 ;
      RECT  8922.5 120502.5 9025.0 120567.5 ;
      RECT  14177.5 120775.0 14242.5 120840.0 ;
      RECT  14177.5 120287.5 14242.5 120352.5 ;
      RECT  11315.0 120775.0 14210.0 120840.0 ;
      RECT  14177.5 120320.0 14242.5 120807.5 ;
      RECT  14210.0 120287.5 17105.0 120352.5 ;
      RECT  8890.0 122210.0 8955.0 122275.0 ;
      RECT  8890.0 122482.5 8955.0 122547.5 ;
      RECT  8820.0 122210.0 8922.5 122275.0 ;
      RECT  8890.0 122242.5 8955.0 122515.0 ;
      RECT  8922.5 122482.5 9025.0 122547.5 ;
      RECT  14177.5 122210.0 14242.5 122275.0 ;
      RECT  14177.5 122697.5 14242.5 122762.5 ;
      RECT  11315.0 122210.0 14210.0 122275.0 ;
      RECT  14177.5 122242.5 14242.5 122730.0 ;
      RECT  14210.0 122697.5 17105.0 122762.5 ;
      RECT  8890.0 123465.0 8955.0 123530.0 ;
      RECT  8890.0 123192.5 8955.0 123257.5 ;
      RECT  8820.0 123465.0 8922.5 123530.0 ;
      RECT  8890.0 123225.0 8955.0 123497.5 ;
      RECT  8922.5 123192.5 9025.0 123257.5 ;
      RECT  14177.5 123465.0 14242.5 123530.0 ;
      RECT  14177.5 122977.5 14242.5 123042.5 ;
      RECT  11315.0 123465.0 14210.0 123530.0 ;
      RECT  14177.5 123010.0 14242.5 123497.5 ;
      RECT  14210.0 122977.5 17105.0 123042.5 ;
      RECT  8890.0 124900.0 8955.0 124965.0 ;
      RECT  8890.0 125172.5 8955.0 125237.5 ;
      RECT  8820.0 124900.0 8922.5 124965.0 ;
      RECT  8890.0 124932.5 8955.0 125205.0 ;
      RECT  8922.5 125172.5 9025.0 125237.5 ;
      RECT  14177.5 124900.0 14242.5 124965.0 ;
      RECT  14177.5 125387.5 14242.5 125452.5 ;
      RECT  11315.0 124900.0 14210.0 124965.0 ;
      RECT  14177.5 124932.5 14242.5 125420.0 ;
      RECT  14210.0 125387.5 17105.0 125452.5 ;
      RECT  8890.0 126155.0 8955.0 126220.0 ;
      RECT  8890.0 125882.5 8955.0 125947.5 ;
      RECT  8820.0 126155.0 8922.5 126220.0 ;
      RECT  8890.0 125915.0 8955.0 126187.5 ;
      RECT  8922.5 125882.5 9025.0 125947.5 ;
      RECT  14177.5 126155.0 14242.5 126220.0 ;
      RECT  14177.5 125667.5 14242.5 125732.5 ;
      RECT  11315.0 126155.0 14210.0 126220.0 ;
      RECT  14177.5 125700.0 14242.5 126187.5 ;
      RECT  14210.0 125667.5 17105.0 125732.5 ;
      RECT  8890.0 127590.0 8955.0 127655.0 ;
      RECT  8890.0 127862.5 8955.0 127927.5 ;
      RECT  8820.0 127590.0 8922.5 127655.0 ;
      RECT  8890.0 127622.5 8955.0 127895.0 ;
      RECT  8922.5 127862.5 9025.0 127927.5 ;
      RECT  14177.5 127590.0 14242.5 127655.0 ;
      RECT  14177.5 128077.5 14242.5 128142.5 ;
      RECT  11315.0 127590.0 14210.0 127655.0 ;
      RECT  14177.5 127622.5 14242.5 128110.0 ;
      RECT  14210.0 128077.5 17105.0 128142.5 ;
      RECT  8890.0 128845.0 8955.0 128910.0 ;
      RECT  8890.0 128572.5 8955.0 128637.5 ;
      RECT  8820.0 128845.0 8922.5 128910.0 ;
      RECT  8890.0 128605.0 8955.0 128877.5 ;
      RECT  8922.5 128572.5 9025.0 128637.5 ;
      RECT  14177.5 128845.0 14242.5 128910.0 ;
      RECT  14177.5 128357.5 14242.5 128422.5 ;
      RECT  11315.0 128845.0 14210.0 128910.0 ;
      RECT  14177.5 128390.0 14242.5 128877.5 ;
      RECT  14210.0 128357.5 17105.0 128422.5 ;
      RECT  8890.0 130280.0 8955.0 130345.0 ;
      RECT  8890.0 130552.5 8955.0 130617.5 ;
      RECT  8820.0 130280.0 8922.5 130345.0 ;
      RECT  8890.0 130312.5 8955.0 130585.0 ;
      RECT  8922.5 130552.5 9025.0 130617.5 ;
      RECT  14177.5 130280.0 14242.5 130345.0 ;
      RECT  14177.5 130767.5 14242.5 130832.5 ;
      RECT  11315.0 130280.0 14210.0 130345.0 ;
      RECT  14177.5 130312.5 14242.5 130800.0 ;
      RECT  14210.0 130767.5 17105.0 130832.5 ;
      RECT  8890.0 131535.0 8955.0 131600.0 ;
      RECT  8890.0 131262.5 8955.0 131327.5 ;
      RECT  8820.0 131535.0 8922.5 131600.0 ;
      RECT  8890.0 131295.0 8955.0 131567.5 ;
      RECT  8922.5 131262.5 9025.0 131327.5 ;
      RECT  14177.5 131535.0 14242.5 131600.0 ;
      RECT  14177.5 131047.5 14242.5 131112.5 ;
      RECT  11315.0 131535.0 14210.0 131600.0 ;
      RECT  14177.5 131080.0 14242.5 131567.5 ;
      RECT  14210.0 131047.5 17105.0 131112.5 ;
      RECT  8890.0 132970.0 8955.0 133035.0 ;
      RECT  8890.0 133242.5 8955.0 133307.5 ;
      RECT  8820.0 132970.0 8922.5 133035.0 ;
      RECT  8890.0 133002.5 8955.0 133275.0 ;
      RECT  8922.5 133242.5 9025.0 133307.5 ;
      RECT  14177.5 132970.0 14242.5 133035.0 ;
      RECT  14177.5 133457.5 14242.5 133522.5 ;
      RECT  11315.0 132970.0 14210.0 133035.0 ;
      RECT  14177.5 133002.5 14242.5 133490.0 ;
      RECT  14210.0 133457.5 17105.0 133522.5 ;
      RECT  8890.0 134225.0 8955.0 134290.0 ;
      RECT  8890.0 133952.5 8955.0 134017.5 ;
      RECT  8820.0 134225.0 8922.5 134290.0 ;
      RECT  8890.0 133985.0 8955.0 134257.5 ;
      RECT  8922.5 133952.5 9025.0 134017.5 ;
      RECT  14177.5 134225.0 14242.5 134290.0 ;
      RECT  14177.5 133737.5 14242.5 133802.5 ;
      RECT  11315.0 134225.0 14210.0 134290.0 ;
      RECT  14177.5 133770.0 14242.5 134257.5 ;
      RECT  14210.0 133737.5 17105.0 133802.5 ;
      RECT  8890.0 135660.0 8955.0 135725.0 ;
      RECT  8890.0 135932.5 8955.0 135997.5 ;
      RECT  8820.0 135660.0 8922.5 135725.0 ;
      RECT  8890.0 135692.5 8955.0 135965.0 ;
      RECT  8922.5 135932.5 9025.0 135997.5 ;
      RECT  14177.5 135660.0 14242.5 135725.0 ;
      RECT  14177.5 136147.5 14242.5 136212.5 ;
      RECT  11315.0 135660.0 14210.0 135725.0 ;
      RECT  14177.5 135692.5 14242.5 136180.0 ;
      RECT  14210.0 136147.5 17105.0 136212.5 ;
      RECT  8890.0 136915.0 8955.0 136980.0 ;
      RECT  8890.0 136642.5 8955.0 136707.5 ;
      RECT  8820.0 136915.0 8922.5 136980.0 ;
      RECT  8890.0 136675.0 8955.0 136947.5 ;
      RECT  8922.5 136642.5 9025.0 136707.5 ;
      RECT  14177.5 136915.0 14242.5 136980.0 ;
      RECT  14177.5 136427.5 14242.5 136492.5 ;
      RECT  11315.0 136915.0 14210.0 136980.0 ;
      RECT  14177.5 136460.0 14242.5 136947.5 ;
      RECT  14210.0 136427.5 17105.0 136492.5 ;
      RECT  8890.0 138350.0 8955.0 138415.0 ;
      RECT  8890.0 138622.5 8955.0 138687.5 ;
      RECT  8820.0 138350.0 8922.5 138415.0 ;
      RECT  8890.0 138382.5 8955.0 138655.0 ;
      RECT  8922.5 138622.5 9025.0 138687.5 ;
      RECT  14177.5 138350.0 14242.5 138415.0 ;
      RECT  14177.5 138837.5 14242.5 138902.5 ;
      RECT  11315.0 138350.0 14210.0 138415.0 ;
      RECT  14177.5 138382.5 14242.5 138870.0 ;
      RECT  14210.0 138837.5 17105.0 138902.5 ;
      RECT  8890.0 139605.0 8955.0 139670.0 ;
      RECT  8890.0 139332.5 8955.0 139397.5 ;
      RECT  8820.0 139605.0 8922.5 139670.0 ;
      RECT  8890.0 139365.0 8955.0 139637.5 ;
      RECT  8922.5 139332.5 9025.0 139397.5 ;
      RECT  14177.5 139605.0 14242.5 139670.0 ;
      RECT  14177.5 139117.5 14242.5 139182.5 ;
      RECT  11315.0 139605.0 14210.0 139670.0 ;
      RECT  14177.5 139150.0 14242.5 139637.5 ;
      RECT  14210.0 139117.5 17105.0 139182.5 ;
      RECT  8890.0 141040.0 8955.0 141105.0 ;
      RECT  8890.0 141312.5 8955.0 141377.5 ;
      RECT  8820.0 141040.0 8922.5 141105.0 ;
      RECT  8890.0 141072.5 8955.0 141345.0 ;
      RECT  8922.5 141312.5 9025.0 141377.5 ;
      RECT  14177.5 141040.0 14242.5 141105.0 ;
      RECT  14177.5 141527.5 14242.5 141592.5 ;
      RECT  11315.0 141040.0 14210.0 141105.0 ;
      RECT  14177.5 141072.5 14242.5 141560.0 ;
      RECT  14210.0 141527.5 17105.0 141592.5 ;
      RECT  8890.0 142295.0 8955.0 142360.0 ;
      RECT  8890.0 142022.5 8955.0 142087.5 ;
      RECT  8820.0 142295.0 8922.5 142360.0 ;
      RECT  8890.0 142055.0 8955.0 142327.5 ;
      RECT  8922.5 142022.5 9025.0 142087.5 ;
      RECT  14177.5 142295.0 14242.5 142360.0 ;
      RECT  14177.5 141807.5 14242.5 141872.5 ;
      RECT  11315.0 142295.0 14210.0 142360.0 ;
      RECT  14177.5 141840.0 14242.5 142327.5 ;
      RECT  14210.0 141807.5 17105.0 141872.5 ;
      RECT  8890.0 143730.0 8955.0 143795.0 ;
      RECT  8890.0 144002.5 8955.0 144067.5 ;
      RECT  8820.0 143730.0 8922.5 143795.0 ;
      RECT  8890.0 143762.5 8955.0 144035.0 ;
      RECT  8922.5 144002.5 9025.0 144067.5 ;
      RECT  14177.5 143730.0 14242.5 143795.0 ;
      RECT  14177.5 144217.5 14242.5 144282.5 ;
      RECT  11315.0 143730.0 14210.0 143795.0 ;
      RECT  14177.5 143762.5 14242.5 144250.0 ;
      RECT  14210.0 144217.5 17105.0 144282.5 ;
      RECT  8890.0 144985.0 8955.0 145050.0 ;
      RECT  8890.0 144712.5 8955.0 144777.5 ;
      RECT  8820.0 144985.0 8922.5 145050.0 ;
      RECT  8890.0 144745.0 8955.0 145017.5 ;
      RECT  8922.5 144712.5 9025.0 144777.5 ;
      RECT  14177.5 144985.0 14242.5 145050.0 ;
      RECT  14177.5 144497.5 14242.5 144562.5 ;
      RECT  11315.0 144985.0 14210.0 145050.0 ;
      RECT  14177.5 144530.0 14242.5 145017.5 ;
      RECT  14210.0 144497.5 17105.0 144562.5 ;
      RECT  8890.0 146420.0 8955.0 146485.0 ;
      RECT  8890.0 146692.5 8955.0 146757.5 ;
      RECT  8820.0 146420.0 8922.5 146485.0 ;
      RECT  8890.0 146452.5 8955.0 146725.0 ;
      RECT  8922.5 146692.5 9025.0 146757.5 ;
      RECT  14177.5 146420.0 14242.5 146485.0 ;
      RECT  14177.5 146907.5 14242.5 146972.5 ;
      RECT  11315.0 146420.0 14210.0 146485.0 ;
      RECT  14177.5 146452.5 14242.5 146940.0 ;
      RECT  14210.0 146907.5 17105.0 146972.5 ;
      RECT  8890.0 147675.0 8955.0 147740.0 ;
      RECT  8890.0 147402.5 8955.0 147467.5 ;
      RECT  8820.0 147675.0 8922.5 147740.0 ;
      RECT  8890.0 147435.0 8955.0 147707.5 ;
      RECT  8922.5 147402.5 9025.0 147467.5 ;
      RECT  14177.5 147675.0 14242.5 147740.0 ;
      RECT  14177.5 147187.5 14242.5 147252.5 ;
      RECT  11315.0 147675.0 14210.0 147740.0 ;
      RECT  14177.5 147220.0 14242.5 147707.5 ;
      RECT  14210.0 147187.5 17105.0 147252.5 ;
      RECT  8890.0 149110.0 8955.0 149175.0 ;
      RECT  8890.0 149382.5 8955.0 149447.5 ;
      RECT  8820.0 149110.0 8922.5 149175.0 ;
      RECT  8890.0 149142.5 8955.0 149415.0 ;
      RECT  8922.5 149382.5 9025.0 149447.5 ;
      RECT  14177.5 149110.0 14242.5 149175.0 ;
      RECT  14177.5 149597.5 14242.5 149662.5 ;
      RECT  11315.0 149110.0 14210.0 149175.0 ;
      RECT  14177.5 149142.5 14242.5 149630.0 ;
      RECT  14210.0 149597.5 17105.0 149662.5 ;
      RECT  8890.0 150365.0 8955.0 150430.0 ;
      RECT  8890.0 150092.5 8955.0 150157.5 ;
      RECT  8820.0 150365.0 8922.5 150430.0 ;
      RECT  8890.0 150125.0 8955.0 150397.5 ;
      RECT  8922.5 150092.5 9025.0 150157.5 ;
      RECT  14177.5 150365.0 14242.5 150430.0 ;
      RECT  14177.5 149877.5 14242.5 149942.5 ;
      RECT  11315.0 150365.0 14210.0 150430.0 ;
      RECT  14177.5 149910.0 14242.5 150397.5 ;
      RECT  14210.0 149877.5 17105.0 149942.5 ;
      RECT  8890.0 151800.0 8955.0 151865.0 ;
      RECT  8890.0 152072.5 8955.0 152137.5 ;
      RECT  8820.0 151800.0 8922.5 151865.0 ;
      RECT  8890.0 151832.5 8955.0 152105.0 ;
      RECT  8922.5 152072.5 9025.0 152137.5 ;
      RECT  14177.5 151800.0 14242.5 151865.0 ;
      RECT  14177.5 152287.5 14242.5 152352.5 ;
      RECT  11315.0 151800.0 14210.0 151865.0 ;
      RECT  14177.5 151832.5 14242.5 152320.0 ;
      RECT  14210.0 152287.5 17105.0 152352.5 ;
      RECT  8890.0 153055.0 8955.0 153120.0 ;
      RECT  8890.0 152782.5 8955.0 152847.5 ;
      RECT  8820.0 153055.0 8922.5 153120.0 ;
      RECT  8890.0 152815.0 8955.0 153087.5 ;
      RECT  8922.5 152782.5 9025.0 152847.5 ;
      RECT  14177.5 153055.0 14242.5 153120.0 ;
      RECT  14177.5 152567.5 14242.5 152632.5 ;
      RECT  11315.0 153055.0 14210.0 153120.0 ;
      RECT  14177.5 152600.0 14242.5 153087.5 ;
      RECT  14210.0 152567.5 17105.0 152632.5 ;
      RECT  8890.0 154490.0 8955.0 154555.0 ;
      RECT  8890.0 154762.5 8955.0 154827.5 ;
      RECT  8820.0 154490.0 8922.5 154555.0 ;
      RECT  8890.0 154522.5 8955.0 154795.0 ;
      RECT  8922.5 154762.5 9025.0 154827.5 ;
      RECT  14177.5 154490.0 14242.5 154555.0 ;
      RECT  14177.5 154977.5 14242.5 155042.5 ;
      RECT  11315.0 154490.0 14210.0 154555.0 ;
      RECT  14177.5 154522.5 14242.5 155010.0 ;
      RECT  14210.0 154977.5 17105.0 155042.5 ;
      RECT  8890.0 155745.0 8955.0 155810.0 ;
      RECT  8890.0 155472.5 8955.0 155537.5 ;
      RECT  8820.0 155745.0 8922.5 155810.0 ;
      RECT  8890.0 155505.0 8955.0 155777.5 ;
      RECT  8922.5 155472.5 9025.0 155537.5 ;
      RECT  14177.5 155745.0 14242.5 155810.0 ;
      RECT  14177.5 155257.5 14242.5 155322.5 ;
      RECT  11315.0 155745.0 14210.0 155810.0 ;
      RECT  14177.5 155290.0 14242.5 155777.5 ;
      RECT  14210.0 155257.5 17105.0 155322.5 ;
      RECT  8890.0 157180.0 8955.0 157245.0 ;
      RECT  8890.0 157452.5 8955.0 157517.5 ;
      RECT  8820.0 157180.0 8922.5 157245.0 ;
      RECT  8890.0 157212.5 8955.0 157485.0 ;
      RECT  8922.5 157452.5 9025.0 157517.5 ;
      RECT  14177.5 157180.0 14242.5 157245.0 ;
      RECT  14177.5 157667.5 14242.5 157732.5 ;
      RECT  11315.0 157180.0 14210.0 157245.0 ;
      RECT  14177.5 157212.5 14242.5 157700.0 ;
      RECT  14210.0 157667.5 17105.0 157732.5 ;
      RECT  8890.0 158435.0 8955.0 158500.0 ;
      RECT  8890.0 158162.5 8955.0 158227.5 ;
      RECT  8820.0 158435.0 8922.5 158500.0 ;
      RECT  8890.0 158195.0 8955.0 158467.5 ;
      RECT  8922.5 158162.5 9025.0 158227.5 ;
      RECT  14177.5 158435.0 14242.5 158500.0 ;
      RECT  14177.5 157947.5 14242.5 158012.5 ;
      RECT  11315.0 158435.0 14210.0 158500.0 ;
      RECT  14177.5 157980.0 14242.5 158467.5 ;
      RECT  14210.0 157947.5 17105.0 158012.5 ;
      RECT  8890.0 159870.0 8955.0 159935.0 ;
      RECT  8890.0 160142.5 8955.0 160207.5 ;
      RECT  8820.0 159870.0 8922.5 159935.0 ;
      RECT  8890.0 159902.5 8955.0 160175.0 ;
      RECT  8922.5 160142.5 9025.0 160207.5 ;
      RECT  14177.5 159870.0 14242.5 159935.0 ;
      RECT  14177.5 160357.5 14242.5 160422.5 ;
      RECT  11315.0 159870.0 14210.0 159935.0 ;
      RECT  14177.5 159902.5 14242.5 160390.0 ;
      RECT  14210.0 160357.5 17105.0 160422.5 ;
      RECT  8890.0 161125.0 8955.0 161190.0 ;
      RECT  8890.0 160852.5 8955.0 160917.5 ;
      RECT  8820.0 161125.0 8922.5 161190.0 ;
      RECT  8890.0 160885.0 8955.0 161157.5 ;
      RECT  8922.5 160852.5 9025.0 160917.5 ;
      RECT  14177.5 161125.0 14242.5 161190.0 ;
      RECT  14177.5 160637.5 14242.5 160702.5 ;
      RECT  11315.0 161125.0 14210.0 161190.0 ;
      RECT  14177.5 160670.0 14242.5 161157.5 ;
      RECT  14210.0 160637.5 17105.0 160702.5 ;
      RECT  8890.0 162560.0 8955.0 162625.0 ;
      RECT  8890.0 162832.5 8955.0 162897.5 ;
      RECT  8820.0 162560.0 8922.5 162625.0 ;
      RECT  8890.0 162592.5 8955.0 162865.0 ;
      RECT  8922.5 162832.5 9025.0 162897.5 ;
      RECT  14177.5 162560.0 14242.5 162625.0 ;
      RECT  14177.5 163047.5 14242.5 163112.5 ;
      RECT  11315.0 162560.0 14210.0 162625.0 ;
      RECT  14177.5 162592.5 14242.5 163080.0 ;
      RECT  14210.0 163047.5 17105.0 163112.5 ;
      RECT  8890.0 163815.0 8955.0 163880.0 ;
      RECT  8890.0 163542.5 8955.0 163607.5 ;
      RECT  8820.0 163815.0 8922.5 163880.0 ;
      RECT  8890.0 163575.0 8955.0 163847.5 ;
      RECT  8922.5 163542.5 9025.0 163607.5 ;
      RECT  14177.5 163815.0 14242.5 163880.0 ;
      RECT  14177.5 163327.5 14242.5 163392.5 ;
      RECT  11315.0 163815.0 14210.0 163880.0 ;
      RECT  14177.5 163360.0 14242.5 163847.5 ;
      RECT  14210.0 163327.5 17105.0 163392.5 ;
      RECT  8890.0 165250.0 8955.0 165315.0 ;
      RECT  8890.0 165522.5 8955.0 165587.5 ;
      RECT  8820.0 165250.0 8922.5 165315.0 ;
      RECT  8890.0 165282.5 8955.0 165555.0 ;
      RECT  8922.5 165522.5 9025.0 165587.5 ;
      RECT  14177.5 165250.0 14242.5 165315.0 ;
      RECT  14177.5 165737.5 14242.5 165802.5 ;
      RECT  11315.0 165250.0 14210.0 165315.0 ;
      RECT  14177.5 165282.5 14242.5 165770.0 ;
      RECT  14210.0 165737.5 17105.0 165802.5 ;
      RECT  8890.0 166505.0 8955.0 166570.0 ;
      RECT  8890.0 166232.5 8955.0 166297.5 ;
      RECT  8820.0 166505.0 8922.5 166570.0 ;
      RECT  8890.0 166265.0 8955.0 166537.5 ;
      RECT  8922.5 166232.5 9025.0 166297.5 ;
      RECT  14177.5 166505.0 14242.5 166570.0 ;
      RECT  14177.5 166017.5 14242.5 166082.5 ;
      RECT  11315.0 166505.0 14210.0 166570.0 ;
      RECT  14177.5 166050.0 14242.5 166537.5 ;
      RECT  14210.0 166017.5 17105.0 166082.5 ;
      RECT  8890.0 167940.0 8955.0 168005.0 ;
      RECT  8890.0 168212.5 8955.0 168277.5 ;
      RECT  8820.0 167940.0 8922.5 168005.0 ;
      RECT  8890.0 167972.5 8955.0 168245.0 ;
      RECT  8922.5 168212.5 9025.0 168277.5 ;
      RECT  14177.5 167940.0 14242.5 168005.0 ;
      RECT  14177.5 168427.5 14242.5 168492.5 ;
      RECT  11315.0 167940.0 14210.0 168005.0 ;
      RECT  14177.5 167972.5 14242.5 168460.0 ;
      RECT  14210.0 168427.5 17105.0 168492.5 ;
      RECT  8890.0 169195.0 8955.0 169260.0 ;
      RECT  8890.0 168922.5 8955.0 168987.5 ;
      RECT  8820.0 169195.0 8922.5 169260.0 ;
      RECT  8890.0 168955.0 8955.0 169227.5 ;
      RECT  8922.5 168922.5 9025.0 168987.5 ;
      RECT  14177.5 169195.0 14242.5 169260.0 ;
      RECT  14177.5 168707.5 14242.5 168772.5 ;
      RECT  11315.0 169195.0 14210.0 169260.0 ;
      RECT  14177.5 168740.0 14242.5 169227.5 ;
      RECT  14210.0 168707.5 17105.0 168772.5 ;
      RECT  8890.0 170630.0 8955.0 170695.0 ;
      RECT  8890.0 170902.5 8955.0 170967.5 ;
      RECT  8820.0 170630.0 8922.5 170695.0 ;
      RECT  8890.0 170662.5 8955.0 170935.0 ;
      RECT  8922.5 170902.5 9025.0 170967.5 ;
      RECT  14177.5 170630.0 14242.5 170695.0 ;
      RECT  14177.5 171117.5 14242.5 171182.5 ;
      RECT  11315.0 170630.0 14210.0 170695.0 ;
      RECT  14177.5 170662.5 14242.5 171150.0 ;
      RECT  14210.0 171117.5 17105.0 171182.5 ;
      RECT  8890.0 171885.0 8955.0 171950.0 ;
      RECT  8890.0 171612.5 8955.0 171677.5 ;
      RECT  8820.0 171885.0 8922.5 171950.0 ;
      RECT  8890.0 171645.0 8955.0 171917.5 ;
      RECT  8922.5 171612.5 9025.0 171677.5 ;
      RECT  14177.5 171885.0 14242.5 171950.0 ;
      RECT  14177.5 171397.5 14242.5 171462.5 ;
      RECT  11315.0 171885.0 14210.0 171950.0 ;
      RECT  14177.5 171430.0 14242.5 171917.5 ;
      RECT  14210.0 171397.5 17105.0 171462.5 ;
      RECT  8890.0 173320.0 8955.0 173385.0 ;
      RECT  8890.0 173592.5 8955.0 173657.5 ;
      RECT  8820.0 173320.0 8922.5 173385.0 ;
      RECT  8890.0 173352.5 8955.0 173625.0 ;
      RECT  8922.5 173592.5 9025.0 173657.5 ;
      RECT  14177.5 173320.0 14242.5 173385.0 ;
      RECT  14177.5 173807.5 14242.5 173872.5 ;
      RECT  11315.0 173320.0 14210.0 173385.0 ;
      RECT  14177.5 173352.5 14242.5 173840.0 ;
      RECT  14210.0 173807.5 17105.0 173872.5 ;
      RECT  8890.0 174575.0 8955.0 174640.0 ;
      RECT  8890.0 174302.5 8955.0 174367.5 ;
      RECT  8820.0 174575.0 8922.5 174640.0 ;
      RECT  8890.0 174335.0 8955.0 174607.5 ;
      RECT  8922.5 174302.5 9025.0 174367.5 ;
      RECT  14177.5 174575.0 14242.5 174640.0 ;
      RECT  14177.5 174087.5 14242.5 174152.5 ;
      RECT  11315.0 174575.0 14210.0 174640.0 ;
      RECT  14177.5 174120.0 14242.5 174607.5 ;
      RECT  14210.0 174087.5 17105.0 174152.5 ;
      RECT  8890.0 176010.0 8955.0 176075.0 ;
      RECT  8890.0 176282.5 8955.0 176347.5 ;
      RECT  8820.0 176010.0 8922.5 176075.0 ;
      RECT  8890.0 176042.5 8955.0 176315.0 ;
      RECT  8922.5 176282.5 9025.0 176347.5 ;
      RECT  14177.5 176010.0 14242.5 176075.0 ;
      RECT  14177.5 176497.5 14242.5 176562.5 ;
      RECT  11315.0 176010.0 14210.0 176075.0 ;
      RECT  14177.5 176042.5 14242.5 176530.0 ;
      RECT  14210.0 176497.5 17105.0 176562.5 ;
      RECT  8890.0 177265.0 8955.0 177330.0 ;
      RECT  8890.0 176992.5 8955.0 177057.5 ;
      RECT  8820.0 177265.0 8922.5 177330.0 ;
      RECT  8890.0 177025.0 8955.0 177297.5 ;
      RECT  8922.5 176992.5 9025.0 177057.5 ;
      RECT  14177.5 177265.0 14242.5 177330.0 ;
      RECT  14177.5 176777.5 14242.5 176842.5 ;
      RECT  11315.0 177265.0 14210.0 177330.0 ;
      RECT  14177.5 176810.0 14242.5 177297.5 ;
      RECT  14210.0 176777.5 17105.0 176842.5 ;
      RECT  8890.0 178700.0 8955.0 178765.0 ;
      RECT  8890.0 178972.5 8955.0 179037.5 ;
      RECT  8820.0 178700.0 8922.5 178765.0 ;
      RECT  8890.0 178732.5 8955.0 179005.0 ;
      RECT  8922.5 178972.5 9025.0 179037.5 ;
      RECT  14177.5 178700.0 14242.5 178765.0 ;
      RECT  14177.5 179187.5 14242.5 179252.5 ;
      RECT  11315.0 178700.0 14210.0 178765.0 ;
      RECT  14177.5 178732.5 14242.5 179220.0 ;
      RECT  14210.0 179187.5 17105.0 179252.5 ;
      RECT  8890.0 179955.0 8955.0 180020.0 ;
      RECT  8890.0 179682.5 8955.0 179747.5 ;
      RECT  8820.0 179955.0 8922.5 180020.0 ;
      RECT  8890.0 179715.0 8955.0 179987.5 ;
      RECT  8922.5 179682.5 9025.0 179747.5 ;
      RECT  14177.5 179955.0 14242.5 180020.0 ;
      RECT  14177.5 179467.5 14242.5 179532.5 ;
      RECT  11315.0 179955.0 14210.0 180020.0 ;
      RECT  14177.5 179500.0 14242.5 179987.5 ;
      RECT  14210.0 179467.5 17105.0 179532.5 ;
      RECT  8890.0 181390.0 8955.0 181455.0 ;
      RECT  8890.0 181662.5 8955.0 181727.5 ;
      RECT  8820.0 181390.0 8922.5 181455.0 ;
      RECT  8890.0 181422.5 8955.0 181695.0 ;
      RECT  8922.5 181662.5 9025.0 181727.5 ;
      RECT  14177.5 181390.0 14242.5 181455.0 ;
      RECT  14177.5 181877.5 14242.5 181942.5 ;
      RECT  11315.0 181390.0 14210.0 181455.0 ;
      RECT  14177.5 181422.5 14242.5 181910.0 ;
      RECT  14210.0 181877.5 17105.0 181942.5 ;
      RECT  8890.0 182645.0 8955.0 182710.0 ;
      RECT  8890.0 182372.5 8955.0 182437.5 ;
      RECT  8820.0 182645.0 8922.5 182710.0 ;
      RECT  8890.0 182405.0 8955.0 182677.5 ;
      RECT  8922.5 182372.5 9025.0 182437.5 ;
      RECT  14177.5 182645.0 14242.5 182710.0 ;
      RECT  14177.5 182157.5 14242.5 182222.5 ;
      RECT  11315.0 182645.0 14210.0 182710.0 ;
      RECT  14177.5 182190.0 14242.5 182677.5 ;
      RECT  14210.0 182157.5 17105.0 182222.5 ;
      RECT  8890.0 184080.0 8955.0 184145.0 ;
      RECT  8890.0 184352.5 8955.0 184417.5 ;
      RECT  8820.0 184080.0 8922.5 184145.0 ;
      RECT  8890.0 184112.5 8955.0 184385.0 ;
      RECT  8922.5 184352.5 9025.0 184417.5 ;
      RECT  14177.5 184080.0 14242.5 184145.0 ;
      RECT  14177.5 184567.5 14242.5 184632.5 ;
      RECT  11315.0 184080.0 14210.0 184145.0 ;
      RECT  14177.5 184112.5 14242.5 184600.0 ;
      RECT  14210.0 184567.5 17105.0 184632.5 ;
      RECT  8890.0 185335.0 8955.0 185400.0 ;
      RECT  8890.0 185062.5 8955.0 185127.5 ;
      RECT  8820.0 185335.0 8922.5 185400.0 ;
      RECT  8890.0 185095.0 8955.0 185367.5 ;
      RECT  8922.5 185062.5 9025.0 185127.5 ;
      RECT  14177.5 185335.0 14242.5 185400.0 ;
      RECT  14177.5 184847.5 14242.5 184912.5 ;
      RECT  11315.0 185335.0 14210.0 185400.0 ;
      RECT  14177.5 184880.0 14242.5 185367.5 ;
      RECT  14210.0 184847.5 17105.0 184912.5 ;
      RECT  8890.0 186770.0 8955.0 186835.0 ;
      RECT  8890.0 187042.5 8955.0 187107.5 ;
      RECT  8820.0 186770.0 8922.5 186835.0 ;
      RECT  8890.0 186802.5 8955.0 187075.0 ;
      RECT  8922.5 187042.5 9025.0 187107.5 ;
      RECT  14177.5 186770.0 14242.5 186835.0 ;
      RECT  14177.5 187257.5 14242.5 187322.5 ;
      RECT  11315.0 186770.0 14210.0 186835.0 ;
      RECT  14177.5 186802.5 14242.5 187290.0 ;
      RECT  14210.0 187257.5 17105.0 187322.5 ;
      RECT  8890.0 188025.0 8955.0 188090.0 ;
      RECT  8890.0 187752.5 8955.0 187817.5 ;
      RECT  8820.0 188025.0 8922.5 188090.0 ;
      RECT  8890.0 187785.0 8955.0 188057.5 ;
      RECT  8922.5 187752.5 9025.0 187817.5 ;
      RECT  14177.5 188025.0 14242.5 188090.0 ;
      RECT  14177.5 187537.5 14242.5 187602.5 ;
      RECT  11315.0 188025.0 14210.0 188090.0 ;
      RECT  14177.5 187570.0 14242.5 188057.5 ;
      RECT  14210.0 187537.5 17105.0 187602.5 ;
      RECT  8890.0 189460.0 8955.0 189525.0 ;
      RECT  8890.0 189732.5 8955.0 189797.5 ;
      RECT  8820.0 189460.0 8922.5 189525.0 ;
      RECT  8890.0 189492.5 8955.0 189765.0 ;
      RECT  8922.5 189732.5 9025.0 189797.5 ;
      RECT  14177.5 189460.0 14242.5 189525.0 ;
      RECT  14177.5 189947.5 14242.5 190012.5 ;
      RECT  11315.0 189460.0 14210.0 189525.0 ;
      RECT  14177.5 189492.5 14242.5 189980.0 ;
      RECT  14210.0 189947.5 17105.0 190012.5 ;
      RECT  8890.0 190715.0 8955.0 190780.0 ;
      RECT  8890.0 190442.5 8955.0 190507.5 ;
      RECT  8820.0 190715.0 8922.5 190780.0 ;
      RECT  8890.0 190475.0 8955.0 190747.5 ;
      RECT  8922.5 190442.5 9025.0 190507.5 ;
      RECT  14177.5 190715.0 14242.5 190780.0 ;
      RECT  14177.5 190227.5 14242.5 190292.5 ;
      RECT  11315.0 190715.0 14210.0 190780.0 ;
      RECT  14177.5 190260.0 14242.5 190747.5 ;
      RECT  14210.0 190227.5 17105.0 190292.5 ;
      RECT  8890.0 192150.0 8955.0 192215.0 ;
      RECT  8890.0 192422.5 8955.0 192487.5 ;
      RECT  8820.0 192150.0 8922.5 192215.0 ;
      RECT  8890.0 192182.5 8955.0 192455.0 ;
      RECT  8922.5 192422.5 9025.0 192487.5 ;
      RECT  14177.5 192150.0 14242.5 192215.0 ;
      RECT  14177.5 192637.5 14242.5 192702.5 ;
      RECT  11315.0 192150.0 14210.0 192215.0 ;
      RECT  14177.5 192182.5 14242.5 192670.0 ;
      RECT  14210.0 192637.5 17105.0 192702.5 ;
      RECT  8890.0 193405.0 8955.0 193470.0 ;
      RECT  8890.0 193132.5 8955.0 193197.5 ;
      RECT  8820.0 193405.0 8922.5 193470.0 ;
      RECT  8890.0 193165.0 8955.0 193437.5 ;
      RECT  8922.5 193132.5 9025.0 193197.5 ;
      RECT  14177.5 193405.0 14242.5 193470.0 ;
      RECT  14177.5 192917.5 14242.5 192982.5 ;
      RECT  11315.0 193405.0 14210.0 193470.0 ;
      RECT  14177.5 192950.0 14242.5 193437.5 ;
      RECT  14210.0 192917.5 17105.0 192982.5 ;
      RECT  8890.0 194840.0 8955.0 194905.0 ;
      RECT  8890.0 195112.5 8955.0 195177.5 ;
      RECT  8820.0 194840.0 8922.5 194905.0 ;
      RECT  8890.0 194872.5 8955.0 195145.0 ;
      RECT  8922.5 195112.5 9025.0 195177.5 ;
      RECT  14177.5 194840.0 14242.5 194905.0 ;
      RECT  14177.5 195327.5 14242.5 195392.5 ;
      RECT  11315.0 194840.0 14210.0 194905.0 ;
      RECT  14177.5 194872.5 14242.5 195360.0 ;
      RECT  14210.0 195327.5 17105.0 195392.5 ;
      RECT  8890.0 196095.0 8955.0 196160.0 ;
      RECT  8890.0 195822.5 8955.0 195887.5 ;
      RECT  8820.0 196095.0 8922.5 196160.0 ;
      RECT  8890.0 195855.0 8955.0 196127.5 ;
      RECT  8922.5 195822.5 9025.0 195887.5 ;
      RECT  14177.5 196095.0 14242.5 196160.0 ;
      RECT  14177.5 195607.5 14242.5 195672.5 ;
      RECT  11315.0 196095.0 14210.0 196160.0 ;
      RECT  14177.5 195640.0 14242.5 196127.5 ;
      RECT  14210.0 195607.5 17105.0 195672.5 ;
      RECT  8890.0 197530.0 8955.0 197595.0 ;
      RECT  8890.0 197802.5 8955.0 197867.5 ;
      RECT  8820.0 197530.0 8922.5 197595.0 ;
      RECT  8890.0 197562.5 8955.0 197835.0 ;
      RECT  8922.5 197802.5 9025.0 197867.5 ;
      RECT  14177.5 197530.0 14242.5 197595.0 ;
      RECT  14177.5 198017.5 14242.5 198082.5 ;
      RECT  11315.0 197530.0 14210.0 197595.0 ;
      RECT  14177.5 197562.5 14242.5 198050.0 ;
      RECT  14210.0 198017.5 17105.0 198082.5 ;
      RECT  8890.0 198785.0 8955.0 198850.0 ;
      RECT  8890.0 198512.5 8955.0 198577.5 ;
      RECT  8820.0 198785.0 8922.5 198850.0 ;
      RECT  8890.0 198545.0 8955.0 198817.5 ;
      RECT  8922.5 198512.5 9025.0 198577.5 ;
      RECT  14177.5 198785.0 14242.5 198850.0 ;
      RECT  14177.5 198297.5 14242.5 198362.5 ;
      RECT  11315.0 198785.0 14210.0 198850.0 ;
      RECT  14177.5 198330.0 14242.5 198817.5 ;
      RECT  14210.0 198297.5 17105.0 198362.5 ;
      RECT  8890.0 200220.0 8955.0 200285.0 ;
      RECT  8890.0 200492.5 8955.0 200557.5 ;
      RECT  8820.0 200220.0 8922.5 200285.0 ;
      RECT  8890.0 200252.5 8955.0 200525.0 ;
      RECT  8922.5 200492.5 9025.0 200557.5 ;
      RECT  14177.5 200220.0 14242.5 200285.0 ;
      RECT  14177.5 200707.5 14242.5 200772.5 ;
      RECT  11315.0 200220.0 14210.0 200285.0 ;
      RECT  14177.5 200252.5 14242.5 200740.0 ;
      RECT  14210.0 200707.5 17105.0 200772.5 ;
      RECT  8890.0 201475.0 8955.0 201540.0 ;
      RECT  8890.0 201202.5 8955.0 201267.5 ;
      RECT  8820.0 201475.0 8922.5 201540.0 ;
      RECT  8890.0 201235.0 8955.0 201507.5 ;
      RECT  8922.5 201202.5 9025.0 201267.5 ;
      RECT  14177.5 201475.0 14242.5 201540.0 ;
      RECT  14177.5 200987.5 14242.5 201052.5 ;
      RECT  11315.0 201475.0 14210.0 201540.0 ;
      RECT  14177.5 201020.0 14242.5 201507.5 ;
      RECT  14210.0 200987.5 17105.0 201052.5 ;
      RECT  8890.0 202910.0 8955.0 202975.0 ;
      RECT  8890.0 203182.5 8955.0 203247.5 ;
      RECT  8820.0 202910.0 8922.5 202975.0 ;
      RECT  8890.0 202942.5 8955.0 203215.0 ;
      RECT  8922.5 203182.5 9025.0 203247.5 ;
      RECT  14177.5 202910.0 14242.5 202975.0 ;
      RECT  14177.5 203397.5 14242.5 203462.5 ;
      RECT  11315.0 202910.0 14210.0 202975.0 ;
      RECT  14177.5 202942.5 14242.5 203430.0 ;
      RECT  14210.0 203397.5 17105.0 203462.5 ;
      RECT  8890.0 204165.0 8955.0 204230.0 ;
      RECT  8890.0 203892.5 8955.0 203957.5 ;
      RECT  8820.0 204165.0 8922.5 204230.0 ;
      RECT  8890.0 203925.0 8955.0 204197.5 ;
      RECT  8922.5 203892.5 9025.0 203957.5 ;
      RECT  14177.5 204165.0 14242.5 204230.0 ;
      RECT  14177.5 203677.5 14242.5 203742.5 ;
      RECT  11315.0 204165.0 14210.0 204230.0 ;
      RECT  14177.5 203710.0 14242.5 204197.5 ;
      RECT  14210.0 203677.5 17105.0 203742.5 ;
      RECT  8890.0 205600.0 8955.0 205665.0 ;
      RECT  8890.0 205872.5 8955.0 205937.5 ;
      RECT  8820.0 205600.0 8922.5 205665.0 ;
      RECT  8890.0 205632.5 8955.0 205905.0 ;
      RECT  8922.5 205872.5 9025.0 205937.5 ;
      RECT  14177.5 205600.0 14242.5 205665.0 ;
      RECT  14177.5 206087.5 14242.5 206152.5 ;
      RECT  11315.0 205600.0 14210.0 205665.0 ;
      RECT  14177.5 205632.5 14242.5 206120.0 ;
      RECT  14210.0 206087.5 17105.0 206152.5 ;
      RECT  9480.0 34067.5 17195.0 34132.5 ;
      RECT  9480.0 36757.5 17195.0 36822.5 ;
      RECT  9480.0 39447.5 17195.0 39512.5 ;
      RECT  9480.0 42137.5 17195.0 42202.5 ;
      RECT  9480.0 44827.5 17195.0 44892.5 ;
      RECT  9480.0 47517.5 17195.0 47582.5 ;
      RECT  9480.0 50207.5 17195.0 50272.5 ;
      RECT  9480.0 52897.5 17195.0 52962.5 ;
      RECT  9480.0 55587.5 17195.0 55652.5 ;
      RECT  9480.0 58277.5 17195.0 58342.5 ;
      RECT  9480.0 60967.5 17195.0 61032.5 ;
      RECT  9480.0 63657.5 17195.0 63722.5 ;
      RECT  9480.0 66347.5 17195.0 66412.5 ;
      RECT  9480.0 69037.5 17195.0 69102.5 ;
      RECT  9480.0 71727.5 17195.0 71792.5 ;
      RECT  9480.0 74417.5 17195.0 74482.5 ;
      RECT  9480.0 77107.5 17195.0 77172.5 ;
      RECT  9480.0 79797.5 17195.0 79862.5 ;
      RECT  9480.0 82487.5 17195.0 82552.5 ;
      RECT  9480.0 85177.5 17195.0 85242.5 ;
      RECT  9480.0 87867.5 17195.0 87932.5 ;
      RECT  9480.0 90557.5 17195.0 90622.5 ;
      RECT  9480.0 93247.5 17195.0 93312.5 ;
      RECT  9480.0 95937.5 17195.0 96002.5 ;
      RECT  9480.0 98627.5 17195.0 98692.5 ;
      RECT  9480.0 101317.5 17195.0 101382.5 ;
      RECT  9480.0 104007.5 17195.0 104072.5 ;
      RECT  9480.0 106697.5 17195.0 106762.5 ;
      RECT  9480.0 109387.5 17195.0 109452.5 ;
      RECT  9480.0 112077.5 17195.0 112142.5 ;
      RECT  9480.0 114767.5 17195.0 114832.5 ;
      RECT  9480.0 117457.5 17195.0 117522.5 ;
      RECT  9480.0 120147.5 17195.0 120212.5 ;
      RECT  9480.0 122837.5 17195.0 122902.5 ;
      RECT  9480.0 125527.5 17195.0 125592.5 ;
      RECT  9480.0 128217.5 17195.0 128282.5 ;
      RECT  9480.0 130907.5 17195.0 130972.5 ;
      RECT  9480.0 133597.5 17195.0 133662.5 ;
      RECT  9480.0 136287.5 17195.0 136352.5 ;
      RECT  9480.0 138977.5 17195.0 139042.5 ;
      RECT  9480.0 141667.5 17195.0 141732.5 ;
      RECT  9480.0 144357.5 17195.0 144422.5 ;
      RECT  9480.0 147047.5 17195.0 147112.5 ;
      RECT  9480.0 149737.5 17195.0 149802.5 ;
      RECT  9480.0 152427.5 17195.0 152492.5 ;
      RECT  9480.0 155117.5 17195.0 155182.5 ;
      RECT  9480.0 157807.5 17195.0 157872.5 ;
      RECT  9480.0 160497.5 17195.0 160562.5 ;
      RECT  9480.0 163187.5 17195.0 163252.5 ;
      RECT  9480.0 165877.5 17195.0 165942.5 ;
      RECT  9480.0 168567.5 17195.0 168632.5 ;
      RECT  9480.0 171257.5 17195.0 171322.5 ;
      RECT  9480.0 173947.5 17195.0 174012.5 ;
      RECT  9480.0 176637.5 17195.0 176702.5 ;
      RECT  9480.0 179327.5 17195.0 179392.5 ;
      RECT  9480.0 182017.5 17195.0 182082.5 ;
      RECT  9480.0 184707.5 17195.0 184772.5 ;
      RECT  9480.0 187397.5 17195.0 187462.5 ;
      RECT  9480.0 190087.5 17195.0 190152.5 ;
      RECT  9480.0 192777.5 17195.0 192842.5 ;
      RECT  9480.0 195467.5 17195.0 195532.5 ;
      RECT  9480.0 198157.5 17195.0 198222.5 ;
      RECT  9480.0 200847.5 17195.0 200912.5 ;
      RECT  9480.0 203537.5 17195.0 203602.5 ;
      RECT  9480.0 206227.5 17195.0 206292.5 ;
      RECT  4175.0 35412.5 107980.0 35477.5 ;
      RECT  4175.0 38102.5 107980.0 38167.5 ;
      RECT  4175.0 40792.5 107980.0 40857.5 ;
      RECT  4175.0 43482.5 107980.0 43547.5 ;
      RECT  4175.0 46172.5 107980.0 46237.5 ;
      RECT  4175.0 48862.5 107980.0 48927.5 ;
      RECT  4175.0 51552.5 107980.0 51617.5 ;
      RECT  4175.0 54242.5 107980.0 54307.5 ;
      RECT  4175.0 56932.5 107980.0 56997.5 ;
      RECT  4175.0 59622.5 107980.0 59687.5 ;
      RECT  4175.0 62312.5 107980.0 62377.5 ;
      RECT  4175.0 65002.5 107980.0 65067.5 ;
      RECT  4175.0 67692.5 107980.0 67757.5 ;
      RECT  4175.0 70382.5 107980.0 70447.5 ;
      RECT  4175.0 73072.5 107980.0 73137.5 ;
      RECT  4175.0 75762.5 107980.0 75827.5 ;
      RECT  4175.0 78452.5 107980.0 78517.5 ;
      RECT  4175.0 81142.5 107980.0 81207.5 ;
      RECT  4175.0 83832.5 107980.0 83897.5 ;
      RECT  4175.0 86522.5 107980.0 86587.5 ;
      RECT  4175.0 89212.5 107980.0 89277.5 ;
      RECT  4175.0 91902.5 107980.0 91967.5 ;
      RECT  4175.0 94592.5 107980.0 94657.5 ;
      RECT  4175.0 97282.5 107980.0 97347.5 ;
      RECT  4175.0 99972.5 107980.0 100037.5 ;
      RECT  4175.0 102662.5 107980.0 102727.5 ;
      RECT  4175.0 105352.5 107980.0 105417.5 ;
      RECT  4175.0 108042.5 107980.0 108107.5 ;
      RECT  4175.0 110732.5 107980.0 110797.5 ;
      RECT  4175.0 113422.5 107980.0 113487.5 ;
      RECT  4175.0 116112.5 107980.0 116177.5 ;
      RECT  4175.0 118802.5 107980.0 118867.5 ;
      RECT  4175.0 121492.5 107980.0 121557.5 ;
      RECT  4175.0 124182.5 107980.0 124247.5 ;
      RECT  4175.0 126872.5 107980.0 126937.5 ;
      RECT  4175.0 129562.5 107980.0 129627.5 ;
      RECT  4175.0 132252.5 107980.0 132317.5 ;
      RECT  4175.0 134942.5 107980.0 135007.5 ;
      RECT  4175.0 137632.5 107980.0 137697.5 ;
      RECT  4175.0 140322.5 107980.0 140387.5 ;
      RECT  4175.0 143012.5 107980.0 143077.5 ;
      RECT  4175.0 145702.5 107980.0 145767.5 ;
      RECT  4175.0 148392.5 107980.0 148457.5 ;
      RECT  4175.0 151082.5 107980.0 151147.5 ;
      RECT  4175.0 153772.5 107980.0 153837.5 ;
      RECT  4175.0 156462.5 107980.0 156527.5 ;
      RECT  4175.0 159152.5 107980.0 159217.5 ;
      RECT  4175.0 161842.5 107980.0 161907.5 ;
      RECT  4175.0 164532.5 107980.0 164597.5 ;
      RECT  4175.0 167222.5 107980.0 167287.5 ;
      RECT  4175.0 169912.5 107980.0 169977.5 ;
      RECT  4175.0 172602.5 107980.0 172667.5 ;
      RECT  4175.0 175292.5 107980.0 175357.5 ;
      RECT  4175.0 177982.5 107980.0 178047.5 ;
      RECT  4175.0 180672.5 107980.0 180737.5 ;
      RECT  4175.0 183362.5 107980.0 183427.5 ;
      RECT  4175.0 186052.5 107980.0 186117.5 ;
      RECT  4175.0 188742.5 107980.0 188807.5 ;
      RECT  4175.0 191432.5 107980.0 191497.5 ;
      RECT  4175.0 194122.5 107980.0 194187.5 ;
      RECT  4175.0 196812.5 107980.0 196877.5 ;
      RECT  4175.0 199502.5 107980.0 199567.5 ;
      RECT  4175.0 202192.5 107980.0 202257.5 ;
      RECT  4175.0 204882.5 107980.0 204947.5 ;
      RECT  11420.0 12752.5 12677.5 12817.5 ;
      RECT  11145.0 14097.5 12882.5 14162.5 ;
      RECT  11420.0 18132.5 13087.5 18197.5 ;
      RECT  11145.0 19477.5 13292.5 19542.5 ;
      RECT  12335.0 23512.5 13497.5 23577.5 ;
      RECT  12060.0 24857.5 13702.5 24922.5 ;
      RECT  11785.0 26202.5 13907.5 26267.5 ;
      RECT  12335.0 12547.5 12472.5 12612.5 ;
      RECT  12335.0 15237.5 12472.5 15302.5 ;
      RECT  12335.0 17927.5 12472.5 17992.5 ;
      RECT  12335.0 20617.5 12472.5 20682.5 ;
      RECT  12335.0 23307.5 12472.5 23372.5 ;
      RECT  12335.0 25997.5 12472.5 26062.5 ;
      RECT  12335.0 28687.5 12472.5 28752.5 ;
      RECT  12335.0 31377.5 12472.5 31442.5 ;
      RECT  4175.0 13892.5 12335.0 13957.5 ;
      RECT  4175.0 16582.5 12335.0 16647.5 ;
      RECT  4175.0 19272.5 12335.0 19337.5 ;
      RECT  4175.0 21962.5 12335.0 22027.5 ;
      RECT  4175.0 24652.5 12335.0 24717.5 ;
      RECT  4175.0 27342.5 12335.0 27407.5 ;
      RECT  4175.0 30032.5 12335.0 30097.5 ;
      RECT  4175.0 32722.5 12335.0 32787.5 ;
      RECT  14112.5 32097.5 17195.0 32162.5 ;
      RECT  14317.5 31957.5 17195.0 32022.5 ;
      RECT  14522.5 31817.5 17195.0 31882.5 ;
      RECT  14727.5 31677.5 17195.0 31742.5 ;
      RECT  11925.0 630.0 14112.5 695.0 ;
      RECT  11925.0 2065.0 14317.5 2130.0 ;
      RECT  11925.0 3320.0 14522.5 3385.0 ;
      RECT  11925.0 4755.0 14727.5 4820.0 ;
      RECT  11925.0 2.5 15102.5 67.5 ;
      RECT  11925.0 2692.5 15102.5 2757.5 ;
      RECT  11925.0 5382.5 15102.5 5447.5 ;
      RECT  4175.0 1347.5 15102.5 1412.5 ;
      RECT  4175.0 4037.5 15102.5 4102.5 ;
      RECT  11095.0 11785.0 12677.5 11850.0 ;
      RECT  11095.0 11080.0 12882.5 11145.0 ;
      RECT  11095.0 10375.0 13087.5 10440.0 ;
      RECT  11095.0 9670.0 13292.5 9735.0 ;
      RECT  11095.0 8965.0 13497.5 9030.0 ;
      RECT  11095.0 8260.0 13702.5 8325.0 ;
      RECT  11095.0 7555.0 13907.5 7620.0 ;
      RECT  11095.0 12137.5 15237.5 12202.5 ;
      RECT  11095.0 11432.5 15237.5 11497.5 ;
      RECT  11095.0 10727.5 15237.5 10792.5 ;
      RECT  11095.0 10022.5 15237.5 10087.5 ;
      RECT  11095.0 9317.5 15237.5 9382.5 ;
      RECT  11095.0 8612.5 15237.5 8677.5 ;
      RECT  11095.0 7907.5 15237.5 7972.5 ;
      RECT  11095.0 7202.5 15237.5 7267.5 ;
      RECT  11095.0 6497.5 15237.5 6562.5 ;
      RECT  11095.0 5792.5 15237.5 5857.5 ;
      RECT  7865.0 5587.5 7930.0 5652.5 ;
      RECT  7865.0 5620.0 7930.0 5825.0 ;
      RECT  4175.0 5587.5 7897.5 5652.5 ;
      RECT  10825.0 5587.5 10890.0 5652.5 ;
      RECT  10825.0 5620.0 10890.0 5825.0 ;
      RECT  4175.0 5587.5 10857.5 5652.5 ;
      RECT  5875.0 5587.5 5940.0 5652.5 ;
      RECT  5875.0 5620.0 5940.0 5825.0 ;
      RECT  4175.0 5587.5 5907.5 5652.5 ;
      RECT  8835.0 5587.5 8900.0 5652.5 ;
      RECT  8835.0 5620.0 8900.0 5825.0 ;
      RECT  4175.0 5587.5 8867.5 5652.5 ;
      RECT  16307.5 15960.0 17195.0 16025.0 ;
      RECT  15897.5 13775.0 17195.0 13840.0 ;
      RECT  16102.5 15322.5 17195.0 15387.5 ;
      RECT  16307.5 207237.5 17195.0 207302.5 ;
      RECT  16512.5 22462.5 17195.0 22527.5 ;
      RECT  16717.5 26487.5 17195.0 26552.5 ;
      RECT  4860.0 12342.5 4925.0 12407.5 ;
      RECT  4860.0 12170.0 4925.0 12375.0 ;
      RECT  4892.5 12342.5 15692.5 12407.5 ;
      RECT  9255.0 206432.5 15757.5 206497.5 ;
      RECT  17195.0 207922.5 107630.0 207987.5 ;
      RECT  17195.0 31060.0 107630.0 31125.0 ;
      RECT  17195.0 22592.5 107630.0 22657.5 ;
      RECT  17195.0 18965.0 107630.0 19030.0 ;
      RECT  17195.0 21925.0 107630.0 21990.0 ;
      RECT  17195.0 16975.0 107630.0 17040.0 ;
      RECT  17195.0 19935.0 107630.0 20000.0 ;
      RECT  17195.0 13905.0 107630.0 13970.0 ;
      RECT  15452.5 15192.5 17195.0 15257.5 ;
      RECT  15452.5 26617.5 17195.0 26682.5 ;
      RECT  15452.5 16120.0 17195.0 16185.0 ;
      RECT  15452.5 23395.0 17195.0 23460.0 ;
      RECT  17195.0 34100.0 17900.0 35445.0 ;
      RECT  17195.0 36790.0 17900.0 35445.0 ;
      RECT  17195.0 36790.0 17900.0 38135.0 ;
      RECT  17195.0 39480.0 17900.0 38135.0 ;
      RECT  17195.0 39480.0 17900.0 40825.0 ;
      RECT  17195.0 42170.0 17900.0 40825.0 ;
      RECT  17195.0 42170.0 17900.0 43515.0 ;
      RECT  17195.0 44860.0 17900.0 43515.0 ;
      RECT  17195.0 44860.0 17900.0 46205.0 ;
      RECT  17195.0 47550.0 17900.0 46205.0 ;
      RECT  17195.0 47550.0 17900.0 48895.0 ;
      RECT  17195.0 50240.0 17900.0 48895.0 ;
      RECT  17195.0 50240.0 17900.0 51585.0 ;
      RECT  17195.0 52930.0 17900.0 51585.0 ;
      RECT  17195.0 52930.0 17900.0 54275.0 ;
      RECT  17195.0 55620.0 17900.0 54275.0 ;
      RECT  17195.0 55620.0 17900.0 56965.0 ;
      RECT  17195.0 58310.0 17900.0 56965.0 ;
      RECT  17195.0 58310.0 17900.0 59655.0 ;
      RECT  17195.0 61000.0 17900.0 59655.0 ;
      RECT  17195.0 61000.0 17900.0 62345.0 ;
      RECT  17195.0 63690.0 17900.0 62345.0 ;
      RECT  17195.0 63690.0 17900.0 65035.0 ;
      RECT  17195.0 66380.0 17900.0 65035.0 ;
      RECT  17195.0 66380.0 17900.0 67725.0 ;
      RECT  17195.0 69070.0 17900.0 67725.0 ;
      RECT  17195.0 69070.0 17900.0 70415.0 ;
      RECT  17195.0 71760.0 17900.0 70415.0 ;
      RECT  17195.0 71760.0 17900.0 73105.0 ;
      RECT  17195.0 74450.0 17900.0 73105.0 ;
      RECT  17195.0 74450.0 17900.0 75795.0 ;
      RECT  17195.0 77140.0 17900.0 75795.0 ;
      RECT  17195.0 77140.0 17900.0 78485.0 ;
      RECT  17195.0 79830.0 17900.0 78485.0 ;
      RECT  17195.0 79830.0 17900.0 81175.0 ;
      RECT  17195.0 82520.0 17900.0 81175.0 ;
      RECT  17195.0 82520.0 17900.0 83865.0 ;
      RECT  17195.0 85210.0 17900.0 83865.0 ;
      RECT  17195.0 85210.0 17900.0 86555.0 ;
      RECT  17195.0 87900.0 17900.0 86555.0 ;
      RECT  17195.0 87900.0 17900.0 89245.0 ;
      RECT  17195.0 90590.0 17900.0 89245.0 ;
      RECT  17195.0 90590.0 17900.0 91935.0 ;
      RECT  17195.0 93280.0 17900.0 91935.0 ;
      RECT  17195.0 93280.0 17900.0 94625.0 ;
      RECT  17195.0 95970.0 17900.0 94625.0 ;
      RECT  17195.0 95970.0 17900.0 97315.0 ;
      RECT  17195.0 98660.0 17900.0 97315.0 ;
      RECT  17195.0 98660.0 17900.0 100005.0 ;
      RECT  17195.0 101350.0 17900.0 100005.0 ;
      RECT  17195.0 101350.0 17900.0 102695.0 ;
      RECT  17195.0 104040.0 17900.0 102695.0 ;
      RECT  17195.0 104040.0 17900.0 105385.0 ;
      RECT  17195.0 106730.0 17900.0 105385.0 ;
      RECT  17195.0 106730.0 17900.0 108075.0 ;
      RECT  17195.0 109420.0 17900.0 108075.0 ;
      RECT  17195.0 109420.0 17900.0 110765.0 ;
      RECT  17195.0 112110.0 17900.0 110765.0 ;
      RECT  17195.0 112110.0 17900.0 113455.0 ;
      RECT  17195.0 114800.0 17900.0 113455.0 ;
      RECT  17195.0 114800.0 17900.0 116145.0 ;
      RECT  17195.0 117490.0 17900.0 116145.0 ;
      RECT  17195.0 117490.0 17900.0 118835.0 ;
      RECT  17195.0 120180.0 17900.0 118835.0 ;
      RECT  17195.0 120180.0 17900.0 121525.0 ;
      RECT  17195.0 122870.0 17900.0 121525.0 ;
      RECT  17195.0 122870.0 17900.0 124215.0 ;
      RECT  17195.0 125560.0 17900.0 124215.0 ;
      RECT  17195.0 125560.0 17900.0 126905.0 ;
      RECT  17195.0 128250.0 17900.0 126905.0 ;
      RECT  17195.0 128250.0 17900.0 129595.0 ;
      RECT  17195.0 130940.0 17900.0 129595.0 ;
      RECT  17195.0 130940.0 17900.0 132285.0 ;
      RECT  17195.0 133630.0 17900.0 132285.0 ;
      RECT  17195.0 133630.0 17900.0 134975.0 ;
      RECT  17195.0 136320.0 17900.0 134975.0 ;
      RECT  17195.0 136320.0 17900.0 137665.0 ;
      RECT  17195.0 139010.0 17900.0 137665.0 ;
      RECT  17195.0 139010.0 17900.0 140355.0 ;
      RECT  17195.0 141700.0 17900.0 140355.0 ;
      RECT  17195.0 141700.0 17900.0 143045.0 ;
      RECT  17195.0 144390.0 17900.0 143045.0 ;
      RECT  17195.0 144390.0 17900.0 145735.0 ;
      RECT  17195.0 147080.0 17900.0 145735.0 ;
      RECT  17195.0 147080.0 17900.0 148425.0 ;
      RECT  17195.0 149770.0 17900.0 148425.0 ;
      RECT  17195.0 149770.0 17900.0 151115.0 ;
      RECT  17195.0 152460.0 17900.0 151115.0 ;
      RECT  17195.0 152460.0 17900.0 153805.0 ;
      RECT  17195.0 155150.0 17900.0 153805.0 ;
      RECT  17195.0 155150.0 17900.0 156495.0 ;
      RECT  17195.0 157840.0 17900.0 156495.0 ;
      RECT  17195.0 157840.0 17900.0 159185.0 ;
      RECT  17195.0 160530.0 17900.0 159185.0 ;
      RECT  17195.0 160530.0 17900.0 161875.0 ;
      RECT  17195.0 163220.0 17900.0 161875.0 ;
      RECT  17195.0 163220.0 17900.0 164565.0 ;
      RECT  17195.0 165910.0 17900.0 164565.0 ;
      RECT  17195.0 165910.0 17900.0 167255.0 ;
      RECT  17195.0 168600.0 17900.0 167255.0 ;
      RECT  17195.0 168600.0 17900.0 169945.0 ;
      RECT  17195.0 171290.0 17900.0 169945.0 ;
      RECT  17195.0 171290.0 17900.0 172635.0 ;
      RECT  17195.0 173980.0 17900.0 172635.0 ;
      RECT  17195.0 173980.0 17900.0 175325.0 ;
      RECT  17195.0 176670.0 17900.0 175325.0 ;
      RECT  17195.0 176670.0 17900.0 178015.0 ;
      RECT  17195.0 179360.0 17900.0 178015.0 ;
      RECT  17195.0 179360.0 17900.0 180705.0 ;
      RECT  17195.0 182050.0 17900.0 180705.0 ;
      RECT  17195.0 182050.0 17900.0 183395.0 ;
      RECT  17195.0 184740.0 17900.0 183395.0 ;
      RECT  17195.0 184740.0 17900.0 186085.0 ;
      RECT  17195.0 187430.0 17900.0 186085.0 ;
      RECT  17195.0 187430.0 17900.0 188775.0 ;
      RECT  17195.0 190120.0 17900.0 188775.0 ;
      RECT  17195.0 190120.0 17900.0 191465.0 ;
      RECT  17195.0 192810.0 17900.0 191465.0 ;
      RECT  17195.0 192810.0 17900.0 194155.0 ;
      RECT  17195.0 195500.0 17900.0 194155.0 ;
      RECT  17195.0 195500.0 17900.0 196845.0 ;
      RECT  17195.0 198190.0 17900.0 196845.0 ;
      RECT  17195.0 198190.0 17900.0 199535.0 ;
      RECT  17195.0 200880.0 17900.0 199535.0 ;
      RECT  17195.0 200880.0 17900.0 202225.0 ;
      RECT  17195.0 203570.0 17900.0 202225.0 ;
      RECT  17195.0 203570.0 17900.0 204915.0 ;
      RECT  17195.0 206260.0 17900.0 204915.0 ;
      RECT  17900.0 34100.0 18605.0 35445.0 ;
      RECT  17900.0 36790.0 18605.0 35445.0 ;
      RECT  17900.0 36790.0 18605.0 38135.0 ;
      RECT  17900.0 39480.0 18605.0 38135.0 ;
      RECT  17900.0 39480.0 18605.0 40825.0 ;
      RECT  17900.0 42170.0 18605.0 40825.0 ;
      RECT  17900.0 42170.0 18605.0 43515.0 ;
      RECT  17900.0 44860.0 18605.0 43515.0 ;
      RECT  17900.0 44860.0 18605.0 46205.0 ;
      RECT  17900.0 47550.0 18605.0 46205.0 ;
      RECT  17900.0 47550.0 18605.0 48895.0 ;
      RECT  17900.0 50240.0 18605.0 48895.0 ;
      RECT  17900.0 50240.0 18605.0 51585.0 ;
      RECT  17900.0 52930.0 18605.0 51585.0 ;
      RECT  17900.0 52930.0 18605.0 54275.0 ;
      RECT  17900.0 55620.0 18605.0 54275.0 ;
      RECT  17900.0 55620.0 18605.0 56965.0 ;
      RECT  17900.0 58310.0 18605.0 56965.0 ;
      RECT  17900.0 58310.0 18605.0 59655.0 ;
      RECT  17900.0 61000.0 18605.0 59655.0 ;
      RECT  17900.0 61000.0 18605.0 62345.0 ;
      RECT  17900.0 63690.0 18605.0 62345.0 ;
      RECT  17900.0 63690.0 18605.0 65035.0 ;
      RECT  17900.0 66380.0 18605.0 65035.0 ;
      RECT  17900.0 66380.0 18605.0 67725.0 ;
      RECT  17900.0 69070.0 18605.0 67725.0 ;
      RECT  17900.0 69070.0 18605.0 70415.0 ;
      RECT  17900.0 71760.0 18605.0 70415.0 ;
      RECT  17900.0 71760.0 18605.0 73105.0 ;
      RECT  17900.0 74450.0 18605.0 73105.0 ;
      RECT  17900.0 74450.0 18605.0 75795.0 ;
      RECT  17900.0 77140.0 18605.0 75795.0 ;
      RECT  17900.0 77140.0 18605.0 78485.0 ;
      RECT  17900.0 79830.0 18605.0 78485.0 ;
      RECT  17900.0 79830.0 18605.0 81175.0 ;
      RECT  17900.0 82520.0 18605.0 81175.0 ;
      RECT  17900.0 82520.0 18605.0 83865.0 ;
      RECT  17900.0 85210.0 18605.0 83865.0 ;
      RECT  17900.0 85210.0 18605.0 86555.0 ;
      RECT  17900.0 87900.0 18605.0 86555.0 ;
      RECT  17900.0 87900.0 18605.0 89245.0 ;
      RECT  17900.0 90590.0 18605.0 89245.0 ;
      RECT  17900.0 90590.0 18605.0 91935.0 ;
      RECT  17900.0 93280.0 18605.0 91935.0 ;
      RECT  17900.0 93280.0 18605.0 94625.0 ;
      RECT  17900.0 95970.0 18605.0 94625.0 ;
      RECT  17900.0 95970.0 18605.0 97315.0 ;
      RECT  17900.0 98660.0 18605.0 97315.0 ;
      RECT  17900.0 98660.0 18605.0 100005.0 ;
      RECT  17900.0 101350.0 18605.0 100005.0 ;
      RECT  17900.0 101350.0 18605.0 102695.0 ;
      RECT  17900.0 104040.0 18605.0 102695.0 ;
      RECT  17900.0 104040.0 18605.0 105385.0 ;
      RECT  17900.0 106730.0 18605.0 105385.0 ;
      RECT  17900.0 106730.0 18605.0 108075.0 ;
      RECT  17900.0 109420.0 18605.0 108075.0 ;
      RECT  17900.0 109420.0 18605.0 110765.0 ;
      RECT  17900.0 112110.0 18605.0 110765.0 ;
      RECT  17900.0 112110.0 18605.0 113455.0 ;
      RECT  17900.0 114800.0 18605.0 113455.0 ;
      RECT  17900.0 114800.0 18605.0 116145.0 ;
      RECT  17900.0 117490.0 18605.0 116145.0 ;
      RECT  17900.0 117490.0 18605.0 118835.0 ;
      RECT  17900.0 120180.0 18605.0 118835.0 ;
      RECT  17900.0 120180.0 18605.0 121525.0 ;
      RECT  17900.0 122870.0 18605.0 121525.0 ;
      RECT  17900.0 122870.0 18605.0 124215.0 ;
      RECT  17900.0 125560.0 18605.0 124215.0 ;
      RECT  17900.0 125560.0 18605.0 126905.0 ;
      RECT  17900.0 128250.0 18605.0 126905.0 ;
      RECT  17900.0 128250.0 18605.0 129595.0 ;
      RECT  17900.0 130940.0 18605.0 129595.0 ;
      RECT  17900.0 130940.0 18605.0 132285.0 ;
      RECT  17900.0 133630.0 18605.0 132285.0 ;
      RECT  17900.0 133630.0 18605.0 134975.0 ;
      RECT  17900.0 136320.0 18605.0 134975.0 ;
      RECT  17900.0 136320.0 18605.0 137665.0 ;
      RECT  17900.0 139010.0 18605.0 137665.0 ;
      RECT  17900.0 139010.0 18605.0 140355.0 ;
      RECT  17900.0 141700.0 18605.0 140355.0 ;
      RECT  17900.0 141700.0 18605.0 143045.0 ;
      RECT  17900.0 144390.0 18605.0 143045.0 ;
      RECT  17900.0 144390.0 18605.0 145735.0 ;
      RECT  17900.0 147080.0 18605.0 145735.0 ;
      RECT  17900.0 147080.0 18605.0 148425.0 ;
      RECT  17900.0 149770.0 18605.0 148425.0 ;
      RECT  17900.0 149770.0 18605.0 151115.0 ;
      RECT  17900.0 152460.0 18605.0 151115.0 ;
      RECT  17900.0 152460.0 18605.0 153805.0 ;
      RECT  17900.0 155150.0 18605.0 153805.0 ;
      RECT  17900.0 155150.0 18605.0 156495.0 ;
      RECT  17900.0 157840.0 18605.0 156495.0 ;
      RECT  17900.0 157840.0 18605.0 159185.0 ;
      RECT  17900.0 160530.0 18605.0 159185.0 ;
      RECT  17900.0 160530.0 18605.0 161875.0 ;
      RECT  17900.0 163220.0 18605.0 161875.0 ;
      RECT  17900.0 163220.0 18605.0 164565.0 ;
      RECT  17900.0 165910.0 18605.0 164565.0 ;
      RECT  17900.0 165910.0 18605.0 167255.0 ;
      RECT  17900.0 168600.0 18605.0 167255.0 ;
      RECT  17900.0 168600.0 18605.0 169945.0 ;
      RECT  17900.0 171290.0 18605.0 169945.0 ;
      RECT  17900.0 171290.0 18605.0 172635.0 ;
      RECT  17900.0 173980.0 18605.0 172635.0 ;
      RECT  17900.0 173980.0 18605.0 175325.0 ;
      RECT  17900.0 176670.0 18605.0 175325.0 ;
      RECT  17900.0 176670.0 18605.0 178015.0 ;
      RECT  17900.0 179360.0 18605.0 178015.0 ;
      RECT  17900.0 179360.0 18605.0 180705.0 ;
      RECT  17900.0 182050.0 18605.0 180705.0 ;
      RECT  17900.0 182050.0 18605.0 183395.0 ;
      RECT  17900.0 184740.0 18605.0 183395.0 ;
      RECT  17900.0 184740.0 18605.0 186085.0 ;
      RECT  17900.0 187430.0 18605.0 186085.0 ;
      RECT  17900.0 187430.0 18605.0 188775.0 ;
      RECT  17900.0 190120.0 18605.0 188775.0 ;
      RECT  17900.0 190120.0 18605.0 191465.0 ;
      RECT  17900.0 192810.0 18605.0 191465.0 ;
      RECT  17900.0 192810.0 18605.0 194155.0 ;
      RECT  17900.0 195500.0 18605.0 194155.0 ;
      RECT  17900.0 195500.0 18605.0 196845.0 ;
      RECT  17900.0 198190.0 18605.0 196845.0 ;
      RECT  17900.0 198190.0 18605.0 199535.0 ;
      RECT  17900.0 200880.0 18605.0 199535.0 ;
      RECT  17900.0 200880.0 18605.0 202225.0 ;
      RECT  17900.0 203570.0 18605.0 202225.0 ;
      RECT  17900.0 203570.0 18605.0 204915.0 ;
      RECT  17900.0 206260.0 18605.0 204915.0 ;
      RECT  18605.0 34100.0 19310.0 35445.0 ;
      RECT  18605.0 36790.0 19310.0 35445.0 ;
      RECT  18605.0 36790.0 19310.0 38135.0 ;
      RECT  18605.0 39480.0 19310.0 38135.0 ;
      RECT  18605.0 39480.0 19310.0 40825.0 ;
      RECT  18605.0 42170.0 19310.0 40825.0 ;
      RECT  18605.0 42170.0 19310.0 43515.0 ;
      RECT  18605.0 44860.0 19310.0 43515.0 ;
      RECT  18605.0 44860.0 19310.0 46205.0 ;
      RECT  18605.0 47550.0 19310.0 46205.0 ;
      RECT  18605.0 47550.0 19310.0 48895.0 ;
      RECT  18605.0 50240.0 19310.0 48895.0 ;
      RECT  18605.0 50240.0 19310.0 51585.0 ;
      RECT  18605.0 52930.0 19310.0 51585.0 ;
      RECT  18605.0 52930.0 19310.0 54275.0 ;
      RECT  18605.0 55620.0 19310.0 54275.0 ;
      RECT  18605.0 55620.0 19310.0 56965.0 ;
      RECT  18605.0 58310.0 19310.0 56965.0 ;
      RECT  18605.0 58310.0 19310.0 59655.0 ;
      RECT  18605.0 61000.0 19310.0 59655.0 ;
      RECT  18605.0 61000.0 19310.0 62345.0 ;
      RECT  18605.0 63690.0 19310.0 62345.0 ;
      RECT  18605.0 63690.0 19310.0 65035.0 ;
      RECT  18605.0 66380.0 19310.0 65035.0 ;
      RECT  18605.0 66380.0 19310.0 67725.0 ;
      RECT  18605.0 69070.0 19310.0 67725.0 ;
      RECT  18605.0 69070.0 19310.0 70415.0 ;
      RECT  18605.0 71760.0 19310.0 70415.0 ;
      RECT  18605.0 71760.0 19310.0 73105.0 ;
      RECT  18605.0 74450.0 19310.0 73105.0 ;
      RECT  18605.0 74450.0 19310.0 75795.0 ;
      RECT  18605.0 77140.0 19310.0 75795.0 ;
      RECT  18605.0 77140.0 19310.0 78485.0 ;
      RECT  18605.0 79830.0 19310.0 78485.0 ;
      RECT  18605.0 79830.0 19310.0 81175.0 ;
      RECT  18605.0 82520.0 19310.0 81175.0 ;
      RECT  18605.0 82520.0 19310.0 83865.0 ;
      RECT  18605.0 85210.0 19310.0 83865.0 ;
      RECT  18605.0 85210.0 19310.0 86555.0 ;
      RECT  18605.0 87900.0 19310.0 86555.0 ;
      RECT  18605.0 87900.0 19310.0 89245.0 ;
      RECT  18605.0 90590.0 19310.0 89245.0 ;
      RECT  18605.0 90590.0 19310.0 91935.0 ;
      RECT  18605.0 93280.0 19310.0 91935.0 ;
      RECT  18605.0 93280.0 19310.0 94625.0 ;
      RECT  18605.0 95970.0 19310.0 94625.0 ;
      RECT  18605.0 95970.0 19310.0 97315.0 ;
      RECT  18605.0 98660.0 19310.0 97315.0 ;
      RECT  18605.0 98660.0 19310.0 100005.0 ;
      RECT  18605.0 101350.0 19310.0 100005.0 ;
      RECT  18605.0 101350.0 19310.0 102695.0 ;
      RECT  18605.0 104040.0 19310.0 102695.0 ;
      RECT  18605.0 104040.0 19310.0 105385.0 ;
      RECT  18605.0 106730.0 19310.0 105385.0 ;
      RECT  18605.0 106730.0 19310.0 108075.0 ;
      RECT  18605.0 109420.0 19310.0 108075.0 ;
      RECT  18605.0 109420.0 19310.0 110765.0 ;
      RECT  18605.0 112110.0 19310.0 110765.0 ;
      RECT  18605.0 112110.0 19310.0 113455.0 ;
      RECT  18605.0 114800.0 19310.0 113455.0 ;
      RECT  18605.0 114800.0 19310.0 116145.0 ;
      RECT  18605.0 117490.0 19310.0 116145.0 ;
      RECT  18605.0 117490.0 19310.0 118835.0 ;
      RECT  18605.0 120180.0 19310.0 118835.0 ;
      RECT  18605.0 120180.0 19310.0 121525.0 ;
      RECT  18605.0 122870.0 19310.0 121525.0 ;
      RECT  18605.0 122870.0 19310.0 124215.0 ;
      RECT  18605.0 125560.0 19310.0 124215.0 ;
      RECT  18605.0 125560.0 19310.0 126905.0 ;
      RECT  18605.0 128250.0 19310.0 126905.0 ;
      RECT  18605.0 128250.0 19310.0 129595.0 ;
      RECT  18605.0 130940.0 19310.0 129595.0 ;
      RECT  18605.0 130940.0 19310.0 132285.0 ;
      RECT  18605.0 133630.0 19310.0 132285.0 ;
      RECT  18605.0 133630.0 19310.0 134975.0 ;
      RECT  18605.0 136320.0 19310.0 134975.0 ;
      RECT  18605.0 136320.0 19310.0 137665.0 ;
      RECT  18605.0 139010.0 19310.0 137665.0 ;
      RECT  18605.0 139010.0 19310.0 140355.0 ;
      RECT  18605.0 141700.0 19310.0 140355.0 ;
      RECT  18605.0 141700.0 19310.0 143045.0 ;
      RECT  18605.0 144390.0 19310.0 143045.0 ;
      RECT  18605.0 144390.0 19310.0 145735.0 ;
      RECT  18605.0 147080.0 19310.0 145735.0 ;
      RECT  18605.0 147080.0 19310.0 148425.0 ;
      RECT  18605.0 149770.0 19310.0 148425.0 ;
      RECT  18605.0 149770.0 19310.0 151115.0 ;
      RECT  18605.0 152460.0 19310.0 151115.0 ;
      RECT  18605.0 152460.0 19310.0 153805.0 ;
      RECT  18605.0 155150.0 19310.0 153805.0 ;
      RECT  18605.0 155150.0 19310.0 156495.0 ;
      RECT  18605.0 157840.0 19310.0 156495.0 ;
      RECT  18605.0 157840.0 19310.0 159185.0 ;
      RECT  18605.0 160530.0 19310.0 159185.0 ;
      RECT  18605.0 160530.0 19310.0 161875.0 ;
      RECT  18605.0 163220.0 19310.0 161875.0 ;
      RECT  18605.0 163220.0 19310.0 164565.0 ;
      RECT  18605.0 165910.0 19310.0 164565.0 ;
      RECT  18605.0 165910.0 19310.0 167255.0 ;
      RECT  18605.0 168600.0 19310.0 167255.0 ;
      RECT  18605.0 168600.0 19310.0 169945.0 ;
      RECT  18605.0 171290.0 19310.0 169945.0 ;
      RECT  18605.0 171290.0 19310.0 172635.0 ;
      RECT  18605.0 173980.0 19310.0 172635.0 ;
      RECT  18605.0 173980.0 19310.0 175325.0 ;
      RECT  18605.0 176670.0 19310.0 175325.0 ;
      RECT  18605.0 176670.0 19310.0 178015.0 ;
      RECT  18605.0 179360.0 19310.0 178015.0 ;
      RECT  18605.0 179360.0 19310.0 180705.0 ;
      RECT  18605.0 182050.0 19310.0 180705.0 ;
      RECT  18605.0 182050.0 19310.0 183395.0 ;
      RECT  18605.0 184740.0 19310.0 183395.0 ;
      RECT  18605.0 184740.0 19310.0 186085.0 ;
      RECT  18605.0 187430.0 19310.0 186085.0 ;
      RECT  18605.0 187430.0 19310.0 188775.0 ;
      RECT  18605.0 190120.0 19310.0 188775.0 ;
      RECT  18605.0 190120.0 19310.0 191465.0 ;
      RECT  18605.0 192810.0 19310.0 191465.0 ;
      RECT  18605.0 192810.0 19310.0 194155.0 ;
      RECT  18605.0 195500.0 19310.0 194155.0 ;
      RECT  18605.0 195500.0 19310.0 196845.0 ;
      RECT  18605.0 198190.0 19310.0 196845.0 ;
      RECT  18605.0 198190.0 19310.0 199535.0 ;
      RECT  18605.0 200880.0 19310.0 199535.0 ;
      RECT  18605.0 200880.0 19310.0 202225.0 ;
      RECT  18605.0 203570.0 19310.0 202225.0 ;
      RECT  18605.0 203570.0 19310.0 204915.0 ;
      RECT  18605.0 206260.0 19310.0 204915.0 ;
      RECT  19310.0 34100.0 20015.0 35445.0 ;
      RECT  19310.0 36790.0 20015.0 35445.0 ;
      RECT  19310.0 36790.0 20015.0 38135.0 ;
      RECT  19310.0 39480.0 20015.0 38135.0 ;
      RECT  19310.0 39480.0 20015.0 40825.0 ;
      RECT  19310.0 42170.0 20015.0 40825.0 ;
      RECT  19310.0 42170.0 20015.0 43515.0 ;
      RECT  19310.0 44860.0 20015.0 43515.0 ;
      RECT  19310.0 44860.0 20015.0 46205.0 ;
      RECT  19310.0 47550.0 20015.0 46205.0 ;
      RECT  19310.0 47550.0 20015.0 48895.0 ;
      RECT  19310.0 50240.0 20015.0 48895.0 ;
      RECT  19310.0 50240.0 20015.0 51585.0 ;
      RECT  19310.0 52930.0 20015.0 51585.0 ;
      RECT  19310.0 52930.0 20015.0 54275.0 ;
      RECT  19310.0 55620.0 20015.0 54275.0 ;
      RECT  19310.0 55620.0 20015.0 56965.0 ;
      RECT  19310.0 58310.0 20015.0 56965.0 ;
      RECT  19310.0 58310.0 20015.0 59655.0 ;
      RECT  19310.0 61000.0 20015.0 59655.0 ;
      RECT  19310.0 61000.0 20015.0 62345.0 ;
      RECT  19310.0 63690.0 20015.0 62345.0 ;
      RECT  19310.0 63690.0 20015.0 65035.0 ;
      RECT  19310.0 66380.0 20015.0 65035.0 ;
      RECT  19310.0 66380.0 20015.0 67725.0 ;
      RECT  19310.0 69070.0 20015.0 67725.0 ;
      RECT  19310.0 69070.0 20015.0 70415.0 ;
      RECT  19310.0 71760.0 20015.0 70415.0 ;
      RECT  19310.0 71760.0 20015.0 73105.0 ;
      RECT  19310.0 74450.0 20015.0 73105.0 ;
      RECT  19310.0 74450.0 20015.0 75795.0 ;
      RECT  19310.0 77140.0 20015.0 75795.0 ;
      RECT  19310.0 77140.0 20015.0 78485.0 ;
      RECT  19310.0 79830.0 20015.0 78485.0 ;
      RECT  19310.0 79830.0 20015.0 81175.0 ;
      RECT  19310.0 82520.0 20015.0 81175.0 ;
      RECT  19310.0 82520.0 20015.0 83865.0 ;
      RECT  19310.0 85210.0 20015.0 83865.0 ;
      RECT  19310.0 85210.0 20015.0 86555.0 ;
      RECT  19310.0 87900.0 20015.0 86555.0 ;
      RECT  19310.0 87900.0 20015.0 89245.0 ;
      RECT  19310.0 90590.0 20015.0 89245.0 ;
      RECT  19310.0 90590.0 20015.0 91935.0 ;
      RECT  19310.0 93280.0 20015.0 91935.0 ;
      RECT  19310.0 93280.0 20015.0 94625.0 ;
      RECT  19310.0 95970.0 20015.0 94625.0 ;
      RECT  19310.0 95970.0 20015.0 97315.0 ;
      RECT  19310.0 98660.0 20015.0 97315.0 ;
      RECT  19310.0 98660.0 20015.0 100005.0 ;
      RECT  19310.0 101350.0 20015.0 100005.0 ;
      RECT  19310.0 101350.0 20015.0 102695.0 ;
      RECT  19310.0 104040.0 20015.0 102695.0 ;
      RECT  19310.0 104040.0 20015.0 105385.0 ;
      RECT  19310.0 106730.0 20015.0 105385.0 ;
      RECT  19310.0 106730.0 20015.0 108075.0 ;
      RECT  19310.0 109420.0 20015.0 108075.0 ;
      RECT  19310.0 109420.0 20015.0 110765.0 ;
      RECT  19310.0 112110.0 20015.0 110765.0 ;
      RECT  19310.0 112110.0 20015.0 113455.0 ;
      RECT  19310.0 114800.0 20015.0 113455.0 ;
      RECT  19310.0 114800.0 20015.0 116145.0 ;
      RECT  19310.0 117490.0 20015.0 116145.0 ;
      RECT  19310.0 117490.0 20015.0 118835.0 ;
      RECT  19310.0 120180.0 20015.0 118835.0 ;
      RECT  19310.0 120180.0 20015.0 121525.0 ;
      RECT  19310.0 122870.0 20015.0 121525.0 ;
      RECT  19310.0 122870.0 20015.0 124215.0 ;
      RECT  19310.0 125560.0 20015.0 124215.0 ;
      RECT  19310.0 125560.0 20015.0 126905.0 ;
      RECT  19310.0 128250.0 20015.0 126905.0 ;
      RECT  19310.0 128250.0 20015.0 129595.0 ;
      RECT  19310.0 130940.0 20015.0 129595.0 ;
      RECT  19310.0 130940.0 20015.0 132285.0 ;
      RECT  19310.0 133630.0 20015.0 132285.0 ;
      RECT  19310.0 133630.0 20015.0 134975.0 ;
      RECT  19310.0 136320.0 20015.0 134975.0 ;
      RECT  19310.0 136320.0 20015.0 137665.0 ;
      RECT  19310.0 139010.0 20015.0 137665.0 ;
      RECT  19310.0 139010.0 20015.0 140355.0 ;
      RECT  19310.0 141700.0 20015.0 140355.0 ;
      RECT  19310.0 141700.0 20015.0 143045.0 ;
      RECT  19310.0 144390.0 20015.0 143045.0 ;
      RECT  19310.0 144390.0 20015.0 145735.0 ;
      RECT  19310.0 147080.0 20015.0 145735.0 ;
      RECT  19310.0 147080.0 20015.0 148425.0 ;
      RECT  19310.0 149770.0 20015.0 148425.0 ;
      RECT  19310.0 149770.0 20015.0 151115.0 ;
      RECT  19310.0 152460.0 20015.0 151115.0 ;
      RECT  19310.0 152460.0 20015.0 153805.0 ;
      RECT  19310.0 155150.0 20015.0 153805.0 ;
      RECT  19310.0 155150.0 20015.0 156495.0 ;
      RECT  19310.0 157840.0 20015.0 156495.0 ;
      RECT  19310.0 157840.0 20015.0 159185.0 ;
      RECT  19310.0 160530.0 20015.0 159185.0 ;
      RECT  19310.0 160530.0 20015.0 161875.0 ;
      RECT  19310.0 163220.0 20015.0 161875.0 ;
      RECT  19310.0 163220.0 20015.0 164565.0 ;
      RECT  19310.0 165910.0 20015.0 164565.0 ;
      RECT  19310.0 165910.0 20015.0 167255.0 ;
      RECT  19310.0 168600.0 20015.0 167255.0 ;
      RECT  19310.0 168600.0 20015.0 169945.0 ;
      RECT  19310.0 171290.0 20015.0 169945.0 ;
      RECT  19310.0 171290.0 20015.0 172635.0 ;
      RECT  19310.0 173980.0 20015.0 172635.0 ;
      RECT  19310.0 173980.0 20015.0 175325.0 ;
      RECT  19310.0 176670.0 20015.0 175325.0 ;
      RECT  19310.0 176670.0 20015.0 178015.0 ;
      RECT  19310.0 179360.0 20015.0 178015.0 ;
      RECT  19310.0 179360.0 20015.0 180705.0 ;
      RECT  19310.0 182050.0 20015.0 180705.0 ;
      RECT  19310.0 182050.0 20015.0 183395.0 ;
      RECT  19310.0 184740.0 20015.0 183395.0 ;
      RECT  19310.0 184740.0 20015.0 186085.0 ;
      RECT  19310.0 187430.0 20015.0 186085.0 ;
      RECT  19310.0 187430.0 20015.0 188775.0 ;
      RECT  19310.0 190120.0 20015.0 188775.0 ;
      RECT  19310.0 190120.0 20015.0 191465.0 ;
      RECT  19310.0 192810.0 20015.0 191465.0 ;
      RECT  19310.0 192810.0 20015.0 194155.0 ;
      RECT  19310.0 195500.0 20015.0 194155.0 ;
      RECT  19310.0 195500.0 20015.0 196845.0 ;
      RECT  19310.0 198190.0 20015.0 196845.0 ;
      RECT  19310.0 198190.0 20015.0 199535.0 ;
      RECT  19310.0 200880.0 20015.0 199535.0 ;
      RECT  19310.0 200880.0 20015.0 202225.0 ;
      RECT  19310.0 203570.0 20015.0 202225.0 ;
      RECT  19310.0 203570.0 20015.0 204915.0 ;
      RECT  19310.0 206260.0 20015.0 204915.0 ;
      RECT  20015.0 34100.0 20720.0 35445.0 ;
      RECT  20015.0 36790.0 20720.0 35445.0 ;
      RECT  20015.0 36790.0 20720.0 38135.0 ;
      RECT  20015.0 39480.0 20720.0 38135.0 ;
      RECT  20015.0 39480.0 20720.0 40825.0 ;
      RECT  20015.0 42170.0 20720.0 40825.0 ;
      RECT  20015.0 42170.0 20720.0 43515.0 ;
      RECT  20015.0 44860.0 20720.0 43515.0 ;
      RECT  20015.0 44860.0 20720.0 46205.0 ;
      RECT  20015.0 47550.0 20720.0 46205.0 ;
      RECT  20015.0 47550.0 20720.0 48895.0 ;
      RECT  20015.0 50240.0 20720.0 48895.0 ;
      RECT  20015.0 50240.0 20720.0 51585.0 ;
      RECT  20015.0 52930.0 20720.0 51585.0 ;
      RECT  20015.0 52930.0 20720.0 54275.0 ;
      RECT  20015.0 55620.0 20720.0 54275.0 ;
      RECT  20015.0 55620.0 20720.0 56965.0 ;
      RECT  20015.0 58310.0 20720.0 56965.0 ;
      RECT  20015.0 58310.0 20720.0 59655.0 ;
      RECT  20015.0 61000.0 20720.0 59655.0 ;
      RECT  20015.0 61000.0 20720.0 62345.0 ;
      RECT  20015.0 63690.0 20720.0 62345.0 ;
      RECT  20015.0 63690.0 20720.0 65035.0 ;
      RECT  20015.0 66380.0 20720.0 65035.0 ;
      RECT  20015.0 66380.0 20720.0 67725.0 ;
      RECT  20015.0 69070.0 20720.0 67725.0 ;
      RECT  20015.0 69070.0 20720.0 70415.0 ;
      RECT  20015.0 71760.0 20720.0 70415.0 ;
      RECT  20015.0 71760.0 20720.0 73105.0 ;
      RECT  20015.0 74450.0 20720.0 73105.0 ;
      RECT  20015.0 74450.0 20720.0 75795.0 ;
      RECT  20015.0 77140.0 20720.0 75795.0 ;
      RECT  20015.0 77140.0 20720.0 78485.0 ;
      RECT  20015.0 79830.0 20720.0 78485.0 ;
      RECT  20015.0 79830.0 20720.0 81175.0 ;
      RECT  20015.0 82520.0 20720.0 81175.0 ;
      RECT  20015.0 82520.0 20720.0 83865.0 ;
      RECT  20015.0 85210.0 20720.0 83865.0 ;
      RECT  20015.0 85210.0 20720.0 86555.0 ;
      RECT  20015.0 87900.0 20720.0 86555.0 ;
      RECT  20015.0 87900.0 20720.0 89245.0 ;
      RECT  20015.0 90590.0 20720.0 89245.0 ;
      RECT  20015.0 90590.0 20720.0 91935.0 ;
      RECT  20015.0 93280.0 20720.0 91935.0 ;
      RECT  20015.0 93280.0 20720.0 94625.0 ;
      RECT  20015.0 95970.0 20720.0 94625.0 ;
      RECT  20015.0 95970.0 20720.0 97315.0 ;
      RECT  20015.0 98660.0 20720.0 97315.0 ;
      RECT  20015.0 98660.0 20720.0 100005.0 ;
      RECT  20015.0 101350.0 20720.0 100005.0 ;
      RECT  20015.0 101350.0 20720.0 102695.0 ;
      RECT  20015.0 104040.0 20720.0 102695.0 ;
      RECT  20015.0 104040.0 20720.0 105385.0 ;
      RECT  20015.0 106730.0 20720.0 105385.0 ;
      RECT  20015.0 106730.0 20720.0 108075.0 ;
      RECT  20015.0 109420.0 20720.0 108075.0 ;
      RECT  20015.0 109420.0 20720.0 110765.0 ;
      RECT  20015.0 112110.0 20720.0 110765.0 ;
      RECT  20015.0 112110.0 20720.0 113455.0 ;
      RECT  20015.0 114800.0 20720.0 113455.0 ;
      RECT  20015.0 114800.0 20720.0 116145.0 ;
      RECT  20015.0 117490.0 20720.0 116145.0 ;
      RECT  20015.0 117490.0 20720.0 118835.0 ;
      RECT  20015.0 120180.0 20720.0 118835.0 ;
      RECT  20015.0 120180.0 20720.0 121525.0 ;
      RECT  20015.0 122870.0 20720.0 121525.0 ;
      RECT  20015.0 122870.0 20720.0 124215.0 ;
      RECT  20015.0 125560.0 20720.0 124215.0 ;
      RECT  20015.0 125560.0 20720.0 126905.0 ;
      RECT  20015.0 128250.0 20720.0 126905.0 ;
      RECT  20015.0 128250.0 20720.0 129595.0 ;
      RECT  20015.0 130940.0 20720.0 129595.0 ;
      RECT  20015.0 130940.0 20720.0 132285.0 ;
      RECT  20015.0 133630.0 20720.0 132285.0 ;
      RECT  20015.0 133630.0 20720.0 134975.0 ;
      RECT  20015.0 136320.0 20720.0 134975.0 ;
      RECT  20015.0 136320.0 20720.0 137665.0 ;
      RECT  20015.0 139010.0 20720.0 137665.0 ;
      RECT  20015.0 139010.0 20720.0 140355.0 ;
      RECT  20015.0 141700.0 20720.0 140355.0 ;
      RECT  20015.0 141700.0 20720.0 143045.0 ;
      RECT  20015.0 144390.0 20720.0 143045.0 ;
      RECT  20015.0 144390.0 20720.0 145735.0 ;
      RECT  20015.0 147080.0 20720.0 145735.0 ;
      RECT  20015.0 147080.0 20720.0 148425.0 ;
      RECT  20015.0 149770.0 20720.0 148425.0 ;
      RECT  20015.0 149770.0 20720.0 151115.0 ;
      RECT  20015.0 152460.0 20720.0 151115.0 ;
      RECT  20015.0 152460.0 20720.0 153805.0 ;
      RECT  20015.0 155150.0 20720.0 153805.0 ;
      RECT  20015.0 155150.0 20720.0 156495.0 ;
      RECT  20015.0 157840.0 20720.0 156495.0 ;
      RECT  20015.0 157840.0 20720.0 159185.0 ;
      RECT  20015.0 160530.0 20720.0 159185.0 ;
      RECT  20015.0 160530.0 20720.0 161875.0 ;
      RECT  20015.0 163220.0 20720.0 161875.0 ;
      RECT  20015.0 163220.0 20720.0 164565.0 ;
      RECT  20015.0 165910.0 20720.0 164565.0 ;
      RECT  20015.0 165910.0 20720.0 167255.0 ;
      RECT  20015.0 168600.0 20720.0 167255.0 ;
      RECT  20015.0 168600.0 20720.0 169945.0 ;
      RECT  20015.0 171290.0 20720.0 169945.0 ;
      RECT  20015.0 171290.0 20720.0 172635.0 ;
      RECT  20015.0 173980.0 20720.0 172635.0 ;
      RECT  20015.0 173980.0 20720.0 175325.0 ;
      RECT  20015.0 176670.0 20720.0 175325.0 ;
      RECT  20015.0 176670.0 20720.0 178015.0 ;
      RECT  20015.0 179360.0 20720.0 178015.0 ;
      RECT  20015.0 179360.0 20720.0 180705.0 ;
      RECT  20015.0 182050.0 20720.0 180705.0 ;
      RECT  20015.0 182050.0 20720.0 183395.0 ;
      RECT  20015.0 184740.0 20720.0 183395.0 ;
      RECT  20015.0 184740.0 20720.0 186085.0 ;
      RECT  20015.0 187430.0 20720.0 186085.0 ;
      RECT  20015.0 187430.0 20720.0 188775.0 ;
      RECT  20015.0 190120.0 20720.0 188775.0 ;
      RECT  20015.0 190120.0 20720.0 191465.0 ;
      RECT  20015.0 192810.0 20720.0 191465.0 ;
      RECT  20015.0 192810.0 20720.0 194155.0 ;
      RECT  20015.0 195500.0 20720.0 194155.0 ;
      RECT  20015.0 195500.0 20720.0 196845.0 ;
      RECT  20015.0 198190.0 20720.0 196845.0 ;
      RECT  20015.0 198190.0 20720.0 199535.0 ;
      RECT  20015.0 200880.0 20720.0 199535.0 ;
      RECT  20015.0 200880.0 20720.0 202225.0 ;
      RECT  20015.0 203570.0 20720.0 202225.0 ;
      RECT  20015.0 203570.0 20720.0 204915.0 ;
      RECT  20015.0 206260.0 20720.0 204915.0 ;
      RECT  20720.0 34100.0 21425.0 35445.0 ;
      RECT  20720.0 36790.0 21425.0 35445.0 ;
      RECT  20720.0 36790.0 21425.0 38135.0 ;
      RECT  20720.0 39480.0 21425.0 38135.0 ;
      RECT  20720.0 39480.0 21425.0 40825.0 ;
      RECT  20720.0 42170.0 21425.0 40825.0 ;
      RECT  20720.0 42170.0 21425.0 43515.0 ;
      RECT  20720.0 44860.0 21425.0 43515.0 ;
      RECT  20720.0 44860.0 21425.0 46205.0 ;
      RECT  20720.0 47550.0 21425.0 46205.0 ;
      RECT  20720.0 47550.0 21425.0 48895.0 ;
      RECT  20720.0 50240.0 21425.0 48895.0 ;
      RECT  20720.0 50240.0 21425.0 51585.0 ;
      RECT  20720.0 52930.0 21425.0 51585.0 ;
      RECT  20720.0 52930.0 21425.0 54275.0 ;
      RECT  20720.0 55620.0 21425.0 54275.0 ;
      RECT  20720.0 55620.0 21425.0 56965.0 ;
      RECT  20720.0 58310.0 21425.0 56965.0 ;
      RECT  20720.0 58310.0 21425.0 59655.0 ;
      RECT  20720.0 61000.0 21425.0 59655.0 ;
      RECT  20720.0 61000.0 21425.0 62345.0 ;
      RECT  20720.0 63690.0 21425.0 62345.0 ;
      RECT  20720.0 63690.0 21425.0 65035.0 ;
      RECT  20720.0 66380.0 21425.0 65035.0 ;
      RECT  20720.0 66380.0 21425.0 67725.0 ;
      RECT  20720.0 69070.0 21425.0 67725.0 ;
      RECT  20720.0 69070.0 21425.0 70415.0 ;
      RECT  20720.0 71760.0 21425.0 70415.0 ;
      RECT  20720.0 71760.0 21425.0 73105.0 ;
      RECT  20720.0 74450.0 21425.0 73105.0 ;
      RECT  20720.0 74450.0 21425.0 75795.0 ;
      RECT  20720.0 77140.0 21425.0 75795.0 ;
      RECT  20720.0 77140.0 21425.0 78485.0 ;
      RECT  20720.0 79830.0 21425.0 78485.0 ;
      RECT  20720.0 79830.0 21425.0 81175.0 ;
      RECT  20720.0 82520.0 21425.0 81175.0 ;
      RECT  20720.0 82520.0 21425.0 83865.0 ;
      RECT  20720.0 85210.0 21425.0 83865.0 ;
      RECT  20720.0 85210.0 21425.0 86555.0 ;
      RECT  20720.0 87900.0 21425.0 86555.0 ;
      RECT  20720.0 87900.0 21425.0 89245.0 ;
      RECT  20720.0 90590.0 21425.0 89245.0 ;
      RECT  20720.0 90590.0 21425.0 91935.0 ;
      RECT  20720.0 93280.0 21425.0 91935.0 ;
      RECT  20720.0 93280.0 21425.0 94625.0 ;
      RECT  20720.0 95970.0 21425.0 94625.0 ;
      RECT  20720.0 95970.0 21425.0 97315.0 ;
      RECT  20720.0 98660.0 21425.0 97315.0 ;
      RECT  20720.0 98660.0 21425.0 100005.0 ;
      RECT  20720.0 101350.0 21425.0 100005.0 ;
      RECT  20720.0 101350.0 21425.0 102695.0 ;
      RECT  20720.0 104040.0 21425.0 102695.0 ;
      RECT  20720.0 104040.0 21425.0 105385.0 ;
      RECT  20720.0 106730.0 21425.0 105385.0 ;
      RECT  20720.0 106730.0 21425.0 108075.0 ;
      RECT  20720.0 109420.0 21425.0 108075.0 ;
      RECT  20720.0 109420.0 21425.0 110765.0 ;
      RECT  20720.0 112110.0 21425.0 110765.0 ;
      RECT  20720.0 112110.0 21425.0 113455.0 ;
      RECT  20720.0 114800.0 21425.0 113455.0 ;
      RECT  20720.0 114800.0 21425.0 116145.0 ;
      RECT  20720.0 117490.0 21425.0 116145.0 ;
      RECT  20720.0 117490.0 21425.0 118835.0 ;
      RECT  20720.0 120180.0 21425.0 118835.0 ;
      RECT  20720.0 120180.0 21425.0 121525.0 ;
      RECT  20720.0 122870.0 21425.0 121525.0 ;
      RECT  20720.0 122870.0 21425.0 124215.0 ;
      RECT  20720.0 125560.0 21425.0 124215.0 ;
      RECT  20720.0 125560.0 21425.0 126905.0 ;
      RECT  20720.0 128250.0 21425.0 126905.0 ;
      RECT  20720.0 128250.0 21425.0 129595.0 ;
      RECT  20720.0 130940.0 21425.0 129595.0 ;
      RECT  20720.0 130940.0 21425.0 132285.0 ;
      RECT  20720.0 133630.0 21425.0 132285.0 ;
      RECT  20720.0 133630.0 21425.0 134975.0 ;
      RECT  20720.0 136320.0 21425.0 134975.0 ;
      RECT  20720.0 136320.0 21425.0 137665.0 ;
      RECT  20720.0 139010.0 21425.0 137665.0 ;
      RECT  20720.0 139010.0 21425.0 140355.0 ;
      RECT  20720.0 141700.0 21425.0 140355.0 ;
      RECT  20720.0 141700.0 21425.0 143045.0 ;
      RECT  20720.0 144390.0 21425.0 143045.0 ;
      RECT  20720.0 144390.0 21425.0 145735.0 ;
      RECT  20720.0 147080.0 21425.0 145735.0 ;
      RECT  20720.0 147080.0 21425.0 148425.0 ;
      RECT  20720.0 149770.0 21425.0 148425.0 ;
      RECT  20720.0 149770.0 21425.0 151115.0 ;
      RECT  20720.0 152460.0 21425.0 151115.0 ;
      RECT  20720.0 152460.0 21425.0 153805.0 ;
      RECT  20720.0 155150.0 21425.0 153805.0 ;
      RECT  20720.0 155150.0 21425.0 156495.0 ;
      RECT  20720.0 157840.0 21425.0 156495.0 ;
      RECT  20720.0 157840.0 21425.0 159185.0 ;
      RECT  20720.0 160530.0 21425.0 159185.0 ;
      RECT  20720.0 160530.0 21425.0 161875.0 ;
      RECT  20720.0 163220.0 21425.0 161875.0 ;
      RECT  20720.0 163220.0 21425.0 164565.0 ;
      RECT  20720.0 165910.0 21425.0 164565.0 ;
      RECT  20720.0 165910.0 21425.0 167255.0 ;
      RECT  20720.0 168600.0 21425.0 167255.0 ;
      RECT  20720.0 168600.0 21425.0 169945.0 ;
      RECT  20720.0 171290.0 21425.0 169945.0 ;
      RECT  20720.0 171290.0 21425.0 172635.0 ;
      RECT  20720.0 173980.0 21425.0 172635.0 ;
      RECT  20720.0 173980.0 21425.0 175325.0 ;
      RECT  20720.0 176670.0 21425.0 175325.0 ;
      RECT  20720.0 176670.0 21425.0 178015.0 ;
      RECT  20720.0 179360.0 21425.0 178015.0 ;
      RECT  20720.0 179360.0 21425.0 180705.0 ;
      RECT  20720.0 182050.0 21425.0 180705.0 ;
      RECT  20720.0 182050.0 21425.0 183395.0 ;
      RECT  20720.0 184740.0 21425.0 183395.0 ;
      RECT  20720.0 184740.0 21425.0 186085.0 ;
      RECT  20720.0 187430.0 21425.0 186085.0 ;
      RECT  20720.0 187430.0 21425.0 188775.0 ;
      RECT  20720.0 190120.0 21425.0 188775.0 ;
      RECT  20720.0 190120.0 21425.0 191465.0 ;
      RECT  20720.0 192810.0 21425.0 191465.0 ;
      RECT  20720.0 192810.0 21425.0 194155.0 ;
      RECT  20720.0 195500.0 21425.0 194155.0 ;
      RECT  20720.0 195500.0 21425.0 196845.0 ;
      RECT  20720.0 198190.0 21425.0 196845.0 ;
      RECT  20720.0 198190.0 21425.0 199535.0 ;
      RECT  20720.0 200880.0 21425.0 199535.0 ;
      RECT  20720.0 200880.0 21425.0 202225.0 ;
      RECT  20720.0 203570.0 21425.0 202225.0 ;
      RECT  20720.0 203570.0 21425.0 204915.0 ;
      RECT  20720.0 206260.0 21425.0 204915.0 ;
      RECT  21425.0 34100.0 22130.0 35445.0 ;
      RECT  21425.0 36790.0 22130.0 35445.0 ;
      RECT  21425.0 36790.0 22130.0 38135.0 ;
      RECT  21425.0 39480.0 22130.0 38135.0 ;
      RECT  21425.0 39480.0 22130.0 40825.0 ;
      RECT  21425.0 42170.0 22130.0 40825.0 ;
      RECT  21425.0 42170.0 22130.0 43515.0 ;
      RECT  21425.0 44860.0 22130.0 43515.0 ;
      RECT  21425.0 44860.0 22130.0 46205.0 ;
      RECT  21425.0 47550.0 22130.0 46205.0 ;
      RECT  21425.0 47550.0 22130.0 48895.0 ;
      RECT  21425.0 50240.0 22130.0 48895.0 ;
      RECT  21425.0 50240.0 22130.0 51585.0 ;
      RECT  21425.0 52930.0 22130.0 51585.0 ;
      RECT  21425.0 52930.0 22130.0 54275.0 ;
      RECT  21425.0 55620.0 22130.0 54275.0 ;
      RECT  21425.0 55620.0 22130.0 56965.0 ;
      RECT  21425.0 58310.0 22130.0 56965.0 ;
      RECT  21425.0 58310.0 22130.0 59655.0 ;
      RECT  21425.0 61000.0 22130.0 59655.0 ;
      RECT  21425.0 61000.0 22130.0 62345.0 ;
      RECT  21425.0 63690.0 22130.0 62345.0 ;
      RECT  21425.0 63690.0 22130.0 65035.0 ;
      RECT  21425.0 66380.0 22130.0 65035.0 ;
      RECT  21425.0 66380.0 22130.0 67725.0 ;
      RECT  21425.0 69070.0 22130.0 67725.0 ;
      RECT  21425.0 69070.0 22130.0 70415.0 ;
      RECT  21425.0 71760.0 22130.0 70415.0 ;
      RECT  21425.0 71760.0 22130.0 73105.0 ;
      RECT  21425.0 74450.0 22130.0 73105.0 ;
      RECT  21425.0 74450.0 22130.0 75795.0 ;
      RECT  21425.0 77140.0 22130.0 75795.0 ;
      RECT  21425.0 77140.0 22130.0 78485.0 ;
      RECT  21425.0 79830.0 22130.0 78485.0 ;
      RECT  21425.0 79830.0 22130.0 81175.0 ;
      RECT  21425.0 82520.0 22130.0 81175.0 ;
      RECT  21425.0 82520.0 22130.0 83865.0 ;
      RECT  21425.0 85210.0 22130.0 83865.0 ;
      RECT  21425.0 85210.0 22130.0 86555.0 ;
      RECT  21425.0 87900.0 22130.0 86555.0 ;
      RECT  21425.0 87900.0 22130.0 89245.0 ;
      RECT  21425.0 90590.0 22130.0 89245.0 ;
      RECT  21425.0 90590.0 22130.0 91935.0 ;
      RECT  21425.0 93280.0 22130.0 91935.0 ;
      RECT  21425.0 93280.0 22130.0 94625.0 ;
      RECT  21425.0 95970.0 22130.0 94625.0 ;
      RECT  21425.0 95970.0 22130.0 97315.0 ;
      RECT  21425.0 98660.0 22130.0 97315.0 ;
      RECT  21425.0 98660.0 22130.0 100005.0 ;
      RECT  21425.0 101350.0 22130.0 100005.0 ;
      RECT  21425.0 101350.0 22130.0 102695.0 ;
      RECT  21425.0 104040.0 22130.0 102695.0 ;
      RECT  21425.0 104040.0 22130.0 105385.0 ;
      RECT  21425.0 106730.0 22130.0 105385.0 ;
      RECT  21425.0 106730.0 22130.0 108075.0 ;
      RECT  21425.0 109420.0 22130.0 108075.0 ;
      RECT  21425.0 109420.0 22130.0 110765.0 ;
      RECT  21425.0 112110.0 22130.0 110765.0 ;
      RECT  21425.0 112110.0 22130.0 113455.0 ;
      RECT  21425.0 114800.0 22130.0 113455.0 ;
      RECT  21425.0 114800.0 22130.0 116145.0 ;
      RECT  21425.0 117490.0 22130.0 116145.0 ;
      RECT  21425.0 117490.0 22130.0 118835.0 ;
      RECT  21425.0 120180.0 22130.0 118835.0 ;
      RECT  21425.0 120180.0 22130.0 121525.0 ;
      RECT  21425.0 122870.0 22130.0 121525.0 ;
      RECT  21425.0 122870.0 22130.0 124215.0 ;
      RECT  21425.0 125560.0 22130.0 124215.0 ;
      RECT  21425.0 125560.0 22130.0 126905.0 ;
      RECT  21425.0 128250.0 22130.0 126905.0 ;
      RECT  21425.0 128250.0 22130.0 129595.0 ;
      RECT  21425.0 130940.0 22130.0 129595.0 ;
      RECT  21425.0 130940.0 22130.0 132285.0 ;
      RECT  21425.0 133630.0 22130.0 132285.0 ;
      RECT  21425.0 133630.0 22130.0 134975.0 ;
      RECT  21425.0 136320.0 22130.0 134975.0 ;
      RECT  21425.0 136320.0 22130.0 137665.0 ;
      RECT  21425.0 139010.0 22130.0 137665.0 ;
      RECT  21425.0 139010.0 22130.0 140355.0 ;
      RECT  21425.0 141700.0 22130.0 140355.0 ;
      RECT  21425.0 141700.0 22130.0 143045.0 ;
      RECT  21425.0 144390.0 22130.0 143045.0 ;
      RECT  21425.0 144390.0 22130.0 145735.0 ;
      RECT  21425.0 147080.0 22130.0 145735.0 ;
      RECT  21425.0 147080.0 22130.0 148425.0 ;
      RECT  21425.0 149770.0 22130.0 148425.0 ;
      RECT  21425.0 149770.0 22130.0 151115.0 ;
      RECT  21425.0 152460.0 22130.0 151115.0 ;
      RECT  21425.0 152460.0 22130.0 153805.0 ;
      RECT  21425.0 155150.0 22130.0 153805.0 ;
      RECT  21425.0 155150.0 22130.0 156495.0 ;
      RECT  21425.0 157840.0 22130.0 156495.0 ;
      RECT  21425.0 157840.0 22130.0 159185.0 ;
      RECT  21425.0 160530.0 22130.0 159185.0 ;
      RECT  21425.0 160530.0 22130.0 161875.0 ;
      RECT  21425.0 163220.0 22130.0 161875.0 ;
      RECT  21425.0 163220.0 22130.0 164565.0 ;
      RECT  21425.0 165910.0 22130.0 164565.0 ;
      RECT  21425.0 165910.0 22130.0 167255.0 ;
      RECT  21425.0 168600.0 22130.0 167255.0 ;
      RECT  21425.0 168600.0 22130.0 169945.0 ;
      RECT  21425.0 171290.0 22130.0 169945.0 ;
      RECT  21425.0 171290.0 22130.0 172635.0 ;
      RECT  21425.0 173980.0 22130.0 172635.0 ;
      RECT  21425.0 173980.0 22130.0 175325.0 ;
      RECT  21425.0 176670.0 22130.0 175325.0 ;
      RECT  21425.0 176670.0 22130.0 178015.0 ;
      RECT  21425.0 179360.0 22130.0 178015.0 ;
      RECT  21425.0 179360.0 22130.0 180705.0 ;
      RECT  21425.0 182050.0 22130.0 180705.0 ;
      RECT  21425.0 182050.0 22130.0 183395.0 ;
      RECT  21425.0 184740.0 22130.0 183395.0 ;
      RECT  21425.0 184740.0 22130.0 186085.0 ;
      RECT  21425.0 187430.0 22130.0 186085.0 ;
      RECT  21425.0 187430.0 22130.0 188775.0 ;
      RECT  21425.0 190120.0 22130.0 188775.0 ;
      RECT  21425.0 190120.0 22130.0 191465.0 ;
      RECT  21425.0 192810.0 22130.0 191465.0 ;
      RECT  21425.0 192810.0 22130.0 194155.0 ;
      RECT  21425.0 195500.0 22130.0 194155.0 ;
      RECT  21425.0 195500.0 22130.0 196845.0 ;
      RECT  21425.0 198190.0 22130.0 196845.0 ;
      RECT  21425.0 198190.0 22130.0 199535.0 ;
      RECT  21425.0 200880.0 22130.0 199535.0 ;
      RECT  21425.0 200880.0 22130.0 202225.0 ;
      RECT  21425.0 203570.0 22130.0 202225.0 ;
      RECT  21425.0 203570.0 22130.0 204915.0 ;
      RECT  21425.0 206260.0 22130.0 204915.0 ;
      RECT  22130.0 34100.0 22835.0 35445.0 ;
      RECT  22130.0 36790.0 22835.0 35445.0 ;
      RECT  22130.0 36790.0 22835.0 38135.0 ;
      RECT  22130.0 39480.0 22835.0 38135.0 ;
      RECT  22130.0 39480.0 22835.0 40825.0 ;
      RECT  22130.0 42170.0 22835.0 40825.0 ;
      RECT  22130.0 42170.0 22835.0 43515.0 ;
      RECT  22130.0 44860.0 22835.0 43515.0 ;
      RECT  22130.0 44860.0 22835.0 46205.0 ;
      RECT  22130.0 47550.0 22835.0 46205.0 ;
      RECT  22130.0 47550.0 22835.0 48895.0 ;
      RECT  22130.0 50240.0 22835.0 48895.0 ;
      RECT  22130.0 50240.0 22835.0 51585.0 ;
      RECT  22130.0 52930.0 22835.0 51585.0 ;
      RECT  22130.0 52930.0 22835.0 54275.0 ;
      RECT  22130.0 55620.0 22835.0 54275.0 ;
      RECT  22130.0 55620.0 22835.0 56965.0 ;
      RECT  22130.0 58310.0 22835.0 56965.0 ;
      RECT  22130.0 58310.0 22835.0 59655.0 ;
      RECT  22130.0 61000.0 22835.0 59655.0 ;
      RECT  22130.0 61000.0 22835.0 62345.0 ;
      RECT  22130.0 63690.0 22835.0 62345.0 ;
      RECT  22130.0 63690.0 22835.0 65035.0 ;
      RECT  22130.0 66380.0 22835.0 65035.0 ;
      RECT  22130.0 66380.0 22835.0 67725.0 ;
      RECT  22130.0 69070.0 22835.0 67725.0 ;
      RECT  22130.0 69070.0 22835.0 70415.0 ;
      RECT  22130.0 71760.0 22835.0 70415.0 ;
      RECT  22130.0 71760.0 22835.0 73105.0 ;
      RECT  22130.0 74450.0 22835.0 73105.0 ;
      RECT  22130.0 74450.0 22835.0 75795.0 ;
      RECT  22130.0 77140.0 22835.0 75795.0 ;
      RECT  22130.0 77140.0 22835.0 78485.0 ;
      RECT  22130.0 79830.0 22835.0 78485.0 ;
      RECT  22130.0 79830.0 22835.0 81175.0 ;
      RECT  22130.0 82520.0 22835.0 81175.0 ;
      RECT  22130.0 82520.0 22835.0 83865.0 ;
      RECT  22130.0 85210.0 22835.0 83865.0 ;
      RECT  22130.0 85210.0 22835.0 86555.0 ;
      RECT  22130.0 87900.0 22835.0 86555.0 ;
      RECT  22130.0 87900.0 22835.0 89245.0 ;
      RECT  22130.0 90590.0 22835.0 89245.0 ;
      RECT  22130.0 90590.0 22835.0 91935.0 ;
      RECT  22130.0 93280.0 22835.0 91935.0 ;
      RECT  22130.0 93280.0 22835.0 94625.0 ;
      RECT  22130.0 95970.0 22835.0 94625.0 ;
      RECT  22130.0 95970.0 22835.0 97315.0 ;
      RECT  22130.0 98660.0 22835.0 97315.0 ;
      RECT  22130.0 98660.0 22835.0 100005.0 ;
      RECT  22130.0 101350.0 22835.0 100005.0 ;
      RECT  22130.0 101350.0 22835.0 102695.0 ;
      RECT  22130.0 104040.0 22835.0 102695.0 ;
      RECT  22130.0 104040.0 22835.0 105385.0 ;
      RECT  22130.0 106730.0 22835.0 105385.0 ;
      RECT  22130.0 106730.0 22835.0 108075.0 ;
      RECT  22130.0 109420.0 22835.0 108075.0 ;
      RECT  22130.0 109420.0 22835.0 110765.0 ;
      RECT  22130.0 112110.0 22835.0 110765.0 ;
      RECT  22130.0 112110.0 22835.0 113455.0 ;
      RECT  22130.0 114800.0 22835.0 113455.0 ;
      RECT  22130.0 114800.0 22835.0 116145.0 ;
      RECT  22130.0 117490.0 22835.0 116145.0 ;
      RECT  22130.0 117490.0 22835.0 118835.0 ;
      RECT  22130.0 120180.0 22835.0 118835.0 ;
      RECT  22130.0 120180.0 22835.0 121525.0 ;
      RECT  22130.0 122870.0 22835.0 121525.0 ;
      RECT  22130.0 122870.0 22835.0 124215.0 ;
      RECT  22130.0 125560.0 22835.0 124215.0 ;
      RECT  22130.0 125560.0 22835.0 126905.0 ;
      RECT  22130.0 128250.0 22835.0 126905.0 ;
      RECT  22130.0 128250.0 22835.0 129595.0 ;
      RECT  22130.0 130940.0 22835.0 129595.0 ;
      RECT  22130.0 130940.0 22835.0 132285.0 ;
      RECT  22130.0 133630.0 22835.0 132285.0 ;
      RECT  22130.0 133630.0 22835.0 134975.0 ;
      RECT  22130.0 136320.0 22835.0 134975.0 ;
      RECT  22130.0 136320.0 22835.0 137665.0 ;
      RECT  22130.0 139010.0 22835.0 137665.0 ;
      RECT  22130.0 139010.0 22835.0 140355.0 ;
      RECT  22130.0 141700.0 22835.0 140355.0 ;
      RECT  22130.0 141700.0 22835.0 143045.0 ;
      RECT  22130.0 144390.0 22835.0 143045.0 ;
      RECT  22130.0 144390.0 22835.0 145735.0 ;
      RECT  22130.0 147080.0 22835.0 145735.0 ;
      RECT  22130.0 147080.0 22835.0 148425.0 ;
      RECT  22130.0 149770.0 22835.0 148425.0 ;
      RECT  22130.0 149770.0 22835.0 151115.0 ;
      RECT  22130.0 152460.0 22835.0 151115.0 ;
      RECT  22130.0 152460.0 22835.0 153805.0 ;
      RECT  22130.0 155150.0 22835.0 153805.0 ;
      RECT  22130.0 155150.0 22835.0 156495.0 ;
      RECT  22130.0 157840.0 22835.0 156495.0 ;
      RECT  22130.0 157840.0 22835.0 159185.0 ;
      RECT  22130.0 160530.0 22835.0 159185.0 ;
      RECT  22130.0 160530.0 22835.0 161875.0 ;
      RECT  22130.0 163220.0 22835.0 161875.0 ;
      RECT  22130.0 163220.0 22835.0 164565.0 ;
      RECT  22130.0 165910.0 22835.0 164565.0 ;
      RECT  22130.0 165910.0 22835.0 167255.0 ;
      RECT  22130.0 168600.0 22835.0 167255.0 ;
      RECT  22130.0 168600.0 22835.0 169945.0 ;
      RECT  22130.0 171290.0 22835.0 169945.0 ;
      RECT  22130.0 171290.0 22835.0 172635.0 ;
      RECT  22130.0 173980.0 22835.0 172635.0 ;
      RECT  22130.0 173980.0 22835.0 175325.0 ;
      RECT  22130.0 176670.0 22835.0 175325.0 ;
      RECT  22130.0 176670.0 22835.0 178015.0 ;
      RECT  22130.0 179360.0 22835.0 178015.0 ;
      RECT  22130.0 179360.0 22835.0 180705.0 ;
      RECT  22130.0 182050.0 22835.0 180705.0 ;
      RECT  22130.0 182050.0 22835.0 183395.0 ;
      RECT  22130.0 184740.0 22835.0 183395.0 ;
      RECT  22130.0 184740.0 22835.0 186085.0 ;
      RECT  22130.0 187430.0 22835.0 186085.0 ;
      RECT  22130.0 187430.0 22835.0 188775.0 ;
      RECT  22130.0 190120.0 22835.0 188775.0 ;
      RECT  22130.0 190120.0 22835.0 191465.0 ;
      RECT  22130.0 192810.0 22835.0 191465.0 ;
      RECT  22130.0 192810.0 22835.0 194155.0 ;
      RECT  22130.0 195500.0 22835.0 194155.0 ;
      RECT  22130.0 195500.0 22835.0 196845.0 ;
      RECT  22130.0 198190.0 22835.0 196845.0 ;
      RECT  22130.0 198190.0 22835.0 199535.0 ;
      RECT  22130.0 200880.0 22835.0 199535.0 ;
      RECT  22130.0 200880.0 22835.0 202225.0 ;
      RECT  22130.0 203570.0 22835.0 202225.0 ;
      RECT  22130.0 203570.0 22835.0 204915.0 ;
      RECT  22130.0 206260.0 22835.0 204915.0 ;
      RECT  22835.0 34100.0 23540.0 35445.0 ;
      RECT  22835.0 36790.0 23540.0 35445.0 ;
      RECT  22835.0 36790.0 23540.0 38135.0 ;
      RECT  22835.0 39480.0 23540.0 38135.0 ;
      RECT  22835.0 39480.0 23540.0 40825.0 ;
      RECT  22835.0 42170.0 23540.0 40825.0 ;
      RECT  22835.0 42170.0 23540.0 43515.0 ;
      RECT  22835.0 44860.0 23540.0 43515.0 ;
      RECT  22835.0 44860.0 23540.0 46205.0 ;
      RECT  22835.0 47550.0 23540.0 46205.0 ;
      RECT  22835.0 47550.0 23540.0 48895.0 ;
      RECT  22835.0 50240.0 23540.0 48895.0 ;
      RECT  22835.0 50240.0 23540.0 51585.0 ;
      RECT  22835.0 52930.0 23540.0 51585.0 ;
      RECT  22835.0 52930.0 23540.0 54275.0 ;
      RECT  22835.0 55620.0 23540.0 54275.0 ;
      RECT  22835.0 55620.0 23540.0 56965.0 ;
      RECT  22835.0 58310.0 23540.0 56965.0 ;
      RECT  22835.0 58310.0 23540.0 59655.0 ;
      RECT  22835.0 61000.0 23540.0 59655.0 ;
      RECT  22835.0 61000.0 23540.0 62345.0 ;
      RECT  22835.0 63690.0 23540.0 62345.0 ;
      RECT  22835.0 63690.0 23540.0 65035.0 ;
      RECT  22835.0 66380.0 23540.0 65035.0 ;
      RECT  22835.0 66380.0 23540.0 67725.0 ;
      RECT  22835.0 69070.0 23540.0 67725.0 ;
      RECT  22835.0 69070.0 23540.0 70415.0 ;
      RECT  22835.0 71760.0 23540.0 70415.0 ;
      RECT  22835.0 71760.0 23540.0 73105.0 ;
      RECT  22835.0 74450.0 23540.0 73105.0 ;
      RECT  22835.0 74450.0 23540.0 75795.0 ;
      RECT  22835.0 77140.0 23540.0 75795.0 ;
      RECT  22835.0 77140.0 23540.0 78485.0 ;
      RECT  22835.0 79830.0 23540.0 78485.0 ;
      RECT  22835.0 79830.0 23540.0 81175.0 ;
      RECT  22835.0 82520.0 23540.0 81175.0 ;
      RECT  22835.0 82520.0 23540.0 83865.0 ;
      RECT  22835.0 85210.0 23540.0 83865.0 ;
      RECT  22835.0 85210.0 23540.0 86555.0 ;
      RECT  22835.0 87900.0 23540.0 86555.0 ;
      RECT  22835.0 87900.0 23540.0 89245.0 ;
      RECT  22835.0 90590.0 23540.0 89245.0 ;
      RECT  22835.0 90590.0 23540.0 91935.0 ;
      RECT  22835.0 93280.0 23540.0 91935.0 ;
      RECT  22835.0 93280.0 23540.0 94625.0 ;
      RECT  22835.0 95970.0 23540.0 94625.0 ;
      RECT  22835.0 95970.0 23540.0 97315.0 ;
      RECT  22835.0 98660.0 23540.0 97315.0 ;
      RECT  22835.0 98660.0 23540.0 100005.0 ;
      RECT  22835.0 101350.0 23540.0 100005.0 ;
      RECT  22835.0 101350.0 23540.0 102695.0 ;
      RECT  22835.0 104040.0 23540.0 102695.0 ;
      RECT  22835.0 104040.0 23540.0 105385.0 ;
      RECT  22835.0 106730.0 23540.0 105385.0 ;
      RECT  22835.0 106730.0 23540.0 108075.0 ;
      RECT  22835.0 109420.0 23540.0 108075.0 ;
      RECT  22835.0 109420.0 23540.0 110765.0 ;
      RECT  22835.0 112110.0 23540.0 110765.0 ;
      RECT  22835.0 112110.0 23540.0 113455.0 ;
      RECT  22835.0 114800.0 23540.0 113455.0 ;
      RECT  22835.0 114800.0 23540.0 116145.0 ;
      RECT  22835.0 117490.0 23540.0 116145.0 ;
      RECT  22835.0 117490.0 23540.0 118835.0 ;
      RECT  22835.0 120180.0 23540.0 118835.0 ;
      RECT  22835.0 120180.0 23540.0 121525.0 ;
      RECT  22835.0 122870.0 23540.0 121525.0 ;
      RECT  22835.0 122870.0 23540.0 124215.0 ;
      RECT  22835.0 125560.0 23540.0 124215.0 ;
      RECT  22835.0 125560.0 23540.0 126905.0 ;
      RECT  22835.0 128250.0 23540.0 126905.0 ;
      RECT  22835.0 128250.0 23540.0 129595.0 ;
      RECT  22835.0 130940.0 23540.0 129595.0 ;
      RECT  22835.0 130940.0 23540.0 132285.0 ;
      RECT  22835.0 133630.0 23540.0 132285.0 ;
      RECT  22835.0 133630.0 23540.0 134975.0 ;
      RECT  22835.0 136320.0 23540.0 134975.0 ;
      RECT  22835.0 136320.0 23540.0 137665.0 ;
      RECT  22835.0 139010.0 23540.0 137665.0 ;
      RECT  22835.0 139010.0 23540.0 140355.0 ;
      RECT  22835.0 141700.0 23540.0 140355.0 ;
      RECT  22835.0 141700.0 23540.0 143045.0 ;
      RECT  22835.0 144390.0 23540.0 143045.0 ;
      RECT  22835.0 144390.0 23540.0 145735.0 ;
      RECT  22835.0 147080.0 23540.0 145735.0 ;
      RECT  22835.0 147080.0 23540.0 148425.0 ;
      RECT  22835.0 149770.0 23540.0 148425.0 ;
      RECT  22835.0 149770.0 23540.0 151115.0 ;
      RECT  22835.0 152460.0 23540.0 151115.0 ;
      RECT  22835.0 152460.0 23540.0 153805.0 ;
      RECT  22835.0 155150.0 23540.0 153805.0 ;
      RECT  22835.0 155150.0 23540.0 156495.0 ;
      RECT  22835.0 157840.0 23540.0 156495.0 ;
      RECT  22835.0 157840.0 23540.0 159185.0 ;
      RECT  22835.0 160530.0 23540.0 159185.0 ;
      RECT  22835.0 160530.0 23540.0 161875.0 ;
      RECT  22835.0 163220.0 23540.0 161875.0 ;
      RECT  22835.0 163220.0 23540.0 164565.0 ;
      RECT  22835.0 165910.0 23540.0 164565.0 ;
      RECT  22835.0 165910.0 23540.0 167255.0 ;
      RECT  22835.0 168600.0 23540.0 167255.0 ;
      RECT  22835.0 168600.0 23540.0 169945.0 ;
      RECT  22835.0 171290.0 23540.0 169945.0 ;
      RECT  22835.0 171290.0 23540.0 172635.0 ;
      RECT  22835.0 173980.0 23540.0 172635.0 ;
      RECT  22835.0 173980.0 23540.0 175325.0 ;
      RECT  22835.0 176670.0 23540.0 175325.0 ;
      RECT  22835.0 176670.0 23540.0 178015.0 ;
      RECT  22835.0 179360.0 23540.0 178015.0 ;
      RECT  22835.0 179360.0 23540.0 180705.0 ;
      RECT  22835.0 182050.0 23540.0 180705.0 ;
      RECT  22835.0 182050.0 23540.0 183395.0 ;
      RECT  22835.0 184740.0 23540.0 183395.0 ;
      RECT  22835.0 184740.0 23540.0 186085.0 ;
      RECT  22835.0 187430.0 23540.0 186085.0 ;
      RECT  22835.0 187430.0 23540.0 188775.0 ;
      RECT  22835.0 190120.0 23540.0 188775.0 ;
      RECT  22835.0 190120.0 23540.0 191465.0 ;
      RECT  22835.0 192810.0 23540.0 191465.0 ;
      RECT  22835.0 192810.0 23540.0 194155.0 ;
      RECT  22835.0 195500.0 23540.0 194155.0 ;
      RECT  22835.0 195500.0 23540.0 196845.0 ;
      RECT  22835.0 198190.0 23540.0 196845.0 ;
      RECT  22835.0 198190.0 23540.0 199535.0 ;
      RECT  22835.0 200880.0 23540.0 199535.0 ;
      RECT  22835.0 200880.0 23540.0 202225.0 ;
      RECT  22835.0 203570.0 23540.0 202225.0 ;
      RECT  22835.0 203570.0 23540.0 204915.0 ;
      RECT  22835.0 206260.0 23540.0 204915.0 ;
      RECT  23540.0 34100.0 24245.0 35445.0 ;
      RECT  23540.0 36790.0 24245.0 35445.0 ;
      RECT  23540.0 36790.0 24245.0 38135.0 ;
      RECT  23540.0 39480.0 24245.0 38135.0 ;
      RECT  23540.0 39480.0 24245.0 40825.0 ;
      RECT  23540.0 42170.0 24245.0 40825.0 ;
      RECT  23540.0 42170.0 24245.0 43515.0 ;
      RECT  23540.0 44860.0 24245.0 43515.0 ;
      RECT  23540.0 44860.0 24245.0 46205.0 ;
      RECT  23540.0 47550.0 24245.0 46205.0 ;
      RECT  23540.0 47550.0 24245.0 48895.0 ;
      RECT  23540.0 50240.0 24245.0 48895.0 ;
      RECT  23540.0 50240.0 24245.0 51585.0 ;
      RECT  23540.0 52930.0 24245.0 51585.0 ;
      RECT  23540.0 52930.0 24245.0 54275.0 ;
      RECT  23540.0 55620.0 24245.0 54275.0 ;
      RECT  23540.0 55620.0 24245.0 56965.0 ;
      RECT  23540.0 58310.0 24245.0 56965.0 ;
      RECT  23540.0 58310.0 24245.0 59655.0 ;
      RECT  23540.0 61000.0 24245.0 59655.0 ;
      RECT  23540.0 61000.0 24245.0 62345.0 ;
      RECT  23540.0 63690.0 24245.0 62345.0 ;
      RECT  23540.0 63690.0 24245.0 65035.0 ;
      RECT  23540.0 66380.0 24245.0 65035.0 ;
      RECT  23540.0 66380.0 24245.0 67725.0 ;
      RECT  23540.0 69070.0 24245.0 67725.0 ;
      RECT  23540.0 69070.0 24245.0 70415.0 ;
      RECT  23540.0 71760.0 24245.0 70415.0 ;
      RECT  23540.0 71760.0 24245.0 73105.0 ;
      RECT  23540.0 74450.0 24245.0 73105.0 ;
      RECT  23540.0 74450.0 24245.0 75795.0 ;
      RECT  23540.0 77140.0 24245.0 75795.0 ;
      RECT  23540.0 77140.0 24245.0 78485.0 ;
      RECT  23540.0 79830.0 24245.0 78485.0 ;
      RECT  23540.0 79830.0 24245.0 81175.0 ;
      RECT  23540.0 82520.0 24245.0 81175.0 ;
      RECT  23540.0 82520.0 24245.0 83865.0 ;
      RECT  23540.0 85210.0 24245.0 83865.0 ;
      RECT  23540.0 85210.0 24245.0 86555.0 ;
      RECT  23540.0 87900.0 24245.0 86555.0 ;
      RECT  23540.0 87900.0 24245.0 89245.0 ;
      RECT  23540.0 90590.0 24245.0 89245.0 ;
      RECT  23540.0 90590.0 24245.0 91935.0 ;
      RECT  23540.0 93280.0 24245.0 91935.0 ;
      RECT  23540.0 93280.0 24245.0 94625.0 ;
      RECT  23540.0 95970.0 24245.0 94625.0 ;
      RECT  23540.0 95970.0 24245.0 97315.0 ;
      RECT  23540.0 98660.0 24245.0 97315.0 ;
      RECT  23540.0 98660.0 24245.0 100005.0 ;
      RECT  23540.0 101350.0 24245.0 100005.0 ;
      RECT  23540.0 101350.0 24245.0 102695.0 ;
      RECT  23540.0 104040.0 24245.0 102695.0 ;
      RECT  23540.0 104040.0 24245.0 105385.0 ;
      RECT  23540.0 106730.0 24245.0 105385.0 ;
      RECT  23540.0 106730.0 24245.0 108075.0 ;
      RECT  23540.0 109420.0 24245.0 108075.0 ;
      RECT  23540.0 109420.0 24245.0 110765.0 ;
      RECT  23540.0 112110.0 24245.0 110765.0 ;
      RECT  23540.0 112110.0 24245.0 113455.0 ;
      RECT  23540.0 114800.0 24245.0 113455.0 ;
      RECT  23540.0 114800.0 24245.0 116145.0 ;
      RECT  23540.0 117490.0 24245.0 116145.0 ;
      RECT  23540.0 117490.0 24245.0 118835.0 ;
      RECT  23540.0 120180.0 24245.0 118835.0 ;
      RECT  23540.0 120180.0 24245.0 121525.0 ;
      RECT  23540.0 122870.0 24245.0 121525.0 ;
      RECT  23540.0 122870.0 24245.0 124215.0 ;
      RECT  23540.0 125560.0 24245.0 124215.0 ;
      RECT  23540.0 125560.0 24245.0 126905.0 ;
      RECT  23540.0 128250.0 24245.0 126905.0 ;
      RECT  23540.0 128250.0 24245.0 129595.0 ;
      RECT  23540.0 130940.0 24245.0 129595.0 ;
      RECT  23540.0 130940.0 24245.0 132285.0 ;
      RECT  23540.0 133630.0 24245.0 132285.0 ;
      RECT  23540.0 133630.0 24245.0 134975.0 ;
      RECT  23540.0 136320.0 24245.0 134975.0 ;
      RECT  23540.0 136320.0 24245.0 137665.0 ;
      RECT  23540.0 139010.0 24245.0 137665.0 ;
      RECT  23540.0 139010.0 24245.0 140355.0 ;
      RECT  23540.0 141700.0 24245.0 140355.0 ;
      RECT  23540.0 141700.0 24245.0 143045.0 ;
      RECT  23540.0 144390.0 24245.0 143045.0 ;
      RECT  23540.0 144390.0 24245.0 145735.0 ;
      RECT  23540.0 147080.0 24245.0 145735.0 ;
      RECT  23540.0 147080.0 24245.0 148425.0 ;
      RECT  23540.0 149770.0 24245.0 148425.0 ;
      RECT  23540.0 149770.0 24245.0 151115.0 ;
      RECT  23540.0 152460.0 24245.0 151115.0 ;
      RECT  23540.0 152460.0 24245.0 153805.0 ;
      RECT  23540.0 155150.0 24245.0 153805.0 ;
      RECT  23540.0 155150.0 24245.0 156495.0 ;
      RECT  23540.0 157840.0 24245.0 156495.0 ;
      RECT  23540.0 157840.0 24245.0 159185.0 ;
      RECT  23540.0 160530.0 24245.0 159185.0 ;
      RECT  23540.0 160530.0 24245.0 161875.0 ;
      RECT  23540.0 163220.0 24245.0 161875.0 ;
      RECT  23540.0 163220.0 24245.0 164565.0 ;
      RECT  23540.0 165910.0 24245.0 164565.0 ;
      RECT  23540.0 165910.0 24245.0 167255.0 ;
      RECT  23540.0 168600.0 24245.0 167255.0 ;
      RECT  23540.0 168600.0 24245.0 169945.0 ;
      RECT  23540.0 171290.0 24245.0 169945.0 ;
      RECT  23540.0 171290.0 24245.0 172635.0 ;
      RECT  23540.0 173980.0 24245.0 172635.0 ;
      RECT  23540.0 173980.0 24245.0 175325.0 ;
      RECT  23540.0 176670.0 24245.0 175325.0 ;
      RECT  23540.0 176670.0 24245.0 178015.0 ;
      RECT  23540.0 179360.0 24245.0 178015.0 ;
      RECT  23540.0 179360.0 24245.0 180705.0 ;
      RECT  23540.0 182050.0 24245.0 180705.0 ;
      RECT  23540.0 182050.0 24245.0 183395.0 ;
      RECT  23540.0 184740.0 24245.0 183395.0 ;
      RECT  23540.0 184740.0 24245.0 186085.0 ;
      RECT  23540.0 187430.0 24245.0 186085.0 ;
      RECT  23540.0 187430.0 24245.0 188775.0 ;
      RECT  23540.0 190120.0 24245.0 188775.0 ;
      RECT  23540.0 190120.0 24245.0 191465.0 ;
      RECT  23540.0 192810.0 24245.0 191465.0 ;
      RECT  23540.0 192810.0 24245.0 194155.0 ;
      RECT  23540.0 195500.0 24245.0 194155.0 ;
      RECT  23540.0 195500.0 24245.0 196845.0 ;
      RECT  23540.0 198190.0 24245.0 196845.0 ;
      RECT  23540.0 198190.0 24245.0 199535.0 ;
      RECT  23540.0 200880.0 24245.0 199535.0 ;
      RECT  23540.0 200880.0 24245.0 202225.0 ;
      RECT  23540.0 203570.0 24245.0 202225.0 ;
      RECT  23540.0 203570.0 24245.0 204915.0 ;
      RECT  23540.0 206260.0 24245.0 204915.0 ;
      RECT  24245.0 34100.0 24950.0 35445.0 ;
      RECT  24245.0 36790.0 24950.0 35445.0 ;
      RECT  24245.0 36790.0 24950.0 38135.0 ;
      RECT  24245.0 39480.0 24950.0 38135.0 ;
      RECT  24245.0 39480.0 24950.0 40825.0 ;
      RECT  24245.0 42170.0 24950.0 40825.0 ;
      RECT  24245.0 42170.0 24950.0 43515.0 ;
      RECT  24245.0 44860.0 24950.0 43515.0 ;
      RECT  24245.0 44860.0 24950.0 46205.0 ;
      RECT  24245.0 47550.0 24950.0 46205.0 ;
      RECT  24245.0 47550.0 24950.0 48895.0 ;
      RECT  24245.0 50240.0 24950.0 48895.0 ;
      RECT  24245.0 50240.0 24950.0 51585.0 ;
      RECT  24245.0 52930.0 24950.0 51585.0 ;
      RECT  24245.0 52930.0 24950.0 54275.0 ;
      RECT  24245.0 55620.0 24950.0 54275.0 ;
      RECT  24245.0 55620.0 24950.0 56965.0 ;
      RECT  24245.0 58310.0 24950.0 56965.0 ;
      RECT  24245.0 58310.0 24950.0 59655.0 ;
      RECT  24245.0 61000.0 24950.0 59655.0 ;
      RECT  24245.0 61000.0 24950.0 62345.0 ;
      RECT  24245.0 63690.0 24950.0 62345.0 ;
      RECT  24245.0 63690.0 24950.0 65035.0 ;
      RECT  24245.0 66380.0 24950.0 65035.0 ;
      RECT  24245.0 66380.0 24950.0 67725.0 ;
      RECT  24245.0 69070.0 24950.0 67725.0 ;
      RECT  24245.0 69070.0 24950.0 70415.0 ;
      RECT  24245.0 71760.0 24950.0 70415.0 ;
      RECT  24245.0 71760.0 24950.0 73105.0 ;
      RECT  24245.0 74450.0 24950.0 73105.0 ;
      RECT  24245.0 74450.0 24950.0 75795.0 ;
      RECT  24245.0 77140.0 24950.0 75795.0 ;
      RECT  24245.0 77140.0 24950.0 78485.0 ;
      RECT  24245.0 79830.0 24950.0 78485.0 ;
      RECT  24245.0 79830.0 24950.0 81175.0 ;
      RECT  24245.0 82520.0 24950.0 81175.0 ;
      RECT  24245.0 82520.0 24950.0 83865.0 ;
      RECT  24245.0 85210.0 24950.0 83865.0 ;
      RECT  24245.0 85210.0 24950.0 86555.0 ;
      RECT  24245.0 87900.0 24950.0 86555.0 ;
      RECT  24245.0 87900.0 24950.0 89245.0 ;
      RECT  24245.0 90590.0 24950.0 89245.0 ;
      RECT  24245.0 90590.0 24950.0 91935.0 ;
      RECT  24245.0 93280.0 24950.0 91935.0 ;
      RECT  24245.0 93280.0 24950.0 94625.0 ;
      RECT  24245.0 95970.0 24950.0 94625.0 ;
      RECT  24245.0 95970.0 24950.0 97315.0 ;
      RECT  24245.0 98660.0 24950.0 97315.0 ;
      RECT  24245.0 98660.0 24950.0 100005.0 ;
      RECT  24245.0 101350.0 24950.0 100005.0 ;
      RECT  24245.0 101350.0 24950.0 102695.0 ;
      RECT  24245.0 104040.0 24950.0 102695.0 ;
      RECT  24245.0 104040.0 24950.0 105385.0 ;
      RECT  24245.0 106730.0 24950.0 105385.0 ;
      RECT  24245.0 106730.0 24950.0 108075.0 ;
      RECT  24245.0 109420.0 24950.0 108075.0 ;
      RECT  24245.0 109420.0 24950.0 110765.0 ;
      RECT  24245.0 112110.0 24950.0 110765.0 ;
      RECT  24245.0 112110.0 24950.0 113455.0 ;
      RECT  24245.0 114800.0 24950.0 113455.0 ;
      RECT  24245.0 114800.0 24950.0 116145.0 ;
      RECT  24245.0 117490.0 24950.0 116145.0 ;
      RECT  24245.0 117490.0 24950.0 118835.0 ;
      RECT  24245.0 120180.0 24950.0 118835.0 ;
      RECT  24245.0 120180.0 24950.0 121525.0 ;
      RECT  24245.0 122870.0 24950.0 121525.0 ;
      RECT  24245.0 122870.0 24950.0 124215.0 ;
      RECT  24245.0 125560.0 24950.0 124215.0 ;
      RECT  24245.0 125560.0 24950.0 126905.0 ;
      RECT  24245.0 128250.0 24950.0 126905.0 ;
      RECT  24245.0 128250.0 24950.0 129595.0 ;
      RECT  24245.0 130940.0 24950.0 129595.0 ;
      RECT  24245.0 130940.0 24950.0 132285.0 ;
      RECT  24245.0 133630.0 24950.0 132285.0 ;
      RECT  24245.0 133630.0 24950.0 134975.0 ;
      RECT  24245.0 136320.0 24950.0 134975.0 ;
      RECT  24245.0 136320.0 24950.0 137665.0 ;
      RECT  24245.0 139010.0 24950.0 137665.0 ;
      RECT  24245.0 139010.0 24950.0 140355.0 ;
      RECT  24245.0 141700.0 24950.0 140355.0 ;
      RECT  24245.0 141700.0 24950.0 143045.0 ;
      RECT  24245.0 144390.0 24950.0 143045.0 ;
      RECT  24245.0 144390.0 24950.0 145735.0 ;
      RECT  24245.0 147080.0 24950.0 145735.0 ;
      RECT  24245.0 147080.0 24950.0 148425.0 ;
      RECT  24245.0 149770.0 24950.0 148425.0 ;
      RECT  24245.0 149770.0 24950.0 151115.0 ;
      RECT  24245.0 152460.0 24950.0 151115.0 ;
      RECT  24245.0 152460.0 24950.0 153805.0 ;
      RECT  24245.0 155150.0 24950.0 153805.0 ;
      RECT  24245.0 155150.0 24950.0 156495.0 ;
      RECT  24245.0 157840.0 24950.0 156495.0 ;
      RECT  24245.0 157840.0 24950.0 159185.0 ;
      RECT  24245.0 160530.0 24950.0 159185.0 ;
      RECT  24245.0 160530.0 24950.0 161875.0 ;
      RECT  24245.0 163220.0 24950.0 161875.0 ;
      RECT  24245.0 163220.0 24950.0 164565.0 ;
      RECT  24245.0 165910.0 24950.0 164565.0 ;
      RECT  24245.0 165910.0 24950.0 167255.0 ;
      RECT  24245.0 168600.0 24950.0 167255.0 ;
      RECT  24245.0 168600.0 24950.0 169945.0 ;
      RECT  24245.0 171290.0 24950.0 169945.0 ;
      RECT  24245.0 171290.0 24950.0 172635.0 ;
      RECT  24245.0 173980.0 24950.0 172635.0 ;
      RECT  24245.0 173980.0 24950.0 175325.0 ;
      RECT  24245.0 176670.0 24950.0 175325.0 ;
      RECT  24245.0 176670.0 24950.0 178015.0 ;
      RECT  24245.0 179360.0 24950.0 178015.0 ;
      RECT  24245.0 179360.0 24950.0 180705.0 ;
      RECT  24245.0 182050.0 24950.0 180705.0 ;
      RECT  24245.0 182050.0 24950.0 183395.0 ;
      RECT  24245.0 184740.0 24950.0 183395.0 ;
      RECT  24245.0 184740.0 24950.0 186085.0 ;
      RECT  24245.0 187430.0 24950.0 186085.0 ;
      RECT  24245.0 187430.0 24950.0 188775.0 ;
      RECT  24245.0 190120.0 24950.0 188775.0 ;
      RECT  24245.0 190120.0 24950.0 191465.0 ;
      RECT  24245.0 192810.0 24950.0 191465.0 ;
      RECT  24245.0 192810.0 24950.0 194155.0 ;
      RECT  24245.0 195500.0 24950.0 194155.0 ;
      RECT  24245.0 195500.0 24950.0 196845.0 ;
      RECT  24245.0 198190.0 24950.0 196845.0 ;
      RECT  24245.0 198190.0 24950.0 199535.0 ;
      RECT  24245.0 200880.0 24950.0 199535.0 ;
      RECT  24245.0 200880.0 24950.0 202225.0 ;
      RECT  24245.0 203570.0 24950.0 202225.0 ;
      RECT  24245.0 203570.0 24950.0 204915.0 ;
      RECT  24245.0 206260.0 24950.0 204915.0 ;
      RECT  24950.0 34100.0 25655.0 35445.0 ;
      RECT  24950.0 36790.0 25655.0 35445.0 ;
      RECT  24950.0 36790.0 25655.0 38135.0 ;
      RECT  24950.0 39480.0 25655.0 38135.0 ;
      RECT  24950.0 39480.0 25655.0 40825.0 ;
      RECT  24950.0 42170.0 25655.0 40825.0 ;
      RECT  24950.0 42170.0 25655.0 43515.0 ;
      RECT  24950.0 44860.0 25655.0 43515.0 ;
      RECT  24950.0 44860.0 25655.0 46205.0 ;
      RECT  24950.0 47550.0 25655.0 46205.0 ;
      RECT  24950.0 47550.0 25655.0 48895.0 ;
      RECT  24950.0 50240.0 25655.0 48895.0 ;
      RECT  24950.0 50240.0 25655.0 51585.0 ;
      RECT  24950.0 52930.0 25655.0 51585.0 ;
      RECT  24950.0 52930.0 25655.0 54275.0 ;
      RECT  24950.0 55620.0 25655.0 54275.0 ;
      RECT  24950.0 55620.0 25655.0 56965.0 ;
      RECT  24950.0 58310.0 25655.0 56965.0 ;
      RECT  24950.0 58310.0 25655.0 59655.0 ;
      RECT  24950.0 61000.0 25655.0 59655.0 ;
      RECT  24950.0 61000.0 25655.0 62345.0 ;
      RECT  24950.0 63690.0 25655.0 62345.0 ;
      RECT  24950.0 63690.0 25655.0 65035.0 ;
      RECT  24950.0 66380.0 25655.0 65035.0 ;
      RECT  24950.0 66380.0 25655.0 67725.0 ;
      RECT  24950.0 69070.0 25655.0 67725.0 ;
      RECT  24950.0 69070.0 25655.0 70415.0 ;
      RECT  24950.0 71760.0 25655.0 70415.0 ;
      RECT  24950.0 71760.0 25655.0 73105.0 ;
      RECT  24950.0 74450.0 25655.0 73105.0 ;
      RECT  24950.0 74450.0 25655.0 75795.0 ;
      RECT  24950.0 77140.0 25655.0 75795.0 ;
      RECT  24950.0 77140.0 25655.0 78485.0 ;
      RECT  24950.0 79830.0 25655.0 78485.0 ;
      RECT  24950.0 79830.0 25655.0 81175.0 ;
      RECT  24950.0 82520.0 25655.0 81175.0 ;
      RECT  24950.0 82520.0 25655.0 83865.0 ;
      RECT  24950.0 85210.0 25655.0 83865.0 ;
      RECT  24950.0 85210.0 25655.0 86555.0 ;
      RECT  24950.0 87900.0 25655.0 86555.0 ;
      RECT  24950.0 87900.0 25655.0 89245.0 ;
      RECT  24950.0 90590.0 25655.0 89245.0 ;
      RECT  24950.0 90590.0 25655.0 91935.0 ;
      RECT  24950.0 93280.0 25655.0 91935.0 ;
      RECT  24950.0 93280.0 25655.0 94625.0 ;
      RECT  24950.0 95970.0 25655.0 94625.0 ;
      RECT  24950.0 95970.0 25655.0 97315.0 ;
      RECT  24950.0 98660.0 25655.0 97315.0 ;
      RECT  24950.0 98660.0 25655.0 100005.0 ;
      RECT  24950.0 101350.0 25655.0 100005.0 ;
      RECT  24950.0 101350.0 25655.0 102695.0 ;
      RECT  24950.0 104040.0 25655.0 102695.0 ;
      RECT  24950.0 104040.0 25655.0 105385.0 ;
      RECT  24950.0 106730.0 25655.0 105385.0 ;
      RECT  24950.0 106730.0 25655.0 108075.0 ;
      RECT  24950.0 109420.0 25655.0 108075.0 ;
      RECT  24950.0 109420.0 25655.0 110765.0 ;
      RECT  24950.0 112110.0 25655.0 110765.0 ;
      RECT  24950.0 112110.0 25655.0 113455.0 ;
      RECT  24950.0 114800.0 25655.0 113455.0 ;
      RECT  24950.0 114800.0 25655.0 116145.0 ;
      RECT  24950.0 117490.0 25655.0 116145.0 ;
      RECT  24950.0 117490.0 25655.0 118835.0 ;
      RECT  24950.0 120180.0 25655.0 118835.0 ;
      RECT  24950.0 120180.0 25655.0 121525.0 ;
      RECT  24950.0 122870.0 25655.0 121525.0 ;
      RECT  24950.0 122870.0 25655.0 124215.0 ;
      RECT  24950.0 125560.0 25655.0 124215.0 ;
      RECT  24950.0 125560.0 25655.0 126905.0 ;
      RECT  24950.0 128250.0 25655.0 126905.0 ;
      RECT  24950.0 128250.0 25655.0 129595.0 ;
      RECT  24950.0 130940.0 25655.0 129595.0 ;
      RECT  24950.0 130940.0 25655.0 132285.0 ;
      RECT  24950.0 133630.0 25655.0 132285.0 ;
      RECT  24950.0 133630.0 25655.0 134975.0 ;
      RECT  24950.0 136320.0 25655.0 134975.0 ;
      RECT  24950.0 136320.0 25655.0 137665.0 ;
      RECT  24950.0 139010.0 25655.0 137665.0 ;
      RECT  24950.0 139010.0 25655.0 140355.0 ;
      RECT  24950.0 141700.0 25655.0 140355.0 ;
      RECT  24950.0 141700.0 25655.0 143045.0 ;
      RECT  24950.0 144390.0 25655.0 143045.0 ;
      RECT  24950.0 144390.0 25655.0 145735.0 ;
      RECT  24950.0 147080.0 25655.0 145735.0 ;
      RECT  24950.0 147080.0 25655.0 148425.0 ;
      RECT  24950.0 149770.0 25655.0 148425.0 ;
      RECT  24950.0 149770.0 25655.0 151115.0 ;
      RECT  24950.0 152460.0 25655.0 151115.0 ;
      RECT  24950.0 152460.0 25655.0 153805.0 ;
      RECT  24950.0 155150.0 25655.0 153805.0 ;
      RECT  24950.0 155150.0 25655.0 156495.0 ;
      RECT  24950.0 157840.0 25655.0 156495.0 ;
      RECT  24950.0 157840.0 25655.0 159185.0 ;
      RECT  24950.0 160530.0 25655.0 159185.0 ;
      RECT  24950.0 160530.0 25655.0 161875.0 ;
      RECT  24950.0 163220.0 25655.0 161875.0 ;
      RECT  24950.0 163220.0 25655.0 164565.0 ;
      RECT  24950.0 165910.0 25655.0 164565.0 ;
      RECT  24950.0 165910.0 25655.0 167255.0 ;
      RECT  24950.0 168600.0 25655.0 167255.0 ;
      RECT  24950.0 168600.0 25655.0 169945.0 ;
      RECT  24950.0 171290.0 25655.0 169945.0 ;
      RECT  24950.0 171290.0 25655.0 172635.0 ;
      RECT  24950.0 173980.0 25655.0 172635.0 ;
      RECT  24950.0 173980.0 25655.0 175325.0 ;
      RECT  24950.0 176670.0 25655.0 175325.0 ;
      RECT  24950.0 176670.0 25655.0 178015.0 ;
      RECT  24950.0 179360.0 25655.0 178015.0 ;
      RECT  24950.0 179360.0 25655.0 180705.0 ;
      RECT  24950.0 182050.0 25655.0 180705.0 ;
      RECT  24950.0 182050.0 25655.0 183395.0 ;
      RECT  24950.0 184740.0 25655.0 183395.0 ;
      RECT  24950.0 184740.0 25655.0 186085.0 ;
      RECT  24950.0 187430.0 25655.0 186085.0 ;
      RECT  24950.0 187430.0 25655.0 188775.0 ;
      RECT  24950.0 190120.0 25655.0 188775.0 ;
      RECT  24950.0 190120.0 25655.0 191465.0 ;
      RECT  24950.0 192810.0 25655.0 191465.0 ;
      RECT  24950.0 192810.0 25655.0 194155.0 ;
      RECT  24950.0 195500.0 25655.0 194155.0 ;
      RECT  24950.0 195500.0 25655.0 196845.0 ;
      RECT  24950.0 198190.0 25655.0 196845.0 ;
      RECT  24950.0 198190.0 25655.0 199535.0 ;
      RECT  24950.0 200880.0 25655.0 199535.0 ;
      RECT  24950.0 200880.0 25655.0 202225.0 ;
      RECT  24950.0 203570.0 25655.0 202225.0 ;
      RECT  24950.0 203570.0 25655.0 204915.0 ;
      RECT  24950.0 206260.0 25655.0 204915.0 ;
      RECT  25655.0 34100.0 26360.0 35445.0 ;
      RECT  25655.0 36790.0 26360.0 35445.0 ;
      RECT  25655.0 36790.0 26360.0 38135.0 ;
      RECT  25655.0 39480.0 26360.0 38135.0 ;
      RECT  25655.0 39480.0 26360.0 40825.0 ;
      RECT  25655.0 42170.0 26360.0 40825.0 ;
      RECT  25655.0 42170.0 26360.0 43515.0 ;
      RECT  25655.0 44860.0 26360.0 43515.0 ;
      RECT  25655.0 44860.0 26360.0 46205.0 ;
      RECT  25655.0 47550.0 26360.0 46205.0 ;
      RECT  25655.0 47550.0 26360.0 48895.0 ;
      RECT  25655.0 50240.0 26360.0 48895.0 ;
      RECT  25655.0 50240.0 26360.0 51585.0 ;
      RECT  25655.0 52930.0 26360.0 51585.0 ;
      RECT  25655.0 52930.0 26360.0 54275.0 ;
      RECT  25655.0 55620.0 26360.0 54275.0 ;
      RECT  25655.0 55620.0 26360.0 56965.0 ;
      RECT  25655.0 58310.0 26360.0 56965.0 ;
      RECT  25655.0 58310.0 26360.0 59655.0 ;
      RECT  25655.0 61000.0 26360.0 59655.0 ;
      RECT  25655.0 61000.0 26360.0 62345.0 ;
      RECT  25655.0 63690.0 26360.0 62345.0 ;
      RECT  25655.0 63690.0 26360.0 65035.0 ;
      RECT  25655.0 66380.0 26360.0 65035.0 ;
      RECT  25655.0 66380.0 26360.0 67725.0 ;
      RECT  25655.0 69070.0 26360.0 67725.0 ;
      RECT  25655.0 69070.0 26360.0 70415.0 ;
      RECT  25655.0 71760.0 26360.0 70415.0 ;
      RECT  25655.0 71760.0 26360.0 73105.0 ;
      RECT  25655.0 74450.0 26360.0 73105.0 ;
      RECT  25655.0 74450.0 26360.0 75795.0 ;
      RECT  25655.0 77140.0 26360.0 75795.0 ;
      RECT  25655.0 77140.0 26360.0 78485.0 ;
      RECT  25655.0 79830.0 26360.0 78485.0 ;
      RECT  25655.0 79830.0 26360.0 81175.0 ;
      RECT  25655.0 82520.0 26360.0 81175.0 ;
      RECT  25655.0 82520.0 26360.0 83865.0 ;
      RECT  25655.0 85210.0 26360.0 83865.0 ;
      RECT  25655.0 85210.0 26360.0 86555.0 ;
      RECT  25655.0 87900.0 26360.0 86555.0 ;
      RECT  25655.0 87900.0 26360.0 89245.0 ;
      RECT  25655.0 90590.0 26360.0 89245.0 ;
      RECT  25655.0 90590.0 26360.0 91935.0 ;
      RECT  25655.0 93280.0 26360.0 91935.0 ;
      RECT  25655.0 93280.0 26360.0 94625.0 ;
      RECT  25655.0 95970.0 26360.0 94625.0 ;
      RECT  25655.0 95970.0 26360.0 97315.0 ;
      RECT  25655.0 98660.0 26360.0 97315.0 ;
      RECT  25655.0 98660.0 26360.0 100005.0 ;
      RECT  25655.0 101350.0 26360.0 100005.0 ;
      RECT  25655.0 101350.0 26360.0 102695.0 ;
      RECT  25655.0 104040.0 26360.0 102695.0 ;
      RECT  25655.0 104040.0 26360.0 105385.0 ;
      RECT  25655.0 106730.0 26360.0 105385.0 ;
      RECT  25655.0 106730.0 26360.0 108075.0 ;
      RECT  25655.0 109420.0 26360.0 108075.0 ;
      RECT  25655.0 109420.0 26360.0 110765.0 ;
      RECT  25655.0 112110.0 26360.0 110765.0 ;
      RECT  25655.0 112110.0 26360.0 113455.0 ;
      RECT  25655.0 114800.0 26360.0 113455.0 ;
      RECT  25655.0 114800.0 26360.0 116145.0 ;
      RECT  25655.0 117490.0 26360.0 116145.0 ;
      RECT  25655.0 117490.0 26360.0 118835.0 ;
      RECT  25655.0 120180.0 26360.0 118835.0 ;
      RECT  25655.0 120180.0 26360.0 121525.0 ;
      RECT  25655.0 122870.0 26360.0 121525.0 ;
      RECT  25655.0 122870.0 26360.0 124215.0 ;
      RECT  25655.0 125560.0 26360.0 124215.0 ;
      RECT  25655.0 125560.0 26360.0 126905.0 ;
      RECT  25655.0 128250.0 26360.0 126905.0 ;
      RECT  25655.0 128250.0 26360.0 129595.0 ;
      RECT  25655.0 130940.0 26360.0 129595.0 ;
      RECT  25655.0 130940.0 26360.0 132285.0 ;
      RECT  25655.0 133630.0 26360.0 132285.0 ;
      RECT  25655.0 133630.0 26360.0 134975.0 ;
      RECT  25655.0 136320.0 26360.0 134975.0 ;
      RECT  25655.0 136320.0 26360.0 137665.0 ;
      RECT  25655.0 139010.0 26360.0 137665.0 ;
      RECT  25655.0 139010.0 26360.0 140355.0 ;
      RECT  25655.0 141700.0 26360.0 140355.0 ;
      RECT  25655.0 141700.0 26360.0 143045.0 ;
      RECT  25655.0 144390.0 26360.0 143045.0 ;
      RECT  25655.0 144390.0 26360.0 145735.0 ;
      RECT  25655.0 147080.0 26360.0 145735.0 ;
      RECT  25655.0 147080.0 26360.0 148425.0 ;
      RECT  25655.0 149770.0 26360.0 148425.0 ;
      RECT  25655.0 149770.0 26360.0 151115.0 ;
      RECT  25655.0 152460.0 26360.0 151115.0 ;
      RECT  25655.0 152460.0 26360.0 153805.0 ;
      RECT  25655.0 155150.0 26360.0 153805.0 ;
      RECT  25655.0 155150.0 26360.0 156495.0 ;
      RECT  25655.0 157840.0 26360.0 156495.0 ;
      RECT  25655.0 157840.0 26360.0 159185.0 ;
      RECT  25655.0 160530.0 26360.0 159185.0 ;
      RECT  25655.0 160530.0 26360.0 161875.0 ;
      RECT  25655.0 163220.0 26360.0 161875.0 ;
      RECT  25655.0 163220.0 26360.0 164565.0 ;
      RECT  25655.0 165910.0 26360.0 164565.0 ;
      RECT  25655.0 165910.0 26360.0 167255.0 ;
      RECT  25655.0 168600.0 26360.0 167255.0 ;
      RECT  25655.0 168600.0 26360.0 169945.0 ;
      RECT  25655.0 171290.0 26360.0 169945.0 ;
      RECT  25655.0 171290.0 26360.0 172635.0 ;
      RECT  25655.0 173980.0 26360.0 172635.0 ;
      RECT  25655.0 173980.0 26360.0 175325.0 ;
      RECT  25655.0 176670.0 26360.0 175325.0 ;
      RECT  25655.0 176670.0 26360.0 178015.0 ;
      RECT  25655.0 179360.0 26360.0 178015.0 ;
      RECT  25655.0 179360.0 26360.0 180705.0 ;
      RECT  25655.0 182050.0 26360.0 180705.0 ;
      RECT  25655.0 182050.0 26360.0 183395.0 ;
      RECT  25655.0 184740.0 26360.0 183395.0 ;
      RECT  25655.0 184740.0 26360.0 186085.0 ;
      RECT  25655.0 187430.0 26360.0 186085.0 ;
      RECT  25655.0 187430.0 26360.0 188775.0 ;
      RECT  25655.0 190120.0 26360.0 188775.0 ;
      RECT  25655.0 190120.0 26360.0 191465.0 ;
      RECT  25655.0 192810.0 26360.0 191465.0 ;
      RECT  25655.0 192810.0 26360.0 194155.0 ;
      RECT  25655.0 195500.0 26360.0 194155.0 ;
      RECT  25655.0 195500.0 26360.0 196845.0 ;
      RECT  25655.0 198190.0 26360.0 196845.0 ;
      RECT  25655.0 198190.0 26360.0 199535.0 ;
      RECT  25655.0 200880.0 26360.0 199535.0 ;
      RECT  25655.0 200880.0 26360.0 202225.0 ;
      RECT  25655.0 203570.0 26360.0 202225.0 ;
      RECT  25655.0 203570.0 26360.0 204915.0 ;
      RECT  25655.0 206260.0 26360.0 204915.0 ;
      RECT  26360.0 34100.0 27065.0 35445.0 ;
      RECT  26360.0 36790.0 27065.0 35445.0 ;
      RECT  26360.0 36790.0 27065.0 38135.0 ;
      RECT  26360.0 39480.0 27065.0 38135.0 ;
      RECT  26360.0 39480.0 27065.0 40825.0 ;
      RECT  26360.0 42170.0 27065.0 40825.0 ;
      RECT  26360.0 42170.0 27065.0 43515.0 ;
      RECT  26360.0 44860.0 27065.0 43515.0 ;
      RECT  26360.0 44860.0 27065.0 46205.0 ;
      RECT  26360.0 47550.0 27065.0 46205.0 ;
      RECT  26360.0 47550.0 27065.0 48895.0 ;
      RECT  26360.0 50240.0 27065.0 48895.0 ;
      RECT  26360.0 50240.0 27065.0 51585.0 ;
      RECT  26360.0 52930.0 27065.0 51585.0 ;
      RECT  26360.0 52930.0 27065.0 54275.0 ;
      RECT  26360.0 55620.0 27065.0 54275.0 ;
      RECT  26360.0 55620.0 27065.0 56965.0 ;
      RECT  26360.0 58310.0 27065.0 56965.0 ;
      RECT  26360.0 58310.0 27065.0 59655.0 ;
      RECT  26360.0 61000.0 27065.0 59655.0 ;
      RECT  26360.0 61000.0 27065.0 62345.0 ;
      RECT  26360.0 63690.0 27065.0 62345.0 ;
      RECT  26360.0 63690.0 27065.0 65035.0 ;
      RECT  26360.0 66380.0 27065.0 65035.0 ;
      RECT  26360.0 66380.0 27065.0 67725.0 ;
      RECT  26360.0 69070.0 27065.0 67725.0 ;
      RECT  26360.0 69070.0 27065.0 70415.0 ;
      RECT  26360.0 71760.0 27065.0 70415.0 ;
      RECT  26360.0 71760.0 27065.0 73105.0 ;
      RECT  26360.0 74450.0 27065.0 73105.0 ;
      RECT  26360.0 74450.0 27065.0 75795.0 ;
      RECT  26360.0 77140.0 27065.0 75795.0 ;
      RECT  26360.0 77140.0 27065.0 78485.0 ;
      RECT  26360.0 79830.0 27065.0 78485.0 ;
      RECT  26360.0 79830.0 27065.0 81175.0 ;
      RECT  26360.0 82520.0 27065.0 81175.0 ;
      RECT  26360.0 82520.0 27065.0 83865.0 ;
      RECT  26360.0 85210.0 27065.0 83865.0 ;
      RECT  26360.0 85210.0 27065.0 86555.0 ;
      RECT  26360.0 87900.0 27065.0 86555.0 ;
      RECT  26360.0 87900.0 27065.0 89245.0 ;
      RECT  26360.0 90590.0 27065.0 89245.0 ;
      RECT  26360.0 90590.0 27065.0 91935.0 ;
      RECT  26360.0 93280.0 27065.0 91935.0 ;
      RECT  26360.0 93280.0 27065.0 94625.0 ;
      RECT  26360.0 95970.0 27065.0 94625.0 ;
      RECT  26360.0 95970.0 27065.0 97315.0 ;
      RECT  26360.0 98660.0 27065.0 97315.0 ;
      RECT  26360.0 98660.0 27065.0 100005.0 ;
      RECT  26360.0 101350.0 27065.0 100005.0 ;
      RECT  26360.0 101350.0 27065.0 102695.0 ;
      RECT  26360.0 104040.0 27065.0 102695.0 ;
      RECT  26360.0 104040.0 27065.0 105385.0 ;
      RECT  26360.0 106730.0 27065.0 105385.0 ;
      RECT  26360.0 106730.0 27065.0 108075.0 ;
      RECT  26360.0 109420.0 27065.0 108075.0 ;
      RECT  26360.0 109420.0 27065.0 110765.0 ;
      RECT  26360.0 112110.0 27065.0 110765.0 ;
      RECT  26360.0 112110.0 27065.0 113455.0 ;
      RECT  26360.0 114800.0 27065.0 113455.0 ;
      RECT  26360.0 114800.0 27065.0 116145.0 ;
      RECT  26360.0 117490.0 27065.0 116145.0 ;
      RECT  26360.0 117490.0 27065.0 118835.0 ;
      RECT  26360.0 120180.0 27065.0 118835.0 ;
      RECT  26360.0 120180.0 27065.0 121525.0 ;
      RECT  26360.0 122870.0 27065.0 121525.0 ;
      RECT  26360.0 122870.0 27065.0 124215.0 ;
      RECT  26360.0 125560.0 27065.0 124215.0 ;
      RECT  26360.0 125560.0 27065.0 126905.0 ;
      RECT  26360.0 128250.0 27065.0 126905.0 ;
      RECT  26360.0 128250.0 27065.0 129595.0 ;
      RECT  26360.0 130940.0 27065.0 129595.0 ;
      RECT  26360.0 130940.0 27065.0 132285.0 ;
      RECT  26360.0 133630.0 27065.0 132285.0 ;
      RECT  26360.0 133630.0 27065.0 134975.0 ;
      RECT  26360.0 136320.0 27065.0 134975.0 ;
      RECT  26360.0 136320.0 27065.0 137665.0 ;
      RECT  26360.0 139010.0 27065.0 137665.0 ;
      RECT  26360.0 139010.0 27065.0 140355.0 ;
      RECT  26360.0 141700.0 27065.0 140355.0 ;
      RECT  26360.0 141700.0 27065.0 143045.0 ;
      RECT  26360.0 144390.0 27065.0 143045.0 ;
      RECT  26360.0 144390.0 27065.0 145735.0 ;
      RECT  26360.0 147080.0 27065.0 145735.0 ;
      RECT  26360.0 147080.0 27065.0 148425.0 ;
      RECT  26360.0 149770.0 27065.0 148425.0 ;
      RECT  26360.0 149770.0 27065.0 151115.0 ;
      RECT  26360.0 152460.0 27065.0 151115.0 ;
      RECT  26360.0 152460.0 27065.0 153805.0 ;
      RECT  26360.0 155150.0 27065.0 153805.0 ;
      RECT  26360.0 155150.0 27065.0 156495.0 ;
      RECT  26360.0 157840.0 27065.0 156495.0 ;
      RECT  26360.0 157840.0 27065.0 159185.0 ;
      RECT  26360.0 160530.0 27065.0 159185.0 ;
      RECT  26360.0 160530.0 27065.0 161875.0 ;
      RECT  26360.0 163220.0 27065.0 161875.0 ;
      RECT  26360.0 163220.0 27065.0 164565.0 ;
      RECT  26360.0 165910.0 27065.0 164565.0 ;
      RECT  26360.0 165910.0 27065.0 167255.0 ;
      RECT  26360.0 168600.0 27065.0 167255.0 ;
      RECT  26360.0 168600.0 27065.0 169945.0 ;
      RECT  26360.0 171290.0 27065.0 169945.0 ;
      RECT  26360.0 171290.0 27065.0 172635.0 ;
      RECT  26360.0 173980.0 27065.0 172635.0 ;
      RECT  26360.0 173980.0 27065.0 175325.0 ;
      RECT  26360.0 176670.0 27065.0 175325.0 ;
      RECT  26360.0 176670.0 27065.0 178015.0 ;
      RECT  26360.0 179360.0 27065.0 178015.0 ;
      RECT  26360.0 179360.0 27065.0 180705.0 ;
      RECT  26360.0 182050.0 27065.0 180705.0 ;
      RECT  26360.0 182050.0 27065.0 183395.0 ;
      RECT  26360.0 184740.0 27065.0 183395.0 ;
      RECT  26360.0 184740.0 27065.0 186085.0 ;
      RECT  26360.0 187430.0 27065.0 186085.0 ;
      RECT  26360.0 187430.0 27065.0 188775.0 ;
      RECT  26360.0 190120.0 27065.0 188775.0 ;
      RECT  26360.0 190120.0 27065.0 191465.0 ;
      RECT  26360.0 192810.0 27065.0 191465.0 ;
      RECT  26360.0 192810.0 27065.0 194155.0 ;
      RECT  26360.0 195500.0 27065.0 194155.0 ;
      RECT  26360.0 195500.0 27065.0 196845.0 ;
      RECT  26360.0 198190.0 27065.0 196845.0 ;
      RECT  26360.0 198190.0 27065.0 199535.0 ;
      RECT  26360.0 200880.0 27065.0 199535.0 ;
      RECT  26360.0 200880.0 27065.0 202225.0 ;
      RECT  26360.0 203570.0 27065.0 202225.0 ;
      RECT  26360.0 203570.0 27065.0 204915.0 ;
      RECT  26360.0 206260.0 27065.0 204915.0 ;
      RECT  27065.0 34100.0 27770.0 35445.0 ;
      RECT  27065.0 36790.0 27770.0 35445.0 ;
      RECT  27065.0 36790.0 27770.0 38135.0 ;
      RECT  27065.0 39480.0 27770.0 38135.0 ;
      RECT  27065.0 39480.0 27770.0 40825.0 ;
      RECT  27065.0 42170.0 27770.0 40825.0 ;
      RECT  27065.0 42170.0 27770.0 43515.0 ;
      RECT  27065.0 44860.0 27770.0 43515.0 ;
      RECT  27065.0 44860.0 27770.0 46205.0 ;
      RECT  27065.0 47550.0 27770.0 46205.0 ;
      RECT  27065.0 47550.0 27770.0 48895.0 ;
      RECT  27065.0 50240.0 27770.0 48895.0 ;
      RECT  27065.0 50240.0 27770.0 51585.0 ;
      RECT  27065.0 52930.0 27770.0 51585.0 ;
      RECT  27065.0 52930.0 27770.0 54275.0 ;
      RECT  27065.0 55620.0 27770.0 54275.0 ;
      RECT  27065.0 55620.0 27770.0 56965.0 ;
      RECT  27065.0 58310.0 27770.0 56965.0 ;
      RECT  27065.0 58310.0 27770.0 59655.0 ;
      RECT  27065.0 61000.0 27770.0 59655.0 ;
      RECT  27065.0 61000.0 27770.0 62345.0 ;
      RECT  27065.0 63690.0 27770.0 62345.0 ;
      RECT  27065.0 63690.0 27770.0 65035.0 ;
      RECT  27065.0 66380.0 27770.0 65035.0 ;
      RECT  27065.0 66380.0 27770.0 67725.0 ;
      RECT  27065.0 69070.0 27770.0 67725.0 ;
      RECT  27065.0 69070.0 27770.0 70415.0 ;
      RECT  27065.0 71760.0 27770.0 70415.0 ;
      RECT  27065.0 71760.0 27770.0 73105.0 ;
      RECT  27065.0 74450.0 27770.0 73105.0 ;
      RECT  27065.0 74450.0 27770.0 75795.0 ;
      RECT  27065.0 77140.0 27770.0 75795.0 ;
      RECT  27065.0 77140.0 27770.0 78485.0 ;
      RECT  27065.0 79830.0 27770.0 78485.0 ;
      RECT  27065.0 79830.0 27770.0 81175.0 ;
      RECT  27065.0 82520.0 27770.0 81175.0 ;
      RECT  27065.0 82520.0 27770.0 83865.0 ;
      RECT  27065.0 85210.0 27770.0 83865.0 ;
      RECT  27065.0 85210.0 27770.0 86555.0 ;
      RECT  27065.0 87900.0 27770.0 86555.0 ;
      RECT  27065.0 87900.0 27770.0 89245.0 ;
      RECT  27065.0 90590.0 27770.0 89245.0 ;
      RECT  27065.0 90590.0 27770.0 91935.0 ;
      RECT  27065.0 93280.0 27770.0 91935.0 ;
      RECT  27065.0 93280.0 27770.0 94625.0 ;
      RECT  27065.0 95970.0 27770.0 94625.0 ;
      RECT  27065.0 95970.0 27770.0 97315.0 ;
      RECT  27065.0 98660.0 27770.0 97315.0 ;
      RECT  27065.0 98660.0 27770.0 100005.0 ;
      RECT  27065.0 101350.0 27770.0 100005.0 ;
      RECT  27065.0 101350.0 27770.0 102695.0 ;
      RECT  27065.0 104040.0 27770.0 102695.0 ;
      RECT  27065.0 104040.0 27770.0 105385.0 ;
      RECT  27065.0 106730.0 27770.0 105385.0 ;
      RECT  27065.0 106730.0 27770.0 108075.0 ;
      RECT  27065.0 109420.0 27770.0 108075.0 ;
      RECT  27065.0 109420.0 27770.0 110765.0 ;
      RECT  27065.0 112110.0 27770.0 110765.0 ;
      RECT  27065.0 112110.0 27770.0 113455.0 ;
      RECT  27065.0 114800.0 27770.0 113455.0 ;
      RECT  27065.0 114800.0 27770.0 116145.0 ;
      RECT  27065.0 117490.0 27770.0 116145.0 ;
      RECT  27065.0 117490.0 27770.0 118835.0 ;
      RECT  27065.0 120180.0 27770.0 118835.0 ;
      RECT  27065.0 120180.0 27770.0 121525.0 ;
      RECT  27065.0 122870.0 27770.0 121525.0 ;
      RECT  27065.0 122870.0 27770.0 124215.0 ;
      RECT  27065.0 125560.0 27770.0 124215.0 ;
      RECT  27065.0 125560.0 27770.0 126905.0 ;
      RECT  27065.0 128250.0 27770.0 126905.0 ;
      RECT  27065.0 128250.0 27770.0 129595.0 ;
      RECT  27065.0 130940.0 27770.0 129595.0 ;
      RECT  27065.0 130940.0 27770.0 132285.0 ;
      RECT  27065.0 133630.0 27770.0 132285.0 ;
      RECT  27065.0 133630.0 27770.0 134975.0 ;
      RECT  27065.0 136320.0 27770.0 134975.0 ;
      RECT  27065.0 136320.0 27770.0 137665.0 ;
      RECT  27065.0 139010.0 27770.0 137665.0 ;
      RECT  27065.0 139010.0 27770.0 140355.0 ;
      RECT  27065.0 141700.0 27770.0 140355.0 ;
      RECT  27065.0 141700.0 27770.0 143045.0 ;
      RECT  27065.0 144390.0 27770.0 143045.0 ;
      RECT  27065.0 144390.0 27770.0 145735.0 ;
      RECT  27065.0 147080.0 27770.0 145735.0 ;
      RECT  27065.0 147080.0 27770.0 148425.0 ;
      RECT  27065.0 149770.0 27770.0 148425.0 ;
      RECT  27065.0 149770.0 27770.0 151115.0 ;
      RECT  27065.0 152460.0 27770.0 151115.0 ;
      RECT  27065.0 152460.0 27770.0 153805.0 ;
      RECT  27065.0 155150.0 27770.0 153805.0 ;
      RECT  27065.0 155150.0 27770.0 156495.0 ;
      RECT  27065.0 157840.0 27770.0 156495.0 ;
      RECT  27065.0 157840.0 27770.0 159185.0 ;
      RECT  27065.0 160530.0 27770.0 159185.0 ;
      RECT  27065.0 160530.0 27770.0 161875.0 ;
      RECT  27065.0 163220.0 27770.0 161875.0 ;
      RECT  27065.0 163220.0 27770.0 164565.0 ;
      RECT  27065.0 165910.0 27770.0 164565.0 ;
      RECT  27065.0 165910.0 27770.0 167255.0 ;
      RECT  27065.0 168600.0 27770.0 167255.0 ;
      RECT  27065.0 168600.0 27770.0 169945.0 ;
      RECT  27065.0 171290.0 27770.0 169945.0 ;
      RECT  27065.0 171290.0 27770.0 172635.0 ;
      RECT  27065.0 173980.0 27770.0 172635.0 ;
      RECT  27065.0 173980.0 27770.0 175325.0 ;
      RECT  27065.0 176670.0 27770.0 175325.0 ;
      RECT  27065.0 176670.0 27770.0 178015.0 ;
      RECT  27065.0 179360.0 27770.0 178015.0 ;
      RECT  27065.0 179360.0 27770.0 180705.0 ;
      RECT  27065.0 182050.0 27770.0 180705.0 ;
      RECT  27065.0 182050.0 27770.0 183395.0 ;
      RECT  27065.0 184740.0 27770.0 183395.0 ;
      RECT  27065.0 184740.0 27770.0 186085.0 ;
      RECT  27065.0 187430.0 27770.0 186085.0 ;
      RECT  27065.0 187430.0 27770.0 188775.0 ;
      RECT  27065.0 190120.0 27770.0 188775.0 ;
      RECT  27065.0 190120.0 27770.0 191465.0 ;
      RECT  27065.0 192810.0 27770.0 191465.0 ;
      RECT  27065.0 192810.0 27770.0 194155.0 ;
      RECT  27065.0 195500.0 27770.0 194155.0 ;
      RECT  27065.0 195500.0 27770.0 196845.0 ;
      RECT  27065.0 198190.0 27770.0 196845.0 ;
      RECT  27065.0 198190.0 27770.0 199535.0 ;
      RECT  27065.0 200880.0 27770.0 199535.0 ;
      RECT  27065.0 200880.0 27770.0 202225.0 ;
      RECT  27065.0 203570.0 27770.0 202225.0 ;
      RECT  27065.0 203570.0 27770.0 204915.0 ;
      RECT  27065.0 206260.0 27770.0 204915.0 ;
      RECT  27770.0 34100.0 28475.0 35445.0 ;
      RECT  27770.0 36790.0 28475.0 35445.0 ;
      RECT  27770.0 36790.0 28475.0 38135.0 ;
      RECT  27770.0 39480.0 28475.0 38135.0 ;
      RECT  27770.0 39480.0 28475.0 40825.0 ;
      RECT  27770.0 42170.0 28475.0 40825.0 ;
      RECT  27770.0 42170.0 28475.0 43515.0 ;
      RECT  27770.0 44860.0 28475.0 43515.0 ;
      RECT  27770.0 44860.0 28475.0 46205.0 ;
      RECT  27770.0 47550.0 28475.0 46205.0 ;
      RECT  27770.0 47550.0 28475.0 48895.0 ;
      RECT  27770.0 50240.0 28475.0 48895.0 ;
      RECT  27770.0 50240.0 28475.0 51585.0 ;
      RECT  27770.0 52930.0 28475.0 51585.0 ;
      RECT  27770.0 52930.0 28475.0 54275.0 ;
      RECT  27770.0 55620.0 28475.0 54275.0 ;
      RECT  27770.0 55620.0 28475.0 56965.0 ;
      RECT  27770.0 58310.0 28475.0 56965.0 ;
      RECT  27770.0 58310.0 28475.0 59655.0 ;
      RECT  27770.0 61000.0 28475.0 59655.0 ;
      RECT  27770.0 61000.0 28475.0 62345.0 ;
      RECT  27770.0 63690.0 28475.0 62345.0 ;
      RECT  27770.0 63690.0 28475.0 65035.0 ;
      RECT  27770.0 66380.0 28475.0 65035.0 ;
      RECT  27770.0 66380.0 28475.0 67725.0 ;
      RECT  27770.0 69070.0 28475.0 67725.0 ;
      RECT  27770.0 69070.0 28475.0 70415.0 ;
      RECT  27770.0 71760.0 28475.0 70415.0 ;
      RECT  27770.0 71760.0 28475.0 73105.0 ;
      RECT  27770.0 74450.0 28475.0 73105.0 ;
      RECT  27770.0 74450.0 28475.0 75795.0 ;
      RECT  27770.0 77140.0 28475.0 75795.0 ;
      RECT  27770.0 77140.0 28475.0 78485.0 ;
      RECT  27770.0 79830.0 28475.0 78485.0 ;
      RECT  27770.0 79830.0 28475.0 81175.0 ;
      RECT  27770.0 82520.0 28475.0 81175.0 ;
      RECT  27770.0 82520.0 28475.0 83865.0 ;
      RECT  27770.0 85210.0 28475.0 83865.0 ;
      RECT  27770.0 85210.0 28475.0 86555.0 ;
      RECT  27770.0 87900.0 28475.0 86555.0 ;
      RECT  27770.0 87900.0 28475.0 89245.0 ;
      RECT  27770.0 90590.0 28475.0 89245.0 ;
      RECT  27770.0 90590.0 28475.0 91935.0 ;
      RECT  27770.0 93280.0 28475.0 91935.0 ;
      RECT  27770.0 93280.0 28475.0 94625.0 ;
      RECT  27770.0 95970.0 28475.0 94625.0 ;
      RECT  27770.0 95970.0 28475.0 97315.0 ;
      RECT  27770.0 98660.0 28475.0 97315.0 ;
      RECT  27770.0 98660.0 28475.0 100005.0 ;
      RECT  27770.0 101350.0 28475.0 100005.0 ;
      RECT  27770.0 101350.0 28475.0 102695.0 ;
      RECT  27770.0 104040.0 28475.0 102695.0 ;
      RECT  27770.0 104040.0 28475.0 105385.0 ;
      RECT  27770.0 106730.0 28475.0 105385.0 ;
      RECT  27770.0 106730.0 28475.0 108075.0 ;
      RECT  27770.0 109420.0 28475.0 108075.0 ;
      RECT  27770.0 109420.0 28475.0 110765.0 ;
      RECT  27770.0 112110.0 28475.0 110765.0 ;
      RECT  27770.0 112110.0 28475.0 113455.0 ;
      RECT  27770.0 114800.0 28475.0 113455.0 ;
      RECT  27770.0 114800.0 28475.0 116145.0 ;
      RECT  27770.0 117490.0 28475.0 116145.0 ;
      RECT  27770.0 117490.0 28475.0 118835.0 ;
      RECT  27770.0 120180.0 28475.0 118835.0 ;
      RECT  27770.0 120180.0 28475.0 121525.0 ;
      RECT  27770.0 122870.0 28475.0 121525.0 ;
      RECT  27770.0 122870.0 28475.0 124215.0 ;
      RECT  27770.0 125560.0 28475.0 124215.0 ;
      RECT  27770.0 125560.0 28475.0 126905.0 ;
      RECT  27770.0 128250.0 28475.0 126905.0 ;
      RECT  27770.0 128250.0 28475.0 129595.0 ;
      RECT  27770.0 130940.0 28475.0 129595.0 ;
      RECT  27770.0 130940.0 28475.0 132285.0 ;
      RECT  27770.0 133630.0 28475.0 132285.0 ;
      RECT  27770.0 133630.0 28475.0 134975.0 ;
      RECT  27770.0 136320.0 28475.0 134975.0 ;
      RECT  27770.0 136320.0 28475.0 137665.0 ;
      RECT  27770.0 139010.0 28475.0 137665.0 ;
      RECT  27770.0 139010.0 28475.0 140355.0 ;
      RECT  27770.0 141700.0 28475.0 140355.0 ;
      RECT  27770.0 141700.0 28475.0 143045.0 ;
      RECT  27770.0 144390.0 28475.0 143045.0 ;
      RECT  27770.0 144390.0 28475.0 145735.0 ;
      RECT  27770.0 147080.0 28475.0 145735.0 ;
      RECT  27770.0 147080.0 28475.0 148425.0 ;
      RECT  27770.0 149770.0 28475.0 148425.0 ;
      RECT  27770.0 149770.0 28475.0 151115.0 ;
      RECT  27770.0 152460.0 28475.0 151115.0 ;
      RECT  27770.0 152460.0 28475.0 153805.0 ;
      RECT  27770.0 155150.0 28475.0 153805.0 ;
      RECT  27770.0 155150.0 28475.0 156495.0 ;
      RECT  27770.0 157840.0 28475.0 156495.0 ;
      RECT  27770.0 157840.0 28475.0 159185.0 ;
      RECT  27770.0 160530.0 28475.0 159185.0 ;
      RECT  27770.0 160530.0 28475.0 161875.0 ;
      RECT  27770.0 163220.0 28475.0 161875.0 ;
      RECT  27770.0 163220.0 28475.0 164565.0 ;
      RECT  27770.0 165910.0 28475.0 164565.0 ;
      RECT  27770.0 165910.0 28475.0 167255.0 ;
      RECT  27770.0 168600.0 28475.0 167255.0 ;
      RECT  27770.0 168600.0 28475.0 169945.0 ;
      RECT  27770.0 171290.0 28475.0 169945.0 ;
      RECT  27770.0 171290.0 28475.0 172635.0 ;
      RECT  27770.0 173980.0 28475.0 172635.0 ;
      RECT  27770.0 173980.0 28475.0 175325.0 ;
      RECT  27770.0 176670.0 28475.0 175325.0 ;
      RECT  27770.0 176670.0 28475.0 178015.0 ;
      RECT  27770.0 179360.0 28475.0 178015.0 ;
      RECT  27770.0 179360.0 28475.0 180705.0 ;
      RECT  27770.0 182050.0 28475.0 180705.0 ;
      RECT  27770.0 182050.0 28475.0 183395.0 ;
      RECT  27770.0 184740.0 28475.0 183395.0 ;
      RECT  27770.0 184740.0 28475.0 186085.0 ;
      RECT  27770.0 187430.0 28475.0 186085.0 ;
      RECT  27770.0 187430.0 28475.0 188775.0 ;
      RECT  27770.0 190120.0 28475.0 188775.0 ;
      RECT  27770.0 190120.0 28475.0 191465.0 ;
      RECT  27770.0 192810.0 28475.0 191465.0 ;
      RECT  27770.0 192810.0 28475.0 194155.0 ;
      RECT  27770.0 195500.0 28475.0 194155.0 ;
      RECT  27770.0 195500.0 28475.0 196845.0 ;
      RECT  27770.0 198190.0 28475.0 196845.0 ;
      RECT  27770.0 198190.0 28475.0 199535.0 ;
      RECT  27770.0 200880.0 28475.0 199535.0 ;
      RECT  27770.0 200880.0 28475.0 202225.0 ;
      RECT  27770.0 203570.0 28475.0 202225.0 ;
      RECT  27770.0 203570.0 28475.0 204915.0 ;
      RECT  27770.0 206260.0 28475.0 204915.0 ;
      RECT  28475.0 34100.0 29180.0 35445.0 ;
      RECT  28475.0 36790.0 29180.0 35445.0 ;
      RECT  28475.0 36790.0 29180.0 38135.0 ;
      RECT  28475.0 39480.0 29180.0 38135.0 ;
      RECT  28475.0 39480.0 29180.0 40825.0 ;
      RECT  28475.0 42170.0 29180.0 40825.0 ;
      RECT  28475.0 42170.0 29180.0 43515.0 ;
      RECT  28475.0 44860.0 29180.0 43515.0 ;
      RECT  28475.0 44860.0 29180.0 46205.0 ;
      RECT  28475.0 47550.0 29180.0 46205.0 ;
      RECT  28475.0 47550.0 29180.0 48895.0 ;
      RECT  28475.0 50240.0 29180.0 48895.0 ;
      RECT  28475.0 50240.0 29180.0 51585.0 ;
      RECT  28475.0 52930.0 29180.0 51585.0 ;
      RECT  28475.0 52930.0 29180.0 54275.0 ;
      RECT  28475.0 55620.0 29180.0 54275.0 ;
      RECT  28475.0 55620.0 29180.0 56965.0 ;
      RECT  28475.0 58310.0 29180.0 56965.0 ;
      RECT  28475.0 58310.0 29180.0 59655.0 ;
      RECT  28475.0 61000.0 29180.0 59655.0 ;
      RECT  28475.0 61000.0 29180.0 62345.0 ;
      RECT  28475.0 63690.0 29180.0 62345.0 ;
      RECT  28475.0 63690.0 29180.0 65035.0 ;
      RECT  28475.0 66380.0 29180.0 65035.0 ;
      RECT  28475.0 66380.0 29180.0 67725.0 ;
      RECT  28475.0 69070.0 29180.0 67725.0 ;
      RECT  28475.0 69070.0 29180.0 70415.0 ;
      RECT  28475.0 71760.0 29180.0 70415.0 ;
      RECT  28475.0 71760.0 29180.0 73105.0 ;
      RECT  28475.0 74450.0 29180.0 73105.0 ;
      RECT  28475.0 74450.0 29180.0 75795.0 ;
      RECT  28475.0 77140.0 29180.0 75795.0 ;
      RECT  28475.0 77140.0 29180.0 78485.0 ;
      RECT  28475.0 79830.0 29180.0 78485.0 ;
      RECT  28475.0 79830.0 29180.0 81175.0 ;
      RECT  28475.0 82520.0 29180.0 81175.0 ;
      RECT  28475.0 82520.0 29180.0 83865.0 ;
      RECT  28475.0 85210.0 29180.0 83865.0 ;
      RECT  28475.0 85210.0 29180.0 86555.0 ;
      RECT  28475.0 87900.0 29180.0 86555.0 ;
      RECT  28475.0 87900.0 29180.0 89245.0 ;
      RECT  28475.0 90590.0 29180.0 89245.0 ;
      RECT  28475.0 90590.0 29180.0 91935.0 ;
      RECT  28475.0 93280.0 29180.0 91935.0 ;
      RECT  28475.0 93280.0 29180.0 94625.0 ;
      RECT  28475.0 95970.0 29180.0 94625.0 ;
      RECT  28475.0 95970.0 29180.0 97315.0 ;
      RECT  28475.0 98660.0 29180.0 97315.0 ;
      RECT  28475.0 98660.0 29180.0 100005.0 ;
      RECT  28475.0 101350.0 29180.0 100005.0 ;
      RECT  28475.0 101350.0 29180.0 102695.0 ;
      RECT  28475.0 104040.0 29180.0 102695.0 ;
      RECT  28475.0 104040.0 29180.0 105385.0 ;
      RECT  28475.0 106730.0 29180.0 105385.0 ;
      RECT  28475.0 106730.0 29180.0 108075.0 ;
      RECT  28475.0 109420.0 29180.0 108075.0 ;
      RECT  28475.0 109420.0 29180.0 110765.0 ;
      RECT  28475.0 112110.0 29180.0 110765.0 ;
      RECT  28475.0 112110.0 29180.0 113455.0 ;
      RECT  28475.0 114800.0 29180.0 113455.0 ;
      RECT  28475.0 114800.0 29180.0 116145.0 ;
      RECT  28475.0 117490.0 29180.0 116145.0 ;
      RECT  28475.0 117490.0 29180.0 118835.0 ;
      RECT  28475.0 120180.0 29180.0 118835.0 ;
      RECT  28475.0 120180.0 29180.0 121525.0 ;
      RECT  28475.0 122870.0 29180.0 121525.0 ;
      RECT  28475.0 122870.0 29180.0 124215.0 ;
      RECT  28475.0 125560.0 29180.0 124215.0 ;
      RECT  28475.0 125560.0 29180.0 126905.0 ;
      RECT  28475.0 128250.0 29180.0 126905.0 ;
      RECT  28475.0 128250.0 29180.0 129595.0 ;
      RECT  28475.0 130940.0 29180.0 129595.0 ;
      RECT  28475.0 130940.0 29180.0 132285.0 ;
      RECT  28475.0 133630.0 29180.0 132285.0 ;
      RECT  28475.0 133630.0 29180.0 134975.0 ;
      RECT  28475.0 136320.0 29180.0 134975.0 ;
      RECT  28475.0 136320.0 29180.0 137665.0 ;
      RECT  28475.0 139010.0 29180.0 137665.0 ;
      RECT  28475.0 139010.0 29180.0 140355.0 ;
      RECT  28475.0 141700.0 29180.0 140355.0 ;
      RECT  28475.0 141700.0 29180.0 143045.0 ;
      RECT  28475.0 144390.0 29180.0 143045.0 ;
      RECT  28475.0 144390.0 29180.0 145735.0 ;
      RECT  28475.0 147080.0 29180.0 145735.0 ;
      RECT  28475.0 147080.0 29180.0 148425.0 ;
      RECT  28475.0 149770.0 29180.0 148425.0 ;
      RECT  28475.0 149770.0 29180.0 151115.0 ;
      RECT  28475.0 152460.0 29180.0 151115.0 ;
      RECT  28475.0 152460.0 29180.0 153805.0 ;
      RECT  28475.0 155150.0 29180.0 153805.0 ;
      RECT  28475.0 155150.0 29180.0 156495.0 ;
      RECT  28475.0 157840.0 29180.0 156495.0 ;
      RECT  28475.0 157840.0 29180.0 159185.0 ;
      RECT  28475.0 160530.0 29180.0 159185.0 ;
      RECT  28475.0 160530.0 29180.0 161875.0 ;
      RECT  28475.0 163220.0 29180.0 161875.0 ;
      RECT  28475.0 163220.0 29180.0 164565.0 ;
      RECT  28475.0 165910.0 29180.0 164565.0 ;
      RECT  28475.0 165910.0 29180.0 167255.0 ;
      RECT  28475.0 168600.0 29180.0 167255.0 ;
      RECT  28475.0 168600.0 29180.0 169945.0 ;
      RECT  28475.0 171290.0 29180.0 169945.0 ;
      RECT  28475.0 171290.0 29180.0 172635.0 ;
      RECT  28475.0 173980.0 29180.0 172635.0 ;
      RECT  28475.0 173980.0 29180.0 175325.0 ;
      RECT  28475.0 176670.0 29180.0 175325.0 ;
      RECT  28475.0 176670.0 29180.0 178015.0 ;
      RECT  28475.0 179360.0 29180.0 178015.0 ;
      RECT  28475.0 179360.0 29180.0 180705.0 ;
      RECT  28475.0 182050.0 29180.0 180705.0 ;
      RECT  28475.0 182050.0 29180.0 183395.0 ;
      RECT  28475.0 184740.0 29180.0 183395.0 ;
      RECT  28475.0 184740.0 29180.0 186085.0 ;
      RECT  28475.0 187430.0 29180.0 186085.0 ;
      RECT  28475.0 187430.0 29180.0 188775.0 ;
      RECT  28475.0 190120.0 29180.0 188775.0 ;
      RECT  28475.0 190120.0 29180.0 191465.0 ;
      RECT  28475.0 192810.0 29180.0 191465.0 ;
      RECT  28475.0 192810.0 29180.0 194155.0 ;
      RECT  28475.0 195500.0 29180.0 194155.0 ;
      RECT  28475.0 195500.0 29180.0 196845.0 ;
      RECT  28475.0 198190.0 29180.0 196845.0 ;
      RECT  28475.0 198190.0 29180.0 199535.0 ;
      RECT  28475.0 200880.0 29180.0 199535.0 ;
      RECT  28475.0 200880.0 29180.0 202225.0 ;
      RECT  28475.0 203570.0 29180.0 202225.0 ;
      RECT  28475.0 203570.0 29180.0 204915.0 ;
      RECT  28475.0 206260.0 29180.0 204915.0 ;
      RECT  29180.0 34100.0 29885.0 35445.0 ;
      RECT  29180.0 36790.0 29885.0 35445.0 ;
      RECT  29180.0 36790.0 29885.0 38135.0 ;
      RECT  29180.0 39480.0 29885.0 38135.0 ;
      RECT  29180.0 39480.0 29885.0 40825.0 ;
      RECT  29180.0 42170.0 29885.0 40825.0 ;
      RECT  29180.0 42170.0 29885.0 43515.0 ;
      RECT  29180.0 44860.0 29885.0 43515.0 ;
      RECT  29180.0 44860.0 29885.0 46205.0 ;
      RECT  29180.0 47550.0 29885.0 46205.0 ;
      RECT  29180.0 47550.0 29885.0 48895.0 ;
      RECT  29180.0 50240.0 29885.0 48895.0 ;
      RECT  29180.0 50240.0 29885.0 51585.0 ;
      RECT  29180.0 52930.0 29885.0 51585.0 ;
      RECT  29180.0 52930.0 29885.0 54275.0 ;
      RECT  29180.0 55620.0 29885.0 54275.0 ;
      RECT  29180.0 55620.0 29885.0 56965.0 ;
      RECT  29180.0 58310.0 29885.0 56965.0 ;
      RECT  29180.0 58310.0 29885.0 59655.0 ;
      RECT  29180.0 61000.0 29885.0 59655.0 ;
      RECT  29180.0 61000.0 29885.0 62345.0 ;
      RECT  29180.0 63690.0 29885.0 62345.0 ;
      RECT  29180.0 63690.0 29885.0 65035.0 ;
      RECT  29180.0 66380.0 29885.0 65035.0 ;
      RECT  29180.0 66380.0 29885.0 67725.0 ;
      RECT  29180.0 69070.0 29885.0 67725.0 ;
      RECT  29180.0 69070.0 29885.0 70415.0 ;
      RECT  29180.0 71760.0 29885.0 70415.0 ;
      RECT  29180.0 71760.0 29885.0 73105.0 ;
      RECT  29180.0 74450.0 29885.0 73105.0 ;
      RECT  29180.0 74450.0 29885.0 75795.0 ;
      RECT  29180.0 77140.0 29885.0 75795.0 ;
      RECT  29180.0 77140.0 29885.0 78485.0 ;
      RECT  29180.0 79830.0 29885.0 78485.0 ;
      RECT  29180.0 79830.0 29885.0 81175.0 ;
      RECT  29180.0 82520.0 29885.0 81175.0 ;
      RECT  29180.0 82520.0 29885.0 83865.0 ;
      RECT  29180.0 85210.0 29885.0 83865.0 ;
      RECT  29180.0 85210.0 29885.0 86555.0 ;
      RECT  29180.0 87900.0 29885.0 86555.0 ;
      RECT  29180.0 87900.0 29885.0 89245.0 ;
      RECT  29180.0 90590.0 29885.0 89245.0 ;
      RECT  29180.0 90590.0 29885.0 91935.0 ;
      RECT  29180.0 93280.0 29885.0 91935.0 ;
      RECT  29180.0 93280.0 29885.0 94625.0 ;
      RECT  29180.0 95970.0 29885.0 94625.0 ;
      RECT  29180.0 95970.0 29885.0 97315.0 ;
      RECT  29180.0 98660.0 29885.0 97315.0 ;
      RECT  29180.0 98660.0 29885.0 100005.0 ;
      RECT  29180.0 101350.0 29885.0 100005.0 ;
      RECT  29180.0 101350.0 29885.0 102695.0 ;
      RECT  29180.0 104040.0 29885.0 102695.0 ;
      RECT  29180.0 104040.0 29885.0 105385.0 ;
      RECT  29180.0 106730.0 29885.0 105385.0 ;
      RECT  29180.0 106730.0 29885.0 108075.0 ;
      RECT  29180.0 109420.0 29885.0 108075.0 ;
      RECT  29180.0 109420.0 29885.0 110765.0 ;
      RECT  29180.0 112110.0 29885.0 110765.0 ;
      RECT  29180.0 112110.0 29885.0 113455.0 ;
      RECT  29180.0 114800.0 29885.0 113455.0 ;
      RECT  29180.0 114800.0 29885.0 116145.0 ;
      RECT  29180.0 117490.0 29885.0 116145.0 ;
      RECT  29180.0 117490.0 29885.0 118835.0 ;
      RECT  29180.0 120180.0 29885.0 118835.0 ;
      RECT  29180.0 120180.0 29885.0 121525.0 ;
      RECT  29180.0 122870.0 29885.0 121525.0 ;
      RECT  29180.0 122870.0 29885.0 124215.0 ;
      RECT  29180.0 125560.0 29885.0 124215.0 ;
      RECT  29180.0 125560.0 29885.0 126905.0 ;
      RECT  29180.0 128250.0 29885.0 126905.0 ;
      RECT  29180.0 128250.0 29885.0 129595.0 ;
      RECT  29180.0 130940.0 29885.0 129595.0 ;
      RECT  29180.0 130940.0 29885.0 132285.0 ;
      RECT  29180.0 133630.0 29885.0 132285.0 ;
      RECT  29180.0 133630.0 29885.0 134975.0 ;
      RECT  29180.0 136320.0 29885.0 134975.0 ;
      RECT  29180.0 136320.0 29885.0 137665.0 ;
      RECT  29180.0 139010.0 29885.0 137665.0 ;
      RECT  29180.0 139010.0 29885.0 140355.0 ;
      RECT  29180.0 141700.0 29885.0 140355.0 ;
      RECT  29180.0 141700.0 29885.0 143045.0 ;
      RECT  29180.0 144390.0 29885.0 143045.0 ;
      RECT  29180.0 144390.0 29885.0 145735.0 ;
      RECT  29180.0 147080.0 29885.0 145735.0 ;
      RECT  29180.0 147080.0 29885.0 148425.0 ;
      RECT  29180.0 149770.0 29885.0 148425.0 ;
      RECT  29180.0 149770.0 29885.0 151115.0 ;
      RECT  29180.0 152460.0 29885.0 151115.0 ;
      RECT  29180.0 152460.0 29885.0 153805.0 ;
      RECT  29180.0 155150.0 29885.0 153805.0 ;
      RECT  29180.0 155150.0 29885.0 156495.0 ;
      RECT  29180.0 157840.0 29885.0 156495.0 ;
      RECT  29180.0 157840.0 29885.0 159185.0 ;
      RECT  29180.0 160530.0 29885.0 159185.0 ;
      RECT  29180.0 160530.0 29885.0 161875.0 ;
      RECT  29180.0 163220.0 29885.0 161875.0 ;
      RECT  29180.0 163220.0 29885.0 164565.0 ;
      RECT  29180.0 165910.0 29885.0 164565.0 ;
      RECT  29180.0 165910.0 29885.0 167255.0 ;
      RECT  29180.0 168600.0 29885.0 167255.0 ;
      RECT  29180.0 168600.0 29885.0 169945.0 ;
      RECT  29180.0 171290.0 29885.0 169945.0 ;
      RECT  29180.0 171290.0 29885.0 172635.0 ;
      RECT  29180.0 173980.0 29885.0 172635.0 ;
      RECT  29180.0 173980.0 29885.0 175325.0 ;
      RECT  29180.0 176670.0 29885.0 175325.0 ;
      RECT  29180.0 176670.0 29885.0 178015.0 ;
      RECT  29180.0 179360.0 29885.0 178015.0 ;
      RECT  29180.0 179360.0 29885.0 180705.0 ;
      RECT  29180.0 182050.0 29885.0 180705.0 ;
      RECT  29180.0 182050.0 29885.0 183395.0 ;
      RECT  29180.0 184740.0 29885.0 183395.0 ;
      RECT  29180.0 184740.0 29885.0 186085.0 ;
      RECT  29180.0 187430.0 29885.0 186085.0 ;
      RECT  29180.0 187430.0 29885.0 188775.0 ;
      RECT  29180.0 190120.0 29885.0 188775.0 ;
      RECT  29180.0 190120.0 29885.0 191465.0 ;
      RECT  29180.0 192810.0 29885.0 191465.0 ;
      RECT  29180.0 192810.0 29885.0 194155.0 ;
      RECT  29180.0 195500.0 29885.0 194155.0 ;
      RECT  29180.0 195500.0 29885.0 196845.0 ;
      RECT  29180.0 198190.0 29885.0 196845.0 ;
      RECT  29180.0 198190.0 29885.0 199535.0 ;
      RECT  29180.0 200880.0 29885.0 199535.0 ;
      RECT  29180.0 200880.0 29885.0 202225.0 ;
      RECT  29180.0 203570.0 29885.0 202225.0 ;
      RECT  29180.0 203570.0 29885.0 204915.0 ;
      RECT  29180.0 206260.0 29885.0 204915.0 ;
      RECT  29885.0 34100.0 30590.0 35445.0 ;
      RECT  29885.0 36790.0 30590.0 35445.0 ;
      RECT  29885.0 36790.0 30590.0 38135.0 ;
      RECT  29885.0 39480.0 30590.0 38135.0 ;
      RECT  29885.0 39480.0 30590.0 40825.0 ;
      RECT  29885.0 42170.0 30590.0 40825.0 ;
      RECT  29885.0 42170.0 30590.0 43515.0 ;
      RECT  29885.0 44860.0 30590.0 43515.0 ;
      RECT  29885.0 44860.0 30590.0 46205.0 ;
      RECT  29885.0 47550.0 30590.0 46205.0 ;
      RECT  29885.0 47550.0 30590.0 48895.0 ;
      RECT  29885.0 50240.0 30590.0 48895.0 ;
      RECT  29885.0 50240.0 30590.0 51585.0 ;
      RECT  29885.0 52930.0 30590.0 51585.0 ;
      RECT  29885.0 52930.0 30590.0 54275.0 ;
      RECT  29885.0 55620.0 30590.0 54275.0 ;
      RECT  29885.0 55620.0 30590.0 56965.0 ;
      RECT  29885.0 58310.0 30590.0 56965.0 ;
      RECT  29885.0 58310.0 30590.0 59655.0 ;
      RECT  29885.0 61000.0 30590.0 59655.0 ;
      RECT  29885.0 61000.0 30590.0 62345.0 ;
      RECT  29885.0 63690.0 30590.0 62345.0 ;
      RECT  29885.0 63690.0 30590.0 65035.0 ;
      RECT  29885.0 66380.0 30590.0 65035.0 ;
      RECT  29885.0 66380.0 30590.0 67725.0 ;
      RECT  29885.0 69070.0 30590.0 67725.0 ;
      RECT  29885.0 69070.0 30590.0 70415.0 ;
      RECT  29885.0 71760.0 30590.0 70415.0 ;
      RECT  29885.0 71760.0 30590.0 73105.0 ;
      RECT  29885.0 74450.0 30590.0 73105.0 ;
      RECT  29885.0 74450.0 30590.0 75795.0 ;
      RECT  29885.0 77140.0 30590.0 75795.0 ;
      RECT  29885.0 77140.0 30590.0 78485.0 ;
      RECT  29885.0 79830.0 30590.0 78485.0 ;
      RECT  29885.0 79830.0 30590.0 81175.0 ;
      RECT  29885.0 82520.0 30590.0 81175.0 ;
      RECT  29885.0 82520.0 30590.0 83865.0 ;
      RECT  29885.0 85210.0 30590.0 83865.0 ;
      RECT  29885.0 85210.0 30590.0 86555.0 ;
      RECT  29885.0 87900.0 30590.0 86555.0 ;
      RECT  29885.0 87900.0 30590.0 89245.0 ;
      RECT  29885.0 90590.0 30590.0 89245.0 ;
      RECT  29885.0 90590.0 30590.0 91935.0 ;
      RECT  29885.0 93280.0 30590.0 91935.0 ;
      RECT  29885.0 93280.0 30590.0 94625.0 ;
      RECT  29885.0 95970.0 30590.0 94625.0 ;
      RECT  29885.0 95970.0 30590.0 97315.0 ;
      RECT  29885.0 98660.0 30590.0 97315.0 ;
      RECT  29885.0 98660.0 30590.0 100005.0 ;
      RECT  29885.0 101350.0 30590.0 100005.0 ;
      RECT  29885.0 101350.0 30590.0 102695.0 ;
      RECT  29885.0 104040.0 30590.0 102695.0 ;
      RECT  29885.0 104040.0 30590.0 105385.0 ;
      RECT  29885.0 106730.0 30590.0 105385.0 ;
      RECT  29885.0 106730.0 30590.0 108075.0 ;
      RECT  29885.0 109420.0 30590.0 108075.0 ;
      RECT  29885.0 109420.0 30590.0 110765.0 ;
      RECT  29885.0 112110.0 30590.0 110765.0 ;
      RECT  29885.0 112110.0 30590.0 113455.0 ;
      RECT  29885.0 114800.0 30590.0 113455.0 ;
      RECT  29885.0 114800.0 30590.0 116145.0 ;
      RECT  29885.0 117490.0 30590.0 116145.0 ;
      RECT  29885.0 117490.0 30590.0 118835.0 ;
      RECT  29885.0 120180.0 30590.0 118835.0 ;
      RECT  29885.0 120180.0 30590.0 121525.0 ;
      RECT  29885.0 122870.0 30590.0 121525.0 ;
      RECT  29885.0 122870.0 30590.0 124215.0 ;
      RECT  29885.0 125560.0 30590.0 124215.0 ;
      RECT  29885.0 125560.0 30590.0 126905.0 ;
      RECT  29885.0 128250.0 30590.0 126905.0 ;
      RECT  29885.0 128250.0 30590.0 129595.0 ;
      RECT  29885.0 130940.0 30590.0 129595.0 ;
      RECT  29885.0 130940.0 30590.0 132285.0 ;
      RECT  29885.0 133630.0 30590.0 132285.0 ;
      RECT  29885.0 133630.0 30590.0 134975.0 ;
      RECT  29885.0 136320.0 30590.0 134975.0 ;
      RECT  29885.0 136320.0 30590.0 137665.0 ;
      RECT  29885.0 139010.0 30590.0 137665.0 ;
      RECT  29885.0 139010.0 30590.0 140355.0 ;
      RECT  29885.0 141700.0 30590.0 140355.0 ;
      RECT  29885.0 141700.0 30590.0 143045.0 ;
      RECT  29885.0 144390.0 30590.0 143045.0 ;
      RECT  29885.0 144390.0 30590.0 145735.0 ;
      RECT  29885.0 147080.0 30590.0 145735.0 ;
      RECT  29885.0 147080.0 30590.0 148425.0 ;
      RECT  29885.0 149770.0 30590.0 148425.0 ;
      RECT  29885.0 149770.0 30590.0 151115.0 ;
      RECT  29885.0 152460.0 30590.0 151115.0 ;
      RECT  29885.0 152460.0 30590.0 153805.0 ;
      RECT  29885.0 155150.0 30590.0 153805.0 ;
      RECT  29885.0 155150.0 30590.0 156495.0 ;
      RECT  29885.0 157840.0 30590.0 156495.0 ;
      RECT  29885.0 157840.0 30590.0 159185.0 ;
      RECT  29885.0 160530.0 30590.0 159185.0 ;
      RECT  29885.0 160530.0 30590.0 161875.0 ;
      RECT  29885.0 163220.0 30590.0 161875.0 ;
      RECT  29885.0 163220.0 30590.0 164565.0 ;
      RECT  29885.0 165910.0 30590.0 164565.0 ;
      RECT  29885.0 165910.0 30590.0 167255.0 ;
      RECT  29885.0 168600.0 30590.0 167255.0 ;
      RECT  29885.0 168600.0 30590.0 169945.0 ;
      RECT  29885.0 171290.0 30590.0 169945.0 ;
      RECT  29885.0 171290.0 30590.0 172635.0 ;
      RECT  29885.0 173980.0 30590.0 172635.0 ;
      RECT  29885.0 173980.0 30590.0 175325.0 ;
      RECT  29885.0 176670.0 30590.0 175325.0 ;
      RECT  29885.0 176670.0 30590.0 178015.0 ;
      RECT  29885.0 179360.0 30590.0 178015.0 ;
      RECT  29885.0 179360.0 30590.0 180705.0 ;
      RECT  29885.0 182050.0 30590.0 180705.0 ;
      RECT  29885.0 182050.0 30590.0 183395.0 ;
      RECT  29885.0 184740.0 30590.0 183395.0 ;
      RECT  29885.0 184740.0 30590.0 186085.0 ;
      RECT  29885.0 187430.0 30590.0 186085.0 ;
      RECT  29885.0 187430.0 30590.0 188775.0 ;
      RECT  29885.0 190120.0 30590.0 188775.0 ;
      RECT  29885.0 190120.0 30590.0 191465.0 ;
      RECT  29885.0 192810.0 30590.0 191465.0 ;
      RECT  29885.0 192810.0 30590.0 194155.0 ;
      RECT  29885.0 195500.0 30590.0 194155.0 ;
      RECT  29885.0 195500.0 30590.0 196845.0 ;
      RECT  29885.0 198190.0 30590.0 196845.0 ;
      RECT  29885.0 198190.0 30590.0 199535.0 ;
      RECT  29885.0 200880.0 30590.0 199535.0 ;
      RECT  29885.0 200880.0 30590.0 202225.0 ;
      RECT  29885.0 203570.0 30590.0 202225.0 ;
      RECT  29885.0 203570.0 30590.0 204915.0 ;
      RECT  29885.0 206260.0 30590.0 204915.0 ;
      RECT  30590.0 34100.0 31295.0 35445.0 ;
      RECT  30590.0 36790.0 31295.0 35445.0 ;
      RECT  30590.0 36790.0 31295.0 38135.0 ;
      RECT  30590.0 39480.0 31295.0 38135.0 ;
      RECT  30590.0 39480.0 31295.0 40825.0 ;
      RECT  30590.0 42170.0 31295.0 40825.0 ;
      RECT  30590.0 42170.0 31295.0 43515.0 ;
      RECT  30590.0 44860.0 31295.0 43515.0 ;
      RECT  30590.0 44860.0 31295.0 46205.0 ;
      RECT  30590.0 47550.0 31295.0 46205.0 ;
      RECT  30590.0 47550.0 31295.0 48895.0 ;
      RECT  30590.0 50240.0 31295.0 48895.0 ;
      RECT  30590.0 50240.0 31295.0 51585.0 ;
      RECT  30590.0 52930.0 31295.0 51585.0 ;
      RECT  30590.0 52930.0 31295.0 54275.0 ;
      RECT  30590.0 55620.0 31295.0 54275.0 ;
      RECT  30590.0 55620.0 31295.0 56965.0 ;
      RECT  30590.0 58310.0 31295.0 56965.0 ;
      RECT  30590.0 58310.0 31295.0 59655.0 ;
      RECT  30590.0 61000.0 31295.0 59655.0 ;
      RECT  30590.0 61000.0 31295.0 62345.0 ;
      RECT  30590.0 63690.0 31295.0 62345.0 ;
      RECT  30590.0 63690.0 31295.0 65035.0 ;
      RECT  30590.0 66380.0 31295.0 65035.0 ;
      RECT  30590.0 66380.0 31295.0 67725.0 ;
      RECT  30590.0 69070.0 31295.0 67725.0 ;
      RECT  30590.0 69070.0 31295.0 70415.0 ;
      RECT  30590.0 71760.0 31295.0 70415.0 ;
      RECT  30590.0 71760.0 31295.0 73105.0 ;
      RECT  30590.0 74450.0 31295.0 73105.0 ;
      RECT  30590.0 74450.0 31295.0 75795.0 ;
      RECT  30590.0 77140.0 31295.0 75795.0 ;
      RECT  30590.0 77140.0 31295.0 78485.0 ;
      RECT  30590.0 79830.0 31295.0 78485.0 ;
      RECT  30590.0 79830.0 31295.0 81175.0 ;
      RECT  30590.0 82520.0 31295.0 81175.0 ;
      RECT  30590.0 82520.0 31295.0 83865.0 ;
      RECT  30590.0 85210.0 31295.0 83865.0 ;
      RECT  30590.0 85210.0 31295.0 86555.0 ;
      RECT  30590.0 87900.0 31295.0 86555.0 ;
      RECT  30590.0 87900.0 31295.0 89245.0 ;
      RECT  30590.0 90590.0 31295.0 89245.0 ;
      RECT  30590.0 90590.0 31295.0 91935.0 ;
      RECT  30590.0 93280.0 31295.0 91935.0 ;
      RECT  30590.0 93280.0 31295.0 94625.0 ;
      RECT  30590.0 95970.0 31295.0 94625.0 ;
      RECT  30590.0 95970.0 31295.0 97315.0 ;
      RECT  30590.0 98660.0 31295.0 97315.0 ;
      RECT  30590.0 98660.0 31295.0 100005.0 ;
      RECT  30590.0 101350.0 31295.0 100005.0 ;
      RECT  30590.0 101350.0 31295.0 102695.0 ;
      RECT  30590.0 104040.0 31295.0 102695.0 ;
      RECT  30590.0 104040.0 31295.0 105385.0 ;
      RECT  30590.0 106730.0 31295.0 105385.0 ;
      RECT  30590.0 106730.0 31295.0 108075.0 ;
      RECT  30590.0 109420.0 31295.0 108075.0 ;
      RECT  30590.0 109420.0 31295.0 110765.0 ;
      RECT  30590.0 112110.0 31295.0 110765.0 ;
      RECT  30590.0 112110.0 31295.0 113455.0 ;
      RECT  30590.0 114800.0 31295.0 113455.0 ;
      RECT  30590.0 114800.0 31295.0 116145.0 ;
      RECT  30590.0 117490.0 31295.0 116145.0 ;
      RECT  30590.0 117490.0 31295.0 118835.0 ;
      RECT  30590.0 120180.0 31295.0 118835.0 ;
      RECT  30590.0 120180.0 31295.0 121525.0 ;
      RECT  30590.0 122870.0 31295.0 121525.0 ;
      RECT  30590.0 122870.0 31295.0 124215.0 ;
      RECT  30590.0 125560.0 31295.0 124215.0 ;
      RECT  30590.0 125560.0 31295.0 126905.0 ;
      RECT  30590.0 128250.0 31295.0 126905.0 ;
      RECT  30590.0 128250.0 31295.0 129595.0 ;
      RECT  30590.0 130940.0 31295.0 129595.0 ;
      RECT  30590.0 130940.0 31295.0 132285.0 ;
      RECT  30590.0 133630.0 31295.0 132285.0 ;
      RECT  30590.0 133630.0 31295.0 134975.0 ;
      RECT  30590.0 136320.0 31295.0 134975.0 ;
      RECT  30590.0 136320.0 31295.0 137665.0 ;
      RECT  30590.0 139010.0 31295.0 137665.0 ;
      RECT  30590.0 139010.0 31295.0 140355.0 ;
      RECT  30590.0 141700.0 31295.0 140355.0 ;
      RECT  30590.0 141700.0 31295.0 143045.0 ;
      RECT  30590.0 144390.0 31295.0 143045.0 ;
      RECT  30590.0 144390.0 31295.0 145735.0 ;
      RECT  30590.0 147080.0 31295.0 145735.0 ;
      RECT  30590.0 147080.0 31295.0 148425.0 ;
      RECT  30590.0 149770.0 31295.0 148425.0 ;
      RECT  30590.0 149770.0 31295.0 151115.0 ;
      RECT  30590.0 152460.0 31295.0 151115.0 ;
      RECT  30590.0 152460.0 31295.0 153805.0 ;
      RECT  30590.0 155150.0 31295.0 153805.0 ;
      RECT  30590.0 155150.0 31295.0 156495.0 ;
      RECT  30590.0 157840.0 31295.0 156495.0 ;
      RECT  30590.0 157840.0 31295.0 159185.0 ;
      RECT  30590.0 160530.0 31295.0 159185.0 ;
      RECT  30590.0 160530.0 31295.0 161875.0 ;
      RECT  30590.0 163220.0 31295.0 161875.0 ;
      RECT  30590.0 163220.0 31295.0 164565.0 ;
      RECT  30590.0 165910.0 31295.0 164565.0 ;
      RECT  30590.0 165910.0 31295.0 167255.0 ;
      RECT  30590.0 168600.0 31295.0 167255.0 ;
      RECT  30590.0 168600.0 31295.0 169945.0 ;
      RECT  30590.0 171290.0 31295.0 169945.0 ;
      RECT  30590.0 171290.0 31295.0 172635.0 ;
      RECT  30590.0 173980.0 31295.0 172635.0 ;
      RECT  30590.0 173980.0 31295.0 175325.0 ;
      RECT  30590.0 176670.0 31295.0 175325.0 ;
      RECT  30590.0 176670.0 31295.0 178015.0 ;
      RECT  30590.0 179360.0 31295.0 178015.0 ;
      RECT  30590.0 179360.0 31295.0 180705.0 ;
      RECT  30590.0 182050.0 31295.0 180705.0 ;
      RECT  30590.0 182050.0 31295.0 183395.0 ;
      RECT  30590.0 184740.0 31295.0 183395.0 ;
      RECT  30590.0 184740.0 31295.0 186085.0 ;
      RECT  30590.0 187430.0 31295.0 186085.0 ;
      RECT  30590.0 187430.0 31295.0 188775.0 ;
      RECT  30590.0 190120.0 31295.0 188775.0 ;
      RECT  30590.0 190120.0 31295.0 191465.0 ;
      RECT  30590.0 192810.0 31295.0 191465.0 ;
      RECT  30590.0 192810.0 31295.0 194155.0 ;
      RECT  30590.0 195500.0 31295.0 194155.0 ;
      RECT  30590.0 195500.0 31295.0 196845.0 ;
      RECT  30590.0 198190.0 31295.0 196845.0 ;
      RECT  30590.0 198190.0 31295.0 199535.0 ;
      RECT  30590.0 200880.0 31295.0 199535.0 ;
      RECT  30590.0 200880.0 31295.0 202225.0 ;
      RECT  30590.0 203570.0 31295.0 202225.0 ;
      RECT  30590.0 203570.0 31295.0 204915.0 ;
      RECT  30590.0 206260.0 31295.0 204915.0 ;
      RECT  31295.0 34100.0 32000.0 35445.0 ;
      RECT  31295.0 36790.0 32000.0 35445.0 ;
      RECT  31295.0 36790.0 32000.0 38135.0 ;
      RECT  31295.0 39480.0 32000.0 38135.0 ;
      RECT  31295.0 39480.0 32000.0 40825.0 ;
      RECT  31295.0 42170.0 32000.0 40825.0 ;
      RECT  31295.0 42170.0 32000.0 43515.0 ;
      RECT  31295.0 44860.0 32000.0 43515.0 ;
      RECT  31295.0 44860.0 32000.0 46205.0 ;
      RECT  31295.0 47550.0 32000.0 46205.0 ;
      RECT  31295.0 47550.0 32000.0 48895.0 ;
      RECT  31295.0 50240.0 32000.0 48895.0 ;
      RECT  31295.0 50240.0 32000.0 51585.0 ;
      RECT  31295.0 52930.0 32000.0 51585.0 ;
      RECT  31295.0 52930.0 32000.0 54275.0 ;
      RECT  31295.0 55620.0 32000.0 54275.0 ;
      RECT  31295.0 55620.0 32000.0 56965.0 ;
      RECT  31295.0 58310.0 32000.0 56965.0 ;
      RECT  31295.0 58310.0 32000.0 59655.0 ;
      RECT  31295.0 61000.0 32000.0 59655.0 ;
      RECT  31295.0 61000.0 32000.0 62345.0 ;
      RECT  31295.0 63690.0 32000.0 62345.0 ;
      RECT  31295.0 63690.0 32000.0 65035.0 ;
      RECT  31295.0 66380.0 32000.0 65035.0 ;
      RECT  31295.0 66380.0 32000.0 67725.0 ;
      RECT  31295.0 69070.0 32000.0 67725.0 ;
      RECT  31295.0 69070.0 32000.0 70415.0 ;
      RECT  31295.0 71760.0 32000.0 70415.0 ;
      RECT  31295.0 71760.0 32000.0 73105.0 ;
      RECT  31295.0 74450.0 32000.0 73105.0 ;
      RECT  31295.0 74450.0 32000.0 75795.0 ;
      RECT  31295.0 77140.0 32000.0 75795.0 ;
      RECT  31295.0 77140.0 32000.0 78485.0 ;
      RECT  31295.0 79830.0 32000.0 78485.0 ;
      RECT  31295.0 79830.0 32000.0 81175.0 ;
      RECT  31295.0 82520.0 32000.0 81175.0 ;
      RECT  31295.0 82520.0 32000.0 83865.0 ;
      RECT  31295.0 85210.0 32000.0 83865.0 ;
      RECT  31295.0 85210.0 32000.0 86555.0 ;
      RECT  31295.0 87900.0 32000.0 86555.0 ;
      RECT  31295.0 87900.0 32000.0 89245.0 ;
      RECT  31295.0 90590.0 32000.0 89245.0 ;
      RECT  31295.0 90590.0 32000.0 91935.0 ;
      RECT  31295.0 93280.0 32000.0 91935.0 ;
      RECT  31295.0 93280.0 32000.0 94625.0 ;
      RECT  31295.0 95970.0 32000.0 94625.0 ;
      RECT  31295.0 95970.0 32000.0 97315.0 ;
      RECT  31295.0 98660.0 32000.0 97315.0 ;
      RECT  31295.0 98660.0 32000.0 100005.0 ;
      RECT  31295.0 101350.0 32000.0 100005.0 ;
      RECT  31295.0 101350.0 32000.0 102695.0 ;
      RECT  31295.0 104040.0 32000.0 102695.0 ;
      RECT  31295.0 104040.0 32000.0 105385.0 ;
      RECT  31295.0 106730.0 32000.0 105385.0 ;
      RECT  31295.0 106730.0 32000.0 108075.0 ;
      RECT  31295.0 109420.0 32000.0 108075.0 ;
      RECT  31295.0 109420.0 32000.0 110765.0 ;
      RECT  31295.0 112110.0 32000.0 110765.0 ;
      RECT  31295.0 112110.0 32000.0 113455.0 ;
      RECT  31295.0 114800.0 32000.0 113455.0 ;
      RECT  31295.0 114800.0 32000.0 116145.0 ;
      RECT  31295.0 117490.0 32000.0 116145.0 ;
      RECT  31295.0 117490.0 32000.0 118835.0 ;
      RECT  31295.0 120180.0 32000.0 118835.0 ;
      RECT  31295.0 120180.0 32000.0 121525.0 ;
      RECT  31295.0 122870.0 32000.0 121525.0 ;
      RECT  31295.0 122870.0 32000.0 124215.0 ;
      RECT  31295.0 125560.0 32000.0 124215.0 ;
      RECT  31295.0 125560.0 32000.0 126905.0 ;
      RECT  31295.0 128250.0 32000.0 126905.0 ;
      RECT  31295.0 128250.0 32000.0 129595.0 ;
      RECT  31295.0 130940.0 32000.0 129595.0 ;
      RECT  31295.0 130940.0 32000.0 132285.0 ;
      RECT  31295.0 133630.0 32000.0 132285.0 ;
      RECT  31295.0 133630.0 32000.0 134975.0 ;
      RECT  31295.0 136320.0 32000.0 134975.0 ;
      RECT  31295.0 136320.0 32000.0 137665.0 ;
      RECT  31295.0 139010.0 32000.0 137665.0 ;
      RECT  31295.0 139010.0 32000.0 140355.0 ;
      RECT  31295.0 141700.0 32000.0 140355.0 ;
      RECT  31295.0 141700.0 32000.0 143045.0 ;
      RECT  31295.0 144390.0 32000.0 143045.0 ;
      RECT  31295.0 144390.0 32000.0 145735.0 ;
      RECT  31295.0 147080.0 32000.0 145735.0 ;
      RECT  31295.0 147080.0 32000.0 148425.0 ;
      RECT  31295.0 149770.0 32000.0 148425.0 ;
      RECT  31295.0 149770.0 32000.0 151115.0 ;
      RECT  31295.0 152460.0 32000.0 151115.0 ;
      RECT  31295.0 152460.0 32000.0 153805.0 ;
      RECT  31295.0 155150.0 32000.0 153805.0 ;
      RECT  31295.0 155150.0 32000.0 156495.0 ;
      RECT  31295.0 157840.0 32000.0 156495.0 ;
      RECT  31295.0 157840.0 32000.0 159185.0 ;
      RECT  31295.0 160530.0 32000.0 159185.0 ;
      RECT  31295.0 160530.0 32000.0 161875.0 ;
      RECT  31295.0 163220.0 32000.0 161875.0 ;
      RECT  31295.0 163220.0 32000.0 164565.0 ;
      RECT  31295.0 165910.0 32000.0 164565.0 ;
      RECT  31295.0 165910.0 32000.0 167255.0 ;
      RECT  31295.0 168600.0 32000.0 167255.0 ;
      RECT  31295.0 168600.0 32000.0 169945.0 ;
      RECT  31295.0 171290.0 32000.0 169945.0 ;
      RECT  31295.0 171290.0 32000.0 172635.0 ;
      RECT  31295.0 173980.0 32000.0 172635.0 ;
      RECT  31295.0 173980.0 32000.0 175325.0 ;
      RECT  31295.0 176670.0 32000.0 175325.0 ;
      RECT  31295.0 176670.0 32000.0 178015.0 ;
      RECT  31295.0 179360.0 32000.0 178015.0 ;
      RECT  31295.0 179360.0 32000.0 180705.0 ;
      RECT  31295.0 182050.0 32000.0 180705.0 ;
      RECT  31295.0 182050.0 32000.0 183395.0 ;
      RECT  31295.0 184740.0 32000.0 183395.0 ;
      RECT  31295.0 184740.0 32000.0 186085.0 ;
      RECT  31295.0 187430.0 32000.0 186085.0 ;
      RECT  31295.0 187430.0 32000.0 188775.0 ;
      RECT  31295.0 190120.0 32000.0 188775.0 ;
      RECT  31295.0 190120.0 32000.0 191465.0 ;
      RECT  31295.0 192810.0 32000.0 191465.0 ;
      RECT  31295.0 192810.0 32000.0 194155.0 ;
      RECT  31295.0 195500.0 32000.0 194155.0 ;
      RECT  31295.0 195500.0 32000.0 196845.0 ;
      RECT  31295.0 198190.0 32000.0 196845.0 ;
      RECT  31295.0 198190.0 32000.0 199535.0 ;
      RECT  31295.0 200880.0 32000.0 199535.0 ;
      RECT  31295.0 200880.0 32000.0 202225.0 ;
      RECT  31295.0 203570.0 32000.0 202225.0 ;
      RECT  31295.0 203570.0 32000.0 204915.0 ;
      RECT  31295.0 206260.0 32000.0 204915.0 ;
      RECT  32000.0 34100.0 32705.0 35445.0 ;
      RECT  32000.0 36790.0 32705.0 35445.0 ;
      RECT  32000.0 36790.0 32705.0 38135.0 ;
      RECT  32000.0 39480.0 32705.0 38135.0 ;
      RECT  32000.0 39480.0 32705.0 40825.0 ;
      RECT  32000.0 42170.0 32705.0 40825.0 ;
      RECT  32000.0 42170.0 32705.0 43515.0 ;
      RECT  32000.0 44860.0 32705.0 43515.0 ;
      RECT  32000.0 44860.0 32705.0 46205.0 ;
      RECT  32000.0 47550.0 32705.0 46205.0 ;
      RECT  32000.0 47550.0 32705.0 48895.0 ;
      RECT  32000.0 50240.0 32705.0 48895.0 ;
      RECT  32000.0 50240.0 32705.0 51585.0 ;
      RECT  32000.0 52930.0 32705.0 51585.0 ;
      RECT  32000.0 52930.0 32705.0 54275.0 ;
      RECT  32000.0 55620.0 32705.0 54275.0 ;
      RECT  32000.0 55620.0 32705.0 56965.0 ;
      RECT  32000.0 58310.0 32705.0 56965.0 ;
      RECT  32000.0 58310.0 32705.0 59655.0 ;
      RECT  32000.0 61000.0 32705.0 59655.0 ;
      RECT  32000.0 61000.0 32705.0 62345.0 ;
      RECT  32000.0 63690.0 32705.0 62345.0 ;
      RECT  32000.0 63690.0 32705.0 65035.0 ;
      RECT  32000.0 66380.0 32705.0 65035.0 ;
      RECT  32000.0 66380.0 32705.0 67725.0 ;
      RECT  32000.0 69070.0 32705.0 67725.0 ;
      RECT  32000.0 69070.0 32705.0 70415.0 ;
      RECT  32000.0 71760.0 32705.0 70415.0 ;
      RECT  32000.0 71760.0 32705.0 73105.0 ;
      RECT  32000.0 74450.0 32705.0 73105.0 ;
      RECT  32000.0 74450.0 32705.0 75795.0 ;
      RECT  32000.0 77140.0 32705.0 75795.0 ;
      RECT  32000.0 77140.0 32705.0 78485.0 ;
      RECT  32000.0 79830.0 32705.0 78485.0 ;
      RECT  32000.0 79830.0 32705.0 81175.0 ;
      RECT  32000.0 82520.0 32705.0 81175.0 ;
      RECT  32000.0 82520.0 32705.0 83865.0 ;
      RECT  32000.0 85210.0 32705.0 83865.0 ;
      RECT  32000.0 85210.0 32705.0 86555.0 ;
      RECT  32000.0 87900.0 32705.0 86555.0 ;
      RECT  32000.0 87900.0 32705.0 89245.0 ;
      RECT  32000.0 90590.0 32705.0 89245.0 ;
      RECT  32000.0 90590.0 32705.0 91935.0 ;
      RECT  32000.0 93280.0 32705.0 91935.0 ;
      RECT  32000.0 93280.0 32705.0 94625.0 ;
      RECT  32000.0 95970.0 32705.0 94625.0 ;
      RECT  32000.0 95970.0 32705.0 97315.0 ;
      RECT  32000.0 98660.0 32705.0 97315.0 ;
      RECT  32000.0 98660.0 32705.0 100005.0 ;
      RECT  32000.0 101350.0 32705.0 100005.0 ;
      RECT  32000.0 101350.0 32705.0 102695.0 ;
      RECT  32000.0 104040.0 32705.0 102695.0 ;
      RECT  32000.0 104040.0 32705.0 105385.0 ;
      RECT  32000.0 106730.0 32705.0 105385.0 ;
      RECT  32000.0 106730.0 32705.0 108075.0 ;
      RECT  32000.0 109420.0 32705.0 108075.0 ;
      RECT  32000.0 109420.0 32705.0 110765.0 ;
      RECT  32000.0 112110.0 32705.0 110765.0 ;
      RECT  32000.0 112110.0 32705.0 113455.0 ;
      RECT  32000.0 114800.0 32705.0 113455.0 ;
      RECT  32000.0 114800.0 32705.0 116145.0 ;
      RECT  32000.0 117490.0 32705.0 116145.0 ;
      RECT  32000.0 117490.0 32705.0 118835.0 ;
      RECT  32000.0 120180.0 32705.0 118835.0 ;
      RECT  32000.0 120180.0 32705.0 121525.0 ;
      RECT  32000.0 122870.0 32705.0 121525.0 ;
      RECT  32000.0 122870.0 32705.0 124215.0 ;
      RECT  32000.0 125560.0 32705.0 124215.0 ;
      RECT  32000.0 125560.0 32705.0 126905.0 ;
      RECT  32000.0 128250.0 32705.0 126905.0 ;
      RECT  32000.0 128250.0 32705.0 129595.0 ;
      RECT  32000.0 130940.0 32705.0 129595.0 ;
      RECT  32000.0 130940.0 32705.0 132285.0 ;
      RECT  32000.0 133630.0 32705.0 132285.0 ;
      RECT  32000.0 133630.0 32705.0 134975.0 ;
      RECT  32000.0 136320.0 32705.0 134975.0 ;
      RECT  32000.0 136320.0 32705.0 137665.0 ;
      RECT  32000.0 139010.0 32705.0 137665.0 ;
      RECT  32000.0 139010.0 32705.0 140355.0 ;
      RECT  32000.0 141700.0 32705.0 140355.0 ;
      RECT  32000.0 141700.0 32705.0 143045.0 ;
      RECT  32000.0 144390.0 32705.0 143045.0 ;
      RECT  32000.0 144390.0 32705.0 145735.0 ;
      RECT  32000.0 147080.0 32705.0 145735.0 ;
      RECT  32000.0 147080.0 32705.0 148425.0 ;
      RECT  32000.0 149770.0 32705.0 148425.0 ;
      RECT  32000.0 149770.0 32705.0 151115.0 ;
      RECT  32000.0 152460.0 32705.0 151115.0 ;
      RECT  32000.0 152460.0 32705.0 153805.0 ;
      RECT  32000.0 155150.0 32705.0 153805.0 ;
      RECT  32000.0 155150.0 32705.0 156495.0 ;
      RECT  32000.0 157840.0 32705.0 156495.0 ;
      RECT  32000.0 157840.0 32705.0 159185.0 ;
      RECT  32000.0 160530.0 32705.0 159185.0 ;
      RECT  32000.0 160530.0 32705.0 161875.0 ;
      RECT  32000.0 163220.0 32705.0 161875.0 ;
      RECT  32000.0 163220.0 32705.0 164565.0 ;
      RECT  32000.0 165910.0 32705.0 164565.0 ;
      RECT  32000.0 165910.0 32705.0 167255.0 ;
      RECT  32000.0 168600.0 32705.0 167255.0 ;
      RECT  32000.0 168600.0 32705.0 169945.0 ;
      RECT  32000.0 171290.0 32705.0 169945.0 ;
      RECT  32000.0 171290.0 32705.0 172635.0 ;
      RECT  32000.0 173980.0 32705.0 172635.0 ;
      RECT  32000.0 173980.0 32705.0 175325.0 ;
      RECT  32000.0 176670.0 32705.0 175325.0 ;
      RECT  32000.0 176670.0 32705.0 178015.0 ;
      RECT  32000.0 179360.0 32705.0 178015.0 ;
      RECT  32000.0 179360.0 32705.0 180705.0 ;
      RECT  32000.0 182050.0 32705.0 180705.0 ;
      RECT  32000.0 182050.0 32705.0 183395.0 ;
      RECT  32000.0 184740.0 32705.0 183395.0 ;
      RECT  32000.0 184740.0 32705.0 186085.0 ;
      RECT  32000.0 187430.0 32705.0 186085.0 ;
      RECT  32000.0 187430.0 32705.0 188775.0 ;
      RECT  32000.0 190120.0 32705.0 188775.0 ;
      RECT  32000.0 190120.0 32705.0 191465.0 ;
      RECT  32000.0 192810.0 32705.0 191465.0 ;
      RECT  32000.0 192810.0 32705.0 194155.0 ;
      RECT  32000.0 195500.0 32705.0 194155.0 ;
      RECT  32000.0 195500.0 32705.0 196845.0 ;
      RECT  32000.0 198190.0 32705.0 196845.0 ;
      RECT  32000.0 198190.0 32705.0 199535.0 ;
      RECT  32000.0 200880.0 32705.0 199535.0 ;
      RECT  32000.0 200880.0 32705.0 202225.0 ;
      RECT  32000.0 203570.0 32705.0 202225.0 ;
      RECT  32000.0 203570.0 32705.0 204915.0 ;
      RECT  32000.0 206260.0 32705.0 204915.0 ;
      RECT  32705.0 34100.0 33410.0 35445.0 ;
      RECT  32705.0 36790.0 33410.0 35445.0 ;
      RECT  32705.0 36790.0 33410.0 38135.0 ;
      RECT  32705.0 39480.0 33410.0 38135.0 ;
      RECT  32705.0 39480.0 33410.0 40825.0 ;
      RECT  32705.0 42170.0 33410.0 40825.0 ;
      RECT  32705.0 42170.0 33410.0 43515.0 ;
      RECT  32705.0 44860.0 33410.0 43515.0 ;
      RECT  32705.0 44860.0 33410.0 46205.0 ;
      RECT  32705.0 47550.0 33410.0 46205.0 ;
      RECT  32705.0 47550.0 33410.0 48895.0 ;
      RECT  32705.0 50240.0 33410.0 48895.0 ;
      RECT  32705.0 50240.0 33410.0 51585.0 ;
      RECT  32705.0 52930.0 33410.0 51585.0 ;
      RECT  32705.0 52930.0 33410.0 54275.0 ;
      RECT  32705.0 55620.0 33410.0 54275.0 ;
      RECT  32705.0 55620.0 33410.0 56965.0 ;
      RECT  32705.0 58310.0 33410.0 56965.0 ;
      RECT  32705.0 58310.0 33410.0 59655.0 ;
      RECT  32705.0 61000.0 33410.0 59655.0 ;
      RECT  32705.0 61000.0 33410.0 62345.0 ;
      RECT  32705.0 63690.0 33410.0 62345.0 ;
      RECT  32705.0 63690.0 33410.0 65035.0 ;
      RECT  32705.0 66380.0 33410.0 65035.0 ;
      RECT  32705.0 66380.0 33410.0 67725.0 ;
      RECT  32705.0 69070.0 33410.0 67725.0 ;
      RECT  32705.0 69070.0 33410.0 70415.0 ;
      RECT  32705.0 71760.0 33410.0 70415.0 ;
      RECT  32705.0 71760.0 33410.0 73105.0 ;
      RECT  32705.0 74450.0 33410.0 73105.0 ;
      RECT  32705.0 74450.0 33410.0 75795.0 ;
      RECT  32705.0 77140.0 33410.0 75795.0 ;
      RECT  32705.0 77140.0 33410.0 78485.0 ;
      RECT  32705.0 79830.0 33410.0 78485.0 ;
      RECT  32705.0 79830.0 33410.0 81175.0 ;
      RECT  32705.0 82520.0 33410.0 81175.0 ;
      RECT  32705.0 82520.0 33410.0 83865.0 ;
      RECT  32705.0 85210.0 33410.0 83865.0 ;
      RECT  32705.0 85210.0 33410.0 86555.0 ;
      RECT  32705.0 87900.0 33410.0 86555.0 ;
      RECT  32705.0 87900.0 33410.0 89245.0 ;
      RECT  32705.0 90590.0 33410.0 89245.0 ;
      RECT  32705.0 90590.0 33410.0 91935.0 ;
      RECT  32705.0 93280.0 33410.0 91935.0 ;
      RECT  32705.0 93280.0 33410.0 94625.0 ;
      RECT  32705.0 95970.0 33410.0 94625.0 ;
      RECT  32705.0 95970.0 33410.0 97315.0 ;
      RECT  32705.0 98660.0 33410.0 97315.0 ;
      RECT  32705.0 98660.0 33410.0 100005.0 ;
      RECT  32705.0 101350.0 33410.0 100005.0 ;
      RECT  32705.0 101350.0 33410.0 102695.0 ;
      RECT  32705.0 104040.0 33410.0 102695.0 ;
      RECT  32705.0 104040.0 33410.0 105385.0 ;
      RECT  32705.0 106730.0 33410.0 105385.0 ;
      RECT  32705.0 106730.0 33410.0 108075.0 ;
      RECT  32705.0 109420.0 33410.0 108075.0 ;
      RECT  32705.0 109420.0 33410.0 110765.0 ;
      RECT  32705.0 112110.0 33410.0 110765.0 ;
      RECT  32705.0 112110.0 33410.0 113455.0 ;
      RECT  32705.0 114800.0 33410.0 113455.0 ;
      RECT  32705.0 114800.0 33410.0 116145.0 ;
      RECT  32705.0 117490.0 33410.0 116145.0 ;
      RECT  32705.0 117490.0 33410.0 118835.0 ;
      RECT  32705.0 120180.0 33410.0 118835.0 ;
      RECT  32705.0 120180.0 33410.0 121525.0 ;
      RECT  32705.0 122870.0 33410.0 121525.0 ;
      RECT  32705.0 122870.0 33410.0 124215.0 ;
      RECT  32705.0 125560.0 33410.0 124215.0 ;
      RECT  32705.0 125560.0 33410.0 126905.0 ;
      RECT  32705.0 128250.0 33410.0 126905.0 ;
      RECT  32705.0 128250.0 33410.0 129595.0 ;
      RECT  32705.0 130940.0 33410.0 129595.0 ;
      RECT  32705.0 130940.0 33410.0 132285.0 ;
      RECT  32705.0 133630.0 33410.0 132285.0 ;
      RECT  32705.0 133630.0 33410.0 134975.0 ;
      RECT  32705.0 136320.0 33410.0 134975.0 ;
      RECT  32705.0 136320.0 33410.0 137665.0 ;
      RECT  32705.0 139010.0 33410.0 137665.0 ;
      RECT  32705.0 139010.0 33410.0 140355.0 ;
      RECT  32705.0 141700.0 33410.0 140355.0 ;
      RECT  32705.0 141700.0 33410.0 143045.0 ;
      RECT  32705.0 144390.0 33410.0 143045.0 ;
      RECT  32705.0 144390.0 33410.0 145735.0 ;
      RECT  32705.0 147080.0 33410.0 145735.0 ;
      RECT  32705.0 147080.0 33410.0 148425.0 ;
      RECT  32705.0 149770.0 33410.0 148425.0 ;
      RECT  32705.0 149770.0 33410.0 151115.0 ;
      RECT  32705.0 152460.0 33410.0 151115.0 ;
      RECT  32705.0 152460.0 33410.0 153805.0 ;
      RECT  32705.0 155150.0 33410.0 153805.0 ;
      RECT  32705.0 155150.0 33410.0 156495.0 ;
      RECT  32705.0 157840.0 33410.0 156495.0 ;
      RECT  32705.0 157840.0 33410.0 159185.0 ;
      RECT  32705.0 160530.0 33410.0 159185.0 ;
      RECT  32705.0 160530.0 33410.0 161875.0 ;
      RECT  32705.0 163220.0 33410.0 161875.0 ;
      RECT  32705.0 163220.0 33410.0 164565.0 ;
      RECT  32705.0 165910.0 33410.0 164565.0 ;
      RECT  32705.0 165910.0 33410.0 167255.0 ;
      RECT  32705.0 168600.0 33410.0 167255.0 ;
      RECT  32705.0 168600.0 33410.0 169945.0 ;
      RECT  32705.0 171290.0 33410.0 169945.0 ;
      RECT  32705.0 171290.0 33410.0 172635.0 ;
      RECT  32705.0 173980.0 33410.0 172635.0 ;
      RECT  32705.0 173980.0 33410.0 175325.0 ;
      RECT  32705.0 176670.0 33410.0 175325.0 ;
      RECT  32705.0 176670.0 33410.0 178015.0 ;
      RECT  32705.0 179360.0 33410.0 178015.0 ;
      RECT  32705.0 179360.0 33410.0 180705.0 ;
      RECT  32705.0 182050.0 33410.0 180705.0 ;
      RECT  32705.0 182050.0 33410.0 183395.0 ;
      RECT  32705.0 184740.0 33410.0 183395.0 ;
      RECT  32705.0 184740.0 33410.0 186085.0 ;
      RECT  32705.0 187430.0 33410.0 186085.0 ;
      RECT  32705.0 187430.0 33410.0 188775.0 ;
      RECT  32705.0 190120.0 33410.0 188775.0 ;
      RECT  32705.0 190120.0 33410.0 191465.0 ;
      RECT  32705.0 192810.0 33410.0 191465.0 ;
      RECT  32705.0 192810.0 33410.0 194155.0 ;
      RECT  32705.0 195500.0 33410.0 194155.0 ;
      RECT  32705.0 195500.0 33410.0 196845.0 ;
      RECT  32705.0 198190.0 33410.0 196845.0 ;
      RECT  32705.0 198190.0 33410.0 199535.0 ;
      RECT  32705.0 200880.0 33410.0 199535.0 ;
      RECT  32705.0 200880.0 33410.0 202225.0 ;
      RECT  32705.0 203570.0 33410.0 202225.0 ;
      RECT  32705.0 203570.0 33410.0 204915.0 ;
      RECT  32705.0 206260.0 33410.0 204915.0 ;
      RECT  33410.0 34100.0 34115.0 35445.0 ;
      RECT  33410.0 36790.0 34115.0 35445.0 ;
      RECT  33410.0 36790.0 34115.0 38135.0 ;
      RECT  33410.0 39480.0 34115.0 38135.0 ;
      RECT  33410.0 39480.0 34115.0 40825.0 ;
      RECT  33410.0 42170.0 34115.0 40825.0 ;
      RECT  33410.0 42170.0 34115.0 43515.0 ;
      RECT  33410.0 44860.0 34115.0 43515.0 ;
      RECT  33410.0 44860.0 34115.0 46205.0 ;
      RECT  33410.0 47550.0 34115.0 46205.0 ;
      RECT  33410.0 47550.0 34115.0 48895.0 ;
      RECT  33410.0 50240.0 34115.0 48895.0 ;
      RECT  33410.0 50240.0 34115.0 51585.0 ;
      RECT  33410.0 52930.0 34115.0 51585.0 ;
      RECT  33410.0 52930.0 34115.0 54275.0 ;
      RECT  33410.0 55620.0 34115.0 54275.0 ;
      RECT  33410.0 55620.0 34115.0 56965.0 ;
      RECT  33410.0 58310.0 34115.0 56965.0 ;
      RECT  33410.0 58310.0 34115.0 59655.0 ;
      RECT  33410.0 61000.0 34115.0 59655.0 ;
      RECT  33410.0 61000.0 34115.0 62345.0 ;
      RECT  33410.0 63690.0 34115.0 62345.0 ;
      RECT  33410.0 63690.0 34115.0 65035.0 ;
      RECT  33410.0 66380.0 34115.0 65035.0 ;
      RECT  33410.0 66380.0 34115.0 67725.0 ;
      RECT  33410.0 69070.0 34115.0 67725.0 ;
      RECT  33410.0 69070.0 34115.0 70415.0 ;
      RECT  33410.0 71760.0 34115.0 70415.0 ;
      RECT  33410.0 71760.0 34115.0 73105.0 ;
      RECT  33410.0 74450.0 34115.0 73105.0 ;
      RECT  33410.0 74450.0 34115.0 75795.0 ;
      RECT  33410.0 77140.0 34115.0 75795.0 ;
      RECT  33410.0 77140.0 34115.0 78485.0 ;
      RECT  33410.0 79830.0 34115.0 78485.0 ;
      RECT  33410.0 79830.0 34115.0 81175.0 ;
      RECT  33410.0 82520.0 34115.0 81175.0 ;
      RECT  33410.0 82520.0 34115.0 83865.0 ;
      RECT  33410.0 85210.0 34115.0 83865.0 ;
      RECT  33410.0 85210.0 34115.0 86555.0 ;
      RECT  33410.0 87900.0 34115.0 86555.0 ;
      RECT  33410.0 87900.0 34115.0 89245.0 ;
      RECT  33410.0 90590.0 34115.0 89245.0 ;
      RECT  33410.0 90590.0 34115.0 91935.0 ;
      RECT  33410.0 93280.0 34115.0 91935.0 ;
      RECT  33410.0 93280.0 34115.0 94625.0 ;
      RECT  33410.0 95970.0 34115.0 94625.0 ;
      RECT  33410.0 95970.0 34115.0 97315.0 ;
      RECT  33410.0 98660.0 34115.0 97315.0 ;
      RECT  33410.0 98660.0 34115.0 100005.0 ;
      RECT  33410.0 101350.0 34115.0 100005.0 ;
      RECT  33410.0 101350.0 34115.0 102695.0 ;
      RECT  33410.0 104040.0 34115.0 102695.0 ;
      RECT  33410.0 104040.0 34115.0 105385.0 ;
      RECT  33410.0 106730.0 34115.0 105385.0 ;
      RECT  33410.0 106730.0 34115.0 108075.0 ;
      RECT  33410.0 109420.0 34115.0 108075.0 ;
      RECT  33410.0 109420.0 34115.0 110765.0 ;
      RECT  33410.0 112110.0 34115.0 110765.0 ;
      RECT  33410.0 112110.0 34115.0 113455.0 ;
      RECT  33410.0 114800.0 34115.0 113455.0 ;
      RECT  33410.0 114800.0 34115.0 116145.0 ;
      RECT  33410.0 117490.0 34115.0 116145.0 ;
      RECT  33410.0 117490.0 34115.0 118835.0 ;
      RECT  33410.0 120180.0 34115.0 118835.0 ;
      RECT  33410.0 120180.0 34115.0 121525.0 ;
      RECT  33410.0 122870.0 34115.0 121525.0 ;
      RECT  33410.0 122870.0 34115.0 124215.0 ;
      RECT  33410.0 125560.0 34115.0 124215.0 ;
      RECT  33410.0 125560.0 34115.0 126905.0 ;
      RECT  33410.0 128250.0 34115.0 126905.0 ;
      RECT  33410.0 128250.0 34115.0 129595.0 ;
      RECT  33410.0 130940.0 34115.0 129595.0 ;
      RECT  33410.0 130940.0 34115.0 132285.0 ;
      RECT  33410.0 133630.0 34115.0 132285.0 ;
      RECT  33410.0 133630.0 34115.0 134975.0 ;
      RECT  33410.0 136320.0 34115.0 134975.0 ;
      RECT  33410.0 136320.0 34115.0 137665.0 ;
      RECT  33410.0 139010.0 34115.0 137665.0 ;
      RECT  33410.0 139010.0 34115.0 140355.0 ;
      RECT  33410.0 141700.0 34115.0 140355.0 ;
      RECT  33410.0 141700.0 34115.0 143045.0 ;
      RECT  33410.0 144390.0 34115.0 143045.0 ;
      RECT  33410.0 144390.0 34115.0 145735.0 ;
      RECT  33410.0 147080.0 34115.0 145735.0 ;
      RECT  33410.0 147080.0 34115.0 148425.0 ;
      RECT  33410.0 149770.0 34115.0 148425.0 ;
      RECT  33410.0 149770.0 34115.0 151115.0 ;
      RECT  33410.0 152460.0 34115.0 151115.0 ;
      RECT  33410.0 152460.0 34115.0 153805.0 ;
      RECT  33410.0 155150.0 34115.0 153805.0 ;
      RECT  33410.0 155150.0 34115.0 156495.0 ;
      RECT  33410.0 157840.0 34115.0 156495.0 ;
      RECT  33410.0 157840.0 34115.0 159185.0 ;
      RECT  33410.0 160530.0 34115.0 159185.0 ;
      RECT  33410.0 160530.0 34115.0 161875.0 ;
      RECT  33410.0 163220.0 34115.0 161875.0 ;
      RECT  33410.0 163220.0 34115.0 164565.0 ;
      RECT  33410.0 165910.0 34115.0 164565.0 ;
      RECT  33410.0 165910.0 34115.0 167255.0 ;
      RECT  33410.0 168600.0 34115.0 167255.0 ;
      RECT  33410.0 168600.0 34115.0 169945.0 ;
      RECT  33410.0 171290.0 34115.0 169945.0 ;
      RECT  33410.0 171290.0 34115.0 172635.0 ;
      RECT  33410.0 173980.0 34115.0 172635.0 ;
      RECT  33410.0 173980.0 34115.0 175325.0 ;
      RECT  33410.0 176670.0 34115.0 175325.0 ;
      RECT  33410.0 176670.0 34115.0 178015.0 ;
      RECT  33410.0 179360.0 34115.0 178015.0 ;
      RECT  33410.0 179360.0 34115.0 180705.0 ;
      RECT  33410.0 182050.0 34115.0 180705.0 ;
      RECT  33410.0 182050.0 34115.0 183395.0 ;
      RECT  33410.0 184740.0 34115.0 183395.0 ;
      RECT  33410.0 184740.0 34115.0 186085.0 ;
      RECT  33410.0 187430.0 34115.0 186085.0 ;
      RECT  33410.0 187430.0 34115.0 188775.0 ;
      RECT  33410.0 190120.0 34115.0 188775.0 ;
      RECT  33410.0 190120.0 34115.0 191465.0 ;
      RECT  33410.0 192810.0 34115.0 191465.0 ;
      RECT  33410.0 192810.0 34115.0 194155.0 ;
      RECT  33410.0 195500.0 34115.0 194155.0 ;
      RECT  33410.0 195500.0 34115.0 196845.0 ;
      RECT  33410.0 198190.0 34115.0 196845.0 ;
      RECT  33410.0 198190.0 34115.0 199535.0 ;
      RECT  33410.0 200880.0 34115.0 199535.0 ;
      RECT  33410.0 200880.0 34115.0 202225.0 ;
      RECT  33410.0 203570.0 34115.0 202225.0 ;
      RECT  33410.0 203570.0 34115.0 204915.0 ;
      RECT  33410.0 206260.0 34115.0 204915.0 ;
      RECT  34115.0 34100.0 34820.0 35445.0 ;
      RECT  34115.0 36790.0 34820.0 35445.0 ;
      RECT  34115.0 36790.0 34820.0 38135.0 ;
      RECT  34115.0 39480.0 34820.0 38135.0 ;
      RECT  34115.0 39480.0 34820.0 40825.0 ;
      RECT  34115.0 42170.0 34820.0 40825.0 ;
      RECT  34115.0 42170.0 34820.0 43515.0 ;
      RECT  34115.0 44860.0 34820.0 43515.0 ;
      RECT  34115.0 44860.0 34820.0 46205.0 ;
      RECT  34115.0 47550.0 34820.0 46205.0 ;
      RECT  34115.0 47550.0 34820.0 48895.0 ;
      RECT  34115.0 50240.0 34820.0 48895.0 ;
      RECT  34115.0 50240.0 34820.0 51585.0 ;
      RECT  34115.0 52930.0 34820.0 51585.0 ;
      RECT  34115.0 52930.0 34820.0 54275.0 ;
      RECT  34115.0 55620.0 34820.0 54275.0 ;
      RECT  34115.0 55620.0 34820.0 56965.0 ;
      RECT  34115.0 58310.0 34820.0 56965.0 ;
      RECT  34115.0 58310.0 34820.0 59655.0 ;
      RECT  34115.0 61000.0 34820.0 59655.0 ;
      RECT  34115.0 61000.0 34820.0 62345.0 ;
      RECT  34115.0 63690.0 34820.0 62345.0 ;
      RECT  34115.0 63690.0 34820.0 65035.0 ;
      RECT  34115.0 66380.0 34820.0 65035.0 ;
      RECT  34115.0 66380.0 34820.0 67725.0 ;
      RECT  34115.0 69070.0 34820.0 67725.0 ;
      RECT  34115.0 69070.0 34820.0 70415.0 ;
      RECT  34115.0 71760.0 34820.0 70415.0 ;
      RECT  34115.0 71760.0 34820.0 73105.0 ;
      RECT  34115.0 74450.0 34820.0 73105.0 ;
      RECT  34115.0 74450.0 34820.0 75795.0 ;
      RECT  34115.0 77140.0 34820.0 75795.0 ;
      RECT  34115.0 77140.0 34820.0 78485.0 ;
      RECT  34115.0 79830.0 34820.0 78485.0 ;
      RECT  34115.0 79830.0 34820.0 81175.0 ;
      RECT  34115.0 82520.0 34820.0 81175.0 ;
      RECT  34115.0 82520.0 34820.0 83865.0 ;
      RECT  34115.0 85210.0 34820.0 83865.0 ;
      RECT  34115.0 85210.0 34820.0 86555.0 ;
      RECT  34115.0 87900.0 34820.0 86555.0 ;
      RECT  34115.0 87900.0 34820.0 89245.0 ;
      RECT  34115.0 90590.0 34820.0 89245.0 ;
      RECT  34115.0 90590.0 34820.0 91935.0 ;
      RECT  34115.0 93280.0 34820.0 91935.0 ;
      RECT  34115.0 93280.0 34820.0 94625.0 ;
      RECT  34115.0 95970.0 34820.0 94625.0 ;
      RECT  34115.0 95970.0 34820.0 97315.0 ;
      RECT  34115.0 98660.0 34820.0 97315.0 ;
      RECT  34115.0 98660.0 34820.0 100005.0 ;
      RECT  34115.0 101350.0 34820.0 100005.0 ;
      RECT  34115.0 101350.0 34820.0 102695.0 ;
      RECT  34115.0 104040.0 34820.0 102695.0 ;
      RECT  34115.0 104040.0 34820.0 105385.0 ;
      RECT  34115.0 106730.0 34820.0 105385.0 ;
      RECT  34115.0 106730.0 34820.0 108075.0 ;
      RECT  34115.0 109420.0 34820.0 108075.0 ;
      RECT  34115.0 109420.0 34820.0 110765.0 ;
      RECT  34115.0 112110.0 34820.0 110765.0 ;
      RECT  34115.0 112110.0 34820.0 113455.0 ;
      RECT  34115.0 114800.0 34820.0 113455.0 ;
      RECT  34115.0 114800.0 34820.0 116145.0 ;
      RECT  34115.0 117490.0 34820.0 116145.0 ;
      RECT  34115.0 117490.0 34820.0 118835.0 ;
      RECT  34115.0 120180.0 34820.0 118835.0 ;
      RECT  34115.0 120180.0 34820.0 121525.0 ;
      RECT  34115.0 122870.0 34820.0 121525.0 ;
      RECT  34115.0 122870.0 34820.0 124215.0 ;
      RECT  34115.0 125560.0 34820.0 124215.0 ;
      RECT  34115.0 125560.0 34820.0 126905.0 ;
      RECT  34115.0 128250.0 34820.0 126905.0 ;
      RECT  34115.0 128250.0 34820.0 129595.0 ;
      RECT  34115.0 130940.0 34820.0 129595.0 ;
      RECT  34115.0 130940.0 34820.0 132285.0 ;
      RECT  34115.0 133630.0 34820.0 132285.0 ;
      RECT  34115.0 133630.0 34820.0 134975.0 ;
      RECT  34115.0 136320.0 34820.0 134975.0 ;
      RECT  34115.0 136320.0 34820.0 137665.0 ;
      RECT  34115.0 139010.0 34820.0 137665.0 ;
      RECT  34115.0 139010.0 34820.0 140355.0 ;
      RECT  34115.0 141700.0 34820.0 140355.0 ;
      RECT  34115.0 141700.0 34820.0 143045.0 ;
      RECT  34115.0 144390.0 34820.0 143045.0 ;
      RECT  34115.0 144390.0 34820.0 145735.0 ;
      RECT  34115.0 147080.0 34820.0 145735.0 ;
      RECT  34115.0 147080.0 34820.0 148425.0 ;
      RECT  34115.0 149770.0 34820.0 148425.0 ;
      RECT  34115.0 149770.0 34820.0 151115.0 ;
      RECT  34115.0 152460.0 34820.0 151115.0 ;
      RECT  34115.0 152460.0 34820.0 153805.0 ;
      RECT  34115.0 155150.0 34820.0 153805.0 ;
      RECT  34115.0 155150.0 34820.0 156495.0 ;
      RECT  34115.0 157840.0 34820.0 156495.0 ;
      RECT  34115.0 157840.0 34820.0 159185.0 ;
      RECT  34115.0 160530.0 34820.0 159185.0 ;
      RECT  34115.0 160530.0 34820.0 161875.0 ;
      RECT  34115.0 163220.0 34820.0 161875.0 ;
      RECT  34115.0 163220.0 34820.0 164565.0 ;
      RECT  34115.0 165910.0 34820.0 164565.0 ;
      RECT  34115.0 165910.0 34820.0 167255.0 ;
      RECT  34115.0 168600.0 34820.0 167255.0 ;
      RECT  34115.0 168600.0 34820.0 169945.0 ;
      RECT  34115.0 171290.0 34820.0 169945.0 ;
      RECT  34115.0 171290.0 34820.0 172635.0 ;
      RECT  34115.0 173980.0 34820.0 172635.0 ;
      RECT  34115.0 173980.0 34820.0 175325.0 ;
      RECT  34115.0 176670.0 34820.0 175325.0 ;
      RECT  34115.0 176670.0 34820.0 178015.0 ;
      RECT  34115.0 179360.0 34820.0 178015.0 ;
      RECT  34115.0 179360.0 34820.0 180705.0 ;
      RECT  34115.0 182050.0 34820.0 180705.0 ;
      RECT  34115.0 182050.0 34820.0 183395.0 ;
      RECT  34115.0 184740.0 34820.0 183395.0 ;
      RECT  34115.0 184740.0 34820.0 186085.0 ;
      RECT  34115.0 187430.0 34820.0 186085.0 ;
      RECT  34115.0 187430.0 34820.0 188775.0 ;
      RECT  34115.0 190120.0 34820.0 188775.0 ;
      RECT  34115.0 190120.0 34820.0 191465.0 ;
      RECT  34115.0 192810.0 34820.0 191465.0 ;
      RECT  34115.0 192810.0 34820.0 194155.0 ;
      RECT  34115.0 195500.0 34820.0 194155.0 ;
      RECT  34115.0 195500.0 34820.0 196845.0 ;
      RECT  34115.0 198190.0 34820.0 196845.0 ;
      RECT  34115.0 198190.0 34820.0 199535.0 ;
      RECT  34115.0 200880.0 34820.0 199535.0 ;
      RECT  34115.0 200880.0 34820.0 202225.0 ;
      RECT  34115.0 203570.0 34820.0 202225.0 ;
      RECT  34115.0 203570.0 34820.0 204915.0 ;
      RECT  34115.0 206260.0 34820.0 204915.0 ;
      RECT  34820.0 34100.0 35525.0 35445.0 ;
      RECT  34820.0 36790.0 35525.0 35445.0 ;
      RECT  34820.0 36790.0 35525.0 38135.0 ;
      RECT  34820.0 39480.0 35525.0 38135.0 ;
      RECT  34820.0 39480.0 35525.0 40825.0 ;
      RECT  34820.0 42170.0 35525.0 40825.0 ;
      RECT  34820.0 42170.0 35525.0 43515.0 ;
      RECT  34820.0 44860.0 35525.0 43515.0 ;
      RECT  34820.0 44860.0 35525.0 46205.0 ;
      RECT  34820.0 47550.0 35525.0 46205.0 ;
      RECT  34820.0 47550.0 35525.0 48895.0 ;
      RECT  34820.0 50240.0 35525.0 48895.0 ;
      RECT  34820.0 50240.0 35525.0 51585.0 ;
      RECT  34820.0 52930.0 35525.0 51585.0 ;
      RECT  34820.0 52930.0 35525.0 54275.0 ;
      RECT  34820.0 55620.0 35525.0 54275.0 ;
      RECT  34820.0 55620.0 35525.0 56965.0 ;
      RECT  34820.0 58310.0 35525.0 56965.0 ;
      RECT  34820.0 58310.0 35525.0 59655.0 ;
      RECT  34820.0 61000.0 35525.0 59655.0 ;
      RECT  34820.0 61000.0 35525.0 62345.0 ;
      RECT  34820.0 63690.0 35525.0 62345.0 ;
      RECT  34820.0 63690.0 35525.0 65035.0 ;
      RECT  34820.0 66380.0 35525.0 65035.0 ;
      RECT  34820.0 66380.0 35525.0 67725.0 ;
      RECT  34820.0 69070.0 35525.0 67725.0 ;
      RECT  34820.0 69070.0 35525.0 70415.0 ;
      RECT  34820.0 71760.0 35525.0 70415.0 ;
      RECT  34820.0 71760.0 35525.0 73105.0 ;
      RECT  34820.0 74450.0 35525.0 73105.0 ;
      RECT  34820.0 74450.0 35525.0 75795.0 ;
      RECT  34820.0 77140.0 35525.0 75795.0 ;
      RECT  34820.0 77140.0 35525.0 78485.0 ;
      RECT  34820.0 79830.0 35525.0 78485.0 ;
      RECT  34820.0 79830.0 35525.0 81175.0 ;
      RECT  34820.0 82520.0 35525.0 81175.0 ;
      RECT  34820.0 82520.0 35525.0 83865.0 ;
      RECT  34820.0 85210.0 35525.0 83865.0 ;
      RECT  34820.0 85210.0 35525.0 86555.0 ;
      RECT  34820.0 87900.0 35525.0 86555.0 ;
      RECT  34820.0 87900.0 35525.0 89245.0 ;
      RECT  34820.0 90590.0 35525.0 89245.0 ;
      RECT  34820.0 90590.0 35525.0 91935.0 ;
      RECT  34820.0 93280.0 35525.0 91935.0 ;
      RECT  34820.0 93280.0 35525.0 94625.0 ;
      RECT  34820.0 95970.0 35525.0 94625.0 ;
      RECT  34820.0 95970.0 35525.0 97315.0 ;
      RECT  34820.0 98660.0 35525.0 97315.0 ;
      RECT  34820.0 98660.0 35525.0 100005.0 ;
      RECT  34820.0 101350.0 35525.0 100005.0 ;
      RECT  34820.0 101350.0 35525.0 102695.0 ;
      RECT  34820.0 104040.0 35525.0 102695.0 ;
      RECT  34820.0 104040.0 35525.0 105385.0 ;
      RECT  34820.0 106730.0 35525.0 105385.0 ;
      RECT  34820.0 106730.0 35525.0 108075.0 ;
      RECT  34820.0 109420.0 35525.0 108075.0 ;
      RECT  34820.0 109420.0 35525.0 110765.0 ;
      RECT  34820.0 112110.0 35525.0 110765.0 ;
      RECT  34820.0 112110.0 35525.0 113455.0 ;
      RECT  34820.0 114800.0 35525.0 113455.0 ;
      RECT  34820.0 114800.0 35525.0 116145.0 ;
      RECT  34820.0 117490.0 35525.0 116145.0 ;
      RECT  34820.0 117490.0 35525.0 118835.0 ;
      RECT  34820.0 120180.0 35525.0 118835.0 ;
      RECT  34820.0 120180.0 35525.0 121525.0 ;
      RECT  34820.0 122870.0 35525.0 121525.0 ;
      RECT  34820.0 122870.0 35525.0 124215.0 ;
      RECT  34820.0 125560.0 35525.0 124215.0 ;
      RECT  34820.0 125560.0 35525.0 126905.0 ;
      RECT  34820.0 128250.0 35525.0 126905.0 ;
      RECT  34820.0 128250.0 35525.0 129595.0 ;
      RECT  34820.0 130940.0 35525.0 129595.0 ;
      RECT  34820.0 130940.0 35525.0 132285.0 ;
      RECT  34820.0 133630.0 35525.0 132285.0 ;
      RECT  34820.0 133630.0 35525.0 134975.0 ;
      RECT  34820.0 136320.0 35525.0 134975.0 ;
      RECT  34820.0 136320.0 35525.0 137665.0 ;
      RECT  34820.0 139010.0 35525.0 137665.0 ;
      RECT  34820.0 139010.0 35525.0 140355.0 ;
      RECT  34820.0 141700.0 35525.0 140355.0 ;
      RECT  34820.0 141700.0 35525.0 143045.0 ;
      RECT  34820.0 144390.0 35525.0 143045.0 ;
      RECT  34820.0 144390.0 35525.0 145735.0 ;
      RECT  34820.0 147080.0 35525.0 145735.0 ;
      RECT  34820.0 147080.0 35525.0 148425.0 ;
      RECT  34820.0 149770.0 35525.0 148425.0 ;
      RECT  34820.0 149770.0 35525.0 151115.0 ;
      RECT  34820.0 152460.0 35525.0 151115.0 ;
      RECT  34820.0 152460.0 35525.0 153805.0 ;
      RECT  34820.0 155150.0 35525.0 153805.0 ;
      RECT  34820.0 155150.0 35525.0 156495.0 ;
      RECT  34820.0 157840.0 35525.0 156495.0 ;
      RECT  34820.0 157840.0 35525.0 159185.0 ;
      RECT  34820.0 160530.0 35525.0 159185.0 ;
      RECT  34820.0 160530.0 35525.0 161875.0 ;
      RECT  34820.0 163220.0 35525.0 161875.0 ;
      RECT  34820.0 163220.0 35525.0 164565.0 ;
      RECT  34820.0 165910.0 35525.0 164565.0 ;
      RECT  34820.0 165910.0 35525.0 167255.0 ;
      RECT  34820.0 168600.0 35525.0 167255.0 ;
      RECT  34820.0 168600.0 35525.0 169945.0 ;
      RECT  34820.0 171290.0 35525.0 169945.0 ;
      RECT  34820.0 171290.0 35525.0 172635.0 ;
      RECT  34820.0 173980.0 35525.0 172635.0 ;
      RECT  34820.0 173980.0 35525.0 175325.0 ;
      RECT  34820.0 176670.0 35525.0 175325.0 ;
      RECT  34820.0 176670.0 35525.0 178015.0 ;
      RECT  34820.0 179360.0 35525.0 178015.0 ;
      RECT  34820.0 179360.0 35525.0 180705.0 ;
      RECT  34820.0 182050.0 35525.0 180705.0 ;
      RECT  34820.0 182050.0 35525.0 183395.0 ;
      RECT  34820.0 184740.0 35525.0 183395.0 ;
      RECT  34820.0 184740.0 35525.0 186085.0 ;
      RECT  34820.0 187430.0 35525.0 186085.0 ;
      RECT  34820.0 187430.0 35525.0 188775.0 ;
      RECT  34820.0 190120.0 35525.0 188775.0 ;
      RECT  34820.0 190120.0 35525.0 191465.0 ;
      RECT  34820.0 192810.0 35525.0 191465.0 ;
      RECT  34820.0 192810.0 35525.0 194155.0 ;
      RECT  34820.0 195500.0 35525.0 194155.0 ;
      RECT  34820.0 195500.0 35525.0 196845.0 ;
      RECT  34820.0 198190.0 35525.0 196845.0 ;
      RECT  34820.0 198190.0 35525.0 199535.0 ;
      RECT  34820.0 200880.0 35525.0 199535.0 ;
      RECT  34820.0 200880.0 35525.0 202225.0 ;
      RECT  34820.0 203570.0 35525.0 202225.0 ;
      RECT  34820.0 203570.0 35525.0 204915.0 ;
      RECT  34820.0 206260.0 35525.0 204915.0 ;
      RECT  35525.0 34100.0 36230.0 35445.0 ;
      RECT  35525.0 36790.0 36230.0 35445.0 ;
      RECT  35525.0 36790.0 36230.0 38135.0 ;
      RECT  35525.0 39480.0 36230.0 38135.0 ;
      RECT  35525.0 39480.0 36230.0 40825.0 ;
      RECT  35525.0 42170.0 36230.0 40825.0 ;
      RECT  35525.0 42170.0 36230.0 43515.0 ;
      RECT  35525.0 44860.0 36230.0 43515.0 ;
      RECT  35525.0 44860.0 36230.0 46205.0 ;
      RECT  35525.0 47550.0 36230.0 46205.0 ;
      RECT  35525.0 47550.0 36230.0 48895.0 ;
      RECT  35525.0 50240.0 36230.0 48895.0 ;
      RECT  35525.0 50240.0 36230.0 51585.0 ;
      RECT  35525.0 52930.0 36230.0 51585.0 ;
      RECT  35525.0 52930.0 36230.0 54275.0 ;
      RECT  35525.0 55620.0 36230.0 54275.0 ;
      RECT  35525.0 55620.0 36230.0 56965.0 ;
      RECT  35525.0 58310.0 36230.0 56965.0 ;
      RECT  35525.0 58310.0 36230.0 59655.0 ;
      RECT  35525.0 61000.0 36230.0 59655.0 ;
      RECT  35525.0 61000.0 36230.0 62345.0 ;
      RECT  35525.0 63690.0 36230.0 62345.0 ;
      RECT  35525.0 63690.0 36230.0 65035.0 ;
      RECT  35525.0 66380.0 36230.0 65035.0 ;
      RECT  35525.0 66380.0 36230.0 67725.0 ;
      RECT  35525.0 69070.0 36230.0 67725.0 ;
      RECT  35525.0 69070.0 36230.0 70415.0 ;
      RECT  35525.0 71760.0 36230.0 70415.0 ;
      RECT  35525.0 71760.0 36230.0 73105.0 ;
      RECT  35525.0 74450.0 36230.0 73105.0 ;
      RECT  35525.0 74450.0 36230.0 75795.0 ;
      RECT  35525.0 77140.0 36230.0 75795.0 ;
      RECT  35525.0 77140.0 36230.0 78485.0 ;
      RECT  35525.0 79830.0 36230.0 78485.0 ;
      RECT  35525.0 79830.0 36230.0 81175.0 ;
      RECT  35525.0 82520.0 36230.0 81175.0 ;
      RECT  35525.0 82520.0 36230.0 83865.0 ;
      RECT  35525.0 85210.0 36230.0 83865.0 ;
      RECT  35525.0 85210.0 36230.0 86555.0 ;
      RECT  35525.0 87900.0 36230.0 86555.0 ;
      RECT  35525.0 87900.0 36230.0 89245.0 ;
      RECT  35525.0 90590.0 36230.0 89245.0 ;
      RECT  35525.0 90590.0 36230.0 91935.0 ;
      RECT  35525.0 93280.0 36230.0 91935.0 ;
      RECT  35525.0 93280.0 36230.0 94625.0 ;
      RECT  35525.0 95970.0 36230.0 94625.0 ;
      RECT  35525.0 95970.0 36230.0 97315.0 ;
      RECT  35525.0 98660.0 36230.0 97315.0 ;
      RECT  35525.0 98660.0 36230.0 100005.0 ;
      RECT  35525.0 101350.0 36230.0 100005.0 ;
      RECT  35525.0 101350.0 36230.0 102695.0 ;
      RECT  35525.0 104040.0 36230.0 102695.0 ;
      RECT  35525.0 104040.0 36230.0 105385.0 ;
      RECT  35525.0 106730.0 36230.0 105385.0 ;
      RECT  35525.0 106730.0 36230.0 108075.0 ;
      RECT  35525.0 109420.0 36230.0 108075.0 ;
      RECT  35525.0 109420.0 36230.0 110765.0 ;
      RECT  35525.0 112110.0 36230.0 110765.0 ;
      RECT  35525.0 112110.0 36230.0 113455.0 ;
      RECT  35525.0 114800.0 36230.0 113455.0 ;
      RECT  35525.0 114800.0 36230.0 116145.0 ;
      RECT  35525.0 117490.0 36230.0 116145.0 ;
      RECT  35525.0 117490.0 36230.0 118835.0 ;
      RECT  35525.0 120180.0 36230.0 118835.0 ;
      RECT  35525.0 120180.0 36230.0 121525.0 ;
      RECT  35525.0 122870.0 36230.0 121525.0 ;
      RECT  35525.0 122870.0 36230.0 124215.0 ;
      RECT  35525.0 125560.0 36230.0 124215.0 ;
      RECT  35525.0 125560.0 36230.0 126905.0 ;
      RECT  35525.0 128250.0 36230.0 126905.0 ;
      RECT  35525.0 128250.0 36230.0 129595.0 ;
      RECT  35525.0 130940.0 36230.0 129595.0 ;
      RECT  35525.0 130940.0 36230.0 132285.0 ;
      RECT  35525.0 133630.0 36230.0 132285.0 ;
      RECT  35525.0 133630.0 36230.0 134975.0 ;
      RECT  35525.0 136320.0 36230.0 134975.0 ;
      RECT  35525.0 136320.0 36230.0 137665.0 ;
      RECT  35525.0 139010.0 36230.0 137665.0 ;
      RECT  35525.0 139010.0 36230.0 140355.0 ;
      RECT  35525.0 141700.0 36230.0 140355.0 ;
      RECT  35525.0 141700.0 36230.0 143045.0 ;
      RECT  35525.0 144390.0 36230.0 143045.0 ;
      RECT  35525.0 144390.0 36230.0 145735.0 ;
      RECT  35525.0 147080.0 36230.0 145735.0 ;
      RECT  35525.0 147080.0 36230.0 148425.0 ;
      RECT  35525.0 149770.0 36230.0 148425.0 ;
      RECT  35525.0 149770.0 36230.0 151115.0 ;
      RECT  35525.0 152460.0 36230.0 151115.0 ;
      RECT  35525.0 152460.0 36230.0 153805.0 ;
      RECT  35525.0 155150.0 36230.0 153805.0 ;
      RECT  35525.0 155150.0 36230.0 156495.0 ;
      RECT  35525.0 157840.0 36230.0 156495.0 ;
      RECT  35525.0 157840.0 36230.0 159185.0 ;
      RECT  35525.0 160530.0 36230.0 159185.0 ;
      RECT  35525.0 160530.0 36230.0 161875.0 ;
      RECT  35525.0 163220.0 36230.0 161875.0 ;
      RECT  35525.0 163220.0 36230.0 164565.0 ;
      RECT  35525.0 165910.0 36230.0 164565.0 ;
      RECT  35525.0 165910.0 36230.0 167255.0 ;
      RECT  35525.0 168600.0 36230.0 167255.0 ;
      RECT  35525.0 168600.0 36230.0 169945.0 ;
      RECT  35525.0 171290.0 36230.0 169945.0 ;
      RECT  35525.0 171290.0 36230.0 172635.0 ;
      RECT  35525.0 173980.0 36230.0 172635.0 ;
      RECT  35525.0 173980.0 36230.0 175325.0 ;
      RECT  35525.0 176670.0 36230.0 175325.0 ;
      RECT  35525.0 176670.0 36230.0 178015.0 ;
      RECT  35525.0 179360.0 36230.0 178015.0 ;
      RECT  35525.0 179360.0 36230.0 180705.0 ;
      RECT  35525.0 182050.0 36230.0 180705.0 ;
      RECT  35525.0 182050.0 36230.0 183395.0 ;
      RECT  35525.0 184740.0 36230.0 183395.0 ;
      RECT  35525.0 184740.0 36230.0 186085.0 ;
      RECT  35525.0 187430.0 36230.0 186085.0 ;
      RECT  35525.0 187430.0 36230.0 188775.0 ;
      RECT  35525.0 190120.0 36230.0 188775.0 ;
      RECT  35525.0 190120.0 36230.0 191465.0 ;
      RECT  35525.0 192810.0 36230.0 191465.0 ;
      RECT  35525.0 192810.0 36230.0 194155.0 ;
      RECT  35525.0 195500.0 36230.0 194155.0 ;
      RECT  35525.0 195500.0 36230.0 196845.0 ;
      RECT  35525.0 198190.0 36230.0 196845.0 ;
      RECT  35525.0 198190.0 36230.0 199535.0 ;
      RECT  35525.0 200880.0 36230.0 199535.0 ;
      RECT  35525.0 200880.0 36230.0 202225.0 ;
      RECT  35525.0 203570.0 36230.0 202225.0 ;
      RECT  35525.0 203570.0 36230.0 204915.0 ;
      RECT  35525.0 206260.0 36230.0 204915.0 ;
      RECT  36230.0 34100.0 36935.0 35445.0 ;
      RECT  36230.0 36790.0 36935.0 35445.0 ;
      RECT  36230.0 36790.0 36935.0 38135.0 ;
      RECT  36230.0 39480.0 36935.0 38135.0 ;
      RECT  36230.0 39480.0 36935.0 40825.0 ;
      RECT  36230.0 42170.0 36935.0 40825.0 ;
      RECT  36230.0 42170.0 36935.0 43515.0 ;
      RECT  36230.0 44860.0 36935.0 43515.0 ;
      RECT  36230.0 44860.0 36935.0 46205.0 ;
      RECT  36230.0 47550.0 36935.0 46205.0 ;
      RECT  36230.0 47550.0 36935.0 48895.0 ;
      RECT  36230.0 50240.0 36935.0 48895.0 ;
      RECT  36230.0 50240.0 36935.0 51585.0 ;
      RECT  36230.0 52930.0 36935.0 51585.0 ;
      RECT  36230.0 52930.0 36935.0 54275.0 ;
      RECT  36230.0 55620.0 36935.0 54275.0 ;
      RECT  36230.0 55620.0 36935.0 56965.0 ;
      RECT  36230.0 58310.0 36935.0 56965.0 ;
      RECT  36230.0 58310.0 36935.0 59655.0 ;
      RECT  36230.0 61000.0 36935.0 59655.0 ;
      RECT  36230.0 61000.0 36935.0 62345.0 ;
      RECT  36230.0 63690.0 36935.0 62345.0 ;
      RECT  36230.0 63690.0 36935.0 65035.0 ;
      RECT  36230.0 66380.0 36935.0 65035.0 ;
      RECT  36230.0 66380.0 36935.0 67725.0 ;
      RECT  36230.0 69070.0 36935.0 67725.0 ;
      RECT  36230.0 69070.0 36935.0 70415.0 ;
      RECT  36230.0 71760.0 36935.0 70415.0 ;
      RECT  36230.0 71760.0 36935.0 73105.0 ;
      RECT  36230.0 74450.0 36935.0 73105.0 ;
      RECT  36230.0 74450.0 36935.0 75795.0 ;
      RECT  36230.0 77140.0 36935.0 75795.0 ;
      RECT  36230.0 77140.0 36935.0 78485.0 ;
      RECT  36230.0 79830.0 36935.0 78485.0 ;
      RECT  36230.0 79830.0 36935.0 81175.0 ;
      RECT  36230.0 82520.0 36935.0 81175.0 ;
      RECT  36230.0 82520.0 36935.0 83865.0 ;
      RECT  36230.0 85210.0 36935.0 83865.0 ;
      RECT  36230.0 85210.0 36935.0 86555.0 ;
      RECT  36230.0 87900.0 36935.0 86555.0 ;
      RECT  36230.0 87900.0 36935.0 89245.0 ;
      RECT  36230.0 90590.0 36935.0 89245.0 ;
      RECT  36230.0 90590.0 36935.0 91935.0 ;
      RECT  36230.0 93280.0 36935.0 91935.0 ;
      RECT  36230.0 93280.0 36935.0 94625.0 ;
      RECT  36230.0 95970.0 36935.0 94625.0 ;
      RECT  36230.0 95970.0 36935.0 97315.0 ;
      RECT  36230.0 98660.0 36935.0 97315.0 ;
      RECT  36230.0 98660.0 36935.0 100005.0 ;
      RECT  36230.0 101350.0 36935.0 100005.0 ;
      RECT  36230.0 101350.0 36935.0 102695.0 ;
      RECT  36230.0 104040.0 36935.0 102695.0 ;
      RECT  36230.0 104040.0 36935.0 105385.0 ;
      RECT  36230.0 106730.0 36935.0 105385.0 ;
      RECT  36230.0 106730.0 36935.0 108075.0 ;
      RECT  36230.0 109420.0 36935.0 108075.0 ;
      RECT  36230.0 109420.0 36935.0 110765.0 ;
      RECT  36230.0 112110.0 36935.0 110765.0 ;
      RECT  36230.0 112110.0 36935.0 113455.0 ;
      RECT  36230.0 114800.0 36935.0 113455.0 ;
      RECT  36230.0 114800.0 36935.0 116145.0 ;
      RECT  36230.0 117490.0 36935.0 116145.0 ;
      RECT  36230.0 117490.0 36935.0 118835.0 ;
      RECT  36230.0 120180.0 36935.0 118835.0 ;
      RECT  36230.0 120180.0 36935.0 121525.0 ;
      RECT  36230.0 122870.0 36935.0 121525.0 ;
      RECT  36230.0 122870.0 36935.0 124215.0 ;
      RECT  36230.0 125560.0 36935.0 124215.0 ;
      RECT  36230.0 125560.0 36935.0 126905.0 ;
      RECT  36230.0 128250.0 36935.0 126905.0 ;
      RECT  36230.0 128250.0 36935.0 129595.0 ;
      RECT  36230.0 130940.0 36935.0 129595.0 ;
      RECT  36230.0 130940.0 36935.0 132285.0 ;
      RECT  36230.0 133630.0 36935.0 132285.0 ;
      RECT  36230.0 133630.0 36935.0 134975.0 ;
      RECT  36230.0 136320.0 36935.0 134975.0 ;
      RECT  36230.0 136320.0 36935.0 137665.0 ;
      RECT  36230.0 139010.0 36935.0 137665.0 ;
      RECT  36230.0 139010.0 36935.0 140355.0 ;
      RECT  36230.0 141700.0 36935.0 140355.0 ;
      RECT  36230.0 141700.0 36935.0 143045.0 ;
      RECT  36230.0 144390.0 36935.0 143045.0 ;
      RECT  36230.0 144390.0 36935.0 145735.0 ;
      RECT  36230.0 147080.0 36935.0 145735.0 ;
      RECT  36230.0 147080.0 36935.0 148425.0 ;
      RECT  36230.0 149770.0 36935.0 148425.0 ;
      RECT  36230.0 149770.0 36935.0 151115.0 ;
      RECT  36230.0 152460.0 36935.0 151115.0 ;
      RECT  36230.0 152460.0 36935.0 153805.0 ;
      RECT  36230.0 155150.0 36935.0 153805.0 ;
      RECT  36230.0 155150.0 36935.0 156495.0 ;
      RECT  36230.0 157840.0 36935.0 156495.0 ;
      RECT  36230.0 157840.0 36935.0 159185.0 ;
      RECT  36230.0 160530.0 36935.0 159185.0 ;
      RECT  36230.0 160530.0 36935.0 161875.0 ;
      RECT  36230.0 163220.0 36935.0 161875.0 ;
      RECT  36230.0 163220.0 36935.0 164565.0 ;
      RECT  36230.0 165910.0 36935.0 164565.0 ;
      RECT  36230.0 165910.0 36935.0 167255.0 ;
      RECT  36230.0 168600.0 36935.0 167255.0 ;
      RECT  36230.0 168600.0 36935.0 169945.0 ;
      RECT  36230.0 171290.0 36935.0 169945.0 ;
      RECT  36230.0 171290.0 36935.0 172635.0 ;
      RECT  36230.0 173980.0 36935.0 172635.0 ;
      RECT  36230.0 173980.0 36935.0 175325.0 ;
      RECT  36230.0 176670.0 36935.0 175325.0 ;
      RECT  36230.0 176670.0 36935.0 178015.0 ;
      RECT  36230.0 179360.0 36935.0 178015.0 ;
      RECT  36230.0 179360.0 36935.0 180705.0 ;
      RECT  36230.0 182050.0 36935.0 180705.0 ;
      RECT  36230.0 182050.0 36935.0 183395.0 ;
      RECT  36230.0 184740.0 36935.0 183395.0 ;
      RECT  36230.0 184740.0 36935.0 186085.0 ;
      RECT  36230.0 187430.0 36935.0 186085.0 ;
      RECT  36230.0 187430.0 36935.0 188775.0 ;
      RECT  36230.0 190120.0 36935.0 188775.0 ;
      RECT  36230.0 190120.0 36935.0 191465.0 ;
      RECT  36230.0 192810.0 36935.0 191465.0 ;
      RECT  36230.0 192810.0 36935.0 194155.0 ;
      RECT  36230.0 195500.0 36935.0 194155.0 ;
      RECT  36230.0 195500.0 36935.0 196845.0 ;
      RECT  36230.0 198190.0 36935.0 196845.0 ;
      RECT  36230.0 198190.0 36935.0 199535.0 ;
      RECT  36230.0 200880.0 36935.0 199535.0 ;
      RECT  36230.0 200880.0 36935.0 202225.0 ;
      RECT  36230.0 203570.0 36935.0 202225.0 ;
      RECT  36230.0 203570.0 36935.0 204915.0 ;
      RECT  36230.0 206260.0 36935.0 204915.0 ;
      RECT  36935.0 34100.0 37640.0 35445.0 ;
      RECT  36935.0 36790.0 37640.0 35445.0 ;
      RECT  36935.0 36790.0 37640.0 38135.0 ;
      RECT  36935.0 39480.0 37640.0 38135.0 ;
      RECT  36935.0 39480.0 37640.0 40825.0 ;
      RECT  36935.0 42170.0 37640.0 40825.0 ;
      RECT  36935.0 42170.0 37640.0 43515.0 ;
      RECT  36935.0 44860.0 37640.0 43515.0 ;
      RECT  36935.0 44860.0 37640.0 46205.0 ;
      RECT  36935.0 47550.0 37640.0 46205.0 ;
      RECT  36935.0 47550.0 37640.0 48895.0 ;
      RECT  36935.0 50240.0 37640.0 48895.0 ;
      RECT  36935.0 50240.0 37640.0 51585.0 ;
      RECT  36935.0 52930.0 37640.0 51585.0 ;
      RECT  36935.0 52930.0 37640.0 54275.0 ;
      RECT  36935.0 55620.0 37640.0 54275.0 ;
      RECT  36935.0 55620.0 37640.0 56965.0 ;
      RECT  36935.0 58310.0 37640.0 56965.0 ;
      RECT  36935.0 58310.0 37640.0 59655.0 ;
      RECT  36935.0 61000.0 37640.0 59655.0 ;
      RECT  36935.0 61000.0 37640.0 62345.0 ;
      RECT  36935.0 63690.0 37640.0 62345.0 ;
      RECT  36935.0 63690.0 37640.0 65035.0 ;
      RECT  36935.0 66380.0 37640.0 65035.0 ;
      RECT  36935.0 66380.0 37640.0 67725.0 ;
      RECT  36935.0 69070.0 37640.0 67725.0 ;
      RECT  36935.0 69070.0 37640.0 70415.0 ;
      RECT  36935.0 71760.0 37640.0 70415.0 ;
      RECT  36935.0 71760.0 37640.0 73105.0 ;
      RECT  36935.0 74450.0 37640.0 73105.0 ;
      RECT  36935.0 74450.0 37640.0 75795.0 ;
      RECT  36935.0 77140.0 37640.0 75795.0 ;
      RECT  36935.0 77140.0 37640.0 78485.0 ;
      RECT  36935.0 79830.0 37640.0 78485.0 ;
      RECT  36935.0 79830.0 37640.0 81175.0 ;
      RECT  36935.0 82520.0 37640.0 81175.0 ;
      RECT  36935.0 82520.0 37640.0 83865.0 ;
      RECT  36935.0 85210.0 37640.0 83865.0 ;
      RECT  36935.0 85210.0 37640.0 86555.0 ;
      RECT  36935.0 87900.0 37640.0 86555.0 ;
      RECT  36935.0 87900.0 37640.0 89245.0 ;
      RECT  36935.0 90590.0 37640.0 89245.0 ;
      RECT  36935.0 90590.0 37640.0 91935.0 ;
      RECT  36935.0 93280.0 37640.0 91935.0 ;
      RECT  36935.0 93280.0 37640.0 94625.0 ;
      RECT  36935.0 95970.0 37640.0 94625.0 ;
      RECT  36935.0 95970.0 37640.0 97315.0 ;
      RECT  36935.0 98660.0 37640.0 97315.0 ;
      RECT  36935.0 98660.0 37640.0 100005.0 ;
      RECT  36935.0 101350.0 37640.0 100005.0 ;
      RECT  36935.0 101350.0 37640.0 102695.0 ;
      RECT  36935.0 104040.0 37640.0 102695.0 ;
      RECT  36935.0 104040.0 37640.0 105385.0 ;
      RECT  36935.0 106730.0 37640.0 105385.0 ;
      RECT  36935.0 106730.0 37640.0 108075.0 ;
      RECT  36935.0 109420.0 37640.0 108075.0 ;
      RECT  36935.0 109420.0 37640.0 110765.0 ;
      RECT  36935.0 112110.0 37640.0 110765.0 ;
      RECT  36935.0 112110.0 37640.0 113455.0 ;
      RECT  36935.0 114800.0 37640.0 113455.0 ;
      RECT  36935.0 114800.0 37640.0 116145.0 ;
      RECT  36935.0 117490.0 37640.0 116145.0 ;
      RECT  36935.0 117490.0 37640.0 118835.0 ;
      RECT  36935.0 120180.0 37640.0 118835.0 ;
      RECT  36935.0 120180.0 37640.0 121525.0 ;
      RECT  36935.0 122870.0 37640.0 121525.0 ;
      RECT  36935.0 122870.0 37640.0 124215.0 ;
      RECT  36935.0 125560.0 37640.0 124215.0 ;
      RECT  36935.0 125560.0 37640.0 126905.0 ;
      RECT  36935.0 128250.0 37640.0 126905.0 ;
      RECT  36935.0 128250.0 37640.0 129595.0 ;
      RECT  36935.0 130940.0 37640.0 129595.0 ;
      RECT  36935.0 130940.0 37640.0 132285.0 ;
      RECT  36935.0 133630.0 37640.0 132285.0 ;
      RECT  36935.0 133630.0 37640.0 134975.0 ;
      RECT  36935.0 136320.0 37640.0 134975.0 ;
      RECT  36935.0 136320.0 37640.0 137665.0 ;
      RECT  36935.0 139010.0 37640.0 137665.0 ;
      RECT  36935.0 139010.0 37640.0 140355.0 ;
      RECT  36935.0 141700.0 37640.0 140355.0 ;
      RECT  36935.0 141700.0 37640.0 143045.0 ;
      RECT  36935.0 144390.0 37640.0 143045.0 ;
      RECT  36935.0 144390.0 37640.0 145735.0 ;
      RECT  36935.0 147080.0 37640.0 145735.0 ;
      RECT  36935.0 147080.0 37640.0 148425.0 ;
      RECT  36935.0 149770.0 37640.0 148425.0 ;
      RECT  36935.0 149770.0 37640.0 151115.0 ;
      RECT  36935.0 152460.0 37640.0 151115.0 ;
      RECT  36935.0 152460.0 37640.0 153805.0 ;
      RECT  36935.0 155150.0 37640.0 153805.0 ;
      RECT  36935.0 155150.0 37640.0 156495.0 ;
      RECT  36935.0 157840.0 37640.0 156495.0 ;
      RECT  36935.0 157840.0 37640.0 159185.0 ;
      RECT  36935.0 160530.0 37640.0 159185.0 ;
      RECT  36935.0 160530.0 37640.0 161875.0 ;
      RECT  36935.0 163220.0 37640.0 161875.0 ;
      RECT  36935.0 163220.0 37640.0 164565.0 ;
      RECT  36935.0 165910.0 37640.0 164565.0 ;
      RECT  36935.0 165910.0 37640.0 167255.0 ;
      RECT  36935.0 168600.0 37640.0 167255.0 ;
      RECT  36935.0 168600.0 37640.0 169945.0 ;
      RECT  36935.0 171290.0 37640.0 169945.0 ;
      RECT  36935.0 171290.0 37640.0 172635.0 ;
      RECT  36935.0 173980.0 37640.0 172635.0 ;
      RECT  36935.0 173980.0 37640.0 175325.0 ;
      RECT  36935.0 176670.0 37640.0 175325.0 ;
      RECT  36935.0 176670.0 37640.0 178015.0 ;
      RECT  36935.0 179360.0 37640.0 178015.0 ;
      RECT  36935.0 179360.0 37640.0 180705.0 ;
      RECT  36935.0 182050.0 37640.0 180705.0 ;
      RECT  36935.0 182050.0 37640.0 183395.0 ;
      RECT  36935.0 184740.0 37640.0 183395.0 ;
      RECT  36935.0 184740.0 37640.0 186085.0 ;
      RECT  36935.0 187430.0 37640.0 186085.0 ;
      RECT  36935.0 187430.0 37640.0 188775.0 ;
      RECT  36935.0 190120.0 37640.0 188775.0 ;
      RECT  36935.0 190120.0 37640.0 191465.0 ;
      RECT  36935.0 192810.0 37640.0 191465.0 ;
      RECT  36935.0 192810.0 37640.0 194155.0 ;
      RECT  36935.0 195500.0 37640.0 194155.0 ;
      RECT  36935.0 195500.0 37640.0 196845.0 ;
      RECT  36935.0 198190.0 37640.0 196845.0 ;
      RECT  36935.0 198190.0 37640.0 199535.0 ;
      RECT  36935.0 200880.0 37640.0 199535.0 ;
      RECT  36935.0 200880.0 37640.0 202225.0 ;
      RECT  36935.0 203570.0 37640.0 202225.0 ;
      RECT  36935.0 203570.0 37640.0 204915.0 ;
      RECT  36935.0 206260.0 37640.0 204915.0 ;
      RECT  37640.0 34100.0 38345.0 35445.0 ;
      RECT  37640.0 36790.0 38345.0 35445.0 ;
      RECT  37640.0 36790.0 38345.0 38135.0 ;
      RECT  37640.0 39480.0 38345.0 38135.0 ;
      RECT  37640.0 39480.0 38345.0 40825.0 ;
      RECT  37640.0 42170.0 38345.0 40825.0 ;
      RECT  37640.0 42170.0 38345.0 43515.0 ;
      RECT  37640.0 44860.0 38345.0 43515.0 ;
      RECT  37640.0 44860.0 38345.0 46205.0 ;
      RECT  37640.0 47550.0 38345.0 46205.0 ;
      RECT  37640.0 47550.0 38345.0 48895.0 ;
      RECT  37640.0 50240.0 38345.0 48895.0 ;
      RECT  37640.0 50240.0 38345.0 51585.0 ;
      RECT  37640.0 52930.0 38345.0 51585.0 ;
      RECT  37640.0 52930.0 38345.0 54275.0 ;
      RECT  37640.0 55620.0 38345.0 54275.0 ;
      RECT  37640.0 55620.0 38345.0 56965.0 ;
      RECT  37640.0 58310.0 38345.0 56965.0 ;
      RECT  37640.0 58310.0 38345.0 59655.0 ;
      RECT  37640.0 61000.0 38345.0 59655.0 ;
      RECT  37640.0 61000.0 38345.0 62345.0 ;
      RECT  37640.0 63690.0 38345.0 62345.0 ;
      RECT  37640.0 63690.0 38345.0 65035.0 ;
      RECT  37640.0 66380.0 38345.0 65035.0 ;
      RECT  37640.0 66380.0 38345.0 67725.0 ;
      RECT  37640.0 69070.0 38345.0 67725.0 ;
      RECT  37640.0 69070.0 38345.0 70415.0 ;
      RECT  37640.0 71760.0 38345.0 70415.0 ;
      RECT  37640.0 71760.0 38345.0 73105.0 ;
      RECT  37640.0 74450.0 38345.0 73105.0 ;
      RECT  37640.0 74450.0 38345.0 75795.0 ;
      RECT  37640.0 77140.0 38345.0 75795.0 ;
      RECT  37640.0 77140.0 38345.0 78485.0 ;
      RECT  37640.0 79830.0 38345.0 78485.0 ;
      RECT  37640.0 79830.0 38345.0 81175.0 ;
      RECT  37640.0 82520.0 38345.0 81175.0 ;
      RECT  37640.0 82520.0 38345.0 83865.0 ;
      RECT  37640.0 85210.0 38345.0 83865.0 ;
      RECT  37640.0 85210.0 38345.0 86555.0 ;
      RECT  37640.0 87900.0 38345.0 86555.0 ;
      RECT  37640.0 87900.0 38345.0 89245.0 ;
      RECT  37640.0 90590.0 38345.0 89245.0 ;
      RECT  37640.0 90590.0 38345.0 91935.0 ;
      RECT  37640.0 93280.0 38345.0 91935.0 ;
      RECT  37640.0 93280.0 38345.0 94625.0 ;
      RECT  37640.0 95970.0 38345.0 94625.0 ;
      RECT  37640.0 95970.0 38345.0 97315.0 ;
      RECT  37640.0 98660.0 38345.0 97315.0 ;
      RECT  37640.0 98660.0 38345.0 100005.0 ;
      RECT  37640.0 101350.0 38345.0 100005.0 ;
      RECT  37640.0 101350.0 38345.0 102695.0 ;
      RECT  37640.0 104040.0 38345.0 102695.0 ;
      RECT  37640.0 104040.0 38345.0 105385.0 ;
      RECT  37640.0 106730.0 38345.0 105385.0 ;
      RECT  37640.0 106730.0 38345.0 108075.0 ;
      RECT  37640.0 109420.0 38345.0 108075.0 ;
      RECT  37640.0 109420.0 38345.0 110765.0 ;
      RECT  37640.0 112110.0 38345.0 110765.0 ;
      RECT  37640.0 112110.0 38345.0 113455.0 ;
      RECT  37640.0 114800.0 38345.0 113455.0 ;
      RECT  37640.0 114800.0 38345.0 116145.0 ;
      RECT  37640.0 117490.0 38345.0 116145.0 ;
      RECT  37640.0 117490.0 38345.0 118835.0 ;
      RECT  37640.0 120180.0 38345.0 118835.0 ;
      RECT  37640.0 120180.0 38345.0 121525.0 ;
      RECT  37640.0 122870.0 38345.0 121525.0 ;
      RECT  37640.0 122870.0 38345.0 124215.0 ;
      RECT  37640.0 125560.0 38345.0 124215.0 ;
      RECT  37640.0 125560.0 38345.0 126905.0 ;
      RECT  37640.0 128250.0 38345.0 126905.0 ;
      RECT  37640.0 128250.0 38345.0 129595.0 ;
      RECT  37640.0 130940.0 38345.0 129595.0 ;
      RECT  37640.0 130940.0 38345.0 132285.0 ;
      RECT  37640.0 133630.0 38345.0 132285.0 ;
      RECT  37640.0 133630.0 38345.0 134975.0 ;
      RECT  37640.0 136320.0 38345.0 134975.0 ;
      RECT  37640.0 136320.0 38345.0 137665.0 ;
      RECT  37640.0 139010.0 38345.0 137665.0 ;
      RECT  37640.0 139010.0 38345.0 140355.0 ;
      RECT  37640.0 141700.0 38345.0 140355.0 ;
      RECT  37640.0 141700.0 38345.0 143045.0 ;
      RECT  37640.0 144390.0 38345.0 143045.0 ;
      RECT  37640.0 144390.0 38345.0 145735.0 ;
      RECT  37640.0 147080.0 38345.0 145735.0 ;
      RECT  37640.0 147080.0 38345.0 148425.0 ;
      RECT  37640.0 149770.0 38345.0 148425.0 ;
      RECT  37640.0 149770.0 38345.0 151115.0 ;
      RECT  37640.0 152460.0 38345.0 151115.0 ;
      RECT  37640.0 152460.0 38345.0 153805.0 ;
      RECT  37640.0 155150.0 38345.0 153805.0 ;
      RECT  37640.0 155150.0 38345.0 156495.0 ;
      RECT  37640.0 157840.0 38345.0 156495.0 ;
      RECT  37640.0 157840.0 38345.0 159185.0 ;
      RECT  37640.0 160530.0 38345.0 159185.0 ;
      RECT  37640.0 160530.0 38345.0 161875.0 ;
      RECT  37640.0 163220.0 38345.0 161875.0 ;
      RECT  37640.0 163220.0 38345.0 164565.0 ;
      RECT  37640.0 165910.0 38345.0 164565.0 ;
      RECT  37640.0 165910.0 38345.0 167255.0 ;
      RECT  37640.0 168600.0 38345.0 167255.0 ;
      RECT  37640.0 168600.0 38345.0 169945.0 ;
      RECT  37640.0 171290.0 38345.0 169945.0 ;
      RECT  37640.0 171290.0 38345.0 172635.0 ;
      RECT  37640.0 173980.0 38345.0 172635.0 ;
      RECT  37640.0 173980.0 38345.0 175325.0 ;
      RECT  37640.0 176670.0 38345.0 175325.0 ;
      RECT  37640.0 176670.0 38345.0 178015.0 ;
      RECT  37640.0 179360.0 38345.0 178015.0 ;
      RECT  37640.0 179360.0 38345.0 180705.0 ;
      RECT  37640.0 182050.0 38345.0 180705.0 ;
      RECT  37640.0 182050.0 38345.0 183395.0 ;
      RECT  37640.0 184740.0 38345.0 183395.0 ;
      RECT  37640.0 184740.0 38345.0 186085.0 ;
      RECT  37640.0 187430.0 38345.0 186085.0 ;
      RECT  37640.0 187430.0 38345.0 188775.0 ;
      RECT  37640.0 190120.0 38345.0 188775.0 ;
      RECT  37640.0 190120.0 38345.0 191465.0 ;
      RECT  37640.0 192810.0 38345.0 191465.0 ;
      RECT  37640.0 192810.0 38345.0 194155.0 ;
      RECT  37640.0 195500.0 38345.0 194155.0 ;
      RECT  37640.0 195500.0 38345.0 196845.0 ;
      RECT  37640.0 198190.0 38345.0 196845.0 ;
      RECT  37640.0 198190.0 38345.0 199535.0 ;
      RECT  37640.0 200880.0 38345.0 199535.0 ;
      RECT  37640.0 200880.0 38345.0 202225.0 ;
      RECT  37640.0 203570.0 38345.0 202225.0 ;
      RECT  37640.0 203570.0 38345.0 204915.0 ;
      RECT  37640.0 206260.0 38345.0 204915.0 ;
      RECT  38345.0 34100.0 39050.0 35445.0 ;
      RECT  38345.0 36790.0 39050.0 35445.0 ;
      RECT  38345.0 36790.0 39050.0 38135.0 ;
      RECT  38345.0 39480.0 39050.0 38135.0 ;
      RECT  38345.0 39480.0 39050.0 40825.0 ;
      RECT  38345.0 42170.0 39050.0 40825.0 ;
      RECT  38345.0 42170.0 39050.0 43515.0 ;
      RECT  38345.0 44860.0 39050.0 43515.0 ;
      RECT  38345.0 44860.0 39050.0 46205.0 ;
      RECT  38345.0 47550.0 39050.0 46205.0 ;
      RECT  38345.0 47550.0 39050.0 48895.0 ;
      RECT  38345.0 50240.0 39050.0 48895.0 ;
      RECT  38345.0 50240.0 39050.0 51585.0 ;
      RECT  38345.0 52930.0 39050.0 51585.0 ;
      RECT  38345.0 52930.0 39050.0 54275.0 ;
      RECT  38345.0 55620.0 39050.0 54275.0 ;
      RECT  38345.0 55620.0 39050.0 56965.0 ;
      RECT  38345.0 58310.0 39050.0 56965.0 ;
      RECT  38345.0 58310.0 39050.0 59655.0 ;
      RECT  38345.0 61000.0 39050.0 59655.0 ;
      RECT  38345.0 61000.0 39050.0 62345.0 ;
      RECT  38345.0 63690.0 39050.0 62345.0 ;
      RECT  38345.0 63690.0 39050.0 65035.0 ;
      RECT  38345.0 66380.0 39050.0 65035.0 ;
      RECT  38345.0 66380.0 39050.0 67725.0 ;
      RECT  38345.0 69070.0 39050.0 67725.0 ;
      RECT  38345.0 69070.0 39050.0 70415.0 ;
      RECT  38345.0 71760.0 39050.0 70415.0 ;
      RECT  38345.0 71760.0 39050.0 73105.0 ;
      RECT  38345.0 74450.0 39050.0 73105.0 ;
      RECT  38345.0 74450.0 39050.0 75795.0 ;
      RECT  38345.0 77140.0 39050.0 75795.0 ;
      RECT  38345.0 77140.0 39050.0 78485.0 ;
      RECT  38345.0 79830.0 39050.0 78485.0 ;
      RECT  38345.0 79830.0 39050.0 81175.0 ;
      RECT  38345.0 82520.0 39050.0 81175.0 ;
      RECT  38345.0 82520.0 39050.0 83865.0 ;
      RECT  38345.0 85210.0 39050.0 83865.0 ;
      RECT  38345.0 85210.0 39050.0 86555.0 ;
      RECT  38345.0 87900.0 39050.0 86555.0 ;
      RECT  38345.0 87900.0 39050.0 89245.0 ;
      RECT  38345.0 90590.0 39050.0 89245.0 ;
      RECT  38345.0 90590.0 39050.0 91935.0 ;
      RECT  38345.0 93280.0 39050.0 91935.0 ;
      RECT  38345.0 93280.0 39050.0 94625.0 ;
      RECT  38345.0 95970.0 39050.0 94625.0 ;
      RECT  38345.0 95970.0 39050.0 97315.0 ;
      RECT  38345.0 98660.0 39050.0 97315.0 ;
      RECT  38345.0 98660.0 39050.0 100005.0 ;
      RECT  38345.0 101350.0 39050.0 100005.0 ;
      RECT  38345.0 101350.0 39050.0 102695.0 ;
      RECT  38345.0 104040.0 39050.0 102695.0 ;
      RECT  38345.0 104040.0 39050.0 105385.0 ;
      RECT  38345.0 106730.0 39050.0 105385.0 ;
      RECT  38345.0 106730.0 39050.0 108075.0 ;
      RECT  38345.0 109420.0 39050.0 108075.0 ;
      RECT  38345.0 109420.0 39050.0 110765.0 ;
      RECT  38345.0 112110.0 39050.0 110765.0 ;
      RECT  38345.0 112110.0 39050.0 113455.0 ;
      RECT  38345.0 114800.0 39050.0 113455.0 ;
      RECT  38345.0 114800.0 39050.0 116145.0 ;
      RECT  38345.0 117490.0 39050.0 116145.0 ;
      RECT  38345.0 117490.0 39050.0 118835.0 ;
      RECT  38345.0 120180.0 39050.0 118835.0 ;
      RECT  38345.0 120180.0 39050.0 121525.0 ;
      RECT  38345.0 122870.0 39050.0 121525.0 ;
      RECT  38345.0 122870.0 39050.0 124215.0 ;
      RECT  38345.0 125560.0 39050.0 124215.0 ;
      RECT  38345.0 125560.0 39050.0 126905.0 ;
      RECT  38345.0 128250.0 39050.0 126905.0 ;
      RECT  38345.0 128250.0 39050.0 129595.0 ;
      RECT  38345.0 130940.0 39050.0 129595.0 ;
      RECT  38345.0 130940.0 39050.0 132285.0 ;
      RECT  38345.0 133630.0 39050.0 132285.0 ;
      RECT  38345.0 133630.0 39050.0 134975.0 ;
      RECT  38345.0 136320.0 39050.0 134975.0 ;
      RECT  38345.0 136320.0 39050.0 137665.0 ;
      RECT  38345.0 139010.0 39050.0 137665.0 ;
      RECT  38345.0 139010.0 39050.0 140355.0 ;
      RECT  38345.0 141700.0 39050.0 140355.0 ;
      RECT  38345.0 141700.0 39050.0 143045.0 ;
      RECT  38345.0 144390.0 39050.0 143045.0 ;
      RECT  38345.0 144390.0 39050.0 145735.0 ;
      RECT  38345.0 147080.0 39050.0 145735.0 ;
      RECT  38345.0 147080.0 39050.0 148425.0 ;
      RECT  38345.0 149770.0 39050.0 148425.0 ;
      RECT  38345.0 149770.0 39050.0 151115.0 ;
      RECT  38345.0 152460.0 39050.0 151115.0 ;
      RECT  38345.0 152460.0 39050.0 153805.0 ;
      RECT  38345.0 155150.0 39050.0 153805.0 ;
      RECT  38345.0 155150.0 39050.0 156495.0 ;
      RECT  38345.0 157840.0 39050.0 156495.0 ;
      RECT  38345.0 157840.0 39050.0 159185.0 ;
      RECT  38345.0 160530.0 39050.0 159185.0 ;
      RECT  38345.0 160530.0 39050.0 161875.0 ;
      RECT  38345.0 163220.0 39050.0 161875.0 ;
      RECT  38345.0 163220.0 39050.0 164565.0 ;
      RECT  38345.0 165910.0 39050.0 164565.0 ;
      RECT  38345.0 165910.0 39050.0 167255.0 ;
      RECT  38345.0 168600.0 39050.0 167255.0 ;
      RECT  38345.0 168600.0 39050.0 169945.0 ;
      RECT  38345.0 171290.0 39050.0 169945.0 ;
      RECT  38345.0 171290.0 39050.0 172635.0 ;
      RECT  38345.0 173980.0 39050.0 172635.0 ;
      RECT  38345.0 173980.0 39050.0 175325.0 ;
      RECT  38345.0 176670.0 39050.0 175325.0 ;
      RECT  38345.0 176670.0 39050.0 178015.0 ;
      RECT  38345.0 179360.0 39050.0 178015.0 ;
      RECT  38345.0 179360.0 39050.0 180705.0 ;
      RECT  38345.0 182050.0 39050.0 180705.0 ;
      RECT  38345.0 182050.0 39050.0 183395.0 ;
      RECT  38345.0 184740.0 39050.0 183395.0 ;
      RECT  38345.0 184740.0 39050.0 186085.0 ;
      RECT  38345.0 187430.0 39050.0 186085.0 ;
      RECT  38345.0 187430.0 39050.0 188775.0 ;
      RECT  38345.0 190120.0 39050.0 188775.0 ;
      RECT  38345.0 190120.0 39050.0 191465.0 ;
      RECT  38345.0 192810.0 39050.0 191465.0 ;
      RECT  38345.0 192810.0 39050.0 194155.0 ;
      RECT  38345.0 195500.0 39050.0 194155.0 ;
      RECT  38345.0 195500.0 39050.0 196845.0 ;
      RECT  38345.0 198190.0 39050.0 196845.0 ;
      RECT  38345.0 198190.0 39050.0 199535.0 ;
      RECT  38345.0 200880.0 39050.0 199535.0 ;
      RECT  38345.0 200880.0 39050.0 202225.0 ;
      RECT  38345.0 203570.0 39050.0 202225.0 ;
      RECT  38345.0 203570.0 39050.0 204915.0 ;
      RECT  38345.0 206260.0 39050.0 204915.0 ;
      RECT  39050.0 34100.0 39755.0 35445.0 ;
      RECT  39050.0 36790.0 39755.0 35445.0 ;
      RECT  39050.0 36790.0 39755.0 38135.0 ;
      RECT  39050.0 39480.0 39755.0 38135.0 ;
      RECT  39050.0 39480.0 39755.0 40825.0 ;
      RECT  39050.0 42170.0 39755.0 40825.0 ;
      RECT  39050.0 42170.0 39755.0 43515.0 ;
      RECT  39050.0 44860.0 39755.0 43515.0 ;
      RECT  39050.0 44860.0 39755.0 46205.0 ;
      RECT  39050.0 47550.0 39755.0 46205.0 ;
      RECT  39050.0 47550.0 39755.0 48895.0 ;
      RECT  39050.0 50240.0 39755.0 48895.0 ;
      RECT  39050.0 50240.0 39755.0 51585.0 ;
      RECT  39050.0 52930.0 39755.0 51585.0 ;
      RECT  39050.0 52930.0 39755.0 54275.0 ;
      RECT  39050.0 55620.0 39755.0 54275.0 ;
      RECT  39050.0 55620.0 39755.0 56965.0 ;
      RECT  39050.0 58310.0 39755.0 56965.0 ;
      RECT  39050.0 58310.0 39755.0 59655.0 ;
      RECT  39050.0 61000.0 39755.0 59655.0 ;
      RECT  39050.0 61000.0 39755.0 62345.0 ;
      RECT  39050.0 63690.0 39755.0 62345.0 ;
      RECT  39050.0 63690.0 39755.0 65035.0 ;
      RECT  39050.0 66380.0 39755.0 65035.0 ;
      RECT  39050.0 66380.0 39755.0 67725.0 ;
      RECT  39050.0 69070.0 39755.0 67725.0 ;
      RECT  39050.0 69070.0 39755.0 70415.0 ;
      RECT  39050.0 71760.0 39755.0 70415.0 ;
      RECT  39050.0 71760.0 39755.0 73105.0 ;
      RECT  39050.0 74450.0 39755.0 73105.0 ;
      RECT  39050.0 74450.0 39755.0 75795.0 ;
      RECT  39050.0 77140.0 39755.0 75795.0 ;
      RECT  39050.0 77140.0 39755.0 78485.0 ;
      RECT  39050.0 79830.0 39755.0 78485.0 ;
      RECT  39050.0 79830.0 39755.0 81175.0 ;
      RECT  39050.0 82520.0 39755.0 81175.0 ;
      RECT  39050.0 82520.0 39755.0 83865.0 ;
      RECT  39050.0 85210.0 39755.0 83865.0 ;
      RECT  39050.0 85210.0 39755.0 86555.0 ;
      RECT  39050.0 87900.0 39755.0 86555.0 ;
      RECT  39050.0 87900.0 39755.0 89245.0 ;
      RECT  39050.0 90590.0 39755.0 89245.0 ;
      RECT  39050.0 90590.0 39755.0 91935.0 ;
      RECT  39050.0 93280.0 39755.0 91935.0 ;
      RECT  39050.0 93280.0 39755.0 94625.0 ;
      RECT  39050.0 95970.0 39755.0 94625.0 ;
      RECT  39050.0 95970.0 39755.0 97315.0 ;
      RECT  39050.0 98660.0 39755.0 97315.0 ;
      RECT  39050.0 98660.0 39755.0 100005.0 ;
      RECT  39050.0 101350.0 39755.0 100005.0 ;
      RECT  39050.0 101350.0 39755.0 102695.0 ;
      RECT  39050.0 104040.0 39755.0 102695.0 ;
      RECT  39050.0 104040.0 39755.0 105385.0 ;
      RECT  39050.0 106730.0 39755.0 105385.0 ;
      RECT  39050.0 106730.0 39755.0 108075.0 ;
      RECT  39050.0 109420.0 39755.0 108075.0 ;
      RECT  39050.0 109420.0 39755.0 110765.0 ;
      RECT  39050.0 112110.0 39755.0 110765.0 ;
      RECT  39050.0 112110.0 39755.0 113455.0 ;
      RECT  39050.0 114800.0 39755.0 113455.0 ;
      RECT  39050.0 114800.0 39755.0 116145.0 ;
      RECT  39050.0 117490.0 39755.0 116145.0 ;
      RECT  39050.0 117490.0 39755.0 118835.0 ;
      RECT  39050.0 120180.0 39755.0 118835.0 ;
      RECT  39050.0 120180.0 39755.0 121525.0 ;
      RECT  39050.0 122870.0 39755.0 121525.0 ;
      RECT  39050.0 122870.0 39755.0 124215.0 ;
      RECT  39050.0 125560.0 39755.0 124215.0 ;
      RECT  39050.0 125560.0 39755.0 126905.0 ;
      RECT  39050.0 128250.0 39755.0 126905.0 ;
      RECT  39050.0 128250.0 39755.0 129595.0 ;
      RECT  39050.0 130940.0 39755.0 129595.0 ;
      RECT  39050.0 130940.0 39755.0 132285.0 ;
      RECT  39050.0 133630.0 39755.0 132285.0 ;
      RECT  39050.0 133630.0 39755.0 134975.0 ;
      RECT  39050.0 136320.0 39755.0 134975.0 ;
      RECT  39050.0 136320.0 39755.0 137665.0 ;
      RECT  39050.0 139010.0 39755.0 137665.0 ;
      RECT  39050.0 139010.0 39755.0 140355.0 ;
      RECT  39050.0 141700.0 39755.0 140355.0 ;
      RECT  39050.0 141700.0 39755.0 143045.0 ;
      RECT  39050.0 144390.0 39755.0 143045.0 ;
      RECT  39050.0 144390.0 39755.0 145735.0 ;
      RECT  39050.0 147080.0 39755.0 145735.0 ;
      RECT  39050.0 147080.0 39755.0 148425.0 ;
      RECT  39050.0 149770.0 39755.0 148425.0 ;
      RECT  39050.0 149770.0 39755.0 151115.0 ;
      RECT  39050.0 152460.0 39755.0 151115.0 ;
      RECT  39050.0 152460.0 39755.0 153805.0 ;
      RECT  39050.0 155150.0 39755.0 153805.0 ;
      RECT  39050.0 155150.0 39755.0 156495.0 ;
      RECT  39050.0 157840.0 39755.0 156495.0 ;
      RECT  39050.0 157840.0 39755.0 159185.0 ;
      RECT  39050.0 160530.0 39755.0 159185.0 ;
      RECT  39050.0 160530.0 39755.0 161875.0 ;
      RECT  39050.0 163220.0 39755.0 161875.0 ;
      RECT  39050.0 163220.0 39755.0 164565.0 ;
      RECT  39050.0 165910.0 39755.0 164565.0 ;
      RECT  39050.0 165910.0 39755.0 167255.0 ;
      RECT  39050.0 168600.0 39755.0 167255.0 ;
      RECT  39050.0 168600.0 39755.0 169945.0 ;
      RECT  39050.0 171290.0 39755.0 169945.0 ;
      RECT  39050.0 171290.0 39755.0 172635.0 ;
      RECT  39050.0 173980.0 39755.0 172635.0 ;
      RECT  39050.0 173980.0 39755.0 175325.0 ;
      RECT  39050.0 176670.0 39755.0 175325.0 ;
      RECT  39050.0 176670.0 39755.0 178015.0 ;
      RECT  39050.0 179360.0 39755.0 178015.0 ;
      RECT  39050.0 179360.0 39755.0 180705.0 ;
      RECT  39050.0 182050.0 39755.0 180705.0 ;
      RECT  39050.0 182050.0 39755.0 183395.0 ;
      RECT  39050.0 184740.0 39755.0 183395.0 ;
      RECT  39050.0 184740.0 39755.0 186085.0 ;
      RECT  39050.0 187430.0 39755.0 186085.0 ;
      RECT  39050.0 187430.0 39755.0 188775.0 ;
      RECT  39050.0 190120.0 39755.0 188775.0 ;
      RECT  39050.0 190120.0 39755.0 191465.0 ;
      RECT  39050.0 192810.0 39755.0 191465.0 ;
      RECT  39050.0 192810.0 39755.0 194155.0 ;
      RECT  39050.0 195500.0 39755.0 194155.0 ;
      RECT  39050.0 195500.0 39755.0 196845.0 ;
      RECT  39050.0 198190.0 39755.0 196845.0 ;
      RECT  39050.0 198190.0 39755.0 199535.0 ;
      RECT  39050.0 200880.0 39755.0 199535.0 ;
      RECT  39050.0 200880.0 39755.0 202225.0 ;
      RECT  39050.0 203570.0 39755.0 202225.0 ;
      RECT  39050.0 203570.0 39755.0 204915.0 ;
      RECT  39050.0 206260.0 39755.0 204915.0 ;
      RECT  39755.0 34100.0 40460.0 35445.0 ;
      RECT  39755.0 36790.0 40460.0 35445.0 ;
      RECT  39755.0 36790.0 40460.0 38135.0 ;
      RECT  39755.0 39480.0 40460.0 38135.0 ;
      RECT  39755.0 39480.0 40460.0 40825.0 ;
      RECT  39755.0 42170.0 40460.0 40825.0 ;
      RECT  39755.0 42170.0 40460.0 43515.0 ;
      RECT  39755.0 44860.0 40460.0 43515.0 ;
      RECT  39755.0 44860.0 40460.0 46205.0 ;
      RECT  39755.0 47550.0 40460.0 46205.0 ;
      RECT  39755.0 47550.0 40460.0 48895.0 ;
      RECT  39755.0 50240.0 40460.0 48895.0 ;
      RECT  39755.0 50240.0 40460.0 51585.0 ;
      RECT  39755.0 52930.0 40460.0 51585.0 ;
      RECT  39755.0 52930.0 40460.0 54275.0 ;
      RECT  39755.0 55620.0 40460.0 54275.0 ;
      RECT  39755.0 55620.0 40460.0 56965.0 ;
      RECT  39755.0 58310.0 40460.0 56965.0 ;
      RECT  39755.0 58310.0 40460.0 59655.0 ;
      RECT  39755.0 61000.0 40460.0 59655.0 ;
      RECT  39755.0 61000.0 40460.0 62345.0 ;
      RECT  39755.0 63690.0 40460.0 62345.0 ;
      RECT  39755.0 63690.0 40460.0 65035.0 ;
      RECT  39755.0 66380.0 40460.0 65035.0 ;
      RECT  39755.0 66380.0 40460.0 67725.0 ;
      RECT  39755.0 69070.0 40460.0 67725.0 ;
      RECT  39755.0 69070.0 40460.0 70415.0 ;
      RECT  39755.0 71760.0 40460.0 70415.0 ;
      RECT  39755.0 71760.0 40460.0 73105.0 ;
      RECT  39755.0 74450.0 40460.0 73105.0 ;
      RECT  39755.0 74450.0 40460.0 75795.0 ;
      RECT  39755.0 77140.0 40460.0 75795.0 ;
      RECT  39755.0 77140.0 40460.0 78485.0 ;
      RECT  39755.0 79830.0 40460.0 78485.0 ;
      RECT  39755.0 79830.0 40460.0 81175.0 ;
      RECT  39755.0 82520.0 40460.0 81175.0 ;
      RECT  39755.0 82520.0 40460.0 83865.0 ;
      RECT  39755.0 85210.0 40460.0 83865.0 ;
      RECT  39755.0 85210.0 40460.0 86555.0 ;
      RECT  39755.0 87900.0 40460.0 86555.0 ;
      RECT  39755.0 87900.0 40460.0 89245.0 ;
      RECT  39755.0 90590.0 40460.0 89245.0 ;
      RECT  39755.0 90590.0 40460.0 91935.0 ;
      RECT  39755.0 93280.0 40460.0 91935.0 ;
      RECT  39755.0 93280.0 40460.0 94625.0 ;
      RECT  39755.0 95970.0 40460.0 94625.0 ;
      RECT  39755.0 95970.0 40460.0 97315.0 ;
      RECT  39755.0 98660.0 40460.0 97315.0 ;
      RECT  39755.0 98660.0 40460.0 100005.0 ;
      RECT  39755.0 101350.0 40460.0 100005.0 ;
      RECT  39755.0 101350.0 40460.0 102695.0 ;
      RECT  39755.0 104040.0 40460.0 102695.0 ;
      RECT  39755.0 104040.0 40460.0 105385.0 ;
      RECT  39755.0 106730.0 40460.0 105385.0 ;
      RECT  39755.0 106730.0 40460.0 108075.0 ;
      RECT  39755.0 109420.0 40460.0 108075.0 ;
      RECT  39755.0 109420.0 40460.0 110765.0 ;
      RECT  39755.0 112110.0 40460.0 110765.0 ;
      RECT  39755.0 112110.0 40460.0 113455.0 ;
      RECT  39755.0 114800.0 40460.0 113455.0 ;
      RECT  39755.0 114800.0 40460.0 116145.0 ;
      RECT  39755.0 117490.0 40460.0 116145.0 ;
      RECT  39755.0 117490.0 40460.0 118835.0 ;
      RECT  39755.0 120180.0 40460.0 118835.0 ;
      RECT  39755.0 120180.0 40460.0 121525.0 ;
      RECT  39755.0 122870.0 40460.0 121525.0 ;
      RECT  39755.0 122870.0 40460.0 124215.0 ;
      RECT  39755.0 125560.0 40460.0 124215.0 ;
      RECT  39755.0 125560.0 40460.0 126905.0 ;
      RECT  39755.0 128250.0 40460.0 126905.0 ;
      RECT  39755.0 128250.0 40460.0 129595.0 ;
      RECT  39755.0 130940.0 40460.0 129595.0 ;
      RECT  39755.0 130940.0 40460.0 132285.0 ;
      RECT  39755.0 133630.0 40460.0 132285.0 ;
      RECT  39755.0 133630.0 40460.0 134975.0 ;
      RECT  39755.0 136320.0 40460.0 134975.0 ;
      RECT  39755.0 136320.0 40460.0 137665.0 ;
      RECT  39755.0 139010.0 40460.0 137665.0 ;
      RECT  39755.0 139010.0 40460.0 140355.0 ;
      RECT  39755.0 141700.0 40460.0 140355.0 ;
      RECT  39755.0 141700.0 40460.0 143045.0 ;
      RECT  39755.0 144390.0 40460.0 143045.0 ;
      RECT  39755.0 144390.0 40460.0 145735.0 ;
      RECT  39755.0 147080.0 40460.0 145735.0 ;
      RECT  39755.0 147080.0 40460.0 148425.0 ;
      RECT  39755.0 149770.0 40460.0 148425.0 ;
      RECT  39755.0 149770.0 40460.0 151115.0 ;
      RECT  39755.0 152460.0 40460.0 151115.0 ;
      RECT  39755.0 152460.0 40460.0 153805.0 ;
      RECT  39755.0 155150.0 40460.0 153805.0 ;
      RECT  39755.0 155150.0 40460.0 156495.0 ;
      RECT  39755.0 157840.0 40460.0 156495.0 ;
      RECT  39755.0 157840.0 40460.0 159185.0 ;
      RECT  39755.0 160530.0 40460.0 159185.0 ;
      RECT  39755.0 160530.0 40460.0 161875.0 ;
      RECT  39755.0 163220.0 40460.0 161875.0 ;
      RECT  39755.0 163220.0 40460.0 164565.0 ;
      RECT  39755.0 165910.0 40460.0 164565.0 ;
      RECT  39755.0 165910.0 40460.0 167255.0 ;
      RECT  39755.0 168600.0 40460.0 167255.0 ;
      RECT  39755.0 168600.0 40460.0 169945.0 ;
      RECT  39755.0 171290.0 40460.0 169945.0 ;
      RECT  39755.0 171290.0 40460.0 172635.0 ;
      RECT  39755.0 173980.0 40460.0 172635.0 ;
      RECT  39755.0 173980.0 40460.0 175325.0 ;
      RECT  39755.0 176670.0 40460.0 175325.0 ;
      RECT  39755.0 176670.0 40460.0 178015.0 ;
      RECT  39755.0 179360.0 40460.0 178015.0 ;
      RECT  39755.0 179360.0 40460.0 180705.0 ;
      RECT  39755.0 182050.0 40460.0 180705.0 ;
      RECT  39755.0 182050.0 40460.0 183395.0 ;
      RECT  39755.0 184740.0 40460.0 183395.0 ;
      RECT  39755.0 184740.0 40460.0 186085.0 ;
      RECT  39755.0 187430.0 40460.0 186085.0 ;
      RECT  39755.0 187430.0 40460.0 188775.0 ;
      RECT  39755.0 190120.0 40460.0 188775.0 ;
      RECT  39755.0 190120.0 40460.0 191465.0 ;
      RECT  39755.0 192810.0 40460.0 191465.0 ;
      RECT  39755.0 192810.0 40460.0 194155.0 ;
      RECT  39755.0 195500.0 40460.0 194155.0 ;
      RECT  39755.0 195500.0 40460.0 196845.0 ;
      RECT  39755.0 198190.0 40460.0 196845.0 ;
      RECT  39755.0 198190.0 40460.0 199535.0 ;
      RECT  39755.0 200880.0 40460.0 199535.0 ;
      RECT  39755.0 200880.0 40460.0 202225.0 ;
      RECT  39755.0 203570.0 40460.0 202225.0 ;
      RECT  39755.0 203570.0 40460.0 204915.0 ;
      RECT  39755.0 206260.0 40460.0 204915.0 ;
      RECT  40460.0 34100.0 41165.0 35445.0 ;
      RECT  40460.0 36790.0 41165.0 35445.0 ;
      RECT  40460.0 36790.0 41165.0 38135.0 ;
      RECT  40460.0 39480.0 41165.0 38135.0 ;
      RECT  40460.0 39480.0 41165.0 40825.0 ;
      RECT  40460.0 42170.0 41165.0 40825.0 ;
      RECT  40460.0 42170.0 41165.0 43515.0 ;
      RECT  40460.0 44860.0 41165.0 43515.0 ;
      RECT  40460.0 44860.0 41165.0 46205.0 ;
      RECT  40460.0 47550.0 41165.0 46205.0 ;
      RECT  40460.0 47550.0 41165.0 48895.0 ;
      RECT  40460.0 50240.0 41165.0 48895.0 ;
      RECT  40460.0 50240.0 41165.0 51585.0 ;
      RECT  40460.0 52930.0 41165.0 51585.0 ;
      RECT  40460.0 52930.0 41165.0 54275.0 ;
      RECT  40460.0 55620.0 41165.0 54275.0 ;
      RECT  40460.0 55620.0 41165.0 56965.0 ;
      RECT  40460.0 58310.0 41165.0 56965.0 ;
      RECT  40460.0 58310.0 41165.0 59655.0 ;
      RECT  40460.0 61000.0 41165.0 59655.0 ;
      RECT  40460.0 61000.0 41165.0 62345.0 ;
      RECT  40460.0 63690.0 41165.0 62345.0 ;
      RECT  40460.0 63690.0 41165.0 65035.0 ;
      RECT  40460.0 66380.0 41165.0 65035.0 ;
      RECT  40460.0 66380.0 41165.0 67725.0 ;
      RECT  40460.0 69070.0 41165.0 67725.0 ;
      RECT  40460.0 69070.0 41165.0 70415.0 ;
      RECT  40460.0 71760.0 41165.0 70415.0 ;
      RECT  40460.0 71760.0 41165.0 73105.0 ;
      RECT  40460.0 74450.0 41165.0 73105.0 ;
      RECT  40460.0 74450.0 41165.0 75795.0 ;
      RECT  40460.0 77140.0 41165.0 75795.0 ;
      RECT  40460.0 77140.0 41165.0 78485.0 ;
      RECT  40460.0 79830.0 41165.0 78485.0 ;
      RECT  40460.0 79830.0 41165.0 81175.0 ;
      RECT  40460.0 82520.0 41165.0 81175.0 ;
      RECT  40460.0 82520.0 41165.0 83865.0 ;
      RECT  40460.0 85210.0 41165.0 83865.0 ;
      RECT  40460.0 85210.0 41165.0 86555.0 ;
      RECT  40460.0 87900.0 41165.0 86555.0 ;
      RECT  40460.0 87900.0 41165.0 89245.0 ;
      RECT  40460.0 90590.0 41165.0 89245.0 ;
      RECT  40460.0 90590.0 41165.0 91935.0 ;
      RECT  40460.0 93280.0 41165.0 91935.0 ;
      RECT  40460.0 93280.0 41165.0 94625.0 ;
      RECT  40460.0 95970.0 41165.0 94625.0 ;
      RECT  40460.0 95970.0 41165.0 97315.0 ;
      RECT  40460.0 98660.0 41165.0 97315.0 ;
      RECT  40460.0 98660.0 41165.0 100005.0 ;
      RECT  40460.0 101350.0 41165.0 100005.0 ;
      RECT  40460.0 101350.0 41165.0 102695.0 ;
      RECT  40460.0 104040.0 41165.0 102695.0 ;
      RECT  40460.0 104040.0 41165.0 105385.0 ;
      RECT  40460.0 106730.0 41165.0 105385.0 ;
      RECT  40460.0 106730.0 41165.0 108075.0 ;
      RECT  40460.0 109420.0 41165.0 108075.0 ;
      RECT  40460.0 109420.0 41165.0 110765.0 ;
      RECT  40460.0 112110.0 41165.0 110765.0 ;
      RECT  40460.0 112110.0 41165.0 113455.0 ;
      RECT  40460.0 114800.0 41165.0 113455.0 ;
      RECT  40460.0 114800.0 41165.0 116145.0 ;
      RECT  40460.0 117490.0 41165.0 116145.0 ;
      RECT  40460.0 117490.0 41165.0 118835.0 ;
      RECT  40460.0 120180.0 41165.0 118835.0 ;
      RECT  40460.0 120180.0 41165.0 121525.0 ;
      RECT  40460.0 122870.0 41165.0 121525.0 ;
      RECT  40460.0 122870.0 41165.0 124215.0 ;
      RECT  40460.0 125560.0 41165.0 124215.0 ;
      RECT  40460.0 125560.0 41165.0 126905.0 ;
      RECT  40460.0 128250.0 41165.0 126905.0 ;
      RECT  40460.0 128250.0 41165.0 129595.0 ;
      RECT  40460.0 130940.0 41165.0 129595.0 ;
      RECT  40460.0 130940.0 41165.0 132285.0 ;
      RECT  40460.0 133630.0 41165.0 132285.0 ;
      RECT  40460.0 133630.0 41165.0 134975.0 ;
      RECT  40460.0 136320.0 41165.0 134975.0 ;
      RECT  40460.0 136320.0 41165.0 137665.0 ;
      RECT  40460.0 139010.0 41165.0 137665.0 ;
      RECT  40460.0 139010.0 41165.0 140355.0 ;
      RECT  40460.0 141700.0 41165.0 140355.0 ;
      RECT  40460.0 141700.0 41165.0 143045.0 ;
      RECT  40460.0 144390.0 41165.0 143045.0 ;
      RECT  40460.0 144390.0 41165.0 145735.0 ;
      RECT  40460.0 147080.0 41165.0 145735.0 ;
      RECT  40460.0 147080.0 41165.0 148425.0 ;
      RECT  40460.0 149770.0 41165.0 148425.0 ;
      RECT  40460.0 149770.0 41165.0 151115.0 ;
      RECT  40460.0 152460.0 41165.0 151115.0 ;
      RECT  40460.0 152460.0 41165.0 153805.0 ;
      RECT  40460.0 155150.0 41165.0 153805.0 ;
      RECT  40460.0 155150.0 41165.0 156495.0 ;
      RECT  40460.0 157840.0 41165.0 156495.0 ;
      RECT  40460.0 157840.0 41165.0 159185.0 ;
      RECT  40460.0 160530.0 41165.0 159185.0 ;
      RECT  40460.0 160530.0 41165.0 161875.0 ;
      RECT  40460.0 163220.0 41165.0 161875.0 ;
      RECT  40460.0 163220.0 41165.0 164565.0 ;
      RECT  40460.0 165910.0 41165.0 164565.0 ;
      RECT  40460.0 165910.0 41165.0 167255.0 ;
      RECT  40460.0 168600.0 41165.0 167255.0 ;
      RECT  40460.0 168600.0 41165.0 169945.0 ;
      RECT  40460.0 171290.0 41165.0 169945.0 ;
      RECT  40460.0 171290.0 41165.0 172635.0 ;
      RECT  40460.0 173980.0 41165.0 172635.0 ;
      RECT  40460.0 173980.0 41165.0 175325.0 ;
      RECT  40460.0 176670.0 41165.0 175325.0 ;
      RECT  40460.0 176670.0 41165.0 178015.0 ;
      RECT  40460.0 179360.0 41165.0 178015.0 ;
      RECT  40460.0 179360.0 41165.0 180705.0 ;
      RECT  40460.0 182050.0 41165.0 180705.0 ;
      RECT  40460.0 182050.0 41165.0 183395.0 ;
      RECT  40460.0 184740.0 41165.0 183395.0 ;
      RECT  40460.0 184740.0 41165.0 186085.0 ;
      RECT  40460.0 187430.0 41165.0 186085.0 ;
      RECT  40460.0 187430.0 41165.0 188775.0 ;
      RECT  40460.0 190120.0 41165.0 188775.0 ;
      RECT  40460.0 190120.0 41165.0 191465.0 ;
      RECT  40460.0 192810.0 41165.0 191465.0 ;
      RECT  40460.0 192810.0 41165.0 194155.0 ;
      RECT  40460.0 195500.0 41165.0 194155.0 ;
      RECT  40460.0 195500.0 41165.0 196845.0 ;
      RECT  40460.0 198190.0 41165.0 196845.0 ;
      RECT  40460.0 198190.0 41165.0 199535.0 ;
      RECT  40460.0 200880.0 41165.0 199535.0 ;
      RECT  40460.0 200880.0 41165.0 202225.0 ;
      RECT  40460.0 203570.0 41165.0 202225.0 ;
      RECT  40460.0 203570.0 41165.0 204915.0 ;
      RECT  40460.0 206260.0 41165.0 204915.0 ;
      RECT  41165.0 34100.0 41870.0 35445.0 ;
      RECT  41165.0 36790.0 41870.0 35445.0 ;
      RECT  41165.0 36790.0 41870.0 38135.0 ;
      RECT  41165.0 39480.0 41870.0 38135.0 ;
      RECT  41165.0 39480.0 41870.0 40825.0 ;
      RECT  41165.0 42170.0 41870.0 40825.0 ;
      RECT  41165.0 42170.0 41870.0 43515.0 ;
      RECT  41165.0 44860.0 41870.0 43515.0 ;
      RECT  41165.0 44860.0 41870.0 46205.0 ;
      RECT  41165.0 47550.0 41870.0 46205.0 ;
      RECT  41165.0 47550.0 41870.0 48895.0 ;
      RECT  41165.0 50240.0 41870.0 48895.0 ;
      RECT  41165.0 50240.0 41870.0 51585.0 ;
      RECT  41165.0 52930.0 41870.0 51585.0 ;
      RECT  41165.0 52930.0 41870.0 54275.0 ;
      RECT  41165.0 55620.0 41870.0 54275.0 ;
      RECT  41165.0 55620.0 41870.0 56965.0 ;
      RECT  41165.0 58310.0 41870.0 56965.0 ;
      RECT  41165.0 58310.0 41870.0 59655.0 ;
      RECT  41165.0 61000.0 41870.0 59655.0 ;
      RECT  41165.0 61000.0 41870.0 62345.0 ;
      RECT  41165.0 63690.0 41870.0 62345.0 ;
      RECT  41165.0 63690.0 41870.0 65035.0 ;
      RECT  41165.0 66380.0 41870.0 65035.0 ;
      RECT  41165.0 66380.0 41870.0 67725.0 ;
      RECT  41165.0 69070.0 41870.0 67725.0 ;
      RECT  41165.0 69070.0 41870.0 70415.0 ;
      RECT  41165.0 71760.0 41870.0 70415.0 ;
      RECT  41165.0 71760.0 41870.0 73105.0 ;
      RECT  41165.0 74450.0 41870.0 73105.0 ;
      RECT  41165.0 74450.0 41870.0 75795.0 ;
      RECT  41165.0 77140.0 41870.0 75795.0 ;
      RECT  41165.0 77140.0 41870.0 78485.0 ;
      RECT  41165.0 79830.0 41870.0 78485.0 ;
      RECT  41165.0 79830.0 41870.0 81175.0 ;
      RECT  41165.0 82520.0 41870.0 81175.0 ;
      RECT  41165.0 82520.0 41870.0 83865.0 ;
      RECT  41165.0 85210.0 41870.0 83865.0 ;
      RECT  41165.0 85210.0 41870.0 86555.0 ;
      RECT  41165.0 87900.0 41870.0 86555.0 ;
      RECT  41165.0 87900.0 41870.0 89245.0 ;
      RECT  41165.0 90590.0 41870.0 89245.0 ;
      RECT  41165.0 90590.0 41870.0 91935.0 ;
      RECT  41165.0 93280.0 41870.0 91935.0 ;
      RECT  41165.0 93280.0 41870.0 94625.0 ;
      RECT  41165.0 95970.0 41870.0 94625.0 ;
      RECT  41165.0 95970.0 41870.0 97315.0 ;
      RECT  41165.0 98660.0 41870.0 97315.0 ;
      RECT  41165.0 98660.0 41870.0 100005.0 ;
      RECT  41165.0 101350.0 41870.0 100005.0 ;
      RECT  41165.0 101350.0 41870.0 102695.0 ;
      RECT  41165.0 104040.0 41870.0 102695.0 ;
      RECT  41165.0 104040.0 41870.0 105385.0 ;
      RECT  41165.0 106730.0 41870.0 105385.0 ;
      RECT  41165.0 106730.0 41870.0 108075.0 ;
      RECT  41165.0 109420.0 41870.0 108075.0 ;
      RECT  41165.0 109420.0 41870.0 110765.0 ;
      RECT  41165.0 112110.0 41870.0 110765.0 ;
      RECT  41165.0 112110.0 41870.0 113455.0 ;
      RECT  41165.0 114800.0 41870.0 113455.0 ;
      RECT  41165.0 114800.0 41870.0 116145.0 ;
      RECT  41165.0 117490.0 41870.0 116145.0 ;
      RECT  41165.0 117490.0 41870.0 118835.0 ;
      RECT  41165.0 120180.0 41870.0 118835.0 ;
      RECT  41165.0 120180.0 41870.0 121525.0 ;
      RECT  41165.0 122870.0 41870.0 121525.0 ;
      RECT  41165.0 122870.0 41870.0 124215.0 ;
      RECT  41165.0 125560.0 41870.0 124215.0 ;
      RECT  41165.0 125560.0 41870.0 126905.0 ;
      RECT  41165.0 128250.0 41870.0 126905.0 ;
      RECT  41165.0 128250.0 41870.0 129595.0 ;
      RECT  41165.0 130940.0 41870.0 129595.0 ;
      RECT  41165.0 130940.0 41870.0 132285.0 ;
      RECT  41165.0 133630.0 41870.0 132285.0 ;
      RECT  41165.0 133630.0 41870.0 134975.0 ;
      RECT  41165.0 136320.0 41870.0 134975.0 ;
      RECT  41165.0 136320.0 41870.0 137665.0 ;
      RECT  41165.0 139010.0 41870.0 137665.0 ;
      RECT  41165.0 139010.0 41870.0 140355.0 ;
      RECT  41165.0 141700.0 41870.0 140355.0 ;
      RECT  41165.0 141700.0 41870.0 143045.0 ;
      RECT  41165.0 144390.0 41870.0 143045.0 ;
      RECT  41165.0 144390.0 41870.0 145735.0 ;
      RECT  41165.0 147080.0 41870.0 145735.0 ;
      RECT  41165.0 147080.0 41870.0 148425.0 ;
      RECT  41165.0 149770.0 41870.0 148425.0 ;
      RECT  41165.0 149770.0 41870.0 151115.0 ;
      RECT  41165.0 152460.0 41870.0 151115.0 ;
      RECT  41165.0 152460.0 41870.0 153805.0 ;
      RECT  41165.0 155150.0 41870.0 153805.0 ;
      RECT  41165.0 155150.0 41870.0 156495.0 ;
      RECT  41165.0 157840.0 41870.0 156495.0 ;
      RECT  41165.0 157840.0 41870.0 159185.0 ;
      RECT  41165.0 160530.0 41870.0 159185.0 ;
      RECT  41165.0 160530.0 41870.0 161875.0 ;
      RECT  41165.0 163220.0 41870.0 161875.0 ;
      RECT  41165.0 163220.0 41870.0 164565.0 ;
      RECT  41165.0 165910.0 41870.0 164565.0 ;
      RECT  41165.0 165910.0 41870.0 167255.0 ;
      RECT  41165.0 168600.0 41870.0 167255.0 ;
      RECT  41165.0 168600.0 41870.0 169945.0 ;
      RECT  41165.0 171290.0 41870.0 169945.0 ;
      RECT  41165.0 171290.0 41870.0 172635.0 ;
      RECT  41165.0 173980.0 41870.0 172635.0 ;
      RECT  41165.0 173980.0 41870.0 175325.0 ;
      RECT  41165.0 176670.0 41870.0 175325.0 ;
      RECT  41165.0 176670.0 41870.0 178015.0 ;
      RECT  41165.0 179360.0 41870.0 178015.0 ;
      RECT  41165.0 179360.0 41870.0 180705.0 ;
      RECT  41165.0 182050.0 41870.0 180705.0 ;
      RECT  41165.0 182050.0 41870.0 183395.0 ;
      RECT  41165.0 184740.0 41870.0 183395.0 ;
      RECT  41165.0 184740.0 41870.0 186085.0 ;
      RECT  41165.0 187430.0 41870.0 186085.0 ;
      RECT  41165.0 187430.0 41870.0 188775.0 ;
      RECT  41165.0 190120.0 41870.0 188775.0 ;
      RECT  41165.0 190120.0 41870.0 191465.0 ;
      RECT  41165.0 192810.0 41870.0 191465.0 ;
      RECT  41165.0 192810.0 41870.0 194155.0 ;
      RECT  41165.0 195500.0 41870.0 194155.0 ;
      RECT  41165.0 195500.0 41870.0 196845.0 ;
      RECT  41165.0 198190.0 41870.0 196845.0 ;
      RECT  41165.0 198190.0 41870.0 199535.0 ;
      RECT  41165.0 200880.0 41870.0 199535.0 ;
      RECT  41165.0 200880.0 41870.0 202225.0 ;
      RECT  41165.0 203570.0 41870.0 202225.0 ;
      RECT  41165.0 203570.0 41870.0 204915.0 ;
      RECT  41165.0 206260.0 41870.0 204915.0 ;
      RECT  41870.0 34100.0 42575.0 35445.0 ;
      RECT  41870.0 36790.0 42575.0 35445.0 ;
      RECT  41870.0 36790.0 42575.0 38135.0 ;
      RECT  41870.0 39480.0 42575.0 38135.0 ;
      RECT  41870.0 39480.0 42575.0 40825.0 ;
      RECT  41870.0 42170.0 42575.0 40825.0 ;
      RECT  41870.0 42170.0 42575.0 43515.0 ;
      RECT  41870.0 44860.0 42575.0 43515.0 ;
      RECT  41870.0 44860.0 42575.0 46205.0 ;
      RECT  41870.0 47550.0 42575.0 46205.0 ;
      RECT  41870.0 47550.0 42575.0 48895.0 ;
      RECT  41870.0 50240.0 42575.0 48895.0 ;
      RECT  41870.0 50240.0 42575.0 51585.0 ;
      RECT  41870.0 52930.0 42575.0 51585.0 ;
      RECT  41870.0 52930.0 42575.0 54275.0 ;
      RECT  41870.0 55620.0 42575.0 54275.0 ;
      RECT  41870.0 55620.0 42575.0 56965.0 ;
      RECT  41870.0 58310.0 42575.0 56965.0 ;
      RECT  41870.0 58310.0 42575.0 59655.0 ;
      RECT  41870.0 61000.0 42575.0 59655.0 ;
      RECT  41870.0 61000.0 42575.0 62345.0 ;
      RECT  41870.0 63690.0 42575.0 62345.0 ;
      RECT  41870.0 63690.0 42575.0 65035.0 ;
      RECT  41870.0 66380.0 42575.0 65035.0 ;
      RECT  41870.0 66380.0 42575.0 67725.0 ;
      RECT  41870.0 69070.0 42575.0 67725.0 ;
      RECT  41870.0 69070.0 42575.0 70415.0 ;
      RECT  41870.0 71760.0 42575.0 70415.0 ;
      RECT  41870.0 71760.0 42575.0 73105.0 ;
      RECT  41870.0 74450.0 42575.0 73105.0 ;
      RECT  41870.0 74450.0 42575.0 75795.0 ;
      RECT  41870.0 77140.0 42575.0 75795.0 ;
      RECT  41870.0 77140.0 42575.0 78485.0 ;
      RECT  41870.0 79830.0 42575.0 78485.0 ;
      RECT  41870.0 79830.0 42575.0 81175.0 ;
      RECT  41870.0 82520.0 42575.0 81175.0 ;
      RECT  41870.0 82520.0 42575.0 83865.0 ;
      RECT  41870.0 85210.0 42575.0 83865.0 ;
      RECT  41870.0 85210.0 42575.0 86555.0 ;
      RECT  41870.0 87900.0 42575.0 86555.0 ;
      RECT  41870.0 87900.0 42575.0 89245.0 ;
      RECT  41870.0 90590.0 42575.0 89245.0 ;
      RECT  41870.0 90590.0 42575.0 91935.0 ;
      RECT  41870.0 93280.0 42575.0 91935.0 ;
      RECT  41870.0 93280.0 42575.0 94625.0 ;
      RECT  41870.0 95970.0 42575.0 94625.0 ;
      RECT  41870.0 95970.0 42575.0 97315.0 ;
      RECT  41870.0 98660.0 42575.0 97315.0 ;
      RECT  41870.0 98660.0 42575.0 100005.0 ;
      RECT  41870.0 101350.0 42575.0 100005.0 ;
      RECT  41870.0 101350.0 42575.0 102695.0 ;
      RECT  41870.0 104040.0 42575.0 102695.0 ;
      RECT  41870.0 104040.0 42575.0 105385.0 ;
      RECT  41870.0 106730.0 42575.0 105385.0 ;
      RECT  41870.0 106730.0 42575.0 108075.0 ;
      RECT  41870.0 109420.0 42575.0 108075.0 ;
      RECT  41870.0 109420.0 42575.0 110765.0 ;
      RECT  41870.0 112110.0 42575.0 110765.0 ;
      RECT  41870.0 112110.0 42575.0 113455.0 ;
      RECT  41870.0 114800.0 42575.0 113455.0 ;
      RECT  41870.0 114800.0 42575.0 116145.0 ;
      RECT  41870.0 117490.0 42575.0 116145.0 ;
      RECT  41870.0 117490.0 42575.0 118835.0 ;
      RECT  41870.0 120180.0 42575.0 118835.0 ;
      RECT  41870.0 120180.0 42575.0 121525.0 ;
      RECT  41870.0 122870.0 42575.0 121525.0 ;
      RECT  41870.0 122870.0 42575.0 124215.0 ;
      RECT  41870.0 125560.0 42575.0 124215.0 ;
      RECT  41870.0 125560.0 42575.0 126905.0 ;
      RECT  41870.0 128250.0 42575.0 126905.0 ;
      RECT  41870.0 128250.0 42575.0 129595.0 ;
      RECT  41870.0 130940.0 42575.0 129595.0 ;
      RECT  41870.0 130940.0 42575.0 132285.0 ;
      RECT  41870.0 133630.0 42575.0 132285.0 ;
      RECT  41870.0 133630.0 42575.0 134975.0 ;
      RECT  41870.0 136320.0 42575.0 134975.0 ;
      RECT  41870.0 136320.0 42575.0 137665.0 ;
      RECT  41870.0 139010.0 42575.0 137665.0 ;
      RECT  41870.0 139010.0 42575.0 140355.0 ;
      RECT  41870.0 141700.0 42575.0 140355.0 ;
      RECT  41870.0 141700.0 42575.0 143045.0 ;
      RECT  41870.0 144390.0 42575.0 143045.0 ;
      RECT  41870.0 144390.0 42575.0 145735.0 ;
      RECT  41870.0 147080.0 42575.0 145735.0 ;
      RECT  41870.0 147080.0 42575.0 148425.0 ;
      RECT  41870.0 149770.0 42575.0 148425.0 ;
      RECT  41870.0 149770.0 42575.0 151115.0 ;
      RECT  41870.0 152460.0 42575.0 151115.0 ;
      RECT  41870.0 152460.0 42575.0 153805.0 ;
      RECT  41870.0 155150.0 42575.0 153805.0 ;
      RECT  41870.0 155150.0 42575.0 156495.0 ;
      RECT  41870.0 157840.0 42575.0 156495.0 ;
      RECT  41870.0 157840.0 42575.0 159185.0 ;
      RECT  41870.0 160530.0 42575.0 159185.0 ;
      RECT  41870.0 160530.0 42575.0 161875.0 ;
      RECT  41870.0 163220.0 42575.0 161875.0 ;
      RECT  41870.0 163220.0 42575.0 164565.0 ;
      RECT  41870.0 165910.0 42575.0 164565.0 ;
      RECT  41870.0 165910.0 42575.0 167255.0 ;
      RECT  41870.0 168600.0 42575.0 167255.0 ;
      RECT  41870.0 168600.0 42575.0 169945.0 ;
      RECT  41870.0 171290.0 42575.0 169945.0 ;
      RECT  41870.0 171290.0 42575.0 172635.0 ;
      RECT  41870.0 173980.0 42575.0 172635.0 ;
      RECT  41870.0 173980.0 42575.0 175325.0 ;
      RECT  41870.0 176670.0 42575.0 175325.0 ;
      RECT  41870.0 176670.0 42575.0 178015.0 ;
      RECT  41870.0 179360.0 42575.0 178015.0 ;
      RECT  41870.0 179360.0 42575.0 180705.0 ;
      RECT  41870.0 182050.0 42575.0 180705.0 ;
      RECT  41870.0 182050.0 42575.0 183395.0 ;
      RECT  41870.0 184740.0 42575.0 183395.0 ;
      RECT  41870.0 184740.0 42575.0 186085.0 ;
      RECT  41870.0 187430.0 42575.0 186085.0 ;
      RECT  41870.0 187430.0 42575.0 188775.0 ;
      RECT  41870.0 190120.0 42575.0 188775.0 ;
      RECT  41870.0 190120.0 42575.0 191465.0 ;
      RECT  41870.0 192810.0 42575.0 191465.0 ;
      RECT  41870.0 192810.0 42575.0 194155.0 ;
      RECT  41870.0 195500.0 42575.0 194155.0 ;
      RECT  41870.0 195500.0 42575.0 196845.0 ;
      RECT  41870.0 198190.0 42575.0 196845.0 ;
      RECT  41870.0 198190.0 42575.0 199535.0 ;
      RECT  41870.0 200880.0 42575.0 199535.0 ;
      RECT  41870.0 200880.0 42575.0 202225.0 ;
      RECT  41870.0 203570.0 42575.0 202225.0 ;
      RECT  41870.0 203570.0 42575.0 204915.0 ;
      RECT  41870.0 206260.0 42575.0 204915.0 ;
      RECT  42575.0 34100.0 43280.0 35445.0 ;
      RECT  42575.0 36790.0 43280.0 35445.0 ;
      RECT  42575.0 36790.0 43280.0 38135.0 ;
      RECT  42575.0 39480.0 43280.0 38135.0 ;
      RECT  42575.0 39480.0 43280.0 40825.0 ;
      RECT  42575.0 42170.0 43280.0 40825.0 ;
      RECT  42575.0 42170.0 43280.0 43515.0 ;
      RECT  42575.0 44860.0 43280.0 43515.0 ;
      RECT  42575.0 44860.0 43280.0 46205.0 ;
      RECT  42575.0 47550.0 43280.0 46205.0 ;
      RECT  42575.0 47550.0 43280.0 48895.0 ;
      RECT  42575.0 50240.0 43280.0 48895.0 ;
      RECT  42575.0 50240.0 43280.0 51585.0 ;
      RECT  42575.0 52930.0 43280.0 51585.0 ;
      RECT  42575.0 52930.0 43280.0 54275.0 ;
      RECT  42575.0 55620.0 43280.0 54275.0 ;
      RECT  42575.0 55620.0 43280.0 56965.0 ;
      RECT  42575.0 58310.0 43280.0 56965.0 ;
      RECT  42575.0 58310.0 43280.0 59655.0 ;
      RECT  42575.0 61000.0 43280.0 59655.0 ;
      RECT  42575.0 61000.0 43280.0 62345.0 ;
      RECT  42575.0 63690.0 43280.0 62345.0 ;
      RECT  42575.0 63690.0 43280.0 65035.0 ;
      RECT  42575.0 66380.0 43280.0 65035.0 ;
      RECT  42575.0 66380.0 43280.0 67725.0 ;
      RECT  42575.0 69070.0 43280.0 67725.0 ;
      RECT  42575.0 69070.0 43280.0 70415.0 ;
      RECT  42575.0 71760.0 43280.0 70415.0 ;
      RECT  42575.0 71760.0 43280.0 73105.0 ;
      RECT  42575.0 74450.0 43280.0 73105.0 ;
      RECT  42575.0 74450.0 43280.0 75795.0 ;
      RECT  42575.0 77140.0 43280.0 75795.0 ;
      RECT  42575.0 77140.0 43280.0 78485.0 ;
      RECT  42575.0 79830.0 43280.0 78485.0 ;
      RECT  42575.0 79830.0 43280.0 81175.0 ;
      RECT  42575.0 82520.0 43280.0 81175.0 ;
      RECT  42575.0 82520.0 43280.0 83865.0 ;
      RECT  42575.0 85210.0 43280.0 83865.0 ;
      RECT  42575.0 85210.0 43280.0 86555.0 ;
      RECT  42575.0 87900.0 43280.0 86555.0 ;
      RECT  42575.0 87900.0 43280.0 89245.0 ;
      RECT  42575.0 90590.0 43280.0 89245.0 ;
      RECT  42575.0 90590.0 43280.0 91935.0 ;
      RECT  42575.0 93280.0 43280.0 91935.0 ;
      RECT  42575.0 93280.0 43280.0 94625.0 ;
      RECT  42575.0 95970.0 43280.0 94625.0 ;
      RECT  42575.0 95970.0 43280.0 97315.0 ;
      RECT  42575.0 98660.0 43280.0 97315.0 ;
      RECT  42575.0 98660.0 43280.0 100005.0 ;
      RECT  42575.0 101350.0 43280.0 100005.0 ;
      RECT  42575.0 101350.0 43280.0 102695.0 ;
      RECT  42575.0 104040.0 43280.0 102695.0 ;
      RECT  42575.0 104040.0 43280.0 105385.0 ;
      RECT  42575.0 106730.0 43280.0 105385.0 ;
      RECT  42575.0 106730.0 43280.0 108075.0 ;
      RECT  42575.0 109420.0 43280.0 108075.0 ;
      RECT  42575.0 109420.0 43280.0 110765.0 ;
      RECT  42575.0 112110.0 43280.0 110765.0 ;
      RECT  42575.0 112110.0 43280.0 113455.0 ;
      RECT  42575.0 114800.0 43280.0 113455.0 ;
      RECT  42575.0 114800.0 43280.0 116145.0 ;
      RECT  42575.0 117490.0 43280.0 116145.0 ;
      RECT  42575.0 117490.0 43280.0 118835.0 ;
      RECT  42575.0 120180.0 43280.0 118835.0 ;
      RECT  42575.0 120180.0 43280.0 121525.0 ;
      RECT  42575.0 122870.0 43280.0 121525.0 ;
      RECT  42575.0 122870.0 43280.0 124215.0 ;
      RECT  42575.0 125560.0 43280.0 124215.0 ;
      RECT  42575.0 125560.0 43280.0 126905.0 ;
      RECT  42575.0 128250.0 43280.0 126905.0 ;
      RECT  42575.0 128250.0 43280.0 129595.0 ;
      RECT  42575.0 130940.0 43280.0 129595.0 ;
      RECT  42575.0 130940.0 43280.0 132285.0 ;
      RECT  42575.0 133630.0 43280.0 132285.0 ;
      RECT  42575.0 133630.0 43280.0 134975.0 ;
      RECT  42575.0 136320.0 43280.0 134975.0 ;
      RECT  42575.0 136320.0 43280.0 137665.0 ;
      RECT  42575.0 139010.0 43280.0 137665.0 ;
      RECT  42575.0 139010.0 43280.0 140355.0 ;
      RECT  42575.0 141700.0 43280.0 140355.0 ;
      RECT  42575.0 141700.0 43280.0 143045.0 ;
      RECT  42575.0 144390.0 43280.0 143045.0 ;
      RECT  42575.0 144390.0 43280.0 145735.0 ;
      RECT  42575.0 147080.0 43280.0 145735.0 ;
      RECT  42575.0 147080.0 43280.0 148425.0 ;
      RECT  42575.0 149770.0 43280.0 148425.0 ;
      RECT  42575.0 149770.0 43280.0 151115.0 ;
      RECT  42575.0 152460.0 43280.0 151115.0 ;
      RECT  42575.0 152460.0 43280.0 153805.0 ;
      RECT  42575.0 155150.0 43280.0 153805.0 ;
      RECT  42575.0 155150.0 43280.0 156495.0 ;
      RECT  42575.0 157840.0 43280.0 156495.0 ;
      RECT  42575.0 157840.0 43280.0 159185.0 ;
      RECT  42575.0 160530.0 43280.0 159185.0 ;
      RECT  42575.0 160530.0 43280.0 161875.0 ;
      RECT  42575.0 163220.0 43280.0 161875.0 ;
      RECT  42575.0 163220.0 43280.0 164565.0 ;
      RECT  42575.0 165910.0 43280.0 164565.0 ;
      RECT  42575.0 165910.0 43280.0 167255.0 ;
      RECT  42575.0 168600.0 43280.0 167255.0 ;
      RECT  42575.0 168600.0 43280.0 169945.0 ;
      RECT  42575.0 171290.0 43280.0 169945.0 ;
      RECT  42575.0 171290.0 43280.0 172635.0 ;
      RECT  42575.0 173980.0 43280.0 172635.0 ;
      RECT  42575.0 173980.0 43280.0 175325.0 ;
      RECT  42575.0 176670.0 43280.0 175325.0 ;
      RECT  42575.0 176670.0 43280.0 178015.0 ;
      RECT  42575.0 179360.0 43280.0 178015.0 ;
      RECT  42575.0 179360.0 43280.0 180705.0 ;
      RECT  42575.0 182050.0 43280.0 180705.0 ;
      RECT  42575.0 182050.0 43280.0 183395.0 ;
      RECT  42575.0 184740.0 43280.0 183395.0 ;
      RECT  42575.0 184740.0 43280.0 186085.0 ;
      RECT  42575.0 187430.0 43280.0 186085.0 ;
      RECT  42575.0 187430.0 43280.0 188775.0 ;
      RECT  42575.0 190120.0 43280.0 188775.0 ;
      RECT  42575.0 190120.0 43280.0 191465.0 ;
      RECT  42575.0 192810.0 43280.0 191465.0 ;
      RECT  42575.0 192810.0 43280.0 194155.0 ;
      RECT  42575.0 195500.0 43280.0 194155.0 ;
      RECT  42575.0 195500.0 43280.0 196845.0 ;
      RECT  42575.0 198190.0 43280.0 196845.0 ;
      RECT  42575.0 198190.0 43280.0 199535.0 ;
      RECT  42575.0 200880.0 43280.0 199535.0 ;
      RECT  42575.0 200880.0 43280.0 202225.0 ;
      RECT  42575.0 203570.0 43280.0 202225.0 ;
      RECT  42575.0 203570.0 43280.0 204915.0 ;
      RECT  42575.0 206260.0 43280.0 204915.0 ;
      RECT  43280.0 34100.0 43985.0 35445.0 ;
      RECT  43280.0 36790.0 43985.0 35445.0 ;
      RECT  43280.0 36790.0 43985.0 38135.0 ;
      RECT  43280.0 39480.0 43985.0 38135.0 ;
      RECT  43280.0 39480.0 43985.0 40825.0 ;
      RECT  43280.0 42170.0 43985.0 40825.0 ;
      RECT  43280.0 42170.0 43985.0 43515.0 ;
      RECT  43280.0 44860.0 43985.0 43515.0 ;
      RECT  43280.0 44860.0 43985.0 46205.0 ;
      RECT  43280.0 47550.0 43985.0 46205.0 ;
      RECT  43280.0 47550.0 43985.0 48895.0 ;
      RECT  43280.0 50240.0 43985.0 48895.0 ;
      RECT  43280.0 50240.0 43985.0 51585.0 ;
      RECT  43280.0 52930.0 43985.0 51585.0 ;
      RECT  43280.0 52930.0 43985.0 54275.0 ;
      RECT  43280.0 55620.0 43985.0 54275.0 ;
      RECT  43280.0 55620.0 43985.0 56965.0 ;
      RECT  43280.0 58310.0 43985.0 56965.0 ;
      RECT  43280.0 58310.0 43985.0 59655.0 ;
      RECT  43280.0 61000.0 43985.0 59655.0 ;
      RECT  43280.0 61000.0 43985.0 62345.0 ;
      RECT  43280.0 63690.0 43985.0 62345.0 ;
      RECT  43280.0 63690.0 43985.0 65035.0 ;
      RECT  43280.0 66380.0 43985.0 65035.0 ;
      RECT  43280.0 66380.0 43985.0 67725.0 ;
      RECT  43280.0 69070.0 43985.0 67725.0 ;
      RECT  43280.0 69070.0 43985.0 70415.0 ;
      RECT  43280.0 71760.0 43985.0 70415.0 ;
      RECT  43280.0 71760.0 43985.0 73105.0 ;
      RECT  43280.0 74450.0 43985.0 73105.0 ;
      RECT  43280.0 74450.0 43985.0 75795.0 ;
      RECT  43280.0 77140.0 43985.0 75795.0 ;
      RECT  43280.0 77140.0 43985.0 78485.0 ;
      RECT  43280.0 79830.0 43985.0 78485.0 ;
      RECT  43280.0 79830.0 43985.0 81175.0 ;
      RECT  43280.0 82520.0 43985.0 81175.0 ;
      RECT  43280.0 82520.0 43985.0 83865.0 ;
      RECT  43280.0 85210.0 43985.0 83865.0 ;
      RECT  43280.0 85210.0 43985.0 86555.0 ;
      RECT  43280.0 87900.0 43985.0 86555.0 ;
      RECT  43280.0 87900.0 43985.0 89245.0 ;
      RECT  43280.0 90590.0 43985.0 89245.0 ;
      RECT  43280.0 90590.0 43985.0 91935.0 ;
      RECT  43280.0 93280.0 43985.0 91935.0 ;
      RECT  43280.0 93280.0 43985.0 94625.0 ;
      RECT  43280.0 95970.0 43985.0 94625.0 ;
      RECT  43280.0 95970.0 43985.0 97315.0 ;
      RECT  43280.0 98660.0 43985.0 97315.0 ;
      RECT  43280.0 98660.0 43985.0 100005.0 ;
      RECT  43280.0 101350.0 43985.0 100005.0 ;
      RECT  43280.0 101350.0 43985.0 102695.0 ;
      RECT  43280.0 104040.0 43985.0 102695.0 ;
      RECT  43280.0 104040.0 43985.0 105385.0 ;
      RECT  43280.0 106730.0 43985.0 105385.0 ;
      RECT  43280.0 106730.0 43985.0 108075.0 ;
      RECT  43280.0 109420.0 43985.0 108075.0 ;
      RECT  43280.0 109420.0 43985.0 110765.0 ;
      RECT  43280.0 112110.0 43985.0 110765.0 ;
      RECT  43280.0 112110.0 43985.0 113455.0 ;
      RECT  43280.0 114800.0 43985.0 113455.0 ;
      RECT  43280.0 114800.0 43985.0 116145.0 ;
      RECT  43280.0 117490.0 43985.0 116145.0 ;
      RECT  43280.0 117490.0 43985.0 118835.0 ;
      RECT  43280.0 120180.0 43985.0 118835.0 ;
      RECT  43280.0 120180.0 43985.0 121525.0 ;
      RECT  43280.0 122870.0 43985.0 121525.0 ;
      RECT  43280.0 122870.0 43985.0 124215.0 ;
      RECT  43280.0 125560.0 43985.0 124215.0 ;
      RECT  43280.0 125560.0 43985.0 126905.0 ;
      RECT  43280.0 128250.0 43985.0 126905.0 ;
      RECT  43280.0 128250.0 43985.0 129595.0 ;
      RECT  43280.0 130940.0 43985.0 129595.0 ;
      RECT  43280.0 130940.0 43985.0 132285.0 ;
      RECT  43280.0 133630.0 43985.0 132285.0 ;
      RECT  43280.0 133630.0 43985.0 134975.0 ;
      RECT  43280.0 136320.0 43985.0 134975.0 ;
      RECT  43280.0 136320.0 43985.0 137665.0 ;
      RECT  43280.0 139010.0 43985.0 137665.0 ;
      RECT  43280.0 139010.0 43985.0 140355.0 ;
      RECT  43280.0 141700.0 43985.0 140355.0 ;
      RECT  43280.0 141700.0 43985.0 143045.0 ;
      RECT  43280.0 144390.0 43985.0 143045.0 ;
      RECT  43280.0 144390.0 43985.0 145735.0 ;
      RECT  43280.0 147080.0 43985.0 145735.0 ;
      RECT  43280.0 147080.0 43985.0 148425.0 ;
      RECT  43280.0 149770.0 43985.0 148425.0 ;
      RECT  43280.0 149770.0 43985.0 151115.0 ;
      RECT  43280.0 152460.0 43985.0 151115.0 ;
      RECT  43280.0 152460.0 43985.0 153805.0 ;
      RECT  43280.0 155150.0 43985.0 153805.0 ;
      RECT  43280.0 155150.0 43985.0 156495.0 ;
      RECT  43280.0 157840.0 43985.0 156495.0 ;
      RECT  43280.0 157840.0 43985.0 159185.0 ;
      RECT  43280.0 160530.0 43985.0 159185.0 ;
      RECT  43280.0 160530.0 43985.0 161875.0 ;
      RECT  43280.0 163220.0 43985.0 161875.0 ;
      RECT  43280.0 163220.0 43985.0 164565.0 ;
      RECT  43280.0 165910.0 43985.0 164565.0 ;
      RECT  43280.0 165910.0 43985.0 167255.0 ;
      RECT  43280.0 168600.0 43985.0 167255.0 ;
      RECT  43280.0 168600.0 43985.0 169945.0 ;
      RECT  43280.0 171290.0 43985.0 169945.0 ;
      RECT  43280.0 171290.0 43985.0 172635.0 ;
      RECT  43280.0 173980.0 43985.0 172635.0 ;
      RECT  43280.0 173980.0 43985.0 175325.0 ;
      RECT  43280.0 176670.0 43985.0 175325.0 ;
      RECT  43280.0 176670.0 43985.0 178015.0 ;
      RECT  43280.0 179360.0 43985.0 178015.0 ;
      RECT  43280.0 179360.0 43985.0 180705.0 ;
      RECT  43280.0 182050.0 43985.0 180705.0 ;
      RECT  43280.0 182050.0 43985.0 183395.0 ;
      RECT  43280.0 184740.0 43985.0 183395.0 ;
      RECT  43280.0 184740.0 43985.0 186085.0 ;
      RECT  43280.0 187430.0 43985.0 186085.0 ;
      RECT  43280.0 187430.0 43985.0 188775.0 ;
      RECT  43280.0 190120.0 43985.0 188775.0 ;
      RECT  43280.0 190120.0 43985.0 191465.0 ;
      RECT  43280.0 192810.0 43985.0 191465.0 ;
      RECT  43280.0 192810.0 43985.0 194155.0 ;
      RECT  43280.0 195500.0 43985.0 194155.0 ;
      RECT  43280.0 195500.0 43985.0 196845.0 ;
      RECT  43280.0 198190.0 43985.0 196845.0 ;
      RECT  43280.0 198190.0 43985.0 199535.0 ;
      RECT  43280.0 200880.0 43985.0 199535.0 ;
      RECT  43280.0 200880.0 43985.0 202225.0 ;
      RECT  43280.0 203570.0 43985.0 202225.0 ;
      RECT  43280.0 203570.0 43985.0 204915.0 ;
      RECT  43280.0 206260.0 43985.0 204915.0 ;
      RECT  43985.0 34100.0 44690.0 35445.0 ;
      RECT  43985.0 36790.0 44690.0 35445.0 ;
      RECT  43985.0 36790.0 44690.0 38135.0 ;
      RECT  43985.0 39480.0 44690.0 38135.0 ;
      RECT  43985.0 39480.0 44690.0 40825.0 ;
      RECT  43985.0 42170.0 44690.0 40825.0 ;
      RECT  43985.0 42170.0 44690.0 43515.0 ;
      RECT  43985.0 44860.0 44690.0 43515.0 ;
      RECT  43985.0 44860.0 44690.0 46205.0 ;
      RECT  43985.0 47550.0 44690.0 46205.0 ;
      RECT  43985.0 47550.0 44690.0 48895.0 ;
      RECT  43985.0 50240.0 44690.0 48895.0 ;
      RECT  43985.0 50240.0 44690.0 51585.0 ;
      RECT  43985.0 52930.0 44690.0 51585.0 ;
      RECT  43985.0 52930.0 44690.0 54275.0 ;
      RECT  43985.0 55620.0 44690.0 54275.0 ;
      RECT  43985.0 55620.0 44690.0 56965.0 ;
      RECT  43985.0 58310.0 44690.0 56965.0 ;
      RECT  43985.0 58310.0 44690.0 59655.0 ;
      RECT  43985.0 61000.0 44690.0 59655.0 ;
      RECT  43985.0 61000.0 44690.0 62345.0 ;
      RECT  43985.0 63690.0 44690.0 62345.0 ;
      RECT  43985.0 63690.0 44690.0 65035.0 ;
      RECT  43985.0 66380.0 44690.0 65035.0 ;
      RECT  43985.0 66380.0 44690.0 67725.0 ;
      RECT  43985.0 69070.0 44690.0 67725.0 ;
      RECT  43985.0 69070.0 44690.0 70415.0 ;
      RECT  43985.0 71760.0 44690.0 70415.0 ;
      RECT  43985.0 71760.0 44690.0 73105.0 ;
      RECT  43985.0 74450.0 44690.0 73105.0 ;
      RECT  43985.0 74450.0 44690.0 75795.0 ;
      RECT  43985.0 77140.0 44690.0 75795.0 ;
      RECT  43985.0 77140.0 44690.0 78485.0 ;
      RECT  43985.0 79830.0 44690.0 78485.0 ;
      RECT  43985.0 79830.0 44690.0 81175.0 ;
      RECT  43985.0 82520.0 44690.0 81175.0 ;
      RECT  43985.0 82520.0 44690.0 83865.0 ;
      RECT  43985.0 85210.0 44690.0 83865.0 ;
      RECT  43985.0 85210.0 44690.0 86555.0 ;
      RECT  43985.0 87900.0 44690.0 86555.0 ;
      RECT  43985.0 87900.0 44690.0 89245.0 ;
      RECT  43985.0 90590.0 44690.0 89245.0 ;
      RECT  43985.0 90590.0 44690.0 91935.0 ;
      RECT  43985.0 93280.0 44690.0 91935.0 ;
      RECT  43985.0 93280.0 44690.0 94625.0 ;
      RECT  43985.0 95970.0 44690.0 94625.0 ;
      RECT  43985.0 95970.0 44690.0 97315.0 ;
      RECT  43985.0 98660.0 44690.0 97315.0 ;
      RECT  43985.0 98660.0 44690.0 100005.0 ;
      RECT  43985.0 101350.0 44690.0 100005.0 ;
      RECT  43985.0 101350.0 44690.0 102695.0 ;
      RECT  43985.0 104040.0 44690.0 102695.0 ;
      RECT  43985.0 104040.0 44690.0 105385.0 ;
      RECT  43985.0 106730.0 44690.0 105385.0 ;
      RECT  43985.0 106730.0 44690.0 108075.0 ;
      RECT  43985.0 109420.0 44690.0 108075.0 ;
      RECT  43985.0 109420.0 44690.0 110765.0 ;
      RECT  43985.0 112110.0 44690.0 110765.0 ;
      RECT  43985.0 112110.0 44690.0 113455.0 ;
      RECT  43985.0 114800.0 44690.0 113455.0 ;
      RECT  43985.0 114800.0 44690.0 116145.0 ;
      RECT  43985.0 117490.0 44690.0 116145.0 ;
      RECT  43985.0 117490.0 44690.0 118835.0 ;
      RECT  43985.0 120180.0 44690.0 118835.0 ;
      RECT  43985.0 120180.0 44690.0 121525.0 ;
      RECT  43985.0 122870.0 44690.0 121525.0 ;
      RECT  43985.0 122870.0 44690.0 124215.0 ;
      RECT  43985.0 125560.0 44690.0 124215.0 ;
      RECT  43985.0 125560.0 44690.0 126905.0 ;
      RECT  43985.0 128250.0 44690.0 126905.0 ;
      RECT  43985.0 128250.0 44690.0 129595.0 ;
      RECT  43985.0 130940.0 44690.0 129595.0 ;
      RECT  43985.0 130940.0 44690.0 132285.0 ;
      RECT  43985.0 133630.0 44690.0 132285.0 ;
      RECT  43985.0 133630.0 44690.0 134975.0 ;
      RECT  43985.0 136320.0 44690.0 134975.0 ;
      RECT  43985.0 136320.0 44690.0 137665.0 ;
      RECT  43985.0 139010.0 44690.0 137665.0 ;
      RECT  43985.0 139010.0 44690.0 140355.0 ;
      RECT  43985.0 141700.0 44690.0 140355.0 ;
      RECT  43985.0 141700.0 44690.0 143045.0 ;
      RECT  43985.0 144390.0 44690.0 143045.0 ;
      RECT  43985.0 144390.0 44690.0 145735.0 ;
      RECT  43985.0 147080.0 44690.0 145735.0 ;
      RECT  43985.0 147080.0 44690.0 148425.0 ;
      RECT  43985.0 149770.0 44690.0 148425.0 ;
      RECT  43985.0 149770.0 44690.0 151115.0 ;
      RECT  43985.0 152460.0 44690.0 151115.0 ;
      RECT  43985.0 152460.0 44690.0 153805.0 ;
      RECT  43985.0 155150.0 44690.0 153805.0 ;
      RECT  43985.0 155150.0 44690.0 156495.0 ;
      RECT  43985.0 157840.0 44690.0 156495.0 ;
      RECT  43985.0 157840.0 44690.0 159185.0 ;
      RECT  43985.0 160530.0 44690.0 159185.0 ;
      RECT  43985.0 160530.0 44690.0 161875.0 ;
      RECT  43985.0 163220.0 44690.0 161875.0 ;
      RECT  43985.0 163220.0 44690.0 164565.0 ;
      RECT  43985.0 165910.0 44690.0 164565.0 ;
      RECT  43985.0 165910.0 44690.0 167255.0 ;
      RECT  43985.0 168600.0 44690.0 167255.0 ;
      RECT  43985.0 168600.0 44690.0 169945.0 ;
      RECT  43985.0 171290.0 44690.0 169945.0 ;
      RECT  43985.0 171290.0 44690.0 172635.0 ;
      RECT  43985.0 173980.0 44690.0 172635.0 ;
      RECT  43985.0 173980.0 44690.0 175325.0 ;
      RECT  43985.0 176670.0 44690.0 175325.0 ;
      RECT  43985.0 176670.0 44690.0 178015.0 ;
      RECT  43985.0 179360.0 44690.0 178015.0 ;
      RECT  43985.0 179360.0 44690.0 180705.0 ;
      RECT  43985.0 182050.0 44690.0 180705.0 ;
      RECT  43985.0 182050.0 44690.0 183395.0 ;
      RECT  43985.0 184740.0 44690.0 183395.0 ;
      RECT  43985.0 184740.0 44690.0 186085.0 ;
      RECT  43985.0 187430.0 44690.0 186085.0 ;
      RECT  43985.0 187430.0 44690.0 188775.0 ;
      RECT  43985.0 190120.0 44690.0 188775.0 ;
      RECT  43985.0 190120.0 44690.0 191465.0 ;
      RECT  43985.0 192810.0 44690.0 191465.0 ;
      RECT  43985.0 192810.0 44690.0 194155.0 ;
      RECT  43985.0 195500.0 44690.0 194155.0 ;
      RECT  43985.0 195500.0 44690.0 196845.0 ;
      RECT  43985.0 198190.0 44690.0 196845.0 ;
      RECT  43985.0 198190.0 44690.0 199535.0 ;
      RECT  43985.0 200880.0 44690.0 199535.0 ;
      RECT  43985.0 200880.0 44690.0 202225.0 ;
      RECT  43985.0 203570.0 44690.0 202225.0 ;
      RECT  43985.0 203570.0 44690.0 204915.0 ;
      RECT  43985.0 206260.0 44690.0 204915.0 ;
      RECT  44690.0 34100.0 45395.0 35445.0 ;
      RECT  44690.0 36790.0 45395.0 35445.0 ;
      RECT  44690.0 36790.0 45395.0 38135.0 ;
      RECT  44690.0 39480.0 45395.0 38135.0 ;
      RECT  44690.0 39480.0 45395.0 40825.0 ;
      RECT  44690.0 42170.0 45395.0 40825.0 ;
      RECT  44690.0 42170.0 45395.0 43515.0 ;
      RECT  44690.0 44860.0 45395.0 43515.0 ;
      RECT  44690.0 44860.0 45395.0 46205.0 ;
      RECT  44690.0 47550.0 45395.0 46205.0 ;
      RECT  44690.0 47550.0 45395.0 48895.0 ;
      RECT  44690.0 50240.0 45395.0 48895.0 ;
      RECT  44690.0 50240.0 45395.0 51585.0 ;
      RECT  44690.0 52930.0 45395.0 51585.0 ;
      RECT  44690.0 52930.0 45395.0 54275.0 ;
      RECT  44690.0 55620.0 45395.0 54275.0 ;
      RECT  44690.0 55620.0 45395.0 56965.0 ;
      RECT  44690.0 58310.0 45395.0 56965.0 ;
      RECT  44690.0 58310.0 45395.0 59655.0 ;
      RECT  44690.0 61000.0 45395.0 59655.0 ;
      RECT  44690.0 61000.0 45395.0 62345.0 ;
      RECT  44690.0 63690.0 45395.0 62345.0 ;
      RECT  44690.0 63690.0 45395.0 65035.0 ;
      RECT  44690.0 66380.0 45395.0 65035.0 ;
      RECT  44690.0 66380.0 45395.0 67725.0 ;
      RECT  44690.0 69070.0 45395.0 67725.0 ;
      RECT  44690.0 69070.0 45395.0 70415.0 ;
      RECT  44690.0 71760.0 45395.0 70415.0 ;
      RECT  44690.0 71760.0 45395.0 73105.0 ;
      RECT  44690.0 74450.0 45395.0 73105.0 ;
      RECT  44690.0 74450.0 45395.0 75795.0 ;
      RECT  44690.0 77140.0 45395.0 75795.0 ;
      RECT  44690.0 77140.0 45395.0 78485.0 ;
      RECT  44690.0 79830.0 45395.0 78485.0 ;
      RECT  44690.0 79830.0 45395.0 81175.0 ;
      RECT  44690.0 82520.0 45395.0 81175.0 ;
      RECT  44690.0 82520.0 45395.0 83865.0 ;
      RECT  44690.0 85210.0 45395.0 83865.0 ;
      RECT  44690.0 85210.0 45395.0 86555.0 ;
      RECT  44690.0 87900.0 45395.0 86555.0 ;
      RECT  44690.0 87900.0 45395.0 89245.0 ;
      RECT  44690.0 90590.0 45395.0 89245.0 ;
      RECT  44690.0 90590.0 45395.0 91935.0 ;
      RECT  44690.0 93280.0 45395.0 91935.0 ;
      RECT  44690.0 93280.0 45395.0 94625.0 ;
      RECT  44690.0 95970.0 45395.0 94625.0 ;
      RECT  44690.0 95970.0 45395.0 97315.0 ;
      RECT  44690.0 98660.0 45395.0 97315.0 ;
      RECT  44690.0 98660.0 45395.0 100005.0 ;
      RECT  44690.0 101350.0 45395.0 100005.0 ;
      RECT  44690.0 101350.0 45395.0 102695.0 ;
      RECT  44690.0 104040.0 45395.0 102695.0 ;
      RECT  44690.0 104040.0 45395.0 105385.0 ;
      RECT  44690.0 106730.0 45395.0 105385.0 ;
      RECT  44690.0 106730.0 45395.0 108075.0 ;
      RECT  44690.0 109420.0 45395.0 108075.0 ;
      RECT  44690.0 109420.0 45395.0 110765.0 ;
      RECT  44690.0 112110.0 45395.0 110765.0 ;
      RECT  44690.0 112110.0 45395.0 113455.0 ;
      RECT  44690.0 114800.0 45395.0 113455.0 ;
      RECT  44690.0 114800.0 45395.0 116145.0 ;
      RECT  44690.0 117490.0 45395.0 116145.0 ;
      RECT  44690.0 117490.0 45395.0 118835.0 ;
      RECT  44690.0 120180.0 45395.0 118835.0 ;
      RECT  44690.0 120180.0 45395.0 121525.0 ;
      RECT  44690.0 122870.0 45395.0 121525.0 ;
      RECT  44690.0 122870.0 45395.0 124215.0 ;
      RECT  44690.0 125560.0 45395.0 124215.0 ;
      RECT  44690.0 125560.0 45395.0 126905.0 ;
      RECT  44690.0 128250.0 45395.0 126905.0 ;
      RECT  44690.0 128250.0 45395.0 129595.0 ;
      RECT  44690.0 130940.0 45395.0 129595.0 ;
      RECT  44690.0 130940.0 45395.0 132285.0 ;
      RECT  44690.0 133630.0 45395.0 132285.0 ;
      RECT  44690.0 133630.0 45395.0 134975.0 ;
      RECT  44690.0 136320.0 45395.0 134975.0 ;
      RECT  44690.0 136320.0 45395.0 137665.0 ;
      RECT  44690.0 139010.0 45395.0 137665.0 ;
      RECT  44690.0 139010.0 45395.0 140355.0 ;
      RECT  44690.0 141700.0 45395.0 140355.0 ;
      RECT  44690.0 141700.0 45395.0 143045.0 ;
      RECT  44690.0 144390.0 45395.0 143045.0 ;
      RECT  44690.0 144390.0 45395.0 145735.0 ;
      RECT  44690.0 147080.0 45395.0 145735.0 ;
      RECT  44690.0 147080.0 45395.0 148425.0 ;
      RECT  44690.0 149770.0 45395.0 148425.0 ;
      RECT  44690.0 149770.0 45395.0 151115.0 ;
      RECT  44690.0 152460.0 45395.0 151115.0 ;
      RECT  44690.0 152460.0 45395.0 153805.0 ;
      RECT  44690.0 155150.0 45395.0 153805.0 ;
      RECT  44690.0 155150.0 45395.0 156495.0 ;
      RECT  44690.0 157840.0 45395.0 156495.0 ;
      RECT  44690.0 157840.0 45395.0 159185.0 ;
      RECT  44690.0 160530.0 45395.0 159185.0 ;
      RECT  44690.0 160530.0 45395.0 161875.0 ;
      RECT  44690.0 163220.0 45395.0 161875.0 ;
      RECT  44690.0 163220.0 45395.0 164565.0 ;
      RECT  44690.0 165910.0 45395.0 164565.0 ;
      RECT  44690.0 165910.0 45395.0 167255.0 ;
      RECT  44690.0 168600.0 45395.0 167255.0 ;
      RECT  44690.0 168600.0 45395.0 169945.0 ;
      RECT  44690.0 171290.0 45395.0 169945.0 ;
      RECT  44690.0 171290.0 45395.0 172635.0 ;
      RECT  44690.0 173980.0 45395.0 172635.0 ;
      RECT  44690.0 173980.0 45395.0 175325.0 ;
      RECT  44690.0 176670.0 45395.0 175325.0 ;
      RECT  44690.0 176670.0 45395.0 178015.0 ;
      RECT  44690.0 179360.0 45395.0 178015.0 ;
      RECT  44690.0 179360.0 45395.0 180705.0 ;
      RECT  44690.0 182050.0 45395.0 180705.0 ;
      RECT  44690.0 182050.0 45395.0 183395.0 ;
      RECT  44690.0 184740.0 45395.0 183395.0 ;
      RECT  44690.0 184740.0 45395.0 186085.0 ;
      RECT  44690.0 187430.0 45395.0 186085.0 ;
      RECT  44690.0 187430.0 45395.0 188775.0 ;
      RECT  44690.0 190120.0 45395.0 188775.0 ;
      RECT  44690.0 190120.0 45395.0 191465.0 ;
      RECT  44690.0 192810.0 45395.0 191465.0 ;
      RECT  44690.0 192810.0 45395.0 194155.0 ;
      RECT  44690.0 195500.0 45395.0 194155.0 ;
      RECT  44690.0 195500.0 45395.0 196845.0 ;
      RECT  44690.0 198190.0 45395.0 196845.0 ;
      RECT  44690.0 198190.0 45395.0 199535.0 ;
      RECT  44690.0 200880.0 45395.0 199535.0 ;
      RECT  44690.0 200880.0 45395.0 202225.0 ;
      RECT  44690.0 203570.0 45395.0 202225.0 ;
      RECT  44690.0 203570.0 45395.0 204915.0 ;
      RECT  44690.0 206260.0 45395.0 204915.0 ;
      RECT  45395.0 34100.0 46100.0 35445.0 ;
      RECT  45395.0 36790.0 46100.0 35445.0 ;
      RECT  45395.0 36790.0 46100.0 38135.0 ;
      RECT  45395.0 39480.0 46100.0 38135.0 ;
      RECT  45395.0 39480.0 46100.0 40825.0 ;
      RECT  45395.0 42170.0 46100.0 40825.0 ;
      RECT  45395.0 42170.0 46100.0 43515.0 ;
      RECT  45395.0 44860.0 46100.0 43515.0 ;
      RECT  45395.0 44860.0 46100.0 46205.0 ;
      RECT  45395.0 47550.0 46100.0 46205.0 ;
      RECT  45395.0 47550.0 46100.0 48895.0 ;
      RECT  45395.0 50240.0 46100.0 48895.0 ;
      RECT  45395.0 50240.0 46100.0 51585.0 ;
      RECT  45395.0 52930.0 46100.0 51585.0 ;
      RECT  45395.0 52930.0 46100.0 54275.0 ;
      RECT  45395.0 55620.0 46100.0 54275.0 ;
      RECT  45395.0 55620.0 46100.0 56965.0 ;
      RECT  45395.0 58310.0 46100.0 56965.0 ;
      RECT  45395.0 58310.0 46100.0 59655.0 ;
      RECT  45395.0 61000.0 46100.0 59655.0 ;
      RECT  45395.0 61000.0 46100.0 62345.0 ;
      RECT  45395.0 63690.0 46100.0 62345.0 ;
      RECT  45395.0 63690.0 46100.0 65035.0 ;
      RECT  45395.0 66380.0 46100.0 65035.0 ;
      RECT  45395.0 66380.0 46100.0 67725.0 ;
      RECT  45395.0 69070.0 46100.0 67725.0 ;
      RECT  45395.0 69070.0 46100.0 70415.0 ;
      RECT  45395.0 71760.0 46100.0 70415.0 ;
      RECT  45395.0 71760.0 46100.0 73105.0 ;
      RECT  45395.0 74450.0 46100.0 73105.0 ;
      RECT  45395.0 74450.0 46100.0 75795.0 ;
      RECT  45395.0 77140.0 46100.0 75795.0 ;
      RECT  45395.0 77140.0 46100.0 78485.0 ;
      RECT  45395.0 79830.0 46100.0 78485.0 ;
      RECT  45395.0 79830.0 46100.0 81175.0 ;
      RECT  45395.0 82520.0 46100.0 81175.0 ;
      RECT  45395.0 82520.0 46100.0 83865.0 ;
      RECT  45395.0 85210.0 46100.0 83865.0 ;
      RECT  45395.0 85210.0 46100.0 86555.0 ;
      RECT  45395.0 87900.0 46100.0 86555.0 ;
      RECT  45395.0 87900.0 46100.0 89245.0 ;
      RECT  45395.0 90590.0 46100.0 89245.0 ;
      RECT  45395.0 90590.0 46100.0 91935.0 ;
      RECT  45395.0 93280.0 46100.0 91935.0 ;
      RECT  45395.0 93280.0 46100.0 94625.0 ;
      RECT  45395.0 95970.0 46100.0 94625.0 ;
      RECT  45395.0 95970.0 46100.0 97315.0 ;
      RECT  45395.0 98660.0 46100.0 97315.0 ;
      RECT  45395.0 98660.0 46100.0 100005.0 ;
      RECT  45395.0 101350.0 46100.0 100005.0 ;
      RECT  45395.0 101350.0 46100.0 102695.0 ;
      RECT  45395.0 104040.0 46100.0 102695.0 ;
      RECT  45395.0 104040.0 46100.0 105385.0 ;
      RECT  45395.0 106730.0 46100.0 105385.0 ;
      RECT  45395.0 106730.0 46100.0 108075.0 ;
      RECT  45395.0 109420.0 46100.0 108075.0 ;
      RECT  45395.0 109420.0 46100.0 110765.0 ;
      RECT  45395.0 112110.0 46100.0 110765.0 ;
      RECT  45395.0 112110.0 46100.0 113455.0 ;
      RECT  45395.0 114800.0 46100.0 113455.0 ;
      RECT  45395.0 114800.0 46100.0 116145.0 ;
      RECT  45395.0 117490.0 46100.0 116145.0 ;
      RECT  45395.0 117490.0 46100.0 118835.0 ;
      RECT  45395.0 120180.0 46100.0 118835.0 ;
      RECT  45395.0 120180.0 46100.0 121525.0 ;
      RECT  45395.0 122870.0 46100.0 121525.0 ;
      RECT  45395.0 122870.0 46100.0 124215.0 ;
      RECT  45395.0 125560.0 46100.0 124215.0 ;
      RECT  45395.0 125560.0 46100.0 126905.0 ;
      RECT  45395.0 128250.0 46100.0 126905.0 ;
      RECT  45395.0 128250.0 46100.0 129595.0 ;
      RECT  45395.0 130940.0 46100.0 129595.0 ;
      RECT  45395.0 130940.0 46100.0 132285.0 ;
      RECT  45395.0 133630.0 46100.0 132285.0 ;
      RECT  45395.0 133630.0 46100.0 134975.0 ;
      RECT  45395.0 136320.0 46100.0 134975.0 ;
      RECT  45395.0 136320.0 46100.0 137665.0 ;
      RECT  45395.0 139010.0 46100.0 137665.0 ;
      RECT  45395.0 139010.0 46100.0 140355.0 ;
      RECT  45395.0 141700.0 46100.0 140355.0 ;
      RECT  45395.0 141700.0 46100.0 143045.0 ;
      RECT  45395.0 144390.0 46100.0 143045.0 ;
      RECT  45395.0 144390.0 46100.0 145735.0 ;
      RECT  45395.0 147080.0 46100.0 145735.0 ;
      RECT  45395.0 147080.0 46100.0 148425.0 ;
      RECT  45395.0 149770.0 46100.0 148425.0 ;
      RECT  45395.0 149770.0 46100.0 151115.0 ;
      RECT  45395.0 152460.0 46100.0 151115.0 ;
      RECT  45395.0 152460.0 46100.0 153805.0 ;
      RECT  45395.0 155150.0 46100.0 153805.0 ;
      RECT  45395.0 155150.0 46100.0 156495.0 ;
      RECT  45395.0 157840.0 46100.0 156495.0 ;
      RECT  45395.0 157840.0 46100.0 159185.0 ;
      RECT  45395.0 160530.0 46100.0 159185.0 ;
      RECT  45395.0 160530.0 46100.0 161875.0 ;
      RECT  45395.0 163220.0 46100.0 161875.0 ;
      RECT  45395.0 163220.0 46100.0 164565.0 ;
      RECT  45395.0 165910.0 46100.0 164565.0 ;
      RECT  45395.0 165910.0 46100.0 167255.0 ;
      RECT  45395.0 168600.0 46100.0 167255.0 ;
      RECT  45395.0 168600.0 46100.0 169945.0 ;
      RECT  45395.0 171290.0 46100.0 169945.0 ;
      RECT  45395.0 171290.0 46100.0 172635.0 ;
      RECT  45395.0 173980.0 46100.0 172635.0 ;
      RECT  45395.0 173980.0 46100.0 175325.0 ;
      RECT  45395.0 176670.0 46100.0 175325.0 ;
      RECT  45395.0 176670.0 46100.0 178015.0 ;
      RECT  45395.0 179360.0 46100.0 178015.0 ;
      RECT  45395.0 179360.0 46100.0 180705.0 ;
      RECT  45395.0 182050.0 46100.0 180705.0 ;
      RECT  45395.0 182050.0 46100.0 183395.0 ;
      RECT  45395.0 184740.0 46100.0 183395.0 ;
      RECT  45395.0 184740.0 46100.0 186085.0 ;
      RECT  45395.0 187430.0 46100.0 186085.0 ;
      RECT  45395.0 187430.0 46100.0 188775.0 ;
      RECT  45395.0 190120.0 46100.0 188775.0 ;
      RECT  45395.0 190120.0 46100.0 191465.0 ;
      RECT  45395.0 192810.0 46100.0 191465.0 ;
      RECT  45395.0 192810.0 46100.0 194155.0 ;
      RECT  45395.0 195500.0 46100.0 194155.0 ;
      RECT  45395.0 195500.0 46100.0 196845.0 ;
      RECT  45395.0 198190.0 46100.0 196845.0 ;
      RECT  45395.0 198190.0 46100.0 199535.0 ;
      RECT  45395.0 200880.0 46100.0 199535.0 ;
      RECT  45395.0 200880.0 46100.0 202225.0 ;
      RECT  45395.0 203570.0 46100.0 202225.0 ;
      RECT  45395.0 203570.0 46100.0 204915.0 ;
      RECT  45395.0 206260.0 46100.0 204915.0 ;
      RECT  46100.0 34100.0 46805.0 35445.0 ;
      RECT  46100.0 36790.0 46805.0 35445.0 ;
      RECT  46100.0 36790.0 46805.0 38135.0 ;
      RECT  46100.0 39480.0 46805.0 38135.0 ;
      RECT  46100.0 39480.0 46805.0 40825.0 ;
      RECT  46100.0 42170.0 46805.0 40825.0 ;
      RECT  46100.0 42170.0 46805.0 43515.0 ;
      RECT  46100.0 44860.0 46805.0 43515.0 ;
      RECT  46100.0 44860.0 46805.0 46205.0 ;
      RECT  46100.0 47550.0 46805.0 46205.0 ;
      RECT  46100.0 47550.0 46805.0 48895.0 ;
      RECT  46100.0 50240.0 46805.0 48895.0 ;
      RECT  46100.0 50240.0 46805.0 51585.0 ;
      RECT  46100.0 52930.0 46805.0 51585.0 ;
      RECT  46100.0 52930.0 46805.0 54275.0 ;
      RECT  46100.0 55620.0 46805.0 54275.0 ;
      RECT  46100.0 55620.0 46805.0 56965.0 ;
      RECT  46100.0 58310.0 46805.0 56965.0 ;
      RECT  46100.0 58310.0 46805.0 59655.0 ;
      RECT  46100.0 61000.0 46805.0 59655.0 ;
      RECT  46100.0 61000.0 46805.0 62345.0 ;
      RECT  46100.0 63690.0 46805.0 62345.0 ;
      RECT  46100.0 63690.0 46805.0 65035.0 ;
      RECT  46100.0 66380.0 46805.0 65035.0 ;
      RECT  46100.0 66380.0 46805.0 67725.0 ;
      RECT  46100.0 69070.0 46805.0 67725.0 ;
      RECT  46100.0 69070.0 46805.0 70415.0 ;
      RECT  46100.0 71760.0 46805.0 70415.0 ;
      RECT  46100.0 71760.0 46805.0 73105.0 ;
      RECT  46100.0 74450.0 46805.0 73105.0 ;
      RECT  46100.0 74450.0 46805.0 75795.0 ;
      RECT  46100.0 77140.0 46805.0 75795.0 ;
      RECT  46100.0 77140.0 46805.0 78485.0 ;
      RECT  46100.0 79830.0 46805.0 78485.0 ;
      RECT  46100.0 79830.0 46805.0 81175.0 ;
      RECT  46100.0 82520.0 46805.0 81175.0 ;
      RECT  46100.0 82520.0 46805.0 83865.0 ;
      RECT  46100.0 85210.0 46805.0 83865.0 ;
      RECT  46100.0 85210.0 46805.0 86555.0 ;
      RECT  46100.0 87900.0 46805.0 86555.0 ;
      RECT  46100.0 87900.0 46805.0 89245.0 ;
      RECT  46100.0 90590.0 46805.0 89245.0 ;
      RECT  46100.0 90590.0 46805.0 91935.0 ;
      RECT  46100.0 93280.0 46805.0 91935.0 ;
      RECT  46100.0 93280.0 46805.0 94625.0 ;
      RECT  46100.0 95970.0 46805.0 94625.0 ;
      RECT  46100.0 95970.0 46805.0 97315.0 ;
      RECT  46100.0 98660.0 46805.0 97315.0 ;
      RECT  46100.0 98660.0 46805.0 100005.0 ;
      RECT  46100.0 101350.0 46805.0 100005.0 ;
      RECT  46100.0 101350.0 46805.0 102695.0 ;
      RECT  46100.0 104040.0 46805.0 102695.0 ;
      RECT  46100.0 104040.0 46805.0 105385.0 ;
      RECT  46100.0 106730.0 46805.0 105385.0 ;
      RECT  46100.0 106730.0 46805.0 108075.0 ;
      RECT  46100.0 109420.0 46805.0 108075.0 ;
      RECT  46100.0 109420.0 46805.0 110765.0 ;
      RECT  46100.0 112110.0 46805.0 110765.0 ;
      RECT  46100.0 112110.0 46805.0 113455.0 ;
      RECT  46100.0 114800.0 46805.0 113455.0 ;
      RECT  46100.0 114800.0 46805.0 116145.0 ;
      RECT  46100.0 117490.0 46805.0 116145.0 ;
      RECT  46100.0 117490.0 46805.0 118835.0 ;
      RECT  46100.0 120180.0 46805.0 118835.0 ;
      RECT  46100.0 120180.0 46805.0 121525.0 ;
      RECT  46100.0 122870.0 46805.0 121525.0 ;
      RECT  46100.0 122870.0 46805.0 124215.0 ;
      RECT  46100.0 125560.0 46805.0 124215.0 ;
      RECT  46100.0 125560.0 46805.0 126905.0 ;
      RECT  46100.0 128250.0 46805.0 126905.0 ;
      RECT  46100.0 128250.0 46805.0 129595.0 ;
      RECT  46100.0 130940.0 46805.0 129595.0 ;
      RECT  46100.0 130940.0 46805.0 132285.0 ;
      RECT  46100.0 133630.0 46805.0 132285.0 ;
      RECT  46100.0 133630.0 46805.0 134975.0 ;
      RECT  46100.0 136320.0 46805.0 134975.0 ;
      RECT  46100.0 136320.0 46805.0 137665.0 ;
      RECT  46100.0 139010.0 46805.0 137665.0 ;
      RECT  46100.0 139010.0 46805.0 140355.0 ;
      RECT  46100.0 141700.0 46805.0 140355.0 ;
      RECT  46100.0 141700.0 46805.0 143045.0 ;
      RECT  46100.0 144390.0 46805.0 143045.0 ;
      RECT  46100.0 144390.0 46805.0 145735.0 ;
      RECT  46100.0 147080.0 46805.0 145735.0 ;
      RECT  46100.0 147080.0 46805.0 148425.0 ;
      RECT  46100.0 149770.0 46805.0 148425.0 ;
      RECT  46100.0 149770.0 46805.0 151115.0 ;
      RECT  46100.0 152460.0 46805.0 151115.0 ;
      RECT  46100.0 152460.0 46805.0 153805.0 ;
      RECT  46100.0 155150.0 46805.0 153805.0 ;
      RECT  46100.0 155150.0 46805.0 156495.0 ;
      RECT  46100.0 157840.0 46805.0 156495.0 ;
      RECT  46100.0 157840.0 46805.0 159185.0 ;
      RECT  46100.0 160530.0 46805.0 159185.0 ;
      RECT  46100.0 160530.0 46805.0 161875.0 ;
      RECT  46100.0 163220.0 46805.0 161875.0 ;
      RECT  46100.0 163220.0 46805.0 164565.0 ;
      RECT  46100.0 165910.0 46805.0 164565.0 ;
      RECT  46100.0 165910.0 46805.0 167255.0 ;
      RECT  46100.0 168600.0 46805.0 167255.0 ;
      RECT  46100.0 168600.0 46805.0 169945.0 ;
      RECT  46100.0 171290.0 46805.0 169945.0 ;
      RECT  46100.0 171290.0 46805.0 172635.0 ;
      RECT  46100.0 173980.0 46805.0 172635.0 ;
      RECT  46100.0 173980.0 46805.0 175325.0 ;
      RECT  46100.0 176670.0 46805.0 175325.0 ;
      RECT  46100.0 176670.0 46805.0 178015.0 ;
      RECT  46100.0 179360.0 46805.0 178015.0 ;
      RECT  46100.0 179360.0 46805.0 180705.0 ;
      RECT  46100.0 182050.0 46805.0 180705.0 ;
      RECT  46100.0 182050.0 46805.0 183395.0 ;
      RECT  46100.0 184740.0 46805.0 183395.0 ;
      RECT  46100.0 184740.0 46805.0 186085.0 ;
      RECT  46100.0 187430.0 46805.0 186085.0 ;
      RECT  46100.0 187430.0 46805.0 188775.0 ;
      RECT  46100.0 190120.0 46805.0 188775.0 ;
      RECT  46100.0 190120.0 46805.0 191465.0 ;
      RECT  46100.0 192810.0 46805.0 191465.0 ;
      RECT  46100.0 192810.0 46805.0 194155.0 ;
      RECT  46100.0 195500.0 46805.0 194155.0 ;
      RECT  46100.0 195500.0 46805.0 196845.0 ;
      RECT  46100.0 198190.0 46805.0 196845.0 ;
      RECT  46100.0 198190.0 46805.0 199535.0 ;
      RECT  46100.0 200880.0 46805.0 199535.0 ;
      RECT  46100.0 200880.0 46805.0 202225.0 ;
      RECT  46100.0 203570.0 46805.0 202225.0 ;
      RECT  46100.0 203570.0 46805.0 204915.0 ;
      RECT  46100.0 206260.0 46805.0 204915.0 ;
      RECT  46805.0 34100.0 47510.0 35445.0 ;
      RECT  46805.0 36790.0 47510.0 35445.0 ;
      RECT  46805.0 36790.0 47510.0 38135.0 ;
      RECT  46805.0 39480.0 47510.0 38135.0 ;
      RECT  46805.0 39480.0 47510.0 40825.0 ;
      RECT  46805.0 42170.0 47510.0 40825.0 ;
      RECT  46805.0 42170.0 47510.0 43515.0 ;
      RECT  46805.0 44860.0 47510.0 43515.0 ;
      RECT  46805.0 44860.0 47510.0 46205.0 ;
      RECT  46805.0 47550.0 47510.0 46205.0 ;
      RECT  46805.0 47550.0 47510.0 48895.0 ;
      RECT  46805.0 50240.0 47510.0 48895.0 ;
      RECT  46805.0 50240.0 47510.0 51585.0 ;
      RECT  46805.0 52930.0 47510.0 51585.0 ;
      RECT  46805.0 52930.0 47510.0 54275.0 ;
      RECT  46805.0 55620.0 47510.0 54275.0 ;
      RECT  46805.0 55620.0 47510.0 56965.0 ;
      RECT  46805.0 58310.0 47510.0 56965.0 ;
      RECT  46805.0 58310.0 47510.0 59655.0 ;
      RECT  46805.0 61000.0 47510.0 59655.0 ;
      RECT  46805.0 61000.0 47510.0 62345.0 ;
      RECT  46805.0 63690.0 47510.0 62345.0 ;
      RECT  46805.0 63690.0 47510.0 65035.0 ;
      RECT  46805.0 66380.0 47510.0 65035.0 ;
      RECT  46805.0 66380.0 47510.0 67725.0 ;
      RECT  46805.0 69070.0 47510.0 67725.0 ;
      RECT  46805.0 69070.0 47510.0 70415.0 ;
      RECT  46805.0 71760.0 47510.0 70415.0 ;
      RECT  46805.0 71760.0 47510.0 73105.0 ;
      RECT  46805.0 74450.0 47510.0 73105.0 ;
      RECT  46805.0 74450.0 47510.0 75795.0 ;
      RECT  46805.0 77140.0 47510.0 75795.0 ;
      RECT  46805.0 77140.0 47510.0 78485.0 ;
      RECT  46805.0 79830.0 47510.0 78485.0 ;
      RECT  46805.0 79830.0 47510.0 81175.0 ;
      RECT  46805.0 82520.0 47510.0 81175.0 ;
      RECT  46805.0 82520.0 47510.0 83865.0 ;
      RECT  46805.0 85210.0 47510.0 83865.0 ;
      RECT  46805.0 85210.0 47510.0 86555.0 ;
      RECT  46805.0 87900.0 47510.0 86555.0 ;
      RECT  46805.0 87900.0 47510.0 89245.0 ;
      RECT  46805.0 90590.0 47510.0 89245.0 ;
      RECT  46805.0 90590.0 47510.0 91935.0 ;
      RECT  46805.0 93280.0 47510.0 91935.0 ;
      RECT  46805.0 93280.0 47510.0 94625.0 ;
      RECT  46805.0 95970.0 47510.0 94625.0 ;
      RECT  46805.0 95970.0 47510.0 97315.0 ;
      RECT  46805.0 98660.0 47510.0 97315.0 ;
      RECT  46805.0 98660.0 47510.0 100005.0 ;
      RECT  46805.0 101350.0 47510.0 100005.0 ;
      RECT  46805.0 101350.0 47510.0 102695.0 ;
      RECT  46805.0 104040.0 47510.0 102695.0 ;
      RECT  46805.0 104040.0 47510.0 105385.0 ;
      RECT  46805.0 106730.0 47510.0 105385.0 ;
      RECT  46805.0 106730.0 47510.0 108075.0 ;
      RECT  46805.0 109420.0 47510.0 108075.0 ;
      RECT  46805.0 109420.0 47510.0 110765.0 ;
      RECT  46805.0 112110.0 47510.0 110765.0 ;
      RECT  46805.0 112110.0 47510.0 113455.0 ;
      RECT  46805.0 114800.0 47510.0 113455.0 ;
      RECT  46805.0 114800.0 47510.0 116145.0 ;
      RECT  46805.0 117490.0 47510.0 116145.0 ;
      RECT  46805.0 117490.0 47510.0 118835.0 ;
      RECT  46805.0 120180.0 47510.0 118835.0 ;
      RECT  46805.0 120180.0 47510.0 121525.0 ;
      RECT  46805.0 122870.0 47510.0 121525.0 ;
      RECT  46805.0 122870.0 47510.0 124215.0 ;
      RECT  46805.0 125560.0 47510.0 124215.0 ;
      RECT  46805.0 125560.0 47510.0 126905.0 ;
      RECT  46805.0 128250.0 47510.0 126905.0 ;
      RECT  46805.0 128250.0 47510.0 129595.0 ;
      RECT  46805.0 130940.0 47510.0 129595.0 ;
      RECT  46805.0 130940.0 47510.0 132285.0 ;
      RECT  46805.0 133630.0 47510.0 132285.0 ;
      RECT  46805.0 133630.0 47510.0 134975.0 ;
      RECT  46805.0 136320.0 47510.0 134975.0 ;
      RECT  46805.0 136320.0 47510.0 137665.0 ;
      RECT  46805.0 139010.0 47510.0 137665.0 ;
      RECT  46805.0 139010.0 47510.0 140355.0 ;
      RECT  46805.0 141700.0 47510.0 140355.0 ;
      RECT  46805.0 141700.0 47510.0 143045.0 ;
      RECT  46805.0 144390.0 47510.0 143045.0 ;
      RECT  46805.0 144390.0 47510.0 145735.0 ;
      RECT  46805.0 147080.0 47510.0 145735.0 ;
      RECT  46805.0 147080.0 47510.0 148425.0 ;
      RECT  46805.0 149770.0 47510.0 148425.0 ;
      RECT  46805.0 149770.0 47510.0 151115.0 ;
      RECT  46805.0 152460.0 47510.0 151115.0 ;
      RECT  46805.0 152460.0 47510.0 153805.0 ;
      RECT  46805.0 155150.0 47510.0 153805.0 ;
      RECT  46805.0 155150.0 47510.0 156495.0 ;
      RECT  46805.0 157840.0 47510.0 156495.0 ;
      RECT  46805.0 157840.0 47510.0 159185.0 ;
      RECT  46805.0 160530.0 47510.0 159185.0 ;
      RECT  46805.0 160530.0 47510.0 161875.0 ;
      RECT  46805.0 163220.0 47510.0 161875.0 ;
      RECT  46805.0 163220.0 47510.0 164565.0 ;
      RECT  46805.0 165910.0 47510.0 164565.0 ;
      RECT  46805.0 165910.0 47510.0 167255.0 ;
      RECT  46805.0 168600.0 47510.0 167255.0 ;
      RECT  46805.0 168600.0 47510.0 169945.0 ;
      RECT  46805.0 171290.0 47510.0 169945.0 ;
      RECT  46805.0 171290.0 47510.0 172635.0 ;
      RECT  46805.0 173980.0 47510.0 172635.0 ;
      RECT  46805.0 173980.0 47510.0 175325.0 ;
      RECT  46805.0 176670.0 47510.0 175325.0 ;
      RECT  46805.0 176670.0 47510.0 178015.0 ;
      RECT  46805.0 179360.0 47510.0 178015.0 ;
      RECT  46805.0 179360.0 47510.0 180705.0 ;
      RECT  46805.0 182050.0 47510.0 180705.0 ;
      RECT  46805.0 182050.0 47510.0 183395.0 ;
      RECT  46805.0 184740.0 47510.0 183395.0 ;
      RECT  46805.0 184740.0 47510.0 186085.0 ;
      RECT  46805.0 187430.0 47510.0 186085.0 ;
      RECT  46805.0 187430.0 47510.0 188775.0 ;
      RECT  46805.0 190120.0 47510.0 188775.0 ;
      RECT  46805.0 190120.0 47510.0 191465.0 ;
      RECT  46805.0 192810.0 47510.0 191465.0 ;
      RECT  46805.0 192810.0 47510.0 194155.0 ;
      RECT  46805.0 195500.0 47510.0 194155.0 ;
      RECT  46805.0 195500.0 47510.0 196845.0 ;
      RECT  46805.0 198190.0 47510.0 196845.0 ;
      RECT  46805.0 198190.0 47510.0 199535.0 ;
      RECT  46805.0 200880.0 47510.0 199535.0 ;
      RECT  46805.0 200880.0 47510.0 202225.0 ;
      RECT  46805.0 203570.0 47510.0 202225.0 ;
      RECT  46805.0 203570.0 47510.0 204915.0 ;
      RECT  46805.0 206260.0 47510.0 204915.0 ;
      RECT  47510.0 34100.0 48215.0 35445.0 ;
      RECT  47510.0 36790.0 48215.0 35445.0 ;
      RECT  47510.0 36790.0 48215.0 38135.0 ;
      RECT  47510.0 39480.0 48215.0 38135.0 ;
      RECT  47510.0 39480.0 48215.0 40825.0 ;
      RECT  47510.0 42170.0 48215.0 40825.0 ;
      RECT  47510.0 42170.0 48215.0 43515.0 ;
      RECT  47510.0 44860.0 48215.0 43515.0 ;
      RECT  47510.0 44860.0 48215.0 46205.0 ;
      RECT  47510.0 47550.0 48215.0 46205.0 ;
      RECT  47510.0 47550.0 48215.0 48895.0 ;
      RECT  47510.0 50240.0 48215.0 48895.0 ;
      RECT  47510.0 50240.0 48215.0 51585.0 ;
      RECT  47510.0 52930.0 48215.0 51585.0 ;
      RECT  47510.0 52930.0 48215.0 54275.0 ;
      RECT  47510.0 55620.0 48215.0 54275.0 ;
      RECT  47510.0 55620.0 48215.0 56965.0 ;
      RECT  47510.0 58310.0 48215.0 56965.0 ;
      RECT  47510.0 58310.0 48215.0 59655.0 ;
      RECT  47510.0 61000.0 48215.0 59655.0 ;
      RECT  47510.0 61000.0 48215.0 62345.0 ;
      RECT  47510.0 63690.0 48215.0 62345.0 ;
      RECT  47510.0 63690.0 48215.0 65035.0 ;
      RECT  47510.0 66380.0 48215.0 65035.0 ;
      RECT  47510.0 66380.0 48215.0 67725.0 ;
      RECT  47510.0 69070.0 48215.0 67725.0 ;
      RECT  47510.0 69070.0 48215.0 70415.0 ;
      RECT  47510.0 71760.0 48215.0 70415.0 ;
      RECT  47510.0 71760.0 48215.0 73105.0 ;
      RECT  47510.0 74450.0 48215.0 73105.0 ;
      RECT  47510.0 74450.0 48215.0 75795.0 ;
      RECT  47510.0 77140.0 48215.0 75795.0 ;
      RECT  47510.0 77140.0 48215.0 78485.0 ;
      RECT  47510.0 79830.0 48215.0 78485.0 ;
      RECT  47510.0 79830.0 48215.0 81175.0 ;
      RECT  47510.0 82520.0 48215.0 81175.0 ;
      RECT  47510.0 82520.0 48215.0 83865.0 ;
      RECT  47510.0 85210.0 48215.0 83865.0 ;
      RECT  47510.0 85210.0 48215.0 86555.0 ;
      RECT  47510.0 87900.0 48215.0 86555.0 ;
      RECT  47510.0 87900.0 48215.0 89245.0 ;
      RECT  47510.0 90590.0 48215.0 89245.0 ;
      RECT  47510.0 90590.0 48215.0 91935.0 ;
      RECT  47510.0 93280.0 48215.0 91935.0 ;
      RECT  47510.0 93280.0 48215.0 94625.0 ;
      RECT  47510.0 95970.0 48215.0 94625.0 ;
      RECT  47510.0 95970.0 48215.0 97315.0 ;
      RECT  47510.0 98660.0 48215.0 97315.0 ;
      RECT  47510.0 98660.0 48215.0 100005.0 ;
      RECT  47510.0 101350.0 48215.0 100005.0 ;
      RECT  47510.0 101350.0 48215.0 102695.0 ;
      RECT  47510.0 104040.0 48215.0 102695.0 ;
      RECT  47510.0 104040.0 48215.0 105385.0 ;
      RECT  47510.0 106730.0 48215.0 105385.0 ;
      RECT  47510.0 106730.0 48215.0 108075.0 ;
      RECT  47510.0 109420.0 48215.0 108075.0 ;
      RECT  47510.0 109420.0 48215.0 110765.0 ;
      RECT  47510.0 112110.0 48215.0 110765.0 ;
      RECT  47510.0 112110.0 48215.0 113455.0 ;
      RECT  47510.0 114800.0 48215.0 113455.0 ;
      RECT  47510.0 114800.0 48215.0 116145.0 ;
      RECT  47510.0 117490.0 48215.0 116145.0 ;
      RECT  47510.0 117490.0 48215.0 118835.0 ;
      RECT  47510.0 120180.0 48215.0 118835.0 ;
      RECT  47510.0 120180.0 48215.0 121525.0 ;
      RECT  47510.0 122870.0 48215.0 121525.0 ;
      RECT  47510.0 122870.0 48215.0 124215.0 ;
      RECT  47510.0 125560.0 48215.0 124215.0 ;
      RECT  47510.0 125560.0 48215.0 126905.0 ;
      RECT  47510.0 128250.0 48215.0 126905.0 ;
      RECT  47510.0 128250.0 48215.0 129595.0 ;
      RECT  47510.0 130940.0 48215.0 129595.0 ;
      RECT  47510.0 130940.0 48215.0 132285.0 ;
      RECT  47510.0 133630.0 48215.0 132285.0 ;
      RECT  47510.0 133630.0 48215.0 134975.0 ;
      RECT  47510.0 136320.0 48215.0 134975.0 ;
      RECT  47510.0 136320.0 48215.0 137665.0 ;
      RECT  47510.0 139010.0 48215.0 137665.0 ;
      RECT  47510.0 139010.0 48215.0 140355.0 ;
      RECT  47510.0 141700.0 48215.0 140355.0 ;
      RECT  47510.0 141700.0 48215.0 143045.0 ;
      RECT  47510.0 144390.0 48215.0 143045.0 ;
      RECT  47510.0 144390.0 48215.0 145735.0 ;
      RECT  47510.0 147080.0 48215.0 145735.0 ;
      RECT  47510.0 147080.0 48215.0 148425.0 ;
      RECT  47510.0 149770.0 48215.0 148425.0 ;
      RECT  47510.0 149770.0 48215.0 151115.0 ;
      RECT  47510.0 152460.0 48215.0 151115.0 ;
      RECT  47510.0 152460.0 48215.0 153805.0 ;
      RECT  47510.0 155150.0 48215.0 153805.0 ;
      RECT  47510.0 155150.0 48215.0 156495.0 ;
      RECT  47510.0 157840.0 48215.0 156495.0 ;
      RECT  47510.0 157840.0 48215.0 159185.0 ;
      RECT  47510.0 160530.0 48215.0 159185.0 ;
      RECT  47510.0 160530.0 48215.0 161875.0 ;
      RECT  47510.0 163220.0 48215.0 161875.0 ;
      RECT  47510.0 163220.0 48215.0 164565.0 ;
      RECT  47510.0 165910.0 48215.0 164565.0 ;
      RECT  47510.0 165910.0 48215.0 167255.0 ;
      RECT  47510.0 168600.0 48215.0 167255.0 ;
      RECT  47510.0 168600.0 48215.0 169945.0 ;
      RECT  47510.0 171290.0 48215.0 169945.0 ;
      RECT  47510.0 171290.0 48215.0 172635.0 ;
      RECT  47510.0 173980.0 48215.0 172635.0 ;
      RECT  47510.0 173980.0 48215.0 175325.0 ;
      RECT  47510.0 176670.0 48215.0 175325.0 ;
      RECT  47510.0 176670.0 48215.0 178015.0 ;
      RECT  47510.0 179360.0 48215.0 178015.0 ;
      RECT  47510.0 179360.0 48215.0 180705.0 ;
      RECT  47510.0 182050.0 48215.0 180705.0 ;
      RECT  47510.0 182050.0 48215.0 183395.0 ;
      RECT  47510.0 184740.0 48215.0 183395.0 ;
      RECT  47510.0 184740.0 48215.0 186085.0 ;
      RECT  47510.0 187430.0 48215.0 186085.0 ;
      RECT  47510.0 187430.0 48215.0 188775.0 ;
      RECT  47510.0 190120.0 48215.0 188775.0 ;
      RECT  47510.0 190120.0 48215.0 191465.0 ;
      RECT  47510.0 192810.0 48215.0 191465.0 ;
      RECT  47510.0 192810.0 48215.0 194155.0 ;
      RECT  47510.0 195500.0 48215.0 194155.0 ;
      RECT  47510.0 195500.0 48215.0 196845.0 ;
      RECT  47510.0 198190.0 48215.0 196845.0 ;
      RECT  47510.0 198190.0 48215.0 199535.0 ;
      RECT  47510.0 200880.0 48215.0 199535.0 ;
      RECT  47510.0 200880.0 48215.0 202225.0 ;
      RECT  47510.0 203570.0 48215.0 202225.0 ;
      RECT  47510.0 203570.0 48215.0 204915.0 ;
      RECT  47510.0 206260.0 48215.0 204915.0 ;
      RECT  48215.0 34100.0 48920.0 35445.0 ;
      RECT  48215.0 36790.0 48920.0 35445.0 ;
      RECT  48215.0 36790.0 48920.0 38135.0 ;
      RECT  48215.0 39480.0 48920.0 38135.0 ;
      RECT  48215.0 39480.0 48920.0 40825.0 ;
      RECT  48215.0 42170.0 48920.0 40825.0 ;
      RECT  48215.0 42170.0 48920.0 43515.0 ;
      RECT  48215.0 44860.0 48920.0 43515.0 ;
      RECT  48215.0 44860.0 48920.0 46205.0 ;
      RECT  48215.0 47550.0 48920.0 46205.0 ;
      RECT  48215.0 47550.0 48920.0 48895.0 ;
      RECT  48215.0 50240.0 48920.0 48895.0 ;
      RECT  48215.0 50240.0 48920.0 51585.0 ;
      RECT  48215.0 52930.0 48920.0 51585.0 ;
      RECT  48215.0 52930.0 48920.0 54275.0 ;
      RECT  48215.0 55620.0 48920.0 54275.0 ;
      RECT  48215.0 55620.0 48920.0 56965.0 ;
      RECT  48215.0 58310.0 48920.0 56965.0 ;
      RECT  48215.0 58310.0 48920.0 59655.0 ;
      RECT  48215.0 61000.0 48920.0 59655.0 ;
      RECT  48215.0 61000.0 48920.0 62345.0 ;
      RECT  48215.0 63690.0 48920.0 62345.0 ;
      RECT  48215.0 63690.0 48920.0 65035.0 ;
      RECT  48215.0 66380.0 48920.0 65035.0 ;
      RECT  48215.0 66380.0 48920.0 67725.0 ;
      RECT  48215.0 69070.0 48920.0 67725.0 ;
      RECT  48215.0 69070.0 48920.0 70415.0 ;
      RECT  48215.0 71760.0 48920.0 70415.0 ;
      RECT  48215.0 71760.0 48920.0 73105.0 ;
      RECT  48215.0 74450.0 48920.0 73105.0 ;
      RECT  48215.0 74450.0 48920.0 75795.0 ;
      RECT  48215.0 77140.0 48920.0 75795.0 ;
      RECT  48215.0 77140.0 48920.0 78485.0 ;
      RECT  48215.0 79830.0 48920.0 78485.0 ;
      RECT  48215.0 79830.0 48920.0 81175.0 ;
      RECT  48215.0 82520.0 48920.0 81175.0 ;
      RECT  48215.0 82520.0 48920.0 83865.0 ;
      RECT  48215.0 85210.0 48920.0 83865.0 ;
      RECT  48215.0 85210.0 48920.0 86555.0 ;
      RECT  48215.0 87900.0 48920.0 86555.0 ;
      RECT  48215.0 87900.0 48920.0 89245.0 ;
      RECT  48215.0 90590.0 48920.0 89245.0 ;
      RECT  48215.0 90590.0 48920.0 91935.0 ;
      RECT  48215.0 93280.0 48920.0 91935.0 ;
      RECT  48215.0 93280.0 48920.0 94625.0 ;
      RECT  48215.0 95970.0 48920.0 94625.0 ;
      RECT  48215.0 95970.0 48920.0 97315.0 ;
      RECT  48215.0 98660.0 48920.0 97315.0 ;
      RECT  48215.0 98660.0 48920.0 100005.0 ;
      RECT  48215.0 101350.0 48920.0 100005.0 ;
      RECT  48215.0 101350.0 48920.0 102695.0 ;
      RECT  48215.0 104040.0 48920.0 102695.0 ;
      RECT  48215.0 104040.0 48920.0 105385.0 ;
      RECT  48215.0 106730.0 48920.0 105385.0 ;
      RECT  48215.0 106730.0 48920.0 108075.0 ;
      RECT  48215.0 109420.0 48920.0 108075.0 ;
      RECT  48215.0 109420.0 48920.0 110765.0 ;
      RECT  48215.0 112110.0 48920.0 110765.0 ;
      RECT  48215.0 112110.0 48920.0 113455.0 ;
      RECT  48215.0 114800.0 48920.0 113455.0 ;
      RECT  48215.0 114800.0 48920.0 116145.0 ;
      RECT  48215.0 117490.0 48920.0 116145.0 ;
      RECT  48215.0 117490.0 48920.0 118835.0 ;
      RECT  48215.0 120180.0 48920.0 118835.0 ;
      RECT  48215.0 120180.0 48920.0 121525.0 ;
      RECT  48215.0 122870.0 48920.0 121525.0 ;
      RECT  48215.0 122870.0 48920.0 124215.0 ;
      RECT  48215.0 125560.0 48920.0 124215.0 ;
      RECT  48215.0 125560.0 48920.0 126905.0 ;
      RECT  48215.0 128250.0 48920.0 126905.0 ;
      RECT  48215.0 128250.0 48920.0 129595.0 ;
      RECT  48215.0 130940.0 48920.0 129595.0 ;
      RECT  48215.0 130940.0 48920.0 132285.0 ;
      RECT  48215.0 133630.0 48920.0 132285.0 ;
      RECT  48215.0 133630.0 48920.0 134975.0 ;
      RECT  48215.0 136320.0 48920.0 134975.0 ;
      RECT  48215.0 136320.0 48920.0 137665.0 ;
      RECT  48215.0 139010.0 48920.0 137665.0 ;
      RECT  48215.0 139010.0 48920.0 140355.0 ;
      RECT  48215.0 141700.0 48920.0 140355.0 ;
      RECT  48215.0 141700.0 48920.0 143045.0 ;
      RECT  48215.0 144390.0 48920.0 143045.0 ;
      RECT  48215.0 144390.0 48920.0 145735.0 ;
      RECT  48215.0 147080.0 48920.0 145735.0 ;
      RECT  48215.0 147080.0 48920.0 148425.0 ;
      RECT  48215.0 149770.0 48920.0 148425.0 ;
      RECT  48215.0 149770.0 48920.0 151115.0 ;
      RECT  48215.0 152460.0 48920.0 151115.0 ;
      RECT  48215.0 152460.0 48920.0 153805.0 ;
      RECT  48215.0 155150.0 48920.0 153805.0 ;
      RECT  48215.0 155150.0 48920.0 156495.0 ;
      RECT  48215.0 157840.0 48920.0 156495.0 ;
      RECT  48215.0 157840.0 48920.0 159185.0 ;
      RECT  48215.0 160530.0 48920.0 159185.0 ;
      RECT  48215.0 160530.0 48920.0 161875.0 ;
      RECT  48215.0 163220.0 48920.0 161875.0 ;
      RECT  48215.0 163220.0 48920.0 164565.0 ;
      RECT  48215.0 165910.0 48920.0 164565.0 ;
      RECT  48215.0 165910.0 48920.0 167255.0 ;
      RECT  48215.0 168600.0 48920.0 167255.0 ;
      RECT  48215.0 168600.0 48920.0 169945.0 ;
      RECT  48215.0 171290.0 48920.0 169945.0 ;
      RECT  48215.0 171290.0 48920.0 172635.0 ;
      RECT  48215.0 173980.0 48920.0 172635.0 ;
      RECT  48215.0 173980.0 48920.0 175325.0 ;
      RECT  48215.0 176670.0 48920.0 175325.0 ;
      RECT  48215.0 176670.0 48920.0 178015.0 ;
      RECT  48215.0 179360.0 48920.0 178015.0 ;
      RECT  48215.0 179360.0 48920.0 180705.0 ;
      RECT  48215.0 182050.0 48920.0 180705.0 ;
      RECT  48215.0 182050.0 48920.0 183395.0 ;
      RECT  48215.0 184740.0 48920.0 183395.0 ;
      RECT  48215.0 184740.0 48920.0 186085.0 ;
      RECT  48215.0 187430.0 48920.0 186085.0 ;
      RECT  48215.0 187430.0 48920.0 188775.0 ;
      RECT  48215.0 190120.0 48920.0 188775.0 ;
      RECT  48215.0 190120.0 48920.0 191465.0 ;
      RECT  48215.0 192810.0 48920.0 191465.0 ;
      RECT  48215.0 192810.0 48920.0 194155.0 ;
      RECT  48215.0 195500.0 48920.0 194155.0 ;
      RECT  48215.0 195500.0 48920.0 196845.0 ;
      RECT  48215.0 198190.0 48920.0 196845.0 ;
      RECT  48215.0 198190.0 48920.0 199535.0 ;
      RECT  48215.0 200880.0 48920.0 199535.0 ;
      RECT  48215.0 200880.0 48920.0 202225.0 ;
      RECT  48215.0 203570.0 48920.0 202225.0 ;
      RECT  48215.0 203570.0 48920.0 204915.0 ;
      RECT  48215.0 206260.0 48920.0 204915.0 ;
      RECT  48920.0 34100.0 49625.0 35445.0 ;
      RECT  48920.0 36790.0 49625.0 35445.0 ;
      RECT  48920.0 36790.0 49625.0 38135.0 ;
      RECT  48920.0 39480.0 49625.0 38135.0 ;
      RECT  48920.0 39480.0 49625.0 40825.0 ;
      RECT  48920.0 42170.0 49625.0 40825.0 ;
      RECT  48920.0 42170.0 49625.0 43515.0 ;
      RECT  48920.0 44860.0 49625.0 43515.0 ;
      RECT  48920.0 44860.0 49625.0 46205.0 ;
      RECT  48920.0 47550.0 49625.0 46205.0 ;
      RECT  48920.0 47550.0 49625.0 48895.0 ;
      RECT  48920.0 50240.0 49625.0 48895.0 ;
      RECT  48920.0 50240.0 49625.0 51585.0 ;
      RECT  48920.0 52930.0 49625.0 51585.0 ;
      RECT  48920.0 52930.0 49625.0 54275.0 ;
      RECT  48920.0 55620.0 49625.0 54275.0 ;
      RECT  48920.0 55620.0 49625.0 56965.0 ;
      RECT  48920.0 58310.0 49625.0 56965.0 ;
      RECT  48920.0 58310.0 49625.0 59655.0 ;
      RECT  48920.0 61000.0 49625.0 59655.0 ;
      RECT  48920.0 61000.0 49625.0 62345.0 ;
      RECT  48920.0 63690.0 49625.0 62345.0 ;
      RECT  48920.0 63690.0 49625.0 65035.0 ;
      RECT  48920.0 66380.0 49625.0 65035.0 ;
      RECT  48920.0 66380.0 49625.0 67725.0 ;
      RECT  48920.0 69070.0 49625.0 67725.0 ;
      RECT  48920.0 69070.0 49625.0 70415.0 ;
      RECT  48920.0 71760.0 49625.0 70415.0 ;
      RECT  48920.0 71760.0 49625.0 73105.0 ;
      RECT  48920.0 74450.0 49625.0 73105.0 ;
      RECT  48920.0 74450.0 49625.0 75795.0 ;
      RECT  48920.0 77140.0 49625.0 75795.0 ;
      RECT  48920.0 77140.0 49625.0 78485.0 ;
      RECT  48920.0 79830.0 49625.0 78485.0 ;
      RECT  48920.0 79830.0 49625.0 81175.0 ;
      RECT  48920.0 82520.0 49625.0 81175.0 ;
      RECT  48920.0 82520.0 49625.0 83865.0 ;
      RECT  48920.0 85210.0 49625.0 83865.0 ;
      RECT  48920.0 85210.0 49625.0 86555.0 ;
      RECT  48920.0 87900.0 49625.0 86555.0 ;
      RECT  48920.0 87900.0 49625.0 89245.0 ;
      RECT  48920.0 90590.0 49625.0 89245.0 ;
      RECT  48920.0 90590.0 49625.0 91935.0 ;
      RECT  48920.0 93280.0 49625.0 91935.0 ;
      RECT  48920.0 93280.0 49625.0 94625.0 ;
      RECT  48920.0 95970.0 49625.0 94625.0 ;
      RECT  48920.0 95970.0 49625.0 97315.0 ;
      RECT  48920.0 98660.0 49625.0 97315.0 ;
      RECT  48920.0 98660.0 49625.0 100005.0 ;
      RECT  48920.0 101350.0 49625.0 100005.0 ;
      RECT  48920.0 101350.0 49625.0 102695.0 ;
      RECT  48920.0 104040.0 49625.0 102695.0 ;
      RECT  48920.0 104040.0 49625.0 105385.0 ;
      RECT  48920.0 106730.0 49625.0 105385.0 ;
      RECT  48920.0 106730.0 49625.0 108075.0 ;
      RECT  48920.0 109420.0 49625.0 108075.0 ;
      RECT  48920.0 109420.0 49625.0 110765.0 ;
      RECT  48920.0 112110.0 49625.0 110765.0 ;
      RECT  48920.0 112110.0 49625.0 113455.0 ;
      RECT  48920.0 114800.0 49625.0 113455.0 ;
      RECT  48920.0 114800.0 49625.0 116145.0 ;
      RECT  48920.0 117490.0 49625.0 116145.0 ;
      RECT  48920.0 117490.0 49625.0 118835.0 ;
      RECT  48920.0 120180.0 49625.0 118835.0 ;
      RECT  48920.0 120180.0 49625.0 121525.0 ;
      RECT  48920.0 122870.0 49625.0 121525.0 ;
      RECT  48920.0 122870.0 49625.0 124215.0 ;
      RECT  48920.0 125560.0 49625.0 124215.0 ;
      RECT  48920.0 125560.0 49625.0 126905.0 ;
      RECT  48920.0 128250.0 49625.0 126905.0 ;
      RECT  48920.0 128250.0 49625.0 129595.0 ;
      RECT  48920.0 130940.0 49625.0 129595.0 ;
      RECT  48920.0 130940.0 49625.0 132285.0 ;
      RECT  48920.0 133630.0 49625.0 132285.0 ;
      RECT  48920.0 133630.0 49625.0 134975.0 ;
      RECT  48920.0 136320.0 49625.0 134975.0 ;
      RECT  48920.0 136320.0 49625.0 137665.0 ;
      RECT  48920.0 139010.0 49625.0 137665.0 ;
      RECT  48920.0 139010.0 49625.0 140355.0 ;
      RECT  48920.0 141700.0 49625.0 140355.0 ;
      RECT  48920.0 141700.0 49625.0 143045.0 ;
      RECT  48920.0 144390.0 49625.0 143045.0 ;
      RECT  48920.0 144390.0 49625.0 145735.0 ;
      RECT  48920.0 147080.0 49625.0 145735.0 ;
      RECT  48920.0 147080.0 49625.0 148425.0 ;
      RECT  48920.0 149770.0 49625.0 148425.0 ;
      RECT  48920.0 149770.0 49625.0 151115.0 ;
      RECT  48920.0 152460.0 49625.0 151115.0 ;
      RECT  48920.0 152460.0 49625.0 153805.0 ;
      RECT  48920.0 155150.0 49625.0 153805.0 ;
      RECT  48920.0 155150.0 49625.0 156495.0 ;
      RECT  48920.0 157840.0 49625.0 156495.0 ;
      RECT  48920.0 157840.0 49625.0 159185.0 ;
      RECT  48920.0 160530.0 49625.0 159185.0 ;
      RECT  48920.0 160530.0 49625.0 161875.0 ;
      RECT  48920.0 163220.0 49625.0 161875.0 ;
      RECT  48920.0 163220.0 49625.0 164565.0 ;
      RECT  48920.0 165910.0 49625.0 164565.0 ;
      RECT  48920.0 165910.0 49625.0 167255.0 ;
      RECT  48920.0 168600.0 49625.0 167255.0 ;
      RECT  48920.0 168600.0 49625.0 169945.0 ;
      RECT  48920.0 171290.0 49625.0 169945.0 ;
      RECT  48920.0 171290.0 49625.0 172635.0 ;
      RECT  48920.0 173980.0 49625.0 172635.0 ;
      RECT  48920.0 173980.0 49625.0 175325.0 ;
      RECT  48920.0 176670.0 49625.0 175325.0 ;
      RECT  48920.0 176670.0 49625.0 178015.0 ;
      RECT  48920.0 179360.0 49625.0 178015.0 ;
      RECT  48920.0 179360.0 49625.0 180705.0 ;
      RECT  48920.0 182050.0 49625.0 180705.0 ;
      RECT  48920.0 182050.0 49625.0 183395.0 ;
      RECT  48920.0 184740.0 49625.0 183395.0 ;
      RECT  48920.0 184740.0 49625.0 186085.0 ;
      RECT  48920.0 187430.0 49625.0 186085.0 ;
      RECT  48920.0 187430.0 49625.0 188775.0 ;
      RECT  48920.0 190120.0 49625.0 188775.0 ;
      RECT  48920.0 190120.0 49625.0 191465.0 ;
      RECT  48920.0 192810.0 49625.0 191465.0 ;
      RECT  48920.0 192810.0 49625.0 194155.0 ;
      RECT  48920.0 195500.0 49625.0 194155.0 ;
      RECT  48920.0 195500.0 49625.0 196845.0 ;
      RECT  48920.0 198190.0 49625.0 196845.0 ;
      RECT  48920.0 198190.0 49625.0 199535.0 ;
      RECT  48920.0 200880.0 49625.0 199535.0 ;
      RECT  48920.0 200880.0 49625.0 202225.0 ;
      RECT  48920.0 203570.0 49625.0 202225.0 ;
      RECT  48920.0 203570.0 49625.0 204915.0 ;
      RECT  48920.0 206260.0 49625.0 204915.0 ;
      RECT  49625.0 34100.0 50330.0 35445.0 ;
      RECT  49625.0 36790.0 50330.0 35445.0 ;
      RECT  49625.0 36790.0 50330.0 38135.0 ;
      RECT  49625.0 39480.0 50330.0 38135.0 ;
      RECT  49625.0 39480.0 50330.0 40825.0 ;
      RECT  49625.0 42170.0 50330.0 40825.0 ;
      RECT  49625.0 42170.0 50330.0 43515.0 ;
      RECT  49625.0 44860.0 50330.0 43515.0 ;
      RECT  49625.0 44860.0 50330.0 46205.0 ;
      RECT  49625.0 47550.0 50330.0 46205.0 ;
      RECT  49625.0 47550.0 50330.0 48895.0 ;
      RECT  49625.0 50240.0 50330.0 48895.0 ;
      RECT  49625.0 50240.0 50330.0 51585.0 ;
      RECT  49625.0 52930.0 50330.0 51585.0 ;
      RECT  49625.0 52930.0 50330.0 54275.0 ;
      RECT  49625.0 55620.0 50330.0 54275.0 ;
      RECT  49625.0 55620.0 50330.0 56965.0 ;
      RECT  49625.0 58310.0 50330.0 56965.0 ;
      RECT  49625.0 58310.0 50330.0 59655.0 ;
      RECT  49625.0 61000.0 50330.0 59655.0 ;
      RECT  49625.0 61000.0 50330.0 62345.0 ;
      RECT  49625.0 63690.0 50330.0 62345.0 ;
      RECT  49625.0 63690.0 50330.0 65035.0 ;
      RECT  49625.0 66380.0 50330.0 65035.0 ;
      RECT  49625.0 66380.0 50330.0 67725.0 ;
      RECT  49625.0 69070.0 50330.0 67725.0 ;
      RECT  49625.0 69070.0 50330.0 70415.0 ;
      RECT  49625.0 71760.0 50330.0 70415.0 ;
      RECT  49625.0 71760.0 50330.0 73105.0 ;
      RECT  49625.0 74450.0 50330.0 73105.0 ;
      RECT  49625.0 74450.0 50330.0 75795.0 ;
      RECT  49625.0 77140.0 50330.0 75795.0 ;
      RECT  49625.0 77140.0 50330.0 78485.0 ;
      RECT  49625.0 79830.0 50330.0 78485.0 ;
      RECT  49625.0 79830.0 50330.0 81175.0 ;
      RECT  49625.0 82520.0 50330.0 81175.0 ;
      RECT  49625.0 82520.0 50330.0 83865.0 ;
      RECT  49625.0 85210.0 50330.0 83865.0 ;
      RECT  49625.0 85210.0 50330.0 86555.0 ;
      RECT  49625.0 87900.0 50330.0 86555.0 ;
      RECT  49625.0 87900.0 50330.0 89245.0 ;
      RECT  49625.0 90590.0 50330.0 89245.0 ;
      RECT  49625.0 90590.0 50330.0 91935.0 ;
      RECT  49625.0 93280.0 50330.0 91935.0 ;
      RECT  49625.0 93280.0 50330.0 94625.0 ;
      RECT  49625.0 95970.0 50330.0 94625.0 ;
      RECT  49625.0 95970.0 50330.0 97315.0 ;
      RECT  49625.0 98660.0 50330.0 97315.0 ;
      RECT  49625.0 98660.0 50330.0 100005.0 ;
      RECT  49625.0 101350.0 50330.0 100005.0 ;
      RECT  49625.0 101350.0 50330.0 102695.0 ;
      RECT  49625.0 104040.0 50330.0 102695.0 ;
      RECT  49625.0 104040.0 50330.0 105385.0 ;
      RECT  49625.0 106730.0 50330.0 105385.0 ;
      RECT  49625.0 106730.0 50330.0 108075.0 ;
      RECT  49625.0 109420.0 50330.0 108075.0 ;
      RECT  49625.0 109420.0 50330.0 110765.0 ;
      RECT  49625.0 112110.0 50330.0 110765.0 ;
      RECT  49625.0 112110.0 50330.0 113455.0 ;
      RECT  49625.0 114800.0 50330.0 113455.0 ;
      RECT  49625.0 114800.0 50330.0 116145.0 ;
      RECT  49625.0 117490.0 50330.0 116145.0 ;
      RECT  49625.0 117490.0 50330.0 118835.0 ;
      RECT  49625.0 120180.0 50330.0 118835.0 ;
      RECT  49625.0 120180.0 50330.0 121525.0 ;
      RECT  49625.0 122870.0 50330.0 121525.0 ;
      RECT  49625.0 122870.0 50330.0 124215.0 ;
      RECT  49625.0 125560.0 50330.0 124215.0 ;
      RECT  49625.0 125560.0 50330.0 126905.0 ;
      RECT  49625.0 128250.0 50330.0 126905.0 ;
      RECT  49625.0 128250.0 50330.0 129595.0 ;
      RECT  49625.0 130940.0 50330.0 129595.0 ;
      RECT  49625.0 130940.0 50330.0 132285.0 ;
      RECT  49625.0 133630.0 50330.0 132285.0 ;
      RECT  49625.0 133630.0 50330.0 134975.0 ;
      RECT  49625.0 136320.0 50330.0 134975.0 ;
      RECT  49625.0 136320.0 50330.0 137665.0 ;
      RECT  49625.0 139010.0 50330.0 137665.0 ;
      RECT  49625.0 139010.0 50330.0 140355.0 ;
      RECT  49625.0 141700.0 50330.0 140355.0 ;
      RECT  49625.0 141700.0 50330.0 143045.0 ;
      RECT  49625.0 144390.0 50330.0 143045.0 ;
      RECT  49625.0 144390.0 50330.0 145735.0 ;
      RECT  49625.0 147080.0 50330.0 145735.0 ;
      RECT  49625.0 147080.0 50330.0 148425.0 ;
      RECT  49625.0 149770.0 50330.0 148425.0 ;
      RECT  49625.0 149770.0 50330.0 151115.0 ;
      RECT  49625.0 152460.0 50330.0 151115.0 ;
      RECT  49625.0 152460.0 50330.0 153805.0 ;
      RECT  49625.0 155150.0 50330.0 153805.0 ;
      RECT  49625.0 155150.0 50330.0 156495.0 ;
      RECT  49625.0 157840.0 50330.0 156495.0 ;
      RECT  49625.0 157840.0 50330.0 159185.0 ;
      RECT  49625.0 160530.0 50330.0 159185.0 ;
      RECT  49625.0 160530.0 50330.0 161875.0 ;
      RECT  49625.0 163220.0 50330.0 161875.0 ;
      RECT  49625.0 163220.0 50330.0 164565.0 ;
      RECT  49625.0 165910.0 50330.0 164565.0 ;
      RECT  49625.0 165910.0 50330.0 167255.0 ;
      RECT  49625.0 168600.0 50330.0 167255.0 ;
      RECT  49625.0 168600.0 50330.0 169945.0 ;
      RECT  49625.0 171290.0 50330.0 169945.0 ;
      RECT  49625.0 171290.0 50330.0 172635.0 ;
      RECT  49625.0 173980.0 50330.0 172635.0 ;
      RECT  49625.0 173980.0 50330.0 175325.0 ;
      RECT  49625.0 176670.0 50330.0 175325.0 ;
      RECT  49625.0 176670.0 50330.0 178015.0 ;
      RECT  49625.0 179360.0 50330.0 178015.0 ;
      RECT  49625.0 179360.0 50330.0 180705.0 ;
      RECT  49625.0 182050.0 50330.0 180705.0 ;
      RECT  49625.0 182050.0 50330.0 183395.0 ;
      RECT  49625.0 184740.0 50330.0 183395.0 ;
      RECT  49625.0 184740.0 50330.0 186085.0 ;
      RECT  49625.0 187430.0 50330.0 186085.0 ;
      RECT  49625.0 187430.0 50330.0 188775.0 ;
      RECT  49625.0 190120.0 50330.0 188775.0 ;
      RECT  49625.0 190120.0 50330.0 191465.0 ;
      RECT  49625.0 192810.0 50330.0 191465.0 ;
      RECT  49625.0 192810.0 50330.0 194155.0 ;
      RECT  49625.0 195500.0 50330.0 194155.0 ;
      RECT  49625.0 195500.0 50330.0 196845.0 ;
      RECT  49625.0 198190.0 50330.0 196845.0 ;
      RECT  49625.0 198190.0 50330.0 199535.0 ;
      RECT  49625.0 200880.0 50330.0 199535.0 ;
      RECT  49625.0 200880.0 50330.0 202225.0 ;
      RECT  49625.0 203570.0 50330.0 202225.0 ;
      RECT  49625.0 203570.0 50330.0 204915.0 ;
      RECT  49625.0 206260.0 50330.0 204915.0 ;
      RECT  50330.0 34100.0 51035.0 35445.0 ;
      RECT  50330.0 36790.0 51035.0 35445.0 ;
      RECT  50330.0 36790.0 51035.0 38135.0 ;
      RECT  50330.0 39480.0 51035.0 38135.0 ;
      RECT  50330.0 39480.0 51035.0 40825.0 ;
      RECT  50330.0 42170.0 51035.0 40825.0 ;
      RECT  50330.0 42170.0 51035.0 43515.0 ;
      RECT  50330.0 44860.0 51035.0 43515.0 ;
      RECT  50330.0 44860.0 51035.0 46205.0 ;
      RECT  50330.0 47550.0 51035.0 46205.0 ;
      RECT  50330.0 47550.0 51035.0 48895.0 ;
      RECT  50330.0 50240.0 51035.0 48895.0 ;
      RECT  50330.0 50240.0 51035.0 51585.0 ;
      RECT  50330.0 52930.0 51035.0 51585.0 ;
      RECT  50330.0 52930.0 51035.0 54275.0 ;
      RECT  50330.0 55620.0 51035.0 54275.0 ;
      RECT  50330.0 55620.0 51035.0 56965.0 ;
      RECT  50330.0 58310.0 51035.0 56965.0 ;
      RECT  50330.0 58310.0 51035.0 59655.0 ;
      RECT  50330.0 61000.0 51035.0 59655.0 ;
      RECT  50330.0 61000.0 51035.0 62345.0 ;
      RECT  50330.0 63690.0 51035.0 62345.0 ;
      RECT  50330.0 63690.0 51035.0 65035.0 ;
      RECT  50330.0 66380.0 51035.0 65035.0 ;
      RECT  50330.0 66380.0 51035.0 67725.0 ;
      RECT  50330.0 69070.0 51035.0 67725.0 ;
      RECT  50330.0 69070.0 51035.0 70415.0 ;
      RECT  50330.0 71760.0 51035.0 70415.0 ;
      RECT  50330.0 71760.0 51035.0 73105.0 ;
      RECT  50330.0 74450.0 51035.0 73105.0 ;
      RECT  50330.0 74450.0 51035.0 75795.0 ;
      RECT  50330.0 77140.0 51035.0 75795.0 ;
      RECT  50330.0 77140.0 51035.0 78485.0 ;
      RECT  50330.0 79830.0 51035.0 78485.0 ;
      RECT  50330.0 79830.0 51035.0 81175.0 ;
      RECT  50330.0 82520.0 51035.0 81175.0 ;
      RECT  50330.0 82520.0 51035.0 83865.0 ;
      RECT  50330.0 85210.0 51035.0 83865.0 ;
      RECT  50330.0 85210.0 51035.0 86555.0 ;
      RECT  50330.0 87900.0 51035.0 86555.0 ;
      RECT  50330.0 87900.0 51035.0 89245.0 ;
      RECT  50330.0 90590.0 51035.0 89245.0 ;
      RECT  50330.0 90590.0 51035.0 91935.0 ;
      RECT  50330.0 93280.0 51035.0 91935.0 ;
      RECT  50330.0 93280.0 51035.0 94625.0 ;
      RECT  50330.0 95970.0 51035.0 94625.0 ;
      RECT  50330.0 95970.0 51035.0 97315.0 ;
      RECT  50330.0 98660.0 51035.0 97315.0 ;
      RECT  50330.0 98660.0 51035.0 100005.0 ;
      RECT  50330.0 101350.0 51035.0 100005.0 ;
      RECT  50330.0 101350.0 51035.0 102695.0 ;
      RECT  50330.0 104040.0 51035.0 102695.0 ;
      RECT  50330.0 104040.0 51035.0 105385.0 ;
      RECT  50330.0 106730.0 51035.0 105385.0 ;
      RECT  50330.0 106730.0 51035.0 108075.0 ;
      RECT  50330.0 109420.0 51035.0 108075.0 ;
      RECT  50330.0 109420.0 51035.0 110765.0 ;
      RECT  50330.0 112110.0 51035.0 110765.0 ;
      RECT  50330.0 112110.0 51035.0 113455.0 ;
      RECT  50330.0 114800.0 51035.0 113455.0 ;
      RECT  50330.0 114800.0 51035.0 116145.0 ;
      RECT  50330.0 117490.0 51035.0 116145.0 ;
      RECT  50330.0 117490.0 51035.0 118835.0 ;
      RECT  50330.0 120180.0 51035.0 118835.0 ;
      RECT  50330.0 120180.0 51035.0 121525.0 ;
      RECT  50330.0 122870.0 51035.0 121525.0 ;
      RECT  50330.0 122870.0 51035.0 124215.0 ;
      RECT  50330.0 125560.0 51035.0 124215.0 ;
      RECT  50330.0 125560.0 51035.0 126905.0 ;
      RECT  50330.0 128250.0 51035.0 126905.0 ;
      RECT  50330.0 128250.0 51035.0 129595.0 ;
      RECT  50330.0 130940.0 51035.0 129595.0 ;
      RECT  50330.0 130940.0 51035.0 132285.0 ;
      RECT  50330.0 133630.0 51035.0 132285.0 ;
      RECT  50330.0 133630.0 51035.0 134975.0 ;
      RECT  50330.0 136320.0 51035.0 134975.0 ;
      RECT  50330.0 136320.0 51035.0 137665.0 ;
      RECT  50330.0 139010.0 51035.0 137665.0 ;
      RECT  50330.0 139010.0 51035.0 140355.0 ;
      RECT  50330.0 141700.0 51035.0 140355.0 ;
      RECT  50330.0 141700.0 51035.0 143045.0 ;
      RECT  50330.0 144390.0 51035.0 143045.0 ;
      RECT  50330.0 144390.0 51035.0 145735.0 ;
      RECT  50330.0 147080.0 51035.0 145735.0 ;
      RECT  50330.0 147080.0 51035.0 148425.0 ;
      RECT  50330.0 149770.0 51035.0 148425.0 ;
      RECT  50330.0 149770.0 51035.0 151115.0 ;
      RECT  50330.0 152460.0 51035.0 151115.0 ;
      RECT  50330.0 152460.0 51035.0 153805.0 ;
      RECT  50330.0 155150.0 51035.0 153805.0 ;
      RECT  50330.0 155150.0 51035.0 156495.0 ;
      RECT  50330.0 157840.0 51035.0 156495.0 ;
      RECT  50330.0 157840.0 51035.0 159185.0 ;
      RECT  50330.0 160530.0 51035.0 159185.0 ;
      RECT  50330.0 160530.0 51035.0 161875.0 ;
      RECT  50330.0 163220.0 51035.0 161875.0 ;
      RECT  50330.0 163220.0 51035.0 164565.0 ;
      RECT  50330.0 165910.0 51035.0 164565.0 ;
      RECT  50330.0 165910.0 51035.0 167255.0 ;
      RECT  50330.0 168600.0 51035.0 167255.0 ;
      RECT  50330.0 168600.0 51035.0 169945.0 ;
      RECT  50330.0 171290.0 51035.0 169945.0 ;
      RECT  50330.0 171290.0 51035.0 172635.0 ;
      RECT  50330.0 173980.0 51035.0 172635.0 ;
      RECT  50330.0 173980.0 51035.0 175325.0 ;
      RECT  50330.0 176670.0 51035.0 175325.0 ;
      RECT  50330.0 176670.0 51035.0 178015.0 ;
      RECT  50330.0 179360.0 51035.0 178015.0 ;
      RECT  50330.0 179360.0 51035.0 180705.0 ;
      RECT  50330.0 182050.0 51035.0 180705.0 ;
      RECT  50330.0 182050.0 51035.0 183395.0 ;
      RECT  50330.0 184740.0 51035.0 183395.0 ;
      RECT  50330.0 184740.0 51035.0 186085.0 ;
      RECT  50330.0 187430.0 51035.0 186085.0 ;
      RECT  50330.0 187430.0 51035.0 188775.0 ;
      RECT  50330.0 190120.0 51035.0 188775.0 ;
      RECT  50330.0 190120.0 51035.0 191465.0 ;
      RECT  50330.0 192810.0 51035.0 191465.0 ;
      RECT  50330.0 192810.0 51035.0 194155.0 ;
      RECT  50330.0 195500.0 51035.0 194155.0 ;
      RECT  50330.0 195500.0 51035.0 196845.0 ;
      RECT  50330.0 198190.0 51035.0 196845.0 ;
      RECT  50330.0 198190.0 51035.0 199535.0 ;
      RECT  50330.0 200880.0 51035.0 199535.0 ;
      RECT  50330.0 200880.0 51035.0 202225.0 ;
      RECT  50330.0 203570.0 51035.0 202225.0 ;
      RECT  50330.0 203570.0 51035.0 204915.0 ;
      RECT  50330.0 206260.0 51035.0 204915.0 ;
      RECT  51035.0 34100.0 51740.0 35445.0 ;
      RECT  51035.0 36790.0 51740.0 35445.0 ;
      RECT  51035.0 36790.0 51740.0 38135.0 ;
      RECT  51035.0 39480.0 51740.0 38135.0 ;
      RECT  51035.0 39480.0 51740.0 40825.0 ;
      RECT  51035.0 42170.0 51740.0 40825.0 ;
      RECT  51035.0 42170.0 51740.0 43515.0 ;
      RECT  51035.0 44860.0 51740.0 43515.0 ;
      RECT  51035.0 44860.0 51740.0 46205.0 ;
      RECT  51035.0 47550.0 51740.0 46205.0 ;
      RECT  51035.0 47550.0 51740.0 48895.0 ;
      RECT  51035.0 50240.0 51740.0 48895.0 ;
      RECT  51035.0 50240.0 51740.0 51585.0 ;
      RECT  51035.0 52930.0 51740.0 51585.0 ;
      RECT  51035.0 52930.0 51740.0 54275.0 ;
      RECT  51035.0 55620.0 51740.0 54275.0 ;
      RECT  51035.0 55620.0 51740.0 56965.0 ;
      RECT  51035.0 58310.0 51740.0 56965.0 ;
      RECT  51035.0 58310.0 51740.0 59655.0 ;
      RECT  51035.0 61000.0 51740.0 59655.0 ;
      RECT  51035.0 61000.0 51740.0 62345.0 ;
      RECT  51035.0 63690.0 51740.0 62345.0 ;
      RECT  51035.0 63690.0 51740.0 65035.0 ;
      RECT  51035.0 66380.0 51740.0 65035.0 ;
      RECT  51035.0 66380.0 51740.0 67725.0 ;
      RECT  51035.0 69070.0 51740.0 67725.0 ;
      RECT  51035.0 69070.0 51740.0 70415.0 ;
      RECT  51035.0 71760.0 51740.0 70415.0 ;
      RECT  51035.0 71760.0 51740.0 73105.0 ;
      RECT  51035.0 74450.0 51740.0 73105.0 ;
      RECT  51035.0 74450.0 51740.0 75795.0 ;
      RECT  51035.0 77140.0 51740.0 75795.0 ;
      RECT  51035.0 77140.0 51740.0 78485.0 ;
      RECT  51035.0 79830.0 51740.0 78485.0 ;
      RECT  51035.0 79830.0 51740.0 81175.0 ;
      RECT  51035.0 82520.0 51740.0 81175.0 ;
      RECT  51035.0 82520.0 51740.0 83865.0 ;
      RECT  51035.0 85210.0 51740.0 83865.0 ;
      RECT  51035.0 85210.0 51740.0 86555.0 ;
      RECT  51035.0 87900.0 51740.0 86555.0 ;
      RECT  51035.0 87900.0 51740.0 89245.0 ;
      RECT  51035.0 90590.0 51740.0 89245.0 ;
      RECT  51035.0 90590.0 51740.0 91935.0 ;
      RECT  51035.0 93280.0 51740.0 91935.0 ;
      RECT  51035.0 93280.0 51740.0 94625.0 ;
      RECT  51035.0 95970.0 51740.0 94625.0 ;
      RECT  51035.0 95970.0 51740.0 97315.0 ;
      RECT  51035.0 98660.0 51740.0 97315.0 ;
      RECT  51035.0 98660.0 51740.0 100005.0 ;
      RECT  51035.0 101350.0 51740.0 100005.0 ;
      RECT  51035.0 101350.0 51740.0 102695.0 ;
      RECT  51035.0 104040.0 51740.0 102695.0 ;
      RECT  51035.0 104040.0 51740.0 105385.0 ;
      RECT  51035.0 106730.0 51740.0 105385.0 ;
      RECT  51035.0 106730.0 51740.0 108075.0 ;
      RECT  51035.0 109420.0 51740.0 108075.0 ;
      RECT  51035.0 109420.0 51740.0 110765.0 ;
      RECT  51035.0 112110.0 51740.0 110765.0 ;
      RECT  51035.0 112110.0 51740.0 113455.0 ;
      RECT  51035.0 114800.0 51740.0 113455.0 ;
      RECT  51035.0 114800.0 51740.0 116145.0 ;
      RECT  51035.0 117490.0 51740.0 116145.0 ;
      RECT  51035.0 117490.0 51740.0 118835.0 ;
      RECT  51035.0 120180.0 51740.0 118835.0 ;
      RECT  51035.0 120180.0 51740.0 121525.0 ;
      RECT  51035.0 122870.0 51740.0 121525.0 ;
      RECT  51035.0 122870.0 51740.0 124215.0 ;
      RECT  51035.0 125560.0 51740.0 124215.0 ;
      RECT  51035.0 125560.0 51740.0 126905.0 ;
      RECT  51035.0 128250.0 51740.0 126905.0 ;
      RECT  51035.0 128250.0 51740.0 129595.0 ;
      RECT  51035.0 130940.0 51740.0 129595.0 ;
      RECT  51035.0 130940.0 51740.0 132285.0 ;
      RECT  51035.0 133630.0 51740.0 132285.0 ;
      RECT  51035.0 133630.0 51740.0 134975.0 ;
      RECT  51035.0 136320.0 51740.0 134975.0 ;
      RECT  51035.0 136320.0 51740.0 137665.0 ;
      RECT  51035.0 139010.0 51740.0 137665.0 ;
      RECT  51035.0 139010.0 51740.0 140355.0 ;
      RECT  51035.0 141700.0 51740.0 140355.0 ;
      RECT  51035.0 141700.0 51740.0 143045.0 ;
      RECT  51035.0 144390.0 51740.0 143045.0 ;
      RECT  51035.0 144390.0 51740.0 145735.0 ;
      RECT  51035.0 147080.0 51740.0 145735.0 ;
      RECT  51035.0 147080.0 51740.0 148425.0 ;
      RECT  51035.0 149770.0 51740.0 148425.0 ;
      RECT  51035.0 149770.0 51740.0 151115.0 ;
      RECT  51035.0 152460.0 51740.0 151115.0 ;
      RECT  51035.0 152460.0 51740.0 153805.0 ;
      RECT  51035.0 155150.0 51740.0 153805.0 ;
      RECT  51035.0 155150.0 51740.0 156495.0 ;
      RECT  51035.0 157840.0 51740.0 156495.0 ;
      RECT  51035.0 157840.0 51740.0 159185.0 ;
      RECT  51035.0 160530.0 51740.0 159185.0 ;
      RECT  51035.0 160530.0 51740.0 161875.0 ;
      RECT  51035.0 163220.0 51740.0 161875.0 ;
      RECT  51035.0 163220.0 51740.0 164565.0 ;
      RECT  51035.0 165910.0 51740.0 164565.0 ;
      RECT  51035.0 165910.0 51740.0 167255.0 ;
      RECT  51035.0 168600.0 51740.0 167255.0 ;
      RECT  51035.0 168600.0 51740.0 169945.0 ;
      RECT  51035.0 171290.0 51740.0 169945.0 ;
      RECT  51035.0 171290.0 51740.0 172635.0 ;
      RECT  51035.0 173980.0 51740.0 172635.0 ;
      RECT  51035.0 173980.0 51740.0 175325.0 ;
      RECT  51035.0 176670.0 51740.0 175325.0 ;
      RECT  51035.0 176670.0 51740.0 178015.0 ;
      RECT  51035.0 179360.0 51740.0 178015.0 ;
      RECT  51035.0 179360.0 51740.0 180705.0 ;
      RECT  51035.0 182050.0 51740.0 180705.0 ;
      RECT  51035.0 182050.0 51740.0 183395.0 ;
      RECT  51035.0 184740.0 51740.0 183395.0 ;
      RECT  51035.0 184740.0 51740.0 186085.0 ;
      RECT  51035.0 187430.0 51740.0 186085.0 ;
      RECT  51035.0 187430.0 51740.0 188775.0 ;
      RECT  51035.0 190120.0 51740.0 188775.0 ;
      RECT  51035.0 190120.0 51740.0 191465.0 ;
      RECT  51035.0 192810.0 51740.0 191465.0 ;
      RECT  51035.0 192810.0 51740.0 194155.0 ;
      RECT  51035.0 195500.0 51740.0 194155.0 ;
      RECT  51035.0 195500.0 51740.0 196845.0 ;
      RECT  51035.0 198190.0 51740.0 196845.0 ;
      RECT  51035.0 198190.0 51740.0 199535.0 ;
      RECT  51035.0 200880.0 51740.0 199535.0 ;
      RECT  51035.0 200880.0 51740.0 202225.0 ;
      RECT  51035.0 203570.0 51740.0 202225.0 ;
      RECT  51035.0 203570.0 51740.0 204915.0 ;
      RECT  51035.0 206260.0 51740.0 204915.0 ;
      RECT  51740.0 34100.0 52445.0 35445.0 ;
      RECT  51740.0 36790.0 52445.0 35445.0 ;
      RECT  51740.0 36790.0 52445.0 38135.0 ;
      RECT  51740.0 39480.0 52445.0 38135.0 ;
      RECT  51740.0 39480.0 52445.0 40825.0 ;
      RECT  51740.0 42170.0 52445.0 40825.0 ;
      RECT  51740.0 42170.0 52445.0 43515.0 ;
      RECT  51740.0 44860.0 52445.0 43515.0 ;
      RECT  51740.0 44860.0 52445.0 46205.0 ;
      RECT  51740.0 47550.0 52445.0 46205.0 ;
      RECT  51740.0 47550.0 52445.0 48895.0 ;
      RECT  51740.0 50240.0 52445.0 48895.0 ;
      RECT  51740.0 50240.0 52445.0 51585.0 ;
      RECT  51740.0 52930.0 52445.0 51585.0 ;
      RECT  51740.0 52930.0 52445.0 54275.0 ;
      RECT  51740.0 55620.0 52445.0 54275.0 ;
      RECT  51740.0 55620.0 52445.0 56965.0 ;
      RECT  51740.0 58310.0 52445.0 56965.0 ;
      RECT  51740.0 58310.0 52445.0 59655.0 ;
      RECT  51740.0 61000.0 52445.0 59655.0 ;
      RECT  51740.0 61000.0 52445.0 62345.0 ;
      RECT  51740.0 63690.0 52445.0 62345.0 ;
      RECT  51740.0 63690.0 52445.0 65035.0 ;
      RECT  51740.0 66380.0 52445.0 65035.0 ;
      RECT  51740.0 66380.0 52445.0 67725.0 ;
      RECT  51740.0 69070.0 52445.0 67725.0 ;
      RECT  51740.0 69070.0 52445.0 70415.0 ;
      RECT  51740.0 71760.0 52445.0 70415.0 ;
      RECT  51740.0 71760.0 52445.0 73105.0 ;
      RECT  51740.0 74450.0 52445.0 73105.0 ;
      RECT  51740.0 74450.0 52445.0 75795.0 ;
      RECT  51740.0 77140.0 52445.0 75795.0 ;
      RECT  51740.0 77140.0 52445.0 78485.0 ;
      RECT  51740.0 79830.0 52445.0 78485.0 ;
      RECT  51740.0 79830.0 52445.0 81175.0 ;
      RECT  51740.0 82520.0 52445.0 81175.0 ;
      RECT  51740.0 82520.0 52445.0 83865.0 ;
      RECT  51740.0 85210.0 52445.0 83865.0 ;
      RECT  51740.0 85210.0 52445.0 86555.0 ;
      RECT  51740.0 87900.0 52445.0 86555.0 ;
      RECT  51740.0 87900.0 52445.0 89245.0 ;
      RECT  51740.0 90590.0 52445.0 89245.0 ;
      RECT  51740.0 90590.0 52445.0 91935.0 ;
      RECT  51740.0 93280.0 52445.0 91935.0 ;
      RECT  51740.0 93280.0 52445.0 94625.0 ;
      RECT  51740.0 95970.0 52445.0 94625.0 ;
      RECT  51740.0 95970.0 52445.0 97315.0 ;
      RECT  51740.0 98660.0 52445.0 97315.0 ;
      RECT  51740.0 98660.0 52445.0 100005.0 ;
      RECT  51740.0 101350.0 52445.0 100005.0 ;
      RECT  51740.0 101350.0 52445.0 102695.0 ;
      RECT  51740.0 104040.0 52445.0 102695.0 ;
      RECT  51740.0 104040.0 52445.0 105385.0 ;
      RECT  51740.0 106730.0 52445.0 105385.0 ;
      RECT  51740.0 106730.0 52445.0 108075.0 ;
      RECT  51740.0 109420.0 52445.0 108075.0 ;
      RECT  51740.0 109420.0 52445.0 110765.0 ;
      RECT  51740.0 112110.0 52445.0 110765.0 ;
      RECT  51740.0 112110.0 52445.0 113455.0 ;
      RECT  51740.0 114800.0 52445.0 113455.0 ;
      RECT  51740.0 114800.0 52445.0 116145.0 ;
      RECT  51740.0 117490.0 52445.0 116145.0 ;
      RECT  51740.0 117490.0 52445.0 118835.0 ;
      RECT  51740.0 120180.0 52445.0 118835.0 ;
      RECT  51740.0 120180.0 52445.0 121525.0 ;
      RECT  51740.0 122870.0 52445.0 121525.0 ;
      RECT  51740.0 122870.0 52445.0 124215.0 ;
      RECT  51740.0 125560.0 52445.0 124215.0 ;
      RECT  51740.0 125560.0 52445.0 126905.0 ;
      RECT  51740.0 128250.0 52445.0 126905.0 ;
      RECT  51740.0 128250.0 52445.0 129595.0 ;
      RECT  51740.0 130940.0 52445.0 129595.0 ;
      RECT  51740.0 130940.0 52445.0 132285.0 ;
      RECT  51740.0 133630.0 52445.0 132285.0 ;
      RECT  51740.0 133630.0 52445.0 134975.0 ;
      RECT  51740.0 136320.0 52445.0 134975.0 ;
      RECT  51740.0 136320.0 52445.0 137665.0 ;
      RECT  51740.0 139010.0 52445.0 137665.0 ;
      RECT  51740.0 139010.0 52445.0 140355.0 ;
      RECT  51740.0 141700.0 52445.0 140355.0 ;
      RECT  51740.0 141700.0 52445.0 143045.0 ;
      RECT  51740.0 144390.0 52445.0 143045.0 ;
      RECT  51740.0 144390.0 52445.0 145735.0 ;
      RECT  51740.0 147080.0 52445.0 145735.0 ;
      RECT  51740.0 147080.0 52445.0 148425.0 ;
      RECT  51740.0 149770.0 52445.0 148425.0 ;
      RECT  51740.0 149770.0 52445.0 151115.0 ;
      RECT  51740.0 152460.0 52445.0 151115.0 ;
      RECT  51740.0 152460.0 52445.0 153805.0 ;
      RECT  51740.0 155150.0 52445.0 153805.0 ;
      RECT  51740.0 155150.0 52445.0 156495.0 ;
      RECT  51740.0 157840.0 52445.0 156495.0 ;
      RECT  51740.0 157840.0 52445.0 159185.0 ;
      RECT  51740.0 160530.0 52445.0 159185.0 ;
      RECT  51740.0 160530.0 52445.0 161875.0 ;
      RECT  51740.0 163220.0 52445.0 161875.0 ;
      RECT  51740.0 163220.0 52445.0 164565.0 ;
      RECT  51740.0 165910.0 52445.0 164565.0 ;
      RECT  51740.0 165910.0 52445.0 167255.0 ;
      RECT  51740.0 168600.0 52445.0 167255.0 ;
      RECT  51740.0 168600.0 52445.0 169945.0 ;
      RECT  51740.0 171290.0 52445.0 169945.0 ;
      RECT  51740.0 171290.0 52445.0 172635.0 ;
      RECT  51740.0 173980.0 52445.0 172635.0 ;
      RECT  51740.0 173980.0 52445.0 175325.0 ;
      RECT  51740.0 176670.0 52445.0 175325.0 ;
      RECT  51740.0 176670.0 52445.0 178015.0 ;
      RECT  51740.0 179360.0 52445.0 178015.0 ;
      RECT  51740.0 179360.0 52445.0 180705.0 ;
      RECT  51740.0 182050.0 52445.0 180705.0 ;
      RECT  51740.0 182050.0 52445.0 183395.0 ;
      RECT  51740.0 184740.0 52445.0 183395.0 ;
      RECT  51740.0 184740.0 52445.0 186085.0 ;
      RECT  51740.0 187430.0 52445.0 186085.0 ;
      RECT  51740.0 187430.0 52445.0 188775.0 ;
      RECT  51740.0 190120.0 52445.0 188775.0 ;
      RECT  51740.0 190120.0 52445.0 191465.0 ;
      RECT  51740.0 192810.0 52445.0 191465.0 ;
      RECT  51740.0 192810.0 52445.0 194155.0 ;
      RECT  51740.0 195500.0 52445.0 194155.0 ;
      RECT  51740.0 195500.0 52445.0 196845.0 ;
      RECT  51740.0 198190.0 52445.0 196845.0 ;
      RECT  51740.0 198190.0 52445.0 199535.0 ;
      RECT  51740.0 200880.0 52445.0 199535.0 ;
      RECT  51740.0 200880.0 52445.0 202225.0 ;
      RECT  51740.0 203570.0 52445.0 202225.0 ;
      RECT  51740.0 203570.0 52445.0 204915.0 ;
      RECT  51740.0 206260.0 52445.0 204915.0 ;
      RECT  52445.0 34100.0 53150.0 35445.0 ;
      RECT  52445.0 36790.0 53150.0 35445.0 ;
      RECT  52445.0 36790.0 53150.0 38135.0 ;
      RECT  52445.0 39480.0 53150.0 38135.0 ;
      RECT  52445.0 39480.0 53150.0 40825.0 ;
      RECT  52445.0 42170.0 53150.0 40825.0 ;
      RECT  52445.0 42170.0 53150.0 43515.0 ;
      RECT  52445.0 44860.0 53150.0 43515.0 ;
      RECT  52445.0 44860.0 53150.0 46205.0 ;
      RECT  52445.0 47550.0 53150.0 46205.0 ;
      RECT  52445.0 47550.0 53150.0 48895.0 ;
      RECT  52445.0 50240.0 53150.0 48895.0 ;
      RECT  52445.0 50240.0 53150.0 51585.0 ;
      RECT  52445.0 52930.0 53150.0 51585.0 ;
      RECT  52445.0 52930.0 53150.0 54275.0 ;
      RECT  52445.0 55620.0 53150.0 54275.0 ;
      RECT  52445.0 55620.0 53150.0 56965.0 ;
      RECT  52445.0 58310.0 53150.0 56965.0 ;
      RECT  52445.0 58310.0 53150.0 59655.0 ;
      RECT  52445.0 61000.0 53150.0 59655.0 ;
      RECT  52445.0 61000.0 53150.0 62345.0 ;
      RECT  52445.0 63690.0 53150.0 62345.0 ;
      RECT  52445.0 63690.0 53150.0 65035.0 ;
      RECT  52445.0 66380.0 53150.0 65035.0 ;
      RECT  52445.0 66380.0 53150.0 67725.0 ;
      RECT  52445.0 69070.0 53150.0 67725.0 ;
      RECT  52445.0 69070.0 53150.0 70415.0 ;
      RECT  52445.0 71760.0 53150.0 70415.0 ;
      RECT  52445.0 71760.0 53150.0 73105.0 ;
      RECT  52445.0 74450.0 53150.0 73105.0 ;
      RECT  52445.0 74450.0 53150.0 75795.0 ;
      RECT  52445.0 77140.0 53150.0 75795.0 ;
      RECT  52445.0 77140.0 53150.0 78485.0 ;
      RECT  52445.0 79830.0 53150.0 78485.0 ;
      RECT  52445.0 79830.0 53150.0 81175.0 ;
      RECT  52445.0 82520.0 53150.0 81175.0 ;
      RECT  52445.0 82520.0 53150.0 83865.0 ;
      RECT  52445.0 85210.0 53150.0 83865.0 ;
      RECT  52445.0 85210.0 53150.0 86555.0 ;
      RECT  52445.0 87900.0 53150.0 86555.0 ;
      RECT  52445.0 87900.0 53150.0 89245.0 ;
      RECT  52445.0 90590.0 53150.0 89245.0 ;
      RECT  52445.0 90590.0 53150.0 91935.0 ;
      RECT  52445.0 93280.0 53150.0 91935.0 ;
      RECT  52445.0 93280.0 53150.0 94625.0 ;
      RECT  52445.0 95970.0 53150.0 94625.0 ;
      RECT  52445.0 95970.0 53150.0 97315.0 ;
      RECT  52445.0 98660.0 53150.0 97315.0 ;
      RECT  52445.0 98660.0 53150.0 100005.0 ;
      RECT  52445.0 101350.0 53150.0 100005.0 ;
      RECT  52445.0 101350.0 53150.0 102695.0 ;
      RECT  52445.0 104040.0 53150.0 102695.0 ;
      RECT  52445.0 104040.0 53150.0 105385.0 ;
      RECT  52445.0 106730.0 53150.0 105385.0 ;
      RECT  52445.0 106730.0 53150.0 108075.0 ;
      RECT  52445.0 109420.0 53150.0 108075.0 ;
      RECT  52445.0 109420.0 53150.0 110765.0 ;
      RECT  52445.0 112110.0 53150.0 110765.0 ;
      RECT  52445.0 112110.0 53150.0 113455.0 ;
      RECT  52445.0 114800.0 53150.0 113455.0 ;
      RECT  52445.0 114800.0 53150.0 116145.0 ;
      RECT  52445.0 117490.0 53150.0 116145.0 ;
      RECT  52445.0 117490.0 53150.0 118835.0 ;
      RECT  52445.0 120180.0 53150.0 118835.0 ;
      RECT  52445.0 120180.0 53150.0 121525.0 ;
      RECT  52445.0 122870.0 53150.0 121525.0 ;
      RECT  52445.0 122870.0 53150.0 124215.0 ;
      RECT  52445.0 125560.0 53150.0 124215.0 ;
      RECT  52445.0 125560.0 53150.0 126905.0 ;
      RECT  52445.0 128250.0 53150.0 126905.0 ;
      RECT  52445.0 128250.0 53150.0 129595.0 ;
      RECT  52445.0 130940.0 53150.0 129595.0 ;
      RECT  52445.0 130940.0 53150.0 132285.0 ;
      RECT  52445.0 133630.0 53150.0 132285.0 ;
      RECT  52445.0 133630.0 53150.0 134975.0 ;
      RECT  52445.0 136320.0 53150.0 134975.0 ;
      RECT  52445.0 136320.0 53150.0 137665.0 ;
      RECT  52445.0 139010.0 53150.0 137665.0 ;
      RECT  52445.0 139010.0 53150.0 140355.0 ;
      RECT  52445.0 141700.0 53150.0 140355.0 ;
      RECT  52445.0 141700.0 53150.0 143045.0 ;
      RECT  52445.0 144390.0 53150.0 143045.0 ;
      RECT  52445.0 144390.0 53150.0 145735.0 ;
      RECT  52445.0 147080.0 53150.0 145735.0 ;
      RECT  52445.0 147080.0 53150.0 148425.0 ;
      RECT  52445.0 149770.0 53150.0 148425.0 ;
      RECT  52445.0 149770.0 53150.0 151115.0 ;
      RECT  52445.0 152460.0 53150.0 151115.0 ;
      RECT  52445.0 152460.0 53150.0 153805.0 ;
      RECT  52445.0 155150.0 53150.0 153805.0 ;
      RECT  52445.0 155150.0 53150.0 156495.0 ;
      RECT  52445.0 157840.0 53150.0 156495.0 ;
      RECT  52445.0 157840.0 53150.0 159185.0 ;
      RECT  52445.0 160530.0 53150.0 159185.0 ;
      RECT  52445.0 160530.0 53150.0 161875.0 ;
      RECT  52445.0 163220.0 53150.0 161875.0 ;
      RECT  52445.0 163220.0 53150.0 164565.0 ;
      RECT  52445.0 165910.0 53150.0 164565.0 ;
      RECT  52445.0 165910.0 53150.0 167255.0 ;
      RECT  52445.0 168600.0 53150.0 167255.0 ;
      RECT  52445.0 168600.0 53150.0 169945.0 ;
      RECT  52445.0 171290.0 53150.0 169945.0 ;
      RECT  52445.0 171290.0 53150.0 172635.0 ;
      RECT  52445.0 173980.0 53150.0 172635.0 ;
      RECT  52445.0 173980.0 53150.0 175325.0 ;
      RECT  52445.0 176670.0 53150.0 175325.0 ;
      RECT  52445.0 176670.0 53150.0 178015.0 ;
      RECT  52445.0 179360.0 53150.0 178015.0 ;
      RECT  52445.0 179360.0 53150.0 180705.0 ;
      RECT  52445.0 182050.0 53150.0 180705.0 ;
      RECT  52445.0 182050.0 53150.0 183395.0 ;
      RECT  52445.0 184740.0 53150.0 183395.0 ;
      RECT  52445.0 184740.0 53150.0 186085.0 ;
      RECT  52445.0 187430.0 53150.0 186085.0 ;
      RECT  52445.0 187430.0 53150.0 188775.0 ;
      RECT  52445.0 190120.0 53150.0 188775.0 ;
      RECT  52445.0 190120.0 53150.0 191465.0 ;
      RECT  52445.0 192810.0 53150.0 191465.0 ;
      RECT  52445.0 192810.0 53150.0 194155.0 ;
      RECT  52445.0 195500.0 53150.0 194155.0 ;
      RECT  52445.0 195500.0 53150.0 196845.0 ;
      RECT  52445.0 198190.0 53150.0 196845.0 ;
      RECT  52445.0 198190.0 53150.0 199535.0 ;
      RECT  52445.0 200880.0 53150.0 199535.0 ;
      RECT  52445.0 200880.0 53150.0 202225.0 ;
      RECT  52445.0 203570.0 53150.0 202225.0 ;
      RECT  52445.0 203570.0 53150.0 204915.0 ;
      RECT  52445.0 206260.0 53150.0 204915.0 ;
      RECT  53150.0 34100.0 53855.0 35445.0 ;
      RECT  53150.0 36790.0 53855.0 35445.0 ;
      RECT  53150.0 36790.0 53855.0 38135.0 ;
      RECT  53150.0 39480.0 53855.0 38135.0 ;
      RECT  53150.0 39480.0 53855.0 40825.0 ;
      RECT  53150.0 42170.0 53855.0 40825.0 ;
      RECT  53150.0 42170.0 53855.0 43515.0 ;
      RECT  53150.0 44860.0 53855.0 43515.0 ;
      RECT  53150.0 44860.0 53855.0 46205.0 ;
      RECT  53150.0 47550.0 53855.0 46205.0 ;
      RECT  53150.0 47550.0 53855.0 48895.0 ;
      RECT  53150.0 50240.0 53855.0 48895.0 ;
      RECT  53150.0 50240.0 53855.0 51585.0 ;
      RECT  53150.0 52930.0 53855.0 51585.0 ;
      RECT  53150.0 52930.0 53855.0 54275.0 ;
      RECT  53150.0 55620.0 53855.0 54275.0 ;
      RECT  53150.0 55620.0 53855.0 56965.0 ;
      RECT  53150.0 58310.0 53855.0 56965.0 ;
      RECT  53150.0 58310.0 53855.0 59655.0 ;
      RECT  53150.0 61000.0 53855.0 59655.0 ;
      RECT  53150.0 61000.0 53855.0 62345.0 ;
      RECT  53150.0 63690.0 53855.0 62345.0 ;
      RECT  53150.0 63690.0 53855.0 65035.0 ;
      RECT  53150.0 66380.0 53855.0 65035.0 ;
      RECT  53150.0 66380.0 53855.0 67725.0 ;
      RECT  53150.0 69070.0 53855.0 67725.0 ;
      RECT  53150.0 69070.0 53855.0 70415.0 ;
      RECT  53150.0 71760.0 53855.0 70415.0 ;
      RECT  53150.0 71760.0 53855.0 73105.0 ;
      RECT  53150.0 74450.0 53855.0 73105.0 ;
      RECT  53150.0 74450.0 53855.0 75795.0 ;
      RECT  53150.0 77140.0 53855.0 75795.0 ;
      RECT  53150.0 77140.0 53855.0 78485.0 ;
      RECT  53150.0 79830.0 53855.0 78485.0 ;
      RECT  53150.0 79830.0 53855.0 81175.0 ;
      RECT  53150.0 82520.0 53855.0 81175.0 ;
      RECT  53150.0 82520.0 53855.0 83865.0 ;
      RECT  53150.0 85210.0 53855.0 83865.0 ;
      RECT  53150.0 85210.0 53855.0 86555.0 ;
      RECT  53150.0 87900.0 53855.0 86555.0 ;
      RECT  53150.0 87900.0 53855.0 89245.0 ;
      RECT  53150.0 90590.0 53855.0 89245.0 ;
      RECT  53150.0 90590.0 53855.0 91935.0 ;
      RECT  53150.0 93280.0 53855.0 91935.0 ;
      RECT  53150.0 93280.0 53855.0 94625.0 ;
      RECT  53150.0 95970.0 53855.0 94625.0 ;
      RECT  53150.0 95970.0 53855.0 97315.0 ;
      RECT  53150.0 98660.0 53855.0 97315.0 ;
      RECT  53150.0 98660.0 53855.0 100005.0 ;
      RECT  53150.0 101350.0 53855.0 100005.0 ;
      RECT  53150.0 101350.0 53855.0 102695.0 ;
      RECT  53150.0 104040.0 53855.0 102695.0 ;
      RECT  53150.0 104040.0 53855.0 105385.0 ;
      RECT  53150.0 106730.0 53855.0 105385.0 ;
      RECT  53150.0 106730.0 53855.0 108075.0 ;
      RECT  53150.0 109420.0 53855.0 108075.0 ;
      RECT  53150.0 109420.0 53855.0 110765.0 ;
      RECT  53150.0 112110.0 53855.0 110765.0 ;
      RECT  53150.0 112110.0 53855.0 113455.0 ;
      RECT  53150.0 114800.0 53855.0 113455.0 ;
      RECT  53150.0 114800.0 53855.0 116145.0 ;
      RECT  53150.0 117490.0 53855.0 116145.0 ;
      RECT  53150.0 117490.0 53855.0 118835.0 ;
      RECT  53150.0 120180.0 53855.0 118835.0 ;
      RECT  53150.0 120180.0 53855.0 121525.0 ;
      RECT  53150.0 122870.0 53855.0 121525.0 ;
      RECT  53150.0 122870.0 53855.0 124215.0 ;
      RECT  53150.0 125560.0 53855.0 124215.0 ;
      RECT  53150.0 125560.0 53855.0 126905.0 ;
      RECT  53150.0 128250.0 53855.0 126905.0 ;
      RECT  53150.0 128250.0 53855.0 129595.0 ;
      RECT  53150.0 130940.0 53855.0 129595.0 ;
      RECT  53150.0 130940.0 53855.0 132285.0 ;
      RECT  53150.0 133630.0 53855.0 132285.0 ;
      RECT  53150.0 133630.0 53855.0 134975.0 ;
      RECT  53150.0 136320.0 53855.0 134975.0 ;
      RECT  53150.0 136320.0 53855.0 137665.0 ;
      RECT  53150.0 139010.0 53855.0 137665.0 ;
      RECT  53150.0 139010.0 53855.0 140355.0 ;
      RECT  53150.0 141700.0 53855.0 140355.0 ;
      RECT  53150.0 141700.0 53855.0 143045.0 ;
      RECT  53150.0 144390.0 53855.0 143045.0 ;
      RECT  53150.0 144390.0 53855.0 145735.0 ;
      RECT  53150.0 147080.0 53855.0 145735.0 ;
      RECT  53150.0 147080.0 53855.0 148425.0 ;
      RECT  53150.0 149770.0 53855.0 148425.0 ;
      RECT  53150.0 149770.0 53855.0 151115.0 ;
      RECT  53150.0 152460.0 53855.0 151115.0 ;
      RECT  53150.0 152460.0 53855.0 153805.0 ;
      RECT  53150.0 155150.0 53855.0 153805.0 ;
      RECT  53150.0 155150.0 53855.0 156495.0 ;
      RECT  53150.0 157840.0 53855.0 156495.0 ;
      RECT  53150.0 157840.0 53855.0 159185.0 ;
      RECT  53150.0 160530.0 53855.0 159185.0 ;
      RECT  53150.0 160530.0 53855.0 161875.0 ;
      RECT  53150.0 163220.0 53855.0 161875.0 ;
      RECT  53150.0 163220.0 53855.0 164565.0 ;
      RECT  53150.0 165910.0 53855.0 164565.0 ;
      RECT  53150.0 165910.0 53855.0 167255.0 ;
      RECT  53150.0 168600.0 53855.0 167255.0 ;
      RECT  53150.0 168600.0 53855.0 169945.0 ;
      RECT  53150.0 171290.0 53855.0 169945.0 ;
      RECT  53150.0 171290.0 53855.0 172635.0 ;
      RECT  53150.0 173980.0 53855.0 172635.0 ;
      RECT  53150.0 173980.0 53855.0 175325.0 ;
      RECT  53150.0 176670.0 53855.0 175325.0 ;
      RECT  53150.0 176670.0 53855.0 178015.0 ;
      RECT  53150.0 179360.0 53855.0 178015.0 ;
      RECT  53150.0 179360.0 53855.0 180705.0 ;
      RECT  53150.0 182050.0 53855.0 180705.0 ;
      RECT  53150.0 182050.0 53855.0 183395.0 ;
      RECT  53150.0 184740.0 53855.0 183395.0 ;
      RECT  53150.0 184740.0 53855.0 186085.0 ;
      RECT  53150.0 187430.0 53855.0 186085.0 ;
      RECT  53150.0 187430.0 53855.0 188775.0 ;
      RECT  53150.0 190120.0 53855.0 188775.0 ;
      RECT  53150.0 190120.0 53855.0 191465.0 ;
      RECT  53150.0 192810.0 53855.0 191465.0 ;
      RECT  53150.0 192810.0 53855.0 194155.0 ;
      RECT  53150.0 195500.0 53855.0 194155.0 ;
      RECT  53150.0 195500.0 53855.0 196845.0 ;
      RECT  53150.0 198190.0 53855.0 196845.0 ;
      RECT  53150.0 198190.0 53855.0 199535.0 ;
      RECT  53150.0 200880.0 53855.0 199535.0 ;
      RECT  53150.0 200880.0 53855.0 202225.0 ;
      RECT  53150.0 203570.0 53855.0 202225.0 ;
      RECT  53150.0 203570.0 53855.0 204915.0 ;
      RECT  53150.0 206260.0 53855.0 204915.0 ;
      RECT  53855.0 34100.0 54560.0 35445.0 ;
      RECT  53855.0 36790.0 54560.0 35445.0 ;
      RECT  53855.0 36790.0 54560.0 38135.0 ;
      RECT  53855.0 39480.0 54560.0 38135.0 ;
      RECT  53855.0 39480.0 54560.0 40825.0 ;
      RECT  53855.0 42170.0 54560.0 40825.0 ;
      RECT  53855.0 42170.0 54560.0 43515.0 ;
      RECT  53855.0 44860.0 54560.0 43515.0 ;
      RECT  53855.0 44860.0 54560.0 46205.0 ;
      RECT  53855.0 47550.0 54560.0 46205.0 ;
      RECT  53855.0 47550.0 54560.0 48895.0 ;
      RECT  53855.0 50240.0 54560.0 48895.0 ;
      RECT  53855.0 50240.0 54560.0 51585.0 ;
      RECT  53855.0 52930.0 54560.0 51585.0 ;
      RECT  53855.0 52930.0 54560.0 54275.0 ;
      RECT  53855.0 55620.0 54560.0 54275.0 ;
      RECT  53855.0 55620.0 54560.0 56965.0 ;
      RECT  53855.0 58310.0 54560.0 56965.0 ;
      RECT  53855.0 58310.0 54560.0 59655.0 ;
      RECT  53855.0 61000.0 54560.0 59655.0 ;
      RECT  53855.0 61000.0 54560.0 62345.0 ;
      RECT  53855.0 63690.0 54560.0 62345.0 ;
      RECT  53855.0 63690.0 54560.0 65035.0 ;
      RECT  53855.0 66380.0 54560.0 65035.0 ;
      RECT  53855.0 66380.0 54560.0 67725.0 ;
      RECT  53855.0 69070.0 54560.0 67725.0 ;
      RECT  53855.0 69070.0 54560.0 70415.0 ;
      RECT  53855.0 71760.0 54560.0 70415.0 ;
      RECT  53855.0 71760.0 54560.0 73105.0 ;
      RECT  53855.0 74450.0 54560.0 73105.0 ;
      RECT  53855.0 74450.0 54560.0 75795.0 ;
      RECT  53855.0 77140.0 54560.0 75795.0 ;
      RECT  53855.0 77140.0 54560.0 78485.0 ;
      RECT  53855.0 79830.0 54560.0 78485.0 ;
      RECT  53855.0 79830.0 54560.0 81175.0 ;
      RECT  53855.0 82520.0 54560.0 81175.0 ;
      RECT  53855.0 82520.0 54560.0 83865.0 ;
      RECT  53855.0 85210.0 54560.0 83865.0 ;
      RECT  53855.0 85210.0 54560.0 86555.0 ;
      RECT  53855.0 87900.0 54560.0 86555.0 ;
      RECT  53855.0 87900.0 54560.0 89245.0 ;
      RECT  53855.0 90590.0 54560.0 89245.0 ;
      RECT  53855.0 90590.0 54560.0 91935.0 ;
      RECT  53855.0 93280.0 54560.0 91935.0 ;
      RECT  53855.0 93280.0 54560.0 94625.0 ;
      RECT  53855.0 95970.0 54560.0 94625.0 ;
      RECT  53855.0 95970.0 54560.0 97315.0 ;
      RECT  53855.0 98660.0 54560.0 97315.0 ;
      RECT  53855.0 98660.0 54560.0 100005.0 ;
      RECT  53855.0 101350.0 54560.0 100005.0 ;
      RECT  53855.0 101350.0 54560.0 102695.0 ;
      RECT  53855.0 104040.0 54560.0 102695.0 ;
      RECT  53855.0 104040.0 54560.0 105385.0 ;
      RECT  53855.0 106730.0 54560.0 105385.0 ;
      RECT  53855.0 106730.0 54560.0 108075.0 ;
      RECT  53855.0 109420.0 54560.0 108075.0 ;
      RECT  53855.0 109420.0 54560.0 110765.0 ;
      RECT  53855.0 112110.0 54560.0 110765.0 ;
      RECT  53855.0 112110.0 54560.0 113455.0 ;
      RECT  53855.0 114800.0 54560.0 113455.0 ;
      RECT  53855.0 114800.0 54560.0 116145.0 ;
      RECT  53855.0 117490.0 54560.0 116145.0 ;
      RECT  53855.0 117490.0 54560.0 118835.0 ;
      RECT  53855.0 120180.0 54560.0 118835.0 ;
      RECT  53855.0 120180.0 54560.0 121525.0 ;
      RECT  53855.0 122870.0 54560.0 121525.0 ;
      RECT  53855.0 122870.0 54560.0 124215.0 ;
      RECT  53855.0 125560.0 54560.0 124215.0 ;
      RECT  53855.0 125560.0 54560.0 126905.0 ;
      RECT  53855.0 128250.0 54560.0 126905.0 ;
      RECT  53855.0 128250.0 54560.0 129595.0 ;
      RECT  53855.0 130940.0 54560.0 129595.0 ;
      RECT  53855.0 130940.0 54560.0 132285.0 ;
      RECT  53855.0 133630.0 54560.0 132285.0 ;
      RECT  53855.0 133630.0 54560.0 134975.0 ;
      RECT  53855.0 136320.0 54560.0 134975.0 ;
      RECT  53855.0 136320.0 54560.0 137665.0 ;
      RECT  53855.0 139010.0 54560.0 137665.0 ;
      RECT  53855.0 139010.0 54560.0 140355.0 ;
      RECT  53855.0 141700.0 54560.0 140355.0 ;
      RECT  53855.0 141700.0 54560.0 143045.0 ;
      RECT  53855.0 144390.0 54560.0 143045.0 ;
      RECT  53855.0 144390.0 54560.0 145735.0 ;
      RECT  53855.0 147080.0 54560.0 145735.0 ;
      RECT  53855.0 147080.0 54560.0 148425.0 ;
      RECT  53855.0 149770.0 54560.0 148425.0 ;
      RECT  53855.0 149770.0 54560.0 151115.0 ;
      RECT  53855.0 152460.0 54560.0 151115.0 ;
      RECT  53855.0 152460.0 54560.0 153805.0 ;
      RECT  53855.0 155150.0 54560.0 153805.0 ;
      RECT  53855.0 155150.0 54560.0 156495.0 ;
      RECT  53855.0 157840.0 54560.0 156495.0 ;
      RECT  53855.0 157840.0 54560.0 159185.0 ;
      RECT  53855.0 160530.0 54560.0 159185.0 ;
      RECT  53855.0 160530.0 54560.0 161875.0 ;
      RECT  53855.0 163220.0 54560.0 161875.0 ;
      RECT  53855.0 163220.0 54560.0 164565.0 ;
      RECT  53855.0 165910.0 54560.0 164565.0 ;
      RECT  53855.0 165910.0 54560.0 167255.0 ;
      RECT  53855.0 168600.0 54560.0 167255.0 ;
      RECT  53855.0 168600.0 54560.0 169945.0 ;
      RECT  53855.0 171290.0 54560.0 169945.0 ;
      RECT  53855.0 171290.0 54560.0 172635.0 ;
      RECT  53855.0 173980.0 54560.0 172635.0 ;
      RECT  53855.0 173980.0 54560.0 175325.0 ;
      RECT  53855.0 176670.0 54560.0 175325.0 ;
      RECT  53855.0 176670.0 54560.0 178015.0 ;
      RECT  53855.0 179360.0 54560.0 178015.0 ;
      RECT  53855.0 179360.0 54560.0 180705.0 ;
      RECT  53855.0 182050.0 54560.0 180705.0 ;
      RECT  53855.0 182050.0 54560.0 183395.0 ;
      RECT  53855.0 184740.0 54560.0 183395.0 ;
      RECT  53855.0 184740.0 54560.0 186085.0 ;
      RECT  53855.0 187430.0 54560.0 186085.0 ;
      RECT  53855.0 187430.0 54560.0 188775.0 ;
      RECT  53855.0 190120.0 54560.0 188775.0 ;
      RECT  53855.0 190120.0 54560.0 191465.0 ;
      RECT  53855.0 192810.0 54560.0 191465.0 ;
      RECT  53855.0 192810.0 54560.0 194155.0 ;
      RECT  53855.0 195500.0 54560.0 194155.0 ;
      RECT  53855.0 195500.0 54560.0 196845.0 ;
      RECT  53855.0 198190.0 54560.0 196845.0 ;
      RECT  53855.0 198190.0 54560.0 199535.0 ;
      RECT  53855.0 200880.0 54560.0 199535.0 ;
      RECT  53855.0 200880.0 54560.0 202225.0 ;
      RECT  53855.0 203570.0 54560.0 202225.0 ;
      RECT  53855.0 203570.0 54560.0 204915.0 ;
      RECT  53855.0 206260.0 54560.0 204915.0 ;
      RECT  54560.0 34100.0 55265.0 35445.0 ;
      RECT  54560.0 36790.0 55265.0 35445.0 ;
      RECT  54560.0 36790.0 55265.0 38135.0 ;
      RECT  54560.0 39480.0 55265.0 38135.0 ;
      RECT  54560.0 39480.0 55265.0 40825.0 ;
      RECT  54560.0 42170.0 55265.0 40825.0 ;
      RECT  54560.0 42170.0 55265.0 43515.0 ;
      RECT  54560.0 44860.0 55265.0 43515.0 ;
      RECT  54560.0 44860.0 55265.0 46205.0 ;
      RECT  54560.0 47550.0 55265.0 46205.0 ;
      RECT  54560.0 47550.0 55265.0 48895.0 ;
      RECT  54560.0 50240.0 55265.0 48895.0 ;
      RECT  54560.0 50240.0 55265.0 51585.0 ;
      RECT  54560.0 52930.0 55265.0 51585.0 ;
      RECT  54560.0 52930.0 55265.0 54275.0 ;
      RECT  54560.0 55620.0 55265.0 54275.0 ;
      RECT  54560.0 55620.0 55265.0 56965.0 ;
      RECT  54560.0 58310.0 55265.0 56965.0 ;
      RECT  54560.0 58310.0 55265.0 59655.0 ;
      RECT  54560.0 61000.0 55265.0 59655.0 ;
      RECT  54560.0 61000.0 55265.0 62345.0 ;
      RECT  54560.0 63690.0 55265.0 62345.0 ;
      RECT  54560.0 63690.0 55265.0 65035.0 ;
      RECT  54560.0 66380.0 55265.0 65035.0 ;
      RECT  54560.0 66380.0 55265.0 67725.0 ;
      RECT  54560.0 69070.0 55265.0 67725.0 ;
      RECT  54560.0 69070.0 55265.0 70415.0 ;
      RECT  54560.0 71760.0 55265.0 70415.0 ;
      RECT  54560.0 71760.0 55265.0 73105.0 ;
      RECT  54560.0 74450.0 55265.0 73105.0 ;
      RECT  54560.0 74450.0 55265.0 75795.0 ;
      RECT  54560.0 77140.0 55265.0 75795.0 ;
      RECT  54560.0 77140.0 55265.0 78485.0 ;
      RECT  54560.0 79830.0 55265.0 78485.0 ;
      RECT  54560.0 79830.0 55265.0 81175.0 ;
      RECT  54560.0 82520.0 55265.0 81175.0 ;
      RECT  54560.0 82520.0 55265.0 83865.0 ;
      RECT  54560.0 85210.0 55265.0 83865.0 ;
      RECT  54560.0 85210.0 55265.0 86555.0 ;
      RECT  54560.0 87900.0 55265.0 86555.0 ;
      RECT  54560.0 87900.0 55265.0 89245.0 ;
      RECT  54560.0 90590.0 55265.0 89245.0 ;
      RECT  54560.0 90590.0 55265.0 91935.0 ;
      RECT  54560.0 93280.0 55265.0 91935.0 ;
      RECT  54560.0 93280.0 55265.0 94625.0 ;
      RECT  54560.0 95970.0 55265.0 94625.0 ;
      RECT  54560.0 95970.0 55265.0 97315.0 ;
      RECT  54560.0 98660.0 55265.0 97315.0 ;
      RECT  54560.0 98660.0 55265.0 100005.0 ;
      RECT  54560.0 101350.0 55265.0 100005.0 ;
      RECT  54560.0 101350.0 55265.0 102695.0 ;
      RECT  54560.0 104040.0 55265.0 102695.0 ;
      RECT  54560.0 104040.0 55265.0 105385.0 ;
      RECT  54560.0 106730.0 55265.0 105385.0 ;
      RECT  54560.0 106730.0 55265.0 108075.0 ;
      RECT  54560.0 109420.0 55265.0 108075.0 ;
      RECT  54560.0 109420.0 55265.0 110765.0 ;
      RECT  54560.0 112110.0 55265.0 110765.0 ;
      RECT  54560.0 112110.0 55265.0 113455.0 ;
      RECT  54560.0 114800.0 55265.0 113455.0 ;
      RECT  54560.0 114800.0 55265.0 116145.0 ;
      RECT  54560.0 117490.0 55265.0 116145.0 ;
      RECT  54560.0 117490.0 55265.0 118835.0 ;
      RECT  54560.0 120180.0 55265.0 118835.0 ;
      RECT  54560.0 120180.0 55265.0 121525.0 ;
      RECT  54560.0 122870.0 55265.0 121525.0 ;
      RECT  54560.0 122870.0 55265.0 124215.0 ;
      RECT  54560.0 125560.0 55265.0 124215.0 ;
      RECT  54560.0 125560.0 55265.0 126905.0 ;
      RECT  54560.0 128250.0 55265.0 126905.0 ;
      RECT  54560.0 128250.0 55265.0 129595.0 ;
      RECT  54560.0 130940.0 55265.0 129595.0 ;
      RECT  54560.0 130940.0 55265.0 132285.0 ;
      RECT  54560.0 133630.0 55265.0 132285.0 ;
      RECT  54560.0 133630.0 55265.0 134975.0 ;
      RECT  54560.0 136320.0 55265.0 134975.0 ;
      RECT  54560.0 136320.0 55265.0 137665.0 ;
      RECT  54560.0 139010.0 55265.0 137665.0 ;
      RECT  54560.0 139010.0 55265.0 140355.0 ;
      RECT  54560.0 141700.0 55265.0 140355.0 ;
      RECT  54560.0 141700.0 55265.0 143045.0 ;
      RECT  54560.0 144390.0 55265.0 143045.0 ;
      RECT  54560.0 144390.0 55265.0 145735.0 ;
      RECT  54560.0 147080.0 55265.0 145735.0 ;
      RECT  54560.0 147080.0 55265.0 148425.0 ;
      RECT  54560.0 149770.0 55265.0 148425.0 ;
      RECT  54560.0 149770.0 55265.0 151115.0 ;
      RECT  54560.0 152460.0 55265.0 151115.0 ;
      RECT  54560.0 152460.0 55265.0 153805.0 ;
      RECT  54560.0 155150.0 55265.0 153805.0 ;
      RECT  54560.0 155150.0 55265.0 156495.0 ;
      RECT  54560.0 157840.0 55265.0 156495.0 ;
      RECT  54560.0 157840.0 55265.0 159185.0 ;
      RECT  54560.0 160530.0 55265.0 159185.0 ;
      RECT  54560.0 160530.0 55265.0 161875.0 ;
      RECT  54560.0 163220.0 55265.0 161875.0 ;
      RECT  54560.0 163220.0 55265.0 164565.0 ;
      RECT  54560.0 165910.0 55265.0 164565.0 ;
      RECT  54560.0 165910.0 55265.0 167255.0 ;
      RECT  54560.0 168600.0 55265.0 167255.0 ;
      RECT  54560.0 168600.0 55265.0 169945.0 ;
      RECT  54560.0 171290.0 55265.0 169945.0 ;
      RECT  54560.0 171290.0 55265.0 172635.0 ;
      RECT  54560.0 173980.0 55265.0 172635.0 ;
      RECT  54560.0 173980.0 55265.0 175325.0 ;
      RECT  54560.0 176670.0 55265.0 175325.0 ;
      RECT  54560.0 176670.0 55265.0 178015.0 ;
      RECT  54560.0 179360.0 55265.0 178015.0 ;
      RECT  54560.0 179360.0 55265.0 180705.0 ;
      RECT  54560.0 182050.0 55265.0 180705.0 ;
      RECT  54560.0 182050.0 55265.0 183395.0 ;
      RECT  54560.0 184740.0 55265.0 183395.0 ;
      RECT  54560.0 184740.0 55265.0 186085.0 ;
      RECT  54560.0 187430.0 55265.0 186085.0 ;
      RECT  54560.0 187430.0 55265.0 188775.0 ;
      RECT  54560.0 190120.0 55265.0 188775.0 ;
      RECT  54560.0 190120.0 55265.0 191465.0 ;
      RECT  54560.0 192810.0 55265.0 191465.0 ;
      RECT  54560.0 192810.0 55265.0 194155.0 ;
      RECT  54560.0 195500.0 55265.0 194155.0 ;
      RECT  54560.0 195500.0 55265.0 196845.0 ;
      RECT  54560.0 198190.0 55265.0 196845.0 ;
      RECT  54560.0 198190.0 55265.0 199535.0 ;
      RECT  54560.0 200880.0 55265.0 199535.0 ;
      RECT  54560.0 200880.0 55265.0 202225.0 ;
      RECT  54560.0 203570.0 55265.0 202225.0 ;
      RECT  54560.0 203570.0 55265.0 204915.0 ;
      RECT  54560.0 206260.0 55265.0 204915.0 ;
      RECT  55265.0 34100.0 55970.0 35445.0 ;
      RECT  55265.0 36790.0 55970.0 35445.0 ;
      RECT  55265.0 36790.0 55970.0 38135.0 ;
      RECT  55265.0 39480.0 55970.0 38135.0 ;
      RECT  55265.0 39480.0 55970.0 40825.0 ;
      RECT  55265.0 42170.0 55970.0 40825.0 ;
      RECT  55265.0 42170.0 55970.0 43515.0 ;
      RECT  55265.0 44860.0 55970.0 43515.0 ;
      RECT  55265.0 44860.0 55970.0 46205.0 ;
      RECT  55265.0 47550.0 55970.0 46205.0 ;
      RECT  55265.0 47550.0 55970.0 48895.0 ;
      RECT  55265.0 50240.0 55970.0 48895.0 ;
      RECT  55265.0 50240.0 55970.0 51585.0 ;
      RECT  55265.0 52930.0 55970.0 51585.0 ;
      RECT  55265.0 52930.0 55970.0 54275.0 ;
      RECT  55265.0 55620.0 55970.0 54275.0 ;
      RECT  55265.0 55620.0 55970.0 56965.0 ;
      RECT  55265.0 58310.0 55970.0 56965.0 ;
      RECT  55265.0 58310.0 55970.0 59655.0 ;
      RECT  55265.0 61000.0 55970.0 59655.0 ;
      RECT  55265.0 61000.0 55970.0 62345.0 ;
      RECT  55265.0 63690.0 55970.0 62345.0 ;
      RECT  55265.0 63690.0 55970.0 65035.0 ;
      RECT  55265.0 66380.0 55970.0 65035.0 ;
      RECT  55265.0 66380.0 55970.0 67725.0 ;
      RECT  55265.0 69070.0 55970.0 67725.0 ;
      RECT  55265.0 69070.0 55970.0 70415.0 ;
      RECT  55265.0 71760.0 55970.0 70415.0 ;
      RECT  55265.0 71760.0 55970.0 73105.0 ;
      RECT  55265.0 74450.0 55970.0 73105.0 ;
      RECT  55265.0 74450.0 55970.0 75795.0 ;
      RECT  55265.0 77140.0 55970.0 75795.0 ;
      RECT  55265.0 77140.0 55970.0 78485.0 ;
      RECT  55265.0 79830.0 55970.0 78485.0 ;
      RECT  55265.0 79830.0 55970.0 81175.0 ;
      RECT  55265.0 82520.0 55970.0 81175.0 ;
      RECT  55265.0 82520.0 55970.0 83865.0 ;
      RECT  55265.0 85210.0 55970.0 83865.0 ;
      RECT  55265.0 85210.0 55970.0 86555.0 ;
      RECT  55265.0 87900.0 55970.0 86555.0 ;
      RECT  55265.0 87900.0 55970.0 89245.0 ;
      RECT  55265.0 90590.0 55970.0 89245.0 ;
      RECT  55265.0 90590.0 55970.0 91935.0 ;
      RECT  55265.0 93280.0 55970.0 91935.0 ;
      RECT  55265.0 93280.0 55970.0 94625.0 ;
      RECT  55265.0 95970.0 55970.0 94625.0 ;
      RECT  55265.0 95970.0 55970.0 97315.0 ;
      RECT  55265.0 98660.0 55970.0 97315.0 ;
      RECT  55265.0 98660.0 55970.0 100005.0 ;
      RECT  55265.0 101350.0 55970.0 100005.0 ;
      RECT  55265.0 101350.0 55970.0 102695.0 ;
      RECT  55265.0 104040.0 55970.0 102695.0 ;
      RECT  55265.0 104040.0 55970.0 105385.0 ;
      RECT  55265.0 106730.0 55970.0 105385.0 ;
      RECT  55265.0 106730.0 55970.0 108075.0 ;
      RECT  55265.0 109420.0 55970.0 108075.0 ;
      RECT  55265.0 109420.0 55970.0 110765.0 ;
      RECT  55265.0 112110.0 55970.0 110765.0 ;
      RECT  55265.0 112110.0 55970.0 113455.0 ;
      RECT  55265.0 114800.0 55970.0 113455.0 ;
      RECT  55265.0 114800.0 55970.0 116145.0 ;
      RECT  55265.0 117490.0 55970.0 116145.0 ;
      RECT  55265.0 117490.0 55970.0 118835.0 ;
      RECT  55265.0 120180.0 55970.0 118835.0 ;
      RECT  55265.0 120180.0 55970.0 121525.0 ;
      RECT  55265.0 122870.0 55970.0 121525.0 ;
      RECT  55265.0 122870.0 55970.0 124215.0 ;
      RECT  55265.0 125560.0 55970.0 124215.0 ;
      RECT  55265.0 125560.0 55970.0 126905.0 ;
      RECT  55265.0 128250.0 55970.0 126905.0 ;
      RECT  55265.0 128250.0 55970.0 129595.0 ;
      RECT  55265.0 130940.0 55970.0 129595.0 ;
      RECT  55265.0 130940.0 55970.0 132285.0 ;
      RECT  55265.0 133630.0 55970.0 132285.0 ;
      RECT  55265.0 133630.0 55970.0 134975.0 ;
      RECT  55265.0 136320.0 55970.0 134975.0 ;
      RECT  55265.0 136320.0 55970.0 137665.0 ;
      RECT  55265.0 139010.0 55970.0 137665.0 ;
      RECT  55265.0 139010.0 55970.0 140355.0 ;
      RECT  55265.0 141700.0 55970.0 140355.0 ;
      RECT  55265.0 141700.0 55970.0 143045.0 ;
      RECT  55265.0 144390.0 55970.0 143045.0 ;
      RECT  55265.0 144390.0 55970.0 145735.0 ;
      RECT  55265.0 147080.0 55970.0 145735.0 ;
      RECT  55265.0 147080.0 55970.0 148425.0 ;
      RECT  55265.0 149770.0 55970.0 148425.0 ;
      RECT  55265.0 149770.0 55970.0 151115.0 ;
      RECT  55265.0 152460.0 55970.0 151115.0 ;
      RECT  55265.0 152460.0 55970.0 153805.0 ;
      RECT  55265.0 155150.0 55970.0 153805.0 ;
      RECT  55265.0 155150.0 55970.0 156495.0 ;
      RECT  55265.0 157840.0 55970.0 156495.0 ;
      RECT  55265.0 157840.0 55970.0 159185.0 ;
      RECT  55265.0 160530.0 55970.0 159185.0 ;
      RECT  55265.0 160530.0 55970.0 161875.0 ;
      RECT  55265.0 163220.0 55970.0 161875.0 ;
      RECT  55265.0 163220.0 55970.0 164565.0 ;
      RECT  55265.0 165910.0 55970.0 164565.0 ;
      RECT  55265.0 165910.0 55970.0 167255.0 ;
      RECT  55265.0 168600.0 55970.0 167255.0 ;
      RECT  55265.0 168600.0 55970.0 169945.0 ;
      RECT  55265.0 171290.0 55970.0 169945.0 ;
      RECT  55265.0 171290.0 55970.0 172635.0 ;
      RECT  55265.0 173980.0 55970.0 172635.0 ;
      RECT  55265.0 173980.0 55970.0 175325.0 ;
      RECT  55265.0 176670.0 55970.0 175325.0 ;
      RECT  55265.0 176670.0 55970.0 178015.0 ;
      RECT  55265.0 179360.0 55970.0 178015.0 ;
      RECT  55265.0 179360.0 55970.0 180705.0 ;
      RECT  55265.0 182050.0 55970.0 180705.0 ;
      RECT  55265.0 182050.0 55970.0 183395.0 ;
      RECT  55265.0 184740.0 55970.0 183395.0 ;
      RECT  55265.0 184740.0 55970.0 186085.0 ;
      RECT  55265.0 187430.0 55970.0 186085.0 ;
      RECT  55265.0 187430.0 55970.0 188775.0 ;
      RECT  55265.0 190120.0 55970.0 188775.0 ;
      RECT  55265.0 190120.0 55970.0 191465.0 ;
      RECT  55265.0 192810.0 55970.0 191465.0 ;
      RECT  55265.0 192810.0 55970.0 194155.0 ;
      RECT  55265.0 195500.0 55970.0 194155.0 ;
      RECT  55265.0 195500.0 55970.0 196845.0 ;
      RECT  55265.0 198190.0 55970.0 196845.0 ;
      RECT  55265.0 198190.0 55970.0 199535.0 ;
      RECT  55265.0 200880.0 55970.0 199535.0 ;
      RECT  55265.0 200880.0 55970.0 202225.0 ;
      RECT  55265.0 203570.0 55970.0 202225.0 ;
      RECT  55265.0 203570.0 55970.0 204915.0 ;
      RECT  55265.0 206260.0 55970.0 204915.0 ;
      RECT  55970.0 34100.0 56675.0 35445.0 ;
      RECT  55970.0 36790.0 56675.0 35445.0 ;
      RECT  55970.0 36790.0 56675.0 38135.0 ;
      RECT  55970.0 39480.0 56675.0 38135.0 ;
      RECT  55970.0 39480.0 56675.0 40825.0 ;
      RECT  55970.0 42170.0 56675.0 40825.0 ;
      RECT  55970.0 42170.0 56675.0 43515.0 ;
      RECT  55970.0 44860.0 56675.0 43515.0 ;
      RECT  55970.0 44860.0 56675.0 46205.0 ;
      RECT  55970.0 47550.0 56675.0 46205.0 ;
      RECT  55970.0 47550.0 56675.0 48895.0 ;
      RECT  55970.0 50240.0 56675.0 48895.0 ;
      RECT  55970.0 50240.0 56675.0 51585.0 ;
      RECT  55970.0 52930.0 56675.0 51585.0 ;
      RECT  55970.0 52930.0 56675.0 54275.0 ;
      RECT  55970.0 55620.0 56675.0 54275.0 ;
      RECT  55970.0 55620.0 56675.0 56965.0 ;
      RECT  55970.0 58310.0 56675.0 56965.0 ;
      RECT  55970.0 58310.0 56675.0 59655.0 ;
      RECT  55970.0 61000.0 56675.0 59655.0 ;
      RECT  55970.0 61000.0 56675.0 62345.0 ;
      RECT  55970.0 63690.0 56675.0 62345.0 ;
      RECT  55970.0 63690.0 56675.0 65035.0 ;
      RECT  55970.0 66380.0 56675.0 65035.0 ;
      RECT  55970.0 66380.0 56675.0 67725.0 ;
      RECT  55970.0 69070.0 56675.0 67725.0 ;
      RECT  55970.0 69070.0 56675.0 70415.0 ;
      RECT  55970.0 71760.0 56675.0 70415.0 ;
      RECT  55970.0 71760.0 56675.0 73105.0 ;
      RECT  55970.0 74450.0 56675.0 73105.0 ;
      RECT  55970.0 74450.0 56675.0 75795.0 ;
      RECT  55970.0 77140.0 56675.0 75795.0 ;
      RECT  55970.0 77140.0 56675.0 78485.0 ;
      RECT  55970.0 79830.0 56675.0 78485.0 ;
      RECT  55970.0 79830.0 56675.0 81175.0 ;
      RECT  55970.0 82520.0 56675.0 81175.0 ;
      RECT  55970.0 82520.0 56675.0 83865.0 ;
      RECT  55970.0 85210.0 56675.0 83865.0 ;
      RECT  55970.0 85210.0 56675.0 86555.0 ;
      RECT  55970.0 87900.0 56675.0 86555.0 ;
      RECT  55970.0 87900.0 56675.0 89245.0 ;
      RECT  55970.0 90590.0 56675.0 89245.0 ;
      RECT  55970.0 90590.0 56675.0 91935.0 ;
      RECT  55970.0 93280.0 56675.0 91935.0 ;
      RECT  55970.0 93280.0 56675.0 94625.0 ;
      RECT  55970.0 95970.0 56675.0 94625.0 ;
      RECT  55970.0 95970.0 56675.0 97315.0 ;
      RECT  55970.0 98660.0 56675.0 97315.0 ;
      RECT  55970.0 98660.0 56675.0 100005.0 ;
      RECT  55970.0 101350.0 56675.0 100005.0 ;
      RECT  55970.0 101350.0 56675.0 102695.0 ;
      RECT  55970.0 104040.0 56675.0 102695.0 ;
      RECT  55970.0 104040.0 56675.0 105385.0 ;
      RECT  55970.0 106730.0 56675.0 105385.0 ;
      RECT  55970.0 106730.0 56675.0 108075.0 ;
      RECT  55970.0 109420.0 56675.0 108075.0 ;
      RECT  55970.0 109420.0 56675.0 110765.0 ;
      RECT  55970.0 112110.0 56675.0 110765.0 ;
      RECT  55970.0 112110.0 56675.0 113455.0 ;
      RECT  55970.0 114800.0 56675.0 113455.0 ;
      RECT  55970.0 114800.0 56675.0 116145.0 ;
      RECT  55970.0 117490.0 56675.0 116145.0 ;
      RECT  55970.0 117490.0 56675.0 118835.0 ;
      RECT  55970.0 120180.0 56675.0 118835.0 ;
      RECT  55970.0 120180.0 56675.0 121525.0 ;
      RECT  55970.0 122870.0 56675.0 121525.0 ;
      RECT  55970.0 122870.0 56675.0 124215.0 ;
      RECT  55970.0 125560.0 56675.0 124215.0 ;
      RECT  55970.0 125560.0 56675.0 126905.0 ;
      RECT  55970.0 128250.0 56675.0 126905.0 ;
      RECT  55970.0 128250.0 56675.0 129595.0 ;
      RECT  55970.0 130940.0 56675.0 129595.0 ;
      RECT  55970.0 130940.0 56675.0 132285.0 ;
      RECT  55970.0 133630.0 56675.0 132285.0 ;
      RECT  55970.0 133630.0 56675.0 134975.0 ;
      RECT  55970.0 136320.0 56675.0 134975.0 ;
      RECT  55970.0 136320.0 56675.0 137665.0 ;
      RECT  55970.0 139010.0 56675.0 137665.0 ;
      RECT  55970.0 139010.0 56675.0 140355.0 ;
      RECT  55970.0 141700.0 56675.0 140355.0 ;
      RECT  55970.0 141700.0 56675.0 143045.0 ;
      RECT  55970.0 144390.0 56675.0 143045.0 ;
      RECT  55970.0 144390.0 56675.0 145735.0 ;
      RECT  55970.0 147080.0 56675.0 145735.0 ;
      RECT  55970.0 147080.0 56675.0 148425.0 ;
      RECT  55970.0 149770.0 56675.0 148425.0 ;
      RECT  55970.0 149770.0 56675.0 151115.0 ;
      RECT  55970.0 152460.0 56675.0 151115.0 ;
      RECT  55970.0 152460.0 56675.0 153805.0 ;
      RECT  55970.0 155150.0 56675.0 153805.0 ;
      RECT  55970.0 155150.0 56675.0 156495.0 ;
      RECT  55970.0 157840.0 56675.0 156495.0 ;
      RECT  55970.0 157840.0 56675.0 159185.0 ;
      RECT  55970.0 160530.0 56675.0 159185.0 ;
      RECT  55970.0 160530.0 56675.0 161875.0 ;
      RECT  55970.0 163220.0 56675.0 161875.0 ;
      RECT  55970.0 163220.0 56675.0 164565.0 ;
      RECT  55970.0 165910.0 56675.0 164565.0 ;
      RECT  55970.0 165910.0 56675.0 167255.0 ;
      RECT  55970.0 168600.0 56675.0 167255.0 ;
      RECT  55970.0 168600.0 56675.0 169945.0 ;
      RECT  55970.0 171290.0 56675.0 169945.0 ;
      RECT  55970.0 171290.0 56675.0 172635.0 ;
      RECT  55970.0 173980.0 56675.0 172635.0 ;
      RECT  55970.0 173980.0 56675.0 175325.0 ;
      RECT  55970.0 176670.0 56675.0 175325.0 ;
      RECT  55970.0 176670.0 56675.0 178015.0 ;
      RECT  55970.0 179360.0 56675.0 178015.0 ;
      RECT  55970.0 179360.0 56675.0 180705.0 ;
      RECT  55970.0 182050.0 56675.0 180705.0 ;
      RECT  55970.0 182050.0 56675.0 183395.0 ;
      RECT  55970.0 184740.0 56675.0 183395.0 ;
      RECT  55970.0 184740.0 56675.0 186085.0 ;
      RECT  55970.0 187430.0 56675.0 186085.0 ;
      RECT  55970.0 187430.0 56675.0 188775.0 ;
      RECT  55970.0 190120.0 56675.0 188775.0 ;
      RECT  55970.0 190120.0 56675.0 191465.0 ;
      RECT  55970.0 192810.0 56675.0 191465.0 ;
      RECT  55970.0 192810.0 56675.0 194155.0 ;
      RECT  55970.0 195500.0 56675.0 194155.0 ;
      RECT  55970.0 195500.0 56675.0 196845.0 ;
      RECT  55970.0 198190.0 56675.0 196845.0 ;
      RECT  55970.0 198190.0 56675.0 199535.0 ;
      RECT  55970.0 200880.0 56675.0 199535.0 ;
      RECT  55970.0 200880.0 56675.0 202225.0 ;
      RECT  55970.0 203570.0 56675.0 202225.0 ;
      RECT  55970.0 203570.0 56675.0 204915.0 ;
      RECT  55970.0 206260.0 56675.0 204915.0 ;
      RECT  56675.0 34100.0 57380.0 35445.0 ;
      RECT  56675.0 36790.0 57380.0 35445.0 ;
      RECT  56675.0 36790.0 57380.0 38135.0 ;
      RECT  56675.0 39480.0 57380.0 38135.0 ;
      RECT  56675.0 39480.0 57380.0 40825.0 ;
      RECT  56675.0 42170.0 57380.0 40825.0 ;
      RECT  56675.0 42170.0 57380.0 43515.0 ;
      RECT  56675.0 44860.0 57380.0 43515.0 ;
      RECT  56675.0 44860.0 57380.0 46205.0 ;
      RECT  56675.0 47550.0 57380.0 46205.0 ;
      RECT  56675.0 47550.0 57380.0 48895.0 ;
      RECT  56675.0 50240.0 57380.0 48895.0 ;
      RECT  56675.0 50240.0 57380.0 51585.0 ;
      RECT  56675.0 52930.0 57380.0 51585.0 ;
      RECT  56675.0 52930.0 57380.0 54275.0 ;
      RECT  56675.0 55620.0 57380.0 54275.0 ;
      RECT  56675.0 55620.0 57380.0 56965.0 ;
      RECT  56675.0 58310.0 57380.0 56965.0 ;
      RECT  56675.0 58310.0 57380.0 59655.0 ;
      RECT  56675.0 61000.0 57380.0 59655.0 ;
      RECT  56675.0 61000.0 57380.0 62345.0 ;
      RECT  56675.0 63690.0 57380.0 62345.0 ;
      RECT  56675.0 63690.0 57380.0 65035.0 ;
      RECT  56675.0 66380.0 57380.0 65035.0 ;
      RECT  56675.0 66380.0 57380.0 67725.0 ;
      RECT  56675.0 69070.0 57380.0 67725.0 ;
      RECT  56675.0 69070.0 57380.0 70415.0 ;
      RECT  56675.0 71760.0 57380.0 70415.0 ;
      RECT  56675.0 71760.0 57380.0 73105.0 ;
      RECT  56675.0 74450.0 57380.0 73105.0 ;
      RECT  56675.0 74450.0 57380.0 75795.0 ;
      RECT  56675.0 77140.0 57380.0 75795.0 ;
      RECT  56675.0 77140.0 57380.0 78485.0 ;
      RECT  56675.0 79830.0 57380.0 78485.0 ;
      RECT  56675.0 79830.0 57380.0 81175.0 ;
      RECT  56675.0 82520.0 57380.0 81175.0 ;
      RECT  56675.0 82520.0 57380.0 83865.0 ;
      RECT  56675.0 85210.0 57380.0 83865.0 ;
      RECT  56675.0 85210.0 57380.0 86555.0 ;
      RECT  56675.0 87900.0 57380.0 86555.0 ;
      RECT  56675.0 87900.0 57380.0 89245.0 ;
      RECT  56675.0 90590.0 57380.0 89245.0 ;
      RECT  56675.0 90590.0 57380.0 91935.0 ;
      RECT  56675.0 93280.0 57380.0 91935.0 ;
      RECT  56675.0 93280.0 57380.0 94625.0 ;
      RECT  56675.0 95970.0 57380.0 94625.0 ;
      RECT  56675.0 95970.0 57380.0 97315.0 ;
      RECT  56675.0 98660.0 57380.0 97315.0 ;
      RECT  56675.0 98660.0 57380.0 100005.0 ;
      RECT  56675.0 101350.0 57380.0 100005.0 ;
      RECT  56675.0 101350.0 57380.0 102695.0 ;
      RECT  56675.0 104040.0 57380.0 102695.0 ;
      RECT  56675.0 104040.0 57380.0 105385.0 ;
      RECT  56675.0 106730.0 57380.0 105385.0 ;
      RECT  56675.0 106730.0 57380.0 108075.0 ;
      RECT  56675.0 109420.0 57380.0 108075.0 ;
      RECT  56675.0 109420.0 57380.0 110765.0 ;
      RECT  56675.0 112110.0 57380.0 110765.0 ;
      RECT  56675.0 112110.0 57380.0 113455.0 ;
      RECT  56675.0 114800.0 57380.0 113455.0 ;
      RECT  56675.0 114800.0 57380.0 116145.0 ;
      RECT  56675.0 117490.0 57380.0 116145.0 ;
      RECT  56675.0 117490.0 57380.0 118835.0 ;
      RECT  56675.0 120180.0 57380.0 118835.0 ;
      RECT  56675.0 120180.0 57380.0 121525.0 ;
      RECT  56675.0 122870.0 57380.0 121525.0 ;
      RECT  56675.0 122870.0 57380.0 124215.0 ;
      RECT  56675.0 125560.0 57380.0 124215.0 ;
      RECT  56675.0 125560.0 57380.0 126905.0 ;
      RECT  56675.0 128250.0 57380.0 126905.0 ;
      RECT  56675.0 128250.0 57380.0 129595.0 ;
      RECT  56675.0 130940.0 57380.0 129595.0 ;
      RECT  56675.0 130940.0 57380.0 132285.0 ;
      RECT  56675.0 133630.0 57380.0 132285.0 ;
      RECT  56675.0 133630.0 57380.0 134975.0 ;
      RECT  56675.0 136320.0 57380.0 134975.0 ;
      RECT  56675.0 136320.0 57380.0 137665.0 ;
      RECT  56675.0 139010.0 57380.0 137665.0 ;
      RECT  56675.0 139010.0 57380.0 140355.0 ;
      RECT  56675.0 141700.0 57380.0 140355.0 ;
      RECT  56675.0 141700.0 57380.0 143045.0 ;
      RECT  56675.0 144390.0 57380.0 143045.0 ;
      RECT  56675.0 144390.0 57380.0 145735.0 ;
      RECT  56675.0 147080.0 57380.0 145735.0 ;
      RECT  56675.0 147080.0 57380.0 148425.0 ;
      RECT  56675.0 149770.0 57380.0 148425.0 ;
      RECT  56675.0 149770.0 57380.0 151115.0 ;
      RECT  56675.0 152460.0 57380.0 151115.0 ;
      RECT  56675.0 152460.0 57380.0 153805.0 ;
      RECT  56675.0 155150.0 57380.0 153805.0 ;
      RECT  56675.0 155150.0 57380.0 156495.0 ;
      RECT  56675.0 157840.0 57380.0 156495.0 ;
      RECT  56675.0 157840.0 57380.0 159185.0 ;
      RECT  56675.0 160530.0 57380.0 159185.0 ;
      RECT  56675.0 160530.0 57380.0 161875.0 ;
      RECT  56675.0 163220.0 57380.0 161875.0 ;
      RECT  56675.0 163220.0 57380.0 164565.0 ;
      RECT  56675.0 165910.0 57380.0 164565.0 ;
      RECT  56675.0 165910.0 57380.0 167255.0 ;
      RECT  56675.0 168600.0 57380.0 167255.0 ;
      RECT  56675.0 168600.0 57380.0 169945.0 ;
      RECT  56675.0 171290.0 57380.0 169945.0 ;
      RECT  56675.0 171290.0 57380.0 172635.0 ;
      RECT  56675.0 173980.0 57380.0 172635.0 ;
      RECT  56675.0 173980.0 57380.0 175325.0 ;
      RECT  56675.0 176670.0 57380.0 175325.0 ;
      RECT  56675.0 176670.0 57380.0 178015.0 ;
      RECT  56675.0 179360.0 57380.0 178015.0 ;
      RECT  56675.0 179360.0 57380.0 180705.0 ;
      RECT  56675.0 182050.0 57380.0 180705.0 ;
      RECT  56675.0 182050.0 57380.0 183395.0 ;
      RECT  56675.0 184740.0 57380.0 183395.0 ;
      RECT  56675.0 184740.0 57380.0 186085.0 ;
      RECT  56675.0 187430.0 57380.0 186085.0 ;
      RECT  56675.0 187430.0 57380.0 188775.0 ;
      RECT  56675.0 190120.0 57380.0 188775.0 ;
      RECT  56675.0 190120.0 57380.0 191465.0 ;
      RECT  56675.0 192810.0 57380.0 191465.0 ;
      RECT  56675.0 192810.0 57380.0 194155.0 ;
      RECT  56675.0 195500.0 57380.0 194155.0 ;
      RECT  56675.0 195500.0 57380.0 196845.0 ;
      RECT  56675.0 198190.0 57380.0 196845.0 ;
      RECT  56675.0 198190.0 57380.0 199535.0 ;
      RECT  56675.0 200880.0 57380.0 199535.0 ;
      RECT  56675.0 200880.0 57380.0 202225.0 ;
      RECT  56675.0 203570.0 57380.0 202225.0 ;
      RECT  56675.0 203570.0 57380.0 204915.0 ;
      RECT  56675.0 206260.0 57380.0 204915.0 ;
      RECT  57380.0 34100.0 58085.0 35445.0 ;
      RECT  57380.0 36790.0 58085.0 35445.0 ;
      RECT  57380.0 36790.0 58085.0 38135.0 ;
      RECT  57380.0 39480.0 58085.0 38135.0 ;
      RECT  57380.0 39480.0 58085.0 40825.0 ;
      RECT  57380.0 42170.0 58085.0 40825.0 ;
      RECT  57380.0 42170.0 58085.0 43515.0 ;
      RECT  57380.0 44860.0 58085.0 43515.0 ;
      RECT  57380.0 44860.0 58085.0 46205.0 ;
      RECT  57380.0 47550.0 58085.0 46205.0 ;
      RECT  57380.0 47550.0 58085.0 48895.0 ;
      RECT  57380.0 50240.0 58085.0 48895.0 ;
      RECT  57380.0 50240.0 58085.0 51585.0 ;
      RECT  57380.0 52930.0 58085.0 51585.0 ;
      RECT  57380.0 52930.0 58085.0 54275.0 ;
      RECT  57380.0 55620.0 58085.0 54275.0 ;
      RECT  57380.0 55620.0 58085.0 56965.0 ;
      RECT  57380.0 58310.0 58085.0 56965.0 ;
      RECT  57380.0 58310.0 58085.0 59655.0 ;
      RECT  57380.0 61000.0 58085.0 59655.0 ;
      RECT  57380.0 61000.0 58085.0 62345.0 ;
      RECT  57380.0 63690.0 58085.0 62345.0 ;
      RECT  57380.0 63690.0 58085.0 65035.0 ;
      RECT  57380.0 66380.0 58085.0 65035.0 ;
      RECT  57380.0 66380.0 58085.0 67725.0 ;
      RECT  57380.0 69070.0 58085.0 67725.0 ;
      RECT  57380.0 69070.0 58085.0 70415.0 ;
      RECT  57380.0 71760.0 58085.0 70415.0 ;
      RECT  57380.0 71760.0 58085.0 73105.0 ;
      RECT  57380.0 74450.0 58085.0 73105.0 ;
      RECT  57380.0 74450.0 58085.0 75795.0 ;
      RECT  57380.0 77140.0 58085.0 75795.0 ;
      RECT  57380.0 77140.0 58085.0 78485.0 ;
      RECT  57380.0 79830.0 58085.0 78485.0 ;
      RECT  57380.0 79830.0 58085.0 81175.0 ;
      RECT  57380.0 82520.0 58085.0 81175.0 ;
      RECT  57380.0 82520.0 58085.0 83865.0 ;
      RECT  57380.0 85210.0 58085.0 83865.0 ;
      RECT  57380.0 85210.0 58085.0 86555.0 ;
      RECT  57380.0 87900.0 58085.0 86555.0 ;
      RECT  57380.0 87900.0 58085.0 89245.0 ;
      RECT  57380.0 90590.0 58085.0 89245.0 ;
      RECT  57380.0 90590.0 58085.0 91935.0 ;
      RECT  57380.0 93280.0 58085.0 91935.0 ;
      RECT  57380.0 93280.0 58085.0 94625.0 ;
      RECT  57380.0 95970.0 58085.0 94625.0 ;
      RECT  57380.0 95970.0 58085.0 97315.0 ;
      RECT  57380.0 98660.0 58085.0 97315.0 ;
      RECT  57380.0 98660.0 58085.0 100005.0 ;
      RECT  57380.0 101350.0 58085.0 100005.0 ;
      RECT  57380.0 101350.0 58085.0 102695.0 ;
      RECT  57380.0 104040.0 58085.0 102695.0 ;
      RECT  57380.0 104040.0 58085.0 105385.0 ;
      RECT  57380.0 106730.0 58085.0 105385.0 ;
      RECT  57380.0 106730.0 58085.0 108075.0 ;
      RECT  57380.0 109420.0 58085.0 108075.0 ;
      RECT  57380.0 109420.0 58085.0 110765.0 ;
      RECT  57380.0 112110.0 58085.0 110765.0 ;
      RECT  57380.0 112110.0 58085.0 113455.0 ;
      RECT  57380.0 114800.0 58085.0 113455.0 ;
      RECT  57380.0 114800.0 58085.0 116145.0 ;
      RECT  57380.0 117490.0 58085.0 116145.0 ;
      RECT  57380.0 117490.0 58085.0 118835.0 ;
      RECT  57380.0 120180.0 58085.0 118835.0 ;
      RECT  57380.0 120180.0 58085.0 121525.0 ;
      RECT  57380.0 122870.0 58085.0 121525.0 ;
      RECT  57380.0 122870.0 58085.0 124215.0 ;
      RECT  57380.0 125560.0 58085.0 124215.0 ;
      RECT  57380.0 125560.0 58085.0 126905.0 ;
      RECT  57380.0 128250.0 58085.0 126905.0 ;
      RECT  57380.0 128250.0 58085.0 129595.0 ;
      RECT  57380.0 130940.0 58085.0 129595.0 ;
      RECT  57380.0 130940.0 58085.0 132285.0 ;
      RECT  57380.0 133630.0 58085.0 132285.0 ;
      RECT  57380.0 133630.0 58085.0 134975.0 ;
      RECT  57380.0 136320.0 58085.0 134975.0 ;
      RECT  57380.0 136320.0 58085.0 137665.0 ;
      RECT  57380.0 139010.0 58085.0 137665.0 ;
      RECT  57380.0 139010.0 58085.0 140355.0 ;
      RECT  57380.0 141700.0 58085.0 140355.0 ;
      RECT  57380.0 141700.0 58085.0 143045.0 ;
      RECT  57380.0 144390.0 58085.0 143045.0 ;
      RECT  57380.0 144390.0 58085.0 145735.0 ;
      RECT  57380.0 147080.0 58085.0 145735.0 ;
      RECT  57380.0 147080.0 58085.0 148425.0 ;
      RECT  57380.0 149770.0 58085.0 148425.0 ;
      RECT  57380.0 149770.0 58085.0 151115.0 ;
      RECT  57380.0 152460.0 58085.0 151115.0 ;
      RECT  57380.0 152460.0 58085.0 153805.0 ;
      RECT  57380.0 155150.0 58085.0 153805.0 ;
      RECT  57380.0 155150.0 58085.0 156495.0 ;
      RECT  57380.0 157840.0 58085.0 156495.0 ;
      RECT  57380.0 157840.0 58085.0 159185.0 ;
      RECT  57380.0 160530.0 58085.0 159185.0 ;
      RECT  57380.0 160530.0 58085.0 161875.0 ;
      RECT  57380.0 163220.0 58085.0 161875.0 ;
      RECT  57380.0 163220.0 58085.0 164565.0 ;
      RECT  57380.0 165910.0 58085.0 164565.0 ;
      RECT  57380.0 165910.0 58085.0 167255.0 ;
      RECT  57380.0 168600.0 58085.0 167255.0 ;
      RECT  57380.0 168600.0 58085.0 169945.0 ;
      RECT  57380.0 171290.0 58085.0 169945.0 ;
      RECT  57380.0 171290.0 58085.0 172635.0 ;
      RECT  57380.0 173980.0 58085.0 172635.0 ;
      RECT  57380.0 173980.0 58085.0 175325.0 ;
      RECT  57380.0 176670.0 58085.0 175325.0 ;
      RECT  57380.0 176670.0 58085.0 178015.0 ;
      RECT  57380.0 179360.0 58085.0 178015.0 ;
      RECT  57380.0 179360.0 58085.0 180705.0 ;
      RECT  57380.0 182050.0 58085.0 180705.0 ;
      RECT  57380.0 182050.0 58085.0 183395.0 ;
      RECT  57380.0 184740.0 58085.0 183395.0 ;
      RECT  57380.0 184740.0 58085.0 186085.0 ;
      RECT  57380.0 187430.0 58085.0 186085.0 ;
      RECT  57380.0 187430.0 58085.0 188775.0 ;
      RECT  57380.0 190120.0 58085.0 188775.0 ;
      RECT  57380.0 190120.0 58085.0 191465.0 ;
      RECT  57380.0 192810.0 58085.0 191465.0 ;
      RECT  57380.0 192810.0 58085.0 194155.0 ;
      RECT  57380.0 195500.0 58085.0 194155.0 ;
      RECT  57380.0 195500.0 58085.0 196845.0 ;
      RECT  57380.0 198190.0 58085.0 196845.0 ;
      RECT  57380.0 198190.0 58085.0 199535.0 ;
      RECT  57380.0 200880.0 58085.0 199535.0 ;
      RECT  57380.0 200880.0 58085.0 202225.0 ;
      RECT  57380.0 203570.0 58085.0 202225.0 ;
      RECT  57380.0 203570.0 58085.0 204915.0 ;
      RECT  57380.0 206260.0 58085.0 204915.0 ;
      RECT  58085.0 34100.0 58790.0 35445.0 ;
      RECT  58085.0 36790.0 58790.0 35445.0 ;
      RECT  58085.0 36790.0 58790.0 38135.0 ;
      RECT  58085.0 39480.0 58790.0 38135.0 ;
      RECT  58085.0 39480.0 58790.0 40825.0 ;
      RECT  58085.0 42170.0 58790.0 40825.0 ;
      RECT  58085.0 42170.0 58790.0 43515.0 ;
      RECT  58085.0 44860.0 58790.0 43515.0 ;
      RECT  58085.0 44860.0 58790.0 46205.0 ;
      RECT  58085.0 47550.0 58790.0 46205.0 ;
      RECT  58085.0 47550.0 58790.0 48895.0 ;
      RECT  58085.0 50240.0 58790.0 48895.0 ;
      RECT  58085.0 50240.0 58790.0 51585.0 ;
      RECT  58085.0 52930.0 58790.0 51585.0 ;
      RECT  58085.0 52930.0 58790.0 54275.0 ;
      RECT  58085.0 55620.0 58790.0 54275.0 ;
      RECT  58085.0 55620.0 58790.0 56965.0 ;
      RECT  58085.0 58310.0 58790.0 56965.0 ;
      RECT  58085.0 58310.0 58790.0 59655.0 ;
      RECT  58085.0 61000.0 58790.0 59655.0 ;
      RECT  58085.0 61000.0 58790.0 62345.0 ;
      RECT  58085.0 63690.0 58790.0 62345.0 ;
      RECT  58085.0 63690.0 58790.0 65035.0 ;
      RECT  58085.0 66380.0 58790.0 65035.0 ;
      RECT  58085.0 66380.0 58790.0 67725.0 ;
      RECT  58085.0 69070.0 58790.0 67725.0 ;
      RECT  58085.0 69070.0 58790.0 70415.0 ;
      RECT  58085.0 71760.0 58790.0 70415.0 ;
      RECT  58085.0 71760.0 58790.0 73105.0 ;
      RECT  58085.0 74450.0 58790.0 73105.0 ;
      RECT  58085.0 74450.0 58790.0 75795.0 ;
      RECT  58085.0 77140.0 58790.0 75795.0 ;
      RECT  58085.0 77140.0 58790.0 78485.0 ;
      RECT  58085.0 79830.0 58790.0 78485.0 ;
      RECT  58085.0 79830.0 58790.0 81175.0 ;
      RECT  58085.0 82520.0 58790.0 81175.0 ;
      RECT  58085.0 82520.0 58790.0 83865.0 ;
      RECT  58085.0 85210.0 58790.0 83865.0 ;
      RECT  58085.0 85210.0 58790.0 86555.0 ;
      RECT  58085.0 87900.0 58790.0 86555.0 ;
      RECT  58085.0 87900.0 58790.0 89245.0 ;
      RECT  58085.0 90590.0 58790.0 89245.0 ;
      RECT  58085.0 90590.0 58790.0 91935.0 ;
      RECT  58085.0 93280.0 58790.0 91935.0 ;
      RECT  58085.0 93280.0 58790.0 94625.0 ;
      RECT  58085.0 95970.0 58790.0 94625.0 ;
      RECT  58085.0 95970.0 58790.0 97315.0 ;
      RECT  58085.0 98660.0 58790.0 97315.0 ;
      RECT  58085.0 98660.0 58790.0 100005.0 ;
      RECT  58085.0 101350.0 58790.0 100005.0 ;
      RECT  58085.0 101350.0 58790.0 102695.0 ;
      RECT  58085.0 104040.0 58790.0 102695.0 ;
      RECT  58085.0 104040.0 58790.0 105385.0 ;
      RECT  58085.0 106730.0 58790.0 105385.0 ;
      RECT  58085.0 106730.0 58790.0 108075.0 ;
      RECT  58085.0 109420.0 58790.0 108075.0 ;
      RECT  58085.0 109420.0 58790.0 110765.0 ;
      RECT  58085.0 112110.0 58790.0 110765.0 ;
      RECT  58085.0 112110.0 58790.0 113455.0 ;
      RECT  58085.0 114800.0 58790.0 113455.0 ;
      RECT  58085.0 114800.0 58790.0 116145.0 ;
      RECT  58085.0 117490.0 58790.0 116145.0 ;
      RECT  58085.0 117490.0 58790.0 118835.0 ;
      RECT  58085.0 120180.0 58790.0 118835.0 ;
      RECT  58085.0 120180.0 58790.0 121525.0 ;
      RECT  58085.0 122870.0 58790.0 121525.0 ;
      RECT  58085.0 122870.0 58790.0 124215.0 ;
      RECT  58085.0 125560.0 58790.0 124215.0 ;
      RECT  58085.0 125560.0 58790.0 126905.0 ;
      RECT  58085.0 128250.0 58790.0 126905.0 ;
      RECT  58085.0 128250.0 58790.0 129595.0 ;
      RECT  58085.0 130940.0 58790.0 129595.0 ;
      RECT  58085.0 130940.0 58790.0 132285.0 ;
      RECT  58085.0 133630.0 58790.0 132285.0 ;
      RECT  58085.0 133630.0 58790.0 134975.0 ;
      RECT  58085.0 136320.0 58790.0 134975.0 ;
      RECT  58085.0 136320.0 58790.0 137665.0 ;
      RECT  58085.0 139010.0 58790.0 137665.0 ;
      RECT  58085.0 139010.0 58790.0 140355.0 ;
      RECT  58085.0 141700.0 58790.0 140355.0 ;
      RECT  58085.0 141700.0 58790.0 143045.0 ;
      RECT  58085.0 144390.0 58790.0 143045.0 ;
      RECT  58085.0 144390.0 58790.0 145735.0 ;
      RECT  58085.0 147080.0 58790.0 145735.0 ;
      RECT  58085.0 147080.0 58790.0 148425.0 ;
      RECT  58085.0 149770.0 58790.0 148425.0 ;
      RECT  58085.0 149770.0 58790.0 151115.0 ;
      RECT  58085.0 152460.0 58790.0 151115.0 ;
      RECT  58085.0 152460.0 58790.0 153805.0 ;
      RECT  58085.0 155150.0 58790.0 153805.0 ;
      RECT  58085.0 155150.0 58790.0 156495.0 ;
      RECT  58085.0 157840.0 58790.0 156495.0 ;
      RECT  58085.0 157840.0 58790.0 159185.0 ;
      RECT  58085.0 160530.0 58790.0 159185.0 ;
      RECT  58085.0 160530.0 58790.0 161875.0 ;
      RECT  58085.0 163220.0 58790.0 161875.0 ;
      RECT  58085.0 163220.0 58790.0 164565.0 ;
      RECT  58085.0 165910.0 58790.0 164565.0 ;
      RECT  58085.0 165910.0 58790.0 167255.0 ;
      RECT  58085.0 168600.0 58790.0 167255.0 ;
      RECT  58085.0 168600.0 58790.0 169945.0 ;
      RECT  58085.0 171290.0 58790.0 169945.0 ;
      RECT  58085.0 171290.0 58790.0 172635.0 ;
      RECT  58085.0 173980.0 58790.0 172635.0 ;
      RECT  58085.0 173980.0 58790.0 175325.0 ;
      RECT  58085.0 176670.0 58790.0 175325.0 ;
      RECT  58085.0 176670.0 58790.0 178015.0 ;
      RECT  58085.0 179360.0 58790.0 178015.0 ;
      RECT  58085.0 179360.0 58790.0 180705.0 ;
      RECT  58085.0 182050.0 58790.0 180705.0 ;
      RECT  58085.0 182050.0 58790.0 183395.0 ;
      RECT  58085.0 184740.0 58790.0 183395.0 ;
      RECT  58085.0 184740.0 58790.0 186085.0 ;
      RECT  58085.0 187430.0 58790.0 186085.0 ;
      RECT  58085.0 187430.0 58790.0 188775.0 ;
      RECT  58085.0 190120.0 58790.0 188775.0 ;
      RECT  58085.0 190120.0 58790.0 191465.0 ;
      RECT  58085.0 192810.0 58790.0 191465.0 ;
      RECT  58085.0 192810.0 58790.0 194155.0 ;
      RECT  58085.0 195500.0 58790.0 194155.0 ;
      RECT  58085.0 195500.0 58790.0 196845.0 ;
      RECT  58085.0 198190.0 58790.0 196845.0 ;
      RECT  58085.0 198190.0 58790.0 199535.0 ;
      RECT  58085.0 200880.0 58790.0 199535.0 ;
      RECT  58085.0 200880.0 58790.0 202225.0 ;
      RECT  58085.0 203570.0 58790.0 202225.0 ;
      RECT  58085.0 203570.0 58790.0 204915.0 ;
      RECT  58085.0 206260.0 58790.0 204915.0 ;
      RECT  58790.0 34100.0 59495.0 35445.0 ;
      RECT  58790.0 36790.0 59495.0 35445.0 ;
      RECT  58790.0 36790.0 59495.0 38135.0 ;
      RECT  58790.0 39480.0 59495.0 38135.0 ;
      RECT  58790.0 39480.0 59495.0 40825.0 ;
      RECT  58790.0 42170.0 59495.0 40825.0 ;
      RECT  58790.0 42170.0 59495.0 43515.0 ;
      RECT  58790.0 44860.0 59495.0 43515.0 ;
      RECT  58790.0 44860.0 59495.0 46205.0 ;
      RECT  58790.0 47550.0 59495.0 46205.0 ;
      RECT  58790.0 47550.0 59495.0 48895.0 ;
      RECT  58790.0 50240.0 59495.0 48895.0 ;
      RECT  58790.0 50240.0 59495.0 51585.0 ;
      RECT  58790.0 52930.0 59495.0 51585.0 ;
      RECT  58790.0 52930.0 59495.0 54275.0 ;
      RECT  58790.0 55620.0 59495.0 54275.0 ;
      RECT  58790.0 55620.0 59495.0 56965.0 ;
      RECT  58790.0 58310.0 59495.0 56965.0 ;
      RECT  58790.0 58310.0 59495.0 59655.0 ;
      RECT  58790.0 61000.0 59495.0 59655.0 ;
      RECT  58790.0 61000.0 59495.0 62345.0 ;
      RECT  58790.0 63690.0 59495.0 62345.0 ;
      RECT  58790.0 63690.0 59495.0 65035.0 ;
      RECT  58790.0 66380.0 59495.0 65035.0 ;
      RECT  58790.0 66380.0 59495.0 67725.0 ;
      RECT  58790.0 69070.0 59495.0 67725.0 ;
      RECT  58790.0 69070.0 59495.0 70415.0 ;
      RECT  58790.0 71760.0 59495.0 70415.0 ;
      RECT  58790.0 71760.0 59495.0 73105.0 ;
      RECT  58790.0 74450.0 59495.0 73105.0 ;
      RECT  58790.0 74450.0 59495.0 75795.0 ;
      RECT  58790.0 77140.0 59495.0 75795.0 ;
      RECT  58790.0 77140.0 59495.0 78485.0 ;
      RECT  58790.0 79830.0 59495.0 78485.0 ;
      RECT  58790.0 79830.0 59495.0 81175.0 ;
      RECT  58790.0 82520.0 59495.0 81175.0 ;
      RECT  58790.0 82520.0 59495.0 83865.0 ;
      RECT  58790.0 85210.0 59495.0 83865.0 ;
      RECT  58790.0 85210.0 59495.0 86555.0 ;
      RECT  58790.0 87900.0 59495.0 86555.0 ;
      RECT  58790.0 87900.0 59495.0 89245.0 ;
      RECT  58790.0 90590.0 59495.0 89245.0 ;
      RECT  58790.0 90590.0 59495.0 91935.0 ;
      RECT  58790.0 93280.0 59495.0 91935.0 ;
      RECT  58790.0 93280.0 59495.0 94625.0 ;
      RECT  58790.0 95970.0 59495.0 94625.0 ;
      RECT  58790.0 95970.0 59495.0 97315.0 ;
      RECT  58790.0 98660.0 59495.0 97315.0 ;
      RECT  58790.0 98660.0 59495.0 100005.0 ;
      RECT  58790.0 101350.0 59495.0 100005.0 ;
      RECT  58790.0 101350.0 59495.0 102695.0 ;
      RECT  58790.0 104040.0 59495.0 102695.0 ;
      RECT  58790.0 104040.0 59495.0 105385.0 ;
      RECT  58790.0 106730.0 59495.0 105385.0 ;
      RECT  58790.0 106730.0 59495.0 108075.0 ;
      RECT  58790.0 109420.0 59495.0 108075.0 ;
      RECT  58790.0 109420.0 59495.0 110765.0 ;
      RECT  58790.0 112110.0 59495.0 110765.0 ;
      RECT  58790.0 112110.0 59495.0 113455.0 ;
      RECT  58790.0 114800.0 59495.0 113455.0 ;
      RECT  58790.0 114800.0 59495.0 116145.0 ;
      RECT  58790.0 117490.0 59495.0 116145.0 ;
      RECT  58790.0 117490.0 59495.0 118835.0 ;
      RECT  58790.0 120180.0 59495.0 118835.0 ;
      RECT  58790.0 120180.0 59495.0 121525.0 ;
      RECT  58790.0 122870.0 59495.0 121525.0 ;
      RECT  58790.0 122870.0 59495.0 124215.0 ;
      RECT  58790.0 125560.0 59495.0 124215.0 ;
      RECT  58790.0 125560.0 59495.0 126905.0 ;
      RECT  58790.0 128250.0 59495.0 126905.0 ;
      RECT  58790.0 128250.0 59495.0 129595.0 ;
      RECT  58790.0 130940.0 59495.0 129595.0 ;
      RECT  58790.0 130940.0 59495.0 132285.0 ;
      RECT  58790.0 133630.0 59495.0 132285.0 ;
      RECT  58790.0 133630.0 59495.0 134975.0 ;
      RECT  58790.0 136320.0 59495.0 134975.0 ;
      RECT  58790.0 136320.0 59495.0 137665.0 ;
      RECT  58790.0 139010.0 59495.0 137665.0 ;
      RECT  58790.0 139010.0 59495.0 140355.0 ;
      RECT  58790.0 141700.0 59495.0 140355.0 ;
      RECT  58790.0 141700.0 59495.0 143045.0 ;
      RECT  58790.0 144390.0 59495.0 143045.0 ;
      RECT  58790.0 144390.0 59495.0 145735.0 ;
      RECT  58790.0 147080.0 59495.0 145735.0 ;
      RECT  58790.0 147080.0 59495.0 148425.0 ;
      RECT  58790.0 149770.0 59495.0 148425.0 ;
      RECT  58790.0 149770.0 59495.0 151115.0 ;
      RECT  58790.0 152460.0 59495.0 151115.0 ;
      RECT  58790.0 152460.0 59495.0 153805.0 ;
      RECT  58790.0 155150.0 59495.0 153805.0 ;
      RECT  58790.0 155150.0 59495.0 156495.0 ;
      RECT  58790.0 157840.0 59495.0 156495.0 ;
      RECT  58790.0 157840.0 59495.0 159185.0 ;
      RECT  58790.0 160530.0 59495.0 159185.0 ;
      RECT  58790.0 160530.0 59495.0 161875.0 ;
      RECT  58790.0 163220.0 59495.0 161875.0 ;
      RECT  58790.0 163220.0 59495.0 164565.0 ;
      RECT  58790.0 165910.0 59495.0 164565.0 ;
      RECT  58790.0 165910.0 59495.0 167255.0 ;
      RECT  58790.0 168600.0 59495.0 167255.0 ;
      RECT  58790.0 168600.0 59495.0 169945.0 ;
      RECT  58790.0 171290.0 59495.0 169945.0 ;
      RECT  58790.0 171290.0 59495.0 172635.0 ;
      RECT  58790.0 173980.0 59495.0 172635.0 ;
      RECT  58790.0 173980.0 59495.0 175325.0 ;
      RECT  58790.0 176670.0 59495.0 175325.0 ;
      RECT  58790.0 176670.0 59495.0 178015.0 ;
      RECT  58790.0 179360.0 59495.0 178015.0 ;
      RECT  58790.0 179360.0 59495.0 180705.0 ;
      RECT  58790.0 182050.0 59495.0 180705.0 ;
      RECT  58790.0 182050.0 59495.0 183395.0 ;
      RECT  58790.0 184740.0 59495.0 183395.0 ;
      RECT  58790.0 184740.0 59495.0 186085.0 ;
      RECT  58790.0 187430.0 59495.0 186085.0 ;
      RECT  58790.0 187430.0 59495.0 188775.0 ;
      RECT  58790.0 190120.0 59495.0 188775.0 ;
      RECT  58790.0 190120.0 59495.0 191465.0 ;
      RECT  58790.0 192810.0 59495.0 191465.0 ;
      RECT  58790.0 192810.0 59495.0 194155.0 ;
      RECT  58790.0 195500.0 59495.0 194155.0 ;
      RECT  58790.0 195500.0 59495.0 196845.0 ;
      RECT  58790.0 198190.0 59495.0 196845.0 ;
      RECT  58790.0 198190.0 59495.0 199535.0 ;
      RECT  58790.0 200880.0 59495.0 199535.0 ;
      RECT  58790.0 200880.0 59495.0 202225.0 ;
      RECT  58790.0 203570.0 59495.0 202225.0 ;
      RECT  58790.0 203570.0 59495.0 204915.0 ;
      RECT  58790.0 206260.0 59495.0 204915.0 ;
      RECT  59495.0 34100.0 60200.0 35445.0 ;
      RECT  59495.0 36790.0 60200.0 35445.0 ;
      RECT  59495.0 36790.0 60200.0 38135.0 ;
      RECT  59495.0 39480.0 60200.0 38135.0 ;
      RECT  59495.0 39480.0 60200.0 40825.0 ;
      RECT  59495.0 42170.0 60200.0 40825.0 ;
      RECT  59495.0 42170.0 60200.0 43515.0 ;
      RECT  59495.0 44860.0 60200.0 43515.0 ;
      RECT  59495.0 44860.0 60200.0 46205.0 ;
      RECT  59495.0 47550.0 60200.0 46205.0 ;
      RECT  59495.0 47550.0 60200.0 48895.0 ;
      RECT  59495.0 50240.0 60200.0 48895.0 ;
      RECT  59495.0 50240.0 60200.0 51585.0 ;
      RECT  59495.0 52930.0 60200.0 51585.0 ;
      RECT  59495.0 52930.0 60200.0 54275.0 ;
      RECT  59495.0 55620.0 60200.0 54275.0 ;
      RECT  59495.0 55620.0 60200.0 56965.0 ;
      RECT  59495.0 58310.0 60200.0 56965.0 ;
      RECT  59495.0 58310.0 60200.0 59655.0 ;
      RECT  59495.0 61000.0 60200.0 59655.0 ;
      RECT  59495.0 61000.0 60200.0 62345.0 ;
      RECT  59495.0 63690.0 60200.0 62345.0 ;
      RECT  59495.0 63690.0 60200.0 65035.0 ;
      RECT  59495.0 66380.0 60200.0 65035.0 ;
      RECT  59495.0 66380.0 60200.0 67725.0 ;
      RECT  59495.0 69070.0 60200.0 67725.0 ;
      RECT  59495.0 69070.0 60200.0 70415.0 ;
      RECT  59495.0 71760.0 60200.0 70415.0 ;
      RECT  59495.0 71760.0 60200.0 73105.0 ;
      RECT  59495.0 74450.0 60200.0 73105.0 ;
      RECT  59495.0 74450.0 60200.0 75795.0 ;
      RECT  59495.0 77140.0 60200.0 75795.0 ;
      RECT  59495.0 77140.0 60200.0 78485.0 ;
      RECT  59495.0 79830.0 60200.0 78485.0 ;
      RECT  59495.0 79830.0 60200.0 81175.0 ;
      RECT  59495.0 82520.0 60200.0 81175.0 ;
      RECT  59495.0 82520.0 60200.0 83865.0 ;
      RECT  59495.0 85210.0 60200.0 83865.0 ;
      RECT  59495.0 85210.0 60200.0 86555.0 ;
      RECT  59495.0 87900.0 60200.0 86555.0 ;
      RECT  59495.0 87900.0 60200.0 89245.0 ;
      RECT  59495.0 90590.0 60200.0 89245.0 ;
      RECT  59495.0 90590.0 60200.0 91935.0 ;
      RECT  59495.0 93280.0 60200.0 91935.0 ;
      RECT  59495.0 93280.0 60200.0 94625.0 ;
      RECT  59495.0 95970.0 60200.0 94625.0 ;
      RECT  59495.0 95970.0 60200.0 97315.0 ;
      RECT  59495.0 98660.0 60200.0 97315.0 ;
      RECT  59495.0 98660.0 60200.0 100005.0 ;
      RECT  59495.0 101350.0 60200.0 100005.0 ;
      RECT  59495.0 101350.0 60200.0 102695.0 ;
      RECT  59495.0 104040.0 60200.0 102695.0 ;
      RECT  59495.0 104040.0 60200.0 105385.0 ;
      RECT  59495.0 106730.0 60200.0 105385.0 ;
      RECT  59495.0 106730.0 60200.0 108075.0 ;
      RECT  59495.0 109420.0 60200.0 108075.0 ;
      RECT  59495.0 109420.0 60200.0 110765.0 ;
      RECT  59495.0 112110.0 60200.0 110765.0 ;
      RECT  59495.0 112110.0 60200.0 113455.0 ;
      RECT  59495.0 114800.0 60200.0 113455.0 ;
      RECT  59495.0 114800.0 60200.0 116145.0 ;
      RECT  59495.0 117490.0 60200.0 116145.0 ;
      RECT  59495.0 117490.0 60200.0 118835.0 ;
      RECT  59495.0 120180.0 60200.0 118835.0 ;
      RECT  59495.0 120180.0 60200.0 121525.0 ;
      RECT  59495.0 122870.0 60200.0 121525.0 ;
      RECT  59495.0 122870.0 60200.0 124215.0 ;
      RECT  59495.0 125560.0 60200.0 124215.0 ;
      RECT  59495.0 125560.0 60200.0 126905.0 ;
      RECT  59495.0 128250.0 60200.0 126905.0 ;
      RECT  59495.0 128250.0 60200.0 129595.0 ;
      RECT  59495.0 130940.0 60200.0 129595.0 ;
      RECT  59495.0 130940.0 60200.0 132285.0 ;
      RECT  59495.0 133630.0 60200.0 132285.0 ;
      RECT  59495.0 133630.0 60200.0 134975.0 ;
      RECT  59495.0 136320.0 60200.0 134975.0 ;
      RECT  59495.0 136320.0 60200.0 137665.0 ;
      RECT  59495.0 139010.0 60200.0 137665.0 ;
      RECT  59495.0 139010.0 60200.0 140355.0 ;
      RECT  59495.0 141700.0 60200.0 140355.0 ;
      RECT  59495.0 141700.0 60200.0 143045.0 ;
      RECT  59495.0 144390.0 60200.0 143045.0 ;
      RECT  59495.0 144390.0 60200.0 145735.0 ;
      RECT  59495.0 147080.0 60200.0 145735.0 ;
      RECT  59495.0 147080.0 60200.0 148425.0 ;
      RECT  59495.0 149770.0 60200.0 148425.0 ;
      RECT  59495.0 149770.0 60200.0 151115.0 ;
      RECT  59495.0 152460.0 60200.0 151115.0 ;
      RECT  59495.0 152460.0 60200.0 153805.0 ;
      RECT  59495.0 155150.0 60200.0 153805.0 ;
      RECT  59495.0 155150.0 60200.0 156495.0 ;
      RECT  59495.0 157840.0 60200.0 156495.0 ;
      RECT  59495.0 157840.0 60200.0 159185.0 ;
      RECT  59495.0 160530.0 60200.0 159185.0 ;
      RECT  59495.0 160530.0 60200.0 161875.0 ;
      RECT  59495.0 163220.0 60200.0 161875.0 ;
      RECT  59495.0 163220.0 60200.0 164565.0 ;
      RECT  59495.0 165910.0 60200.0 164565.0 ;
      RECT  59495.0 165910.0 60200.0 167255.0 ;
      RECT  59495.0 168600.0 60200.0 167255.0 ;
      RECT  59495.0 168600.0 60200.0 169945.0 ;
      RECT  59495.0 171290.0 60200.0 169945.0 ;
      RECT  59495.0 171290.0 60200.0 172635.0 ;
      RECT  59495.0 173980.0 60200.0 172635.0 ;
      RECT  59495.0 173980.0 60200.0 175325.0 ;
      RECT  59495.0 176670.0 60200.0 175325.0 ;
      RECT  59495.0 176670.0 60200.0 178015.0 ;
      RECT  59495.0 179360.0 60200.0 178015.0 ;
      RECT  59495.0 179360.0 60200.0 180705.0 ;
      RECT  59495.0 182050.0 60200.0 180705.0 ;
      RECT  59495.0 182050.0 60200.0 183395.0 ;
      RECT  59495.0 184740.0 60200.0 183395.0 ;
      RECT  59495.0 184740.0 60200.0 186085.0 ;
      RECT  59495.0 187430.0 60200.0 186085.0 ;
      RECT  59495.0 187430.0 60200.0 188775.0 ;
      RECT  59495.0 190120.0 60200.0 188775.0 ;
      RECT  59495.0 190120.0 60200.0 191465.0 ;
      RECT  59495.0 192810.0 60200.0 191465.0 ;
      RECT  59495.0 192810.0 60200.0 194155.0 ;
      RECT  59495.0 195500.0 60200.0 194155.0 ;
      RECT  59495.0 195500.0 60200.0 196845.0 ;
      RECT  59495.0 198190.0 60200.0 196845.0 ;
      RECT  59495.0 198190.0 60200.0 199535.0 ;
      RECT  59495.0 200880.0 60200.0 199535.0 ;
      RECT  59495.0 200880.0 60200.0 202225.0 ;
      RECT  59495.0 203570.0 60200.0 202225.0 ;
      RECT  59495.0 203570.0 60200.0 204915.0 ;
      RECT  59495.0 206260.0 60200.0 204915.0 ;
      RECT  60200.0 34100.0 60905.0 35445.0 ;
      RECT  60200.0 36790.0 60905.0 35445.0 ;
      RECT  60200.0 36790.0 60905.0 38135.0 ;
      RECT  60200.0 39480.0 60905.0 38135.0 ;
      RECT  60200.0 39480.0 60905.0 40825.0 ;
      RECT  60200.0 42170.0 60905.0 40825.0 ;
      RECT  60200.0 42170.0 60905.0 43515.0 ;
      RECT  60200.0 44860.0 60905.0 43515.0 ;
      RECT  60200.0 44860.0 60905.0 46205.0 ;
      RECT  60200.0 47550.0 60905.0 46205.0 ;
      RECT  60200.0 47550.0 60905.0 48895.0 ;
      RECT  60200.0 50240.0 60905.0 48895.0 ;
      RECT  60200.0 50240.0 60905.0 51585.0 ;
      RECT  60200.0 52930.0 60905.0 51585.0 ;
      RECT  60200.0 52930.0 60905.0 54275.0 ;
      RECT  60200.0 55620.0 60905.0 54275.0 ;
      RECT  60200.0 55620.0 60905.0 56965.0 ;
      RECT  60200.0 58310.0 60905.0 56965.0 ;
      RECT  60200.0 58310.0 60905.0 59655.0 ;
      RECT  60200.0 61000.0 60905.0 59655.0 ;
      RECT  60200.0 61000.0 60905.0 62345.0 ;
      RECT  60200.0 63690.0 60905.0 62345.0 ;
      RECT  60200.0 63690.0 60905.0 65035.0 ;
      RECT  60200.0 66380.0 60905.0 65035.0 ;
      RECT  60200.0 66380.0 60905.0 67725.0 ;
      RECT  60200.0 69070.0 60905.0 67725.0 ;
      RECT  60200.0 69070.0 60905.0 70415.0 ;
      RECT  60200.0 71760.0 60905.0 70415.0 ;
      RECT  60200.0 71760.0 60905.0 73105.0 ;
      RECT  60200.0 74450.0 60905.0 73105.0 ;
      RECT  60200.0 74450.0 60905.0 75795.0 ;
      RECT  60200.0 77140.0 60905.0 75795.0 ;
      RECT  60200.0 77140.0 60905.0 78485.0 ;
      RECT  60200.0 79830.0 60905.0 78485.0 ;
      RECT  60200.0 79830.0 60905.0 81175.0 ;
      RECT  60200.0 82520.0 60905.0 81175.0 ;
      RECT  60200.0 82520.0 60905.0 83865.0 ;
      RECT  60200.0 85210.0 60905.0 83865.0 ;
      RECT  60200.0 85210.0 60905.0 86555.0 ;
      RECT  60200.0 87900.0 60905.0 86555.0 ;
      RECT  60200.0 87900.0 60905.0 89245.0 ;
      RECT  60200.0 90590.0 60905.0 89245.0 ;
      RECT  60200.0 90590.0 60905.0 91935.0 ;
      RECT  60200.0 93280.0 60905.0 91935.0 ;
      RECT  60200.0 93280.0 60905.0 94625.0 ;
      RECT  60200.0 95970.0 60905.0 94625.0 ;
      RECT  60200.0 95970.0 60905.0 97315.0 ;
      RECT  60200.0 98660.0 60905.0 97315.0 ;
      RECT  60200.0 98660.0 60905.0 100005.0 ;
      RECT  60200.0 101350.0 60905.0 100005.0 ;
      RECT  60200.0 101350.0 60905.0 102695.0 ;
      RECT  60200.0 104040.0 60905.0 102695.0 ;
      RECT  60200.0 104040.0 60905.0 105385.0 ;
      RECT  60200.0 106730.0 60905.0 105385.0 ;
      RECT  60200.0 106730.0 60905.0 108075.0 ;
      RECT  60200.0 109420.0 60905.0 108075.0 ;
      RECT  60200.0 109420.0 60905.0 110765.0 ;
      RECT  60200.0 112110.0 60905.0 110765.0 ;
      RECT  60200.0 112110.0 60905.0 113455.0 ;
      RECT  60200.0 114800.0 60905.0 113455.0 ;
      RECT  60200.0 114800.0 60905.0 116145.0 ;
      RECT  60200.0 117490.0 60905.0 116145.0 ;
      RECT  60200.0 117490.0 60905.0 118835.0 ;
      RECT  60200.0 120180.0 60905.0 118835.0 ;
      RECT  60200.0 120180.0 60905.0 121525.0 ;
      RECT  60200.0 122870.0 60905.0 121525.0 ;
      RECT  60200.0 122870.0 60905.0 124215.0 ;
      RECT  60200.0 125560.0 60905.0 124215.0 ;
      RECT  60200.0 125560.0 60905.0 126905.0 ;
      RECT  60200.0 128250.0 60905.0 126905.0 ;
      RECT  60200.0 128250.0 60905.0 129595.0 ;
      RECT  60200.0 130940.0 60905.0 129595.0 ;
      RECT  60200.0 130940.0 60905.0 132285.0 ;
      RECT  60200.0 133630.0 60905.0 132285.0 ;
      RECT  60200.0 133630.0 60905.0 134975.0 ;
      RECT  60200.0 136320.0 60905.0 134975.0 ;
      RECT  60200.0 136320.0 60905.0 137665.0 ;
      RECT  60200.0 139010.0 60905.0 137665.0 ;
      RECT  60200.0 139010.0 60905.0 140355.0 ;
      RECT  60200.0 141700.0 60905.0 140355.0 ;
      RECT  60200.0 141700.0 60905.0 143045.0 ;
      RECT  60200.0 144390.0 60905.0 143045.0 ;
      RECT  60200.0 144390.0 60905.0 145735.0 ;
      RECT  60200.0 147080.0 60905.0 145735.0 ;
      RECT  60200.0 147080.0 60905.0 148425.0 ;
      RECT  60200.0 149770.0 60905.0 148425.0 ;
      RECT  60200.0 149770.0 60905.0 151115.0 ;
      RECT  60200.0 152460.0 60905.0 151115.0 ;
      RECT  60200.0 152460.0 60905.0 153805.0 ;
      RECT  60200.0 155150.0 60905.0 153805.0 ;
      RECT  60200.0 155150.0 60905.0 156495.0 ;
      RECT  60200.0 157840.0 60905.0 156495.0 ;
      RECT  60200.0 157840.0 60905.0 159185.0 ;
      RECT  60200.0 160530.0 60905.0 159185.0 ;
      RECT  60200.0 160530.0 60905.0 161875.0 ;
      RECT  60200.0 163220.0 60905.0 161875.0 ;
      RECT  60200.0 163220.0 60905.0 164565.0 ;
      RECT  60200.0 165910.0 60905.0 164565.0 ;
      RECT  60200.0 165910.0 60905.0 167255.0 ;
      RECT  60200.0 168600.0 60905.0 167255.0 ;
      RECT  60200.0 168600.0 60905.0 169945.0 ;
      RECT  60200.0 171290.0 60905.0 169945.0 ;
      RECT  60200.0 171290.0 60905.0 172635.0 ;
      RECT  60200.0 173980.0 60905.0 172635.0 ;
      RECT  60200.0 173980.0 60905.0 175325.0 ;
      RECT  60200.0 176670.0 60905.0 175325.0 ;
      RECT  60200.0 176670.0 60905.0 178015.0 ;
      RECT  60200.0 179360.0 60905.0 178015.0 ;
      RECT  60200.0 179360.0 60905.0 180705.0 ;
      RECT  60200.0 182050.0 60905.0 180705.0 ;
      RECT  60200.0 182050.0 60905.0 183395.0 ;
      RECT  60200.0 184740.0 60905.0 183395.0 ;
      RECT  60200.0 184740.0 60905.0 186085.0 ;
      RECT  60200.0 187430.0 60905.0 186085.0 ;
      RECT  60200.0 187430.0 60905.0 188775.0 ;
      RECT  60200.0 190120.0 60905.0 188775.0 ;
      RECT  60200.0 190120.0 60905.0 191465.0 ;
      RECT  60200.0 192810.0 60905.0 191465.0 ;
      RECT  60200.0 192810.0 60905.0 194155.0 ;
      RECT  60200.0 195500.0 60905.0 194155.0 ;
      RECT  60200.0 195500.0 60905.0 196845.0 ;
      RECT  60200.0 198190.0 60905.0 196845.0 ;
      RECT  60200.0 198190.0 60905.0 199535.0 ;
      RECT  60200.0 200880.0 60905.0 199535.0 ;
      RECT  60200.0 200880.0 60905.0 202225.0 ;
      RECT  60200.0 203570.0 60905.0 202225.0 ;
      RECT  60200.0 203570.0 60905.0 204915.0 ;
      RECT  60200.0 206260.0 60905.0 204915.0 ;
      RECT  60905.0 34100.0 61610.0 35445.0 ;
      RECT  60905.0 36790.0 61610.0 35445.0 ;
      RECT  60905.0 36790.0 61610.0 38135.0 ;
      RECT  60905.0 39480.0 61610.0 38135.0 ;
      RECT  60905.0 39480.0 61610.0 40825.0 ;
      RECT  60905.0 42170.0 61610.0 40825.0 ;
      RECT  60905.0 42170.0 61610.0 43515.0 ;
      RECT  60905.0 44860.0 61610.0 43515.0 ;
      RECT  60905.0 44860.0 61610.0 46205.0 ;
      RECT  60905.0 47550.0 61610.0 46205.0 ;
      RECT  60905.0 47550.0 61610.0 48895.0 ;
      RECT  60905.0 50240.0 61610.0 48895.0 ;
      RECT  60905.0 50240.0 61610.0 51585.0 ;
      RECT  60905.0 52930.0 61610.0 51585.0 ;
      RECT  60905.0 52930.0 61610.0 54275.0 ;
      RECT  60905.0 55620.0 61610.0 54275.0 ;
      RECT  60905.0 55620.0 61610.0 56965.0 ;
      RECT  60905.0 58310.0 61610.0 56965.0 ;
      RECT  60905.0 58310.0 61610.0 59655.0 ;
      RECT  60905.0 61000.0 61610.0 59655.0 ;
      RECT  60905.0 61000.0 61610.0 62345.0 ;
      RECT  60905.0 63690.0 61610.0 62345.0 ;
      RECT  60905.0 63690.0 61610.0 65035.0 ;
      RECT  60905.0 66380.0 61610.0 65035.0 ;
      RECT  60905.0 66380.0 61610.0 67725.0 ;
      RECT  60905.0 69070.0 61610.0 67725.0 ;
      RECT  60905.0 69070.0 61610.0 70415.0 ;
      RECT  60905.0 71760.0 61610.0 70415.0 ;
      RECT  60905.0 71760.0 61610.0 73105.0 ;
      RECT  60905.0 74450.0 61610.0 73105.0 ;
      RECT  60905.0 74450.0 61610.0 75795.0 ;
      RECT  60905.0 77140.0 61610.0 75795.0 ;
      RECT  60905.0 77140.0 61610.0 78485.0 ;
      RECT  60905.0 79830.0 61610.0 78485.0 ;
      RECT  60905.0 79830.0 61610.0 81175.0 ;
      RECT  60905.0 82520.0 61610.0 81175.0 ;
      RECT  60905.0 82520.0 61610.0 83865.0 ;
      RECT  60905.0 85210.0 61610.0 83865.0 ;
      RECT  60905.0 85210.0 61610.0 86555.0 ;
      RECT  60905.0 87900.0 61610.0 86555.0 ;
      RECT  60905.0 87900.0 61610.0 89245.0 ;
      RECT  60905.0 90590.0 61610.0 89245.0 ;
      RECT  60905.0 90590.0 61610.0 91935.0 ;
      RECT  60905.0 93280.0 61610.0 91935.0 ;
      RECT  60905.0 93280.0 61610.0 94625.0 ;
      RECT  60905.0 95970.0 61610.0 94625.0 ;
      RECT  60905.0 95970.0 61610.0 97315.0 ;
      RECT  60905.0 98660.0 61610.0 97315.0 ;
      RECT  60905.0 98660.0 61610.0 100005.0 ;
      RECT  60905.0 101350.0 61610.0 100005.0 ;
      RECT  60905.0 101350.0 61610.0 102695.0 ;
      RECT  60905.0 104040.0 61610.0 102695.0 ;
      RECT  60905.0 104040.0 61610.0 105385.0 ;
      RECT  60905.0 106730.0 61610.0 105385.0 ;
      RECT  60905.0 106730.0 61610.0 108075.0 ;
      RECT  60905.0 109420.0 61610.0 108075.0 ;
      RECT  60905.0 109420.0 61610.0 110765.0 ;
      RECT  60905.0 112110.0 61610.0 110765.0 ;
      RECT  60905.0 112110.0 61610.0 113455.0 ;
      RECT  60905.0 114800.0 61610.0 113455.0 ;
      RECT  60905.0 114800.0 61610.0 116145.0 ;
      RECT  60905.0 117490.0 61610.0 116145.0 ;
      RECT  60905.0 117490.0 61610.0 118835.0 ;
      RECT  60905.0 120180.0 61610.0 118835.0 ;
      RECT  60905.0 120180.0 61610.0 121525.0 ;
      RECT  60905.0 122870.0 61610.0 121525.0 ;
      RECT  60905.0 122870.0 61610.0 124215.0 ;
      RECT  60905.0 125560.0 61610.0 124215.0 ;
      RECT  60905.0 125560.0 61610.0 126905.0 ;
      RECT  60905.0 128250.0 61610.0 126905.0 ;
      RECT  60905.0 128250.0 61610.0 129595.0 ;
      RECT  60905.0 130940.0 61610.0 129595.0 ;
      RECT  60905.0 130940.0 61610.0 132285.0 ;
      RECT  60905.0 133630.0 61610.0 132285.0 ;
      RECT  60905.0 133630.0 61610.0 134975.0 ;
      RECT  60905.0 136320.0 61610.0 134975.0 ;
      RECT  60905.0 136320.0 61610.0 137665.0 ;
      RECT  60905.0 139010.0 61610.0 137665.0 ;
      RECT  60905.0 139010.0 61610.0 140355.0 ;
      RECT  60905.0 141700.0 61610.0 140355.0 ;
      RECT  60905.0 141700.0 61610.0 143045.0 ;
      RECT  60905.0 144390.0 61610.0 143045.0 ;
      RECT  60905.0 144390.0 61610.0 145735.0 ;
      RECT  60905.0 147080.0 61610.0 145735.0 ;
      RECT  60905.0 147080.0 61610.0 148425.0 ;
      RECT  60905.0 149770.0 61610.0 148425.0 ;
      RECT  60905.0 149770.0 61610.0 151115.0 ;
      RECT  60905.0 152460.0 61610.0 151115.0 ;
      RECT  60905.0 152460.0 61610.0 153805.0 ;
      RECT  60905.0 155150.0 61610.0 153805.0 ;
      RECT  60905.0 155150.0 61610.0 156495.0 ;
      RECT  60905.0 157840.0 61610.0 156495.0 ;
      RECT  60905.0 157840.0 61610.0 159185.0 ;
      RECT  60905.0 160530.0 61610.0 159185.0 ;
      RECT  60905.0 160530.0 61610.0 161875.0 ;
      RECT  60905.0 163220.0 61610.0 161875.0 ;
      RECT  60905.0 163220.0 61610.0 164565.0 ;
      RECT  60905.0 165910.0 61610.0 164565.0 ;
      RECT  60905.0 165910.0 61610.0 167255.0 ;
      RECT  60905.0 168600.0 61610.0 167255.0 ;
      RECT  60905.0 168600.0 61610.0 169945.0 ;
      RECT  60905.0 171290.0 61610.0 169945.0 ;
      RECT  60905.0 171290.0 61610.0 172635.0 ;
      RECT  60905.0 173980.0 61610.0 172635.0 ;
      RECT  60905.0 173980.0 61610.0 175325.0 ;
      RECT  60905.0 176670.0 61610.0 175325.0 ;
      RECT  60905.0 176670.0 61610.0 178015.0 ;
      RECT  60905.0 179360.0 61610.0 178015.0 ;
      RECT  60905.0 179360.0 61610.0 180705.0 ;
      RECT  60905.0 182050.0 61610.0 180705.0 ;
      RECT  60905.0 182050.0 61610.0 183395.0 ;
      RECT  60905.0 184740.0 61610.0 183395.0 ;
      RECT  60905.0 184740.0 61610.0 186085.0 ;
      RECT  60905.0 187430.0 61610.0 186085.0 ;
      RECT  60905.0 187430.0 61610.0 188775.0 ;
      RECT  60905.0 190120.0 61610.0 188775.0 ;
      RECT  60905.0 190120.0 61610.0 191465.0 ;
      RECT  60905.0 192810.0 61610.0 191465.0 ;
      RECT  60905.0 192810.0 61610.0 194155.0 ;
      RECT  60905.0 195500.0 61610.0 194155.0 ;
      RECT  60905.0 195500.0 61610.0 196845.0 ;
      RECT  60905.0 198190.0 61610.0 196845.0 ;
      RECT  60905.0 198190.0 61610.0 199535.0 ;
      RECT  60905.0 200880.0 61610.0 199535.0 ;
      RECT  60905.0 200880.0 61610.0 202225.0 ;
      RECT  60905.0 203570.0 61610.0 202225.0 ;
      RECT  60905.0 203570.0 61610.0 204915.0 ;
      RECT  60905.0 206260.0 61610.0 204915.0 ;
      RECT  61610.0 34100.0 62315.0 35445.0 ;
      RECT  61610.0 36790.0 62315.0 35445.0 ;
      RECT  61610.0 36790.0 62315.0 38135.0 ;
      RECT  61610.0 39480.0 62315.0 38135.0 ;
      RECT  61610.0 39480.0 62315.0 40825.0 ;
      RECT  61610.0 42170.0 62315.0 40825.0 ;
      RECT  61610.0 42170.0 62315.0 43515.0 ;
      RECT  61610.0 44860.0 62315.0 43515.0 ;
      RECT  61610.0 44860.0 62315.0 46205.0 ;
      RECT  61610.0 47550.0 62315.0 46205.0 ;
      RECT  61610.0 47550.0 62315.0 48895.0 ;
      RECT  61610.0 50240.0 62315.0 48895.0 ;
      RECT  61610.0 50240.0 62315.0 51585.0 ;
      RECT  61610.0 52930.0 62315.0 51585.0 ;
      RECT  61610.0 52930.0 62315.0 54275.0 ;
      RECT  61610.0 55620.0 62315.0 54275.0 ;
      RECT  61610.0 55620.0 62315.0 56965.0 ;
      RECT  61610.0 58310.0 62315.0 56965.0 ;
      RECT  61610.0 58310.0 62315.0 59655.0 ;
      RECT  61610.0 61000.0 62315.0 59655.0 ;
      RECT  61610.0 61000.0 62315.0 62345.0 ;
      RECT  61610.0 63690.0 62315.0 62345.0 ;
      RECT  61610.0 63690.0 62315.0 65035.0 ;
      RECT  61610.0 66380.0 62315.0 65035.0 ;
      RECT  61610.0 66380.0 62315.0 67725.0 ;
      RECT  61610.0 69070.0 62315.0 67725.0 ;
      RECT  61610.0 69070.0 62315.0 70415.0 ;
      RECT  61610.0 71760.0 62315.0 70415.0 ;
      RECT  61610.0 71760.0 62315.0 73105.0 ;
      RECT  61610.0 74450.0 62315.0 73105.0 ;
      RECT  61610.0 74450.0 62315.0 75795.0 ;
      RECT  61610.0 77140.0 62315.0 75795.0 ;
      RECT  61610.0 77140.0 62315.0 78485.0 ;
      RECT  61610.0 79830.0 62315.0 78485.0 ;
      RECT  61610.0 79830.0 62315.0 81175.0 ;
      RECT  61610.0 82520.0 62315.0 81175.0 ;
      RECT  61610.0 82520.0 62315.0 83865.0 ;
      RECT  61610.0 85210.0 62315.0 83865.0 ;
      RECT  61610.0 85210.0 62315.0 86555.0 ;
      RECT  61610.0 87900.0 62315.0 86555.0 ;
      RECT  61610.0 87900.0 62315.0 89245.0 ;
      RECT  61610.0 90590.0 62315.0 89245.0 ;
      RECT  61610.0 90590.0 62315.0 91935.0 ;
      RECT  61610.0 93280.0 62315.0 91935.0 ;
      RECT  61610.0 93280.0 62315.0 94625.0 ;
      RECT  61610.0 95970.0 62315.0 94625.0 ;
      RECT  61610.0 95970.0 62315.0 97315.0 ;
      RECT  61610.0 98660.0 62315.0 97315.0 ;
      RECT  61610.0 98660.0 62315.0 100005.0 ;
      RECT  61610.0 101350.0 62315.0 100005.0 ;
      RECT  61610.0 101350.0 62315.0 102695.0 ;
      RECT  61610.0 104040.0 62315.0 102695.0 ;
      RECT  61610.0 104040.0 62315.0 105385.0 ;
      RECT  61610.0 106730.0 62315.0 105385.0 ;
      RECT  61610.0 106730.0 62315.0 108075.0 ;
      RECT  61610.0 109420.0 62315.0 108075.0 ;
      RECT  61610.0 109420.0 62315.0 110765.0 ;
      RECT  61610.0 112110.0 62315.0 110765.0 ;
      RECT  61610.0 112110.0 62315.0 113455.0 ;
      RECT  61610.0 114800.0 62315.0 113455.0 ;
      RECT  61610.0 114800.0 62315.0 116145.0 ;
      RECT  61610.0 117490.0 62315.0 116145.0 ;
      RECT  61610.0 117490.0 62315.0 118835.0 ;
      RECT  61610.0 120180.0 62315.0 118835.0 ;
      RECT  61610.0 120180.0 62315.0 121525.0 ;
      RECT  61610.0 122870.0 62315.0 121525.0 ;
      RECT  61610.0 122870.0 62315.0 124215.0 ;
      RECT  61610.0 125560.0 62315.0 124215.0 ;
      RECT  61610.0 125560.0 62315.0 126905.0 ;
      RECT  61610.0 128250.0 62315.0 126905.0 ;
      RECT  61610.0 128250.0 62315.0 129595.0 ;
      RECT  61610.0 130940.0 62315.0 129595.0 ;
      RECT  61610.0 130940.0 62315.0 132285.0 ;
      RECT  61610.0 133630.0 62315.0 132285.0 ;
      RECT  61610.0 133630.0 62315.0 134975.0 ;
      RECT  61610.0 136320.0 62315.0 134975.0 ;
      RECT  61610.0 136320.0 62315.0 137665.0 ;
      RECT  61610.0 139010.0 62315.0 137665.0 ;
      RECT  61610.0 139010.0 62315.0 140355.0 ;
      RECT  61610.0 141700.0 62315.0 140355.0 ;
      RECT  61610.0 141700.0 62315.0 143045.0 ;
      RECT  61610.0 144390.0 62315.0 143045.0 ;
      RECT  61610.0 144390.0 62315.0 145735.0 ;
      RECT  61610.0 147080.0 62315.0 145735.0 ;
      RECT  61610.0 147080.0 62315.0 148425.0 ;
      RECT  61610.0 149770.0 62315.0 148425.0 ;
      RECT  61610.0 149770.0 62315.0 151115.0 ;
      RECT  61610.0 152460.0 62315.0 151115.0 ;
      RECT  61610.0 152460.0 62315.0 153805.0 ;
      RECT  61610.0 155150.0 62315.0 153805.0 ;
      RECT  61610.0 155150.0 62315.0 156495.0 ;
      RECT  61610.0 157840.0 62315.0 156495.0 ;
      RECT  61610.0 157840.0 62315.0 159185.0 ;
      RECT  61610.0 160530.0 62315.0 159185.0 ;
      RECT  61610.0 160530.0 62315.0 161875.0 ;
      RECT  61610.0 163220.0 62315.0 161875.0 ;
      RECT  61610.0 163220.0 62315.0 164565.0 ;
      RECT  61610.0 165910.0 62315.0 164565.0 ;
      RECT  61610.0 165910.0 62315.0 167255.0 ;
      RECT  61610.0 168600.0 62315.0 167255.0 ;
      RECT  61610.0 168600.0 62315.0 169945.0 ;
      RECT  61610.0 171290.0 62315.0 169945.0 ;
      RECT  61610.0 171290.0 62315.0 172635.0 ;
      RECT  61610.0 173980.0 62315.0 172635.0 ;
      RECT  61610.0 173980.0 62315.0 175325.0 ;
      RECT  61610.0 176670.0 62315.0 175325.0 ;
      RECT  61610.0 176670.0 62315.0 178015.0 ;
      RECT  61610.0 179360.0 62315.0 178015.0 ;
      RECT  61610.0 179360.0 62315.0 180705.0 ;
      RECT  61610.0 182050.0 62315.0 180705.0 ;
      RECT  61610.0 182050.0 62315.0 183395.0 ;
      RECT  61610.0 184740.0 62315.0 183395.0 ;
      RECT  61610.0 184740.0 62315.0 186085.0 ;
      RECT  61610.0 187430.0 62315.0 186085.0 ;
      RECT  61610.0 187430.0 62315.0 188775.0 ;
      RECT  61610.0 190120.0 62315.0 188775.0 ;
      RECT  61610.0 190120.0 62315.0 191465.0 ;
      RECT  61610.0 192810.0 62315.0 191465.0 ;
      RECT  61610.0 192810.0 62315.0 194155.0 ;
      RECT  61610.0 195500.0 62315.0 194155.0 ;
      RECT  61610.0 195500.0 62315.0 196845.0 ;
      RECT  61610.0 198190.0 62315.0 196845.0 ;
      RECT  61610.0 198190.0 62315.0 199535.0 ;
      RECT  61610.0 200880.0 62315.0 199535.0 ;
      RECT  61610.0 200880.0 62315.0 202225.0 ;
      RECT  61610.0 203570.0 62315.0 202225.0 ;
      RECT  61610.0 203570.0 62315.0 204915.0 ;
      RECT  61610.0 206260.0 62315.0 204915.0 ;
      RECT  62315.0 34100.0 63020.0 35445.0 ;
      RECT  62315.0 36790.0 63020.0 35445.0 ;
      RECT  62315.0 36790.0 63020.0 38135.0 ;
      RECT  62315.0 39480.0 63020.0 38135.0 ;
      RECT  62315.0 39480.0 63020.0 40825.0 ;
      RECT  62315.0 42170.0 63020.0 40825.0 ;
      RECT  62315.0 42170.0 63020.0 43515.0 ;
      RECT  62315.0 44860.0 63020.0 43515.0 ;
      RECT  62315.0 44860.0 63020.0 46205.0 ;
      RECT  62315.0 47550.0 63020.0 46205.0 ;
      RECT  62315.0 47550.0 63020.0 48895.0 ;
      RECT  62315.0 50240.0 63020.0 48895.0 ;
      RECT  62315.0 50240.0 63020.0 51585.0 ;
      RECT  62315.0 52930.0 63020.0 51585.0 ;
      RECT  62315.0 52930.0 63020.0 54275.0 ;
      RECT  62315.0 55620.0 63020.0 54275.0 ;
      RECT  62315.0 55620.0 63020.0 56965.0 ;
      RECT  62315.0 58310.0 63020.0 56965.0 ;
      RECT  62315.0 58310.0 63020.0 59655.0 ;
      RECT  62315.0 61000.0 63020.0 59655.0 ;
      RECT  62315.0 61000.0 63020.0 62345.0 ;
      RECT  62315.0 63690.0 63020.0 62345.0 ;
      RECT  62315.0 63690.0 63020.0 65035.0 ;
      RECT  62315.0 66380.0 63020.0 65035.0 ;
      RECT  62315.0 66380.0 63020.0 67725.0 ;
      RECT  62315.0 69070.0 63020.0 67725.0 ;
      RECT  62315.0 69070.0 63020.0 70415.0 ;
      RECT  62315.0 71760.0 63020.0 70415.0 ;
      RECT  62315.0 71760.0 63020.0 73105.0 ;
      RECT  62315.0 74450.0 63020.0 73105.0 ;
      RECT  62315.0 74450.0 63020.0 75795.0 ;
      RECT  62315.0 77140.0 63020.0 75795.0 ;
      RECT  62315.0 77140.0 63020.0 78485.0 ;
      RECT  62315.0 79830.0 63020.0 78485.0 ;
      RECT  62315.0 79830.0 63020.0 81175.0 ;
      RECT  62315.0 82520.0 63020.0 81175.0 ;
      RECT  62315.0 82520.0 63020.0 83865.0 ;
      RECT  62315.0 85210.0 63020.0 83865.0 ;
      RECT  62315.0 85210.0 63020.0 86555.0 ;
      RECT  62315.0 87900.0 63020.0 86555.0 ;
      RECT  62315.0 87900.0 63020.0 89245.0 ;
      RECT  62315.0 90590.0 63020.0 89245.0 ;
      RECT  62315.0 90590.0 63020.0 91935.0 ;
      RECT  62315.0 93280.0 63020.0 91935.0 ;
      RECT  62315.0 93280.0 63020.0 94625.0 ;
      RECT  62315.0 95970.0 63020.0 94625.0 ;
      RECT  62315.0 95970.0 63020.0 97315.0 ;
      RECT  62315.0 98660.0 63020.0 97315.0 ;
      RECT  62315.0 98660.0 63020.0 100005.0 ;
      RECT  62315.0 101350.0 63020.0 100005.0 ;
      RECT  62315.0 101350.0 63020.0 102695.0 ;
      RECT  62315.0 104040.0 63020.0 102695.0 ;
      RECT  62315.0 104040.0 63020.0 105385.0 ;
      RECT  62315.0 106730.0 63020.0 105385.0 ;
      RECT  62315.0 106730.0 63020.0 108075.0 ;
      RECT  62315.0 109420.0 63020.0 108075.0 ;
      RECT  62315.0 109420.0 63020.0 110765.0 ;
      RECT  62315.0 112110.0 63020.0 110765.0 ;
      RECT  62315.0 112110.0 63020.0 113455.0 ;
      RECT  62315.0 114800.0 63020.0 113455.0 ;
      RECT  62315.0 114800.0 63020.0 116145.0 ;
      RECT  62315.0 117490.0 63020.0 116145.0 ;
      RECT  62315.0 117490.0 63020.0 118835.0 ;
      RECT  62315.0 120180.0 63020.0 118835.0 ;
      RECT  62315.0 120180.0 63020.0 121525.0 ;
      RECT  62315.0 122870.0 63020.0 121525.0 ;
      RECT  62315.0 122870.0 63020.0 124215.0 ;
      RECT  62315.0 125560.0 63020.0 124215.0 ;
      RECT  62315.0 125560.0 63020.0 126905.0 ;
      RECT  62315.0 128250.0 63020.0 126905.0 ;
      RECT  62315.0 128250.0 63020.0 129595.0 ;
      RECT  62315.0 130940.0 63020.0 129595.0 ;
      RECT  62315.0 130940.0 63020.0 132285.0 ;
      RECT  62315.0 133630.0 63020.0 132285.0 ;
      RECT  62315.0 133630.0 63020.0 134975.0 ;
      RECT  62315.0 136320.0 63020.0 134975.0 ;
      RECT  62315.0 136320.0 63020.0 137665.0 ;
      RECT  62315.0 139010.0 63020.0 137665.0 ;
      RECT  62315.0 139010.0 63020.0 140355.0 ;
      RECT  62315.0 141700.0 63020.0 140355.0 ;
      RECT  62315.0 141700.0 63020.0 143045.0 ;
      RECT  62315.0 144390.0 63020.0 143045.0 ;
      RECT  62315.0 144390.0 63020.0 145735.0 ;
      RECT  62315.0 147080.0 63020.0 145735.0 ;
      RECT  62315.0 147080.0 63020.0 148425.0 ;
      RECT  62315.0 149770.0 63020.0 148425.0 ;
      RECT  62315.0 149770.0 63020.0 151115.0 ;
      RECT  62315.0 152460.0 63020.0 151115.0 ;
      RECT  62315.0 152460.0 63020.0 153805.0 ;
      RECT  62315.0 155150.0 63020.0 153805.0 ;
      RECT  62315.0 155150.0 63020.0 156495.0 ;
      RECT  62315.0 157840.0 63020.0 156495.0 ;
      RECT  62315.0 157840.0 63020.0 159185.0 ;
      RECT  62315.0 160530.0 63020.0 159185.0 ;
      RECT  62315.0 160530.0 63020.0 161875.0 ;
      RECT  62315.0 163220.0 63020.0 161875.0 ;
      RECT  62315.0 163220.0 63020.0 164565.0 ;
      RECT  62315.0 165910.0 63020.0 164565.0 ;
      RECT  62315.0 165910.0 63020.0 167255.0 ;
      RECT  62315.0 168600.0 63020.0 167255.0 ;
      RECT  62315.0 168600.0 63020.0 169945.0 ;
      RECT  62315.0 171290.0 63020.0 169945.0 ;
      RECT  62315.0 171290.0 63020.0 172635.0 ;
      RECT  62315.0 173980.0 63020.0 172635.0 ;
      RECT  62315.0 173980.0 63020.0 175325.0 ;
      RECT  62315.0 176670.0 63020.0 175325.0 ;
      RECT  62315.0 176670.0 63020.0 178015.0 ;
      RECT  62315.0 179360.0 63020.0 178015.0 ;
      RECT  62315.0 179360.0 63020.0 180705.0 ;
      RECT  62315.0 182050.0 63020.0 180705.0 ;
      RECT  62315.0 182050.0 63020.0 183395.0 ;
      RECT  62315.0 184740.0 63020.0 183395.0 ;
      RECT  62315.0 184740.0 63020.0 186085.0 ;
      RECT  62315.0 187430.0 63020.0 186085.0 ;
      RECT  62315.0 187430.0 63020.0 188775.0 ;
      RECT  62315.0 190120.0 63020.0 188775.0 ;
      RECT  62315.0 190120.0 63020.0 191465.0 ;
      RECT  62315.0 192810.0 63020.0 191465.0 ;
      RECT  62315.0 192810.0 63020.0 194155.0 ;
      RECT  62315.0 195500.0 63020.0 194155.0 ;
      RECT  62315.0 195500.0 63020.0 196845.0 ;
      RECT  62315.0 198190.0 63020.0 196845.0 ;
      RECT  62315.0 198190.0 63020.0 199535.0 ;
      RECT  62315.0 200880.0 63020.0 199535.0 ;
      RECT  62315.0 200880.0 63020.0 202225.0 ;
      RECT  62315.0 203570.0 63020.0 202225.0 ;
      RECT  62315.0 203570.0 63020.0 204915.0 ;
      RECT  62315.0 206260.0 63020.0 204915.0 ;
      RECT  63020.0 34100.0 63725.0 35445.0 ;
      RECT  63020.0 36790.0 63725.0 35445.0 ;
      RECT  63020.0 36790.0 63725.0 38135.0 ;
      RECT  63020.0 39480.0 63725.0 38135.0 ;
      RECT  63020.0 39480.0 63725.0 40825.0 ;
      RECT  63020.0 42170.0 63725.0 40825.0 ;
      RECT  63020.0 42170.0 63725.0 43515.0 ;
      RECT  63020.0 44860.0 63725.0 43515.0 ;
      RECT  63020.0 44860.0 63725.0 46205.0 ;
      RECT  63020.0 47550.0 63725.0 46205.0 ;
      RECT  63020.0 47550.0 63725.0 48895.0 ;
      RECT  63020.0 50240.0 63725.0 48895.0 ;
      RECT  63020.0 50240.0 63725.0 51585.0 ;
      RECT  63020.0 52930.0 63725.0 51585.0 ;
      RECT  63020.0 52930.0 63725.0 54275.0 ;
      RECT  63020.0 55620.0 63725.0 54275.0 ;
      RECT  63020.0 55620.0 63725.0 56965.0 ;
      RECT  63020.0 58310.0 63725.0 56965.0 ;
      RECT  63020.0 58310.0 63725.0 59655.0 ;
      RECT  63020.0 61000.0 63725.0 59655.0 ;
      RECT  63020.0 61000.0 63725.0 62345.0 ;
      RECT  63020.0 63690.0 63725.0 62345.0 ;
      RECT  63020.0 63690.0 63725.0 65035.0 ;
      RECT  63020.0 66380.0 63725.0 65035.0 ;
      RECT  63020.0 66380.0 63725.0 67725.0 ;
      RECT  63020.0 69070.0 63725.0 67725.0 ;
      RECT  63020.0 69070.0 63725.0 70415.0 ;
      RECT  63020.0 71760.0 63725.0 70415.0 ;
      RECT  63020.0 71760.0 63725.0 73105.0 ;
      RECT  63020.0 74450.0 63725.0 73105.0 ;
      RECT  63020.0 74450.0 63725.0 75795.0 ;
      RECT  63020.0 77140.0 63725.0 75795.0 ;
      RECT  63020.0 77140.0 63725.0 78485.0 ;
      RECT  63020.0 79830.0 63725.0 78485.0 ;
      RECT  63020.0 79830.0 63725.0 81175.0 ;
      RECT  63020.0 82520.0 63725.0 81175.0 ;
      RECT  63020.0 82520.0 63725.0 83865.0 ;
      RECT  63020.0 85210.0 63725.0 83865.0 ;
      RECT  63020.0 85210.0 63725.0 86555.0 ;
      RECT  63020.0 87900.0 63725.0 86555.0 ;
      RECT  63020.0 87900.0 63725.0 89245.0 ;
      RECT  63020.0 90590.0 63725.0 89245.0 ;
      RECT  63020.0 90590.0 63725.0 91935.0 ;
      RECT  63020.0 93280.0 63725.0 91935.0 ;
      RECT  63020.0 93280.0 63725.0 94625.0 ;
      RECT  63020.0 95970.0 63725.0 94625.0 ;
      RECT  63020.0 95970.0 63725.0 97315.0 ;
      RECT  63020.0 98660.0 63725.0 97315.0 ;
      RECT  63020.0 98660.0 63725.0 100005.0 ;
      RECT  63020.0 101350.0 63725.0 100005.0 ;
      RECT  63020.0 101350.0 63725.0 102695.0 ;
      RECT  63020.0 104040.0 63725.0 102695.0 ;
      RECT  63020.0 104040.0 63725.0 105385.0 ;
      RECT  63020.0 106730.0 63725.0 105385.0 ;
      RECT  63020.0 106730.0 63725.0 108075.0 ;
      RECT  63020.0 109420.0 63725.0 108075.0 ;
      RECT  63020.0 109420.0 63725.0 110765.0 ;
      RECT  63020.0 112110.0 63725.0 110765.0 ;
      RECT  63020.0 112110.0 63725.0 113455.0 ;
      RECT  63020.0 114800.0 63725.0 113455.0 ;
      RECT  63020.0 114800.0 63725.0 116145.0 ;
      RECT  63020.0 117490.0 63725.0 116145.0 ;
      RECT  63020.0 117490.0 63725.0 118835.0 ;
      RECT  63020.0 120180.0 63725.0 118835.0 ;
      RECT  63020.0 120180.0 63725.0 121525.0 ;
      RECT  63020.0 122870.0 63725.0 121525.0 ;
      RECT  63020.0 122870.0 63725.0 124215.0 ;
      RECT  63020.0 125560.0 63725.0 124215.0 ;
      RECT  63020.0 125560.0 63725.0 126905.0 ;
      RECT  63020.0 128250.0 63725.0 126905.0 ;
      RECT  63020.0 128250.0 63725.0 129595.0 ;
      RECT  63020.0 130940.0 63725.0 129595.0 ;
      RECT  63020.0 130940.0 63725.0 132285.0 ;
      RECT  63020.0 133630.0 63725.0 132285.0 ;
      RECT  63020.0 133630.0 63725.0 134975.0 ;
      RECT  63020.0 136320.0 63725.0 134975.0 ;
      RECT  63020.0 136320.0 63725.0 137665.0 ;
      RECT  63020.0 139010.0 63725.0 137665.0 ;
      RECT  63020.0 139010.0 63725.0 140355.0 ;
      RECT  63020.0 141700.0 63725.0 140355.0 ;
      RECT  63020.0 141700.0 63725.0 143045.0 ;
      RECT  63020.0 144390.0 63725.0 143045.0 ;
      RECT  63020.0 144390.0 63725.0 145735.0 ;
      RECT  63020.0 147080.0 63725.0 145735.0 ;
      RECT  63020.0 147080.0 63725.0 148425.0 ;
      RECT  63020.0 149770.0 63725.0 148425.0 ;
      RECT  63020.0 149770.0 63725.0 151115.0 ;
      RECT  63020.0 152460.0 63725.0 151115.0 ;
      RECT  63020.0 152460.0 63725.0 153805.0 ;
      RECT  63020.0 155150.0 63725.0 153805.0 ;
      RECT  63020.0 155150.0 63725.0 156495.0 ;
      RECT  63020.0 157840.0 63725.0 156495.0 ;
      RECT  63020.0 157840.0 63725.0 159185.0 ;
      RECT  63020.0 160530.0 63725.0 159185.0 ;
      RECT  63020.0 160530.0 63725.0 161875.0 ;
      RECT  63020.0 163220.0 63725.0 161875.0 ;
      RECT  63020.0 163220.0 63725.0 164565.0 ;
      RECT  63020.0 165910.0 63725.0 164565.0 ;
      RECT  63020.0 165910.0 63725.0 167255.0 ;
      RECT  63020.0 168600.0 63725.0 167255.0 ;
      RECT  63020.0 168600.0 63725.0 169945.0 ;
      RECT  63020.0 171290.0 63725.0 169945.0 ;
      RECT  63020.0 171290.0 63725.0 172635.0 ;
      RECT  63020.0 173980.0 63725.0 172635.0 ;
      RECT  63020.0 173980.0 63725.0 175325.0 ;
      RECT  63020.0 176670.0 63725.0 175325.0 ;
      RECT  63020.0 176670.0 63725.0 178015.0 ;
      RECT  63020.0 179360.0 63725.0 178015.0 ;
      RECT  63020.0 179360.0 63725.0 180705.0 ;
      RECT  63020.0 182050.0 63725.0 180705.0 ;
      RECT  63020.0 182050.0 63725.0 183395.0 ;
      RECT  63020.0 184740.0 63725.0 183395.0 ;
      RECT  63020.0 184740.0 63725.0 186085.0 ;
      RECT  63020.0 187430.0 63725.0 186085.0 ;
      RECT  63020.0 187430.0 63725.0 188775.0 ;
      RECT  63020.0 190120.0 63725.0 188775.0 ;
      RECT  63020.0 190120.0 63725.0 191465.0 ;
      RECT  63020.0 192810.0 63725.0 191465.0 ;
      RECT  63020.0 192810.0 63725.0 194155.0 ;
      RECT  63020.0 195500.0 63725.0 194155.0 ;
      RECT  63020.0 195500.0 63725.0 196845.0 ;
      RECT  63020.0 198190.0 63725.0 196845.0 ;
      RECT  63020.0 198190.0 63725.0 199535.0 ;
      RECT  63020.0 200880.0 63725.0 199535.0 ;
      RECT  63020.0 200880.0 63725.0 202225.0 ;
      RECT  63020.0 203570.0 63725.0 202225.0 ;
      RECT  63020.0 203570.0 63725.0 204915.0 ;
      RECT  63020.0 206260.0 63725.0 204915.0 ;
      RECT  63725.0 34100.0 64430.0 35445.0 ;
      RECT  63725.0 36790.0 64430.0 35445.0 ;
      RECT  63725.0 36790.0 64430.0 38135.0 ;
      RECT  63725.0 39480.0 64430.0 38135.0 ;
      RECT  63725.0 39480.0 64430.0 40825.0 ;
      RECT  63725.0 42170.0 64430.0 40825.0 ;
      RECT  63725.0 42170.0 64430.0 43515.0 ;
      RECT  63725.0 44860.0 64430.0 43515.0 ;
      RECT  63725.0 44860.0 64430.0 46205.0 ;
      RECT  63725.0 47550.0 64430.0 46205.0 ;
      RECT  63725.0 47550.0 64430.0 48895.0 ;
      RECT  63725.0 50240.0 64430.0 48895.0 ;
      RECT  63725.0 50240.0 64430.0 51585.0 ;
      RECT  63725.0 52930.0 64430.0 51585.0 ;
      RECT  63725.0 52930.0 64430.0 54275.0 ;
      RECT  63725.0 55620.0 64430.0 54275.0 ;
      RECT  63725.0 55620.0 64430.0 56965.0 ;
      RECT  63725.0 58310.0 64430.0 56965.0 ;
      RECT  63725.0 58310.0 64430.0 59655.0 ;
      RECT  63725.0 61000.0 64430.0 59655.0 ;
      RECT  63725.0 61000.0 64430.0 62345.0 ;
      RECT  63725.0 63690.0 64430.0 62345.0 ;
      RECT  63725.0 63690.0 64430.0 65035.0 ;
      RECT  63725.0 66380.0 64430.0 65035.0 ;
      RECT  63725.0 66380.0 64430.0 67725.0 ;
      RECT  63725.0 69070.0 64430.0 67725.0 ;
      RECT  63725.0 69070.0 64430.0 70415.0 ;
      RECT  63725.0 71760.0 64430.0 70415.0 ;
      RECT  63725.0 71760.0 64430.0 73105.0 ;
      RECT  63725.0 74450.0 64430.0 73105.0 ;
      RECT  63725.0 74450.0 64430.0 75795.0 ;
      RECT  63725.0 77140.0 64430.0 75795.0 ;
      RECT  63725.0 77140.0 64430.0 78485.0 ;
      RECT  63725.0 79830.0 64430.0 78485.0 ;
      RECT  63725.0 79830.0 64430.0 81175.0 ;
      RECT  63725.0 82520.0 64430.0 81175.0 ;
      RECT  63725.0 82520.0 64430.0 83865.0 ;
      RECT  63725.0 85210.0 64430.0 83865.0 ;
      RECT  63725.0 85210.0 64430.0 86555.0 ;
      RECT  63725.0 87900.0 64430.0 86555.0 ;
      RECT  63725.0 87900.0 64430.0 89245.0 ;
      RECT  63725.0 90590.0 64430.0 89245.0 ;
      RECT  63725.0 90590.0 64430.0 91935.0 ;
      RECT  63725.0 93280.0 64430.0 91935.0 ;
      RECT  63725.0 93280.0 64430.0 94625.0 ;
      RECT  63725.0 95970.0 64430.0 94625.0 ;
      RECT  63725.0 95970.0 64430.0 97315.0 ;
      RECT  63725.0 98660.0 64430.0 97315.0 ;
      RECT  63725.0 98660.0 64430.0 100005.0 ;
      RECT  63725.0 101350.0 64430.0 100005.0 ;
      RECT  63725.0 101350.0 64430.0 102695.0 ;
      RECT  63725.0 104040.0 64430.0 102695.0 ;
      RECT  63725.0 104040.0 64430.0 105385.0 ;
      RECT  63725.0 106730.0 64430.0 105385.0 ;
      RECT  63725.0 106730.0 64430.0 108075.0 ;
      RECT  63725.0 109420.0 64430.0 108075.0 ;
      RECT  63725.0 109420.0 64430.0 110765.0 ;
      RECT  63725.0 112110.0 64430.0 110765.0 ;
      RECT  63725.0 112110.0 64430.0 113455.0 ;
      RECT  63725.0 114800.0 64430.0 113455.0 ;
      RECT  63725.0 114800.0 64430.0 116145.0 ;
      RECT  63725.0 117490.0 64430.0 116145.0 ;
      RECT  63725.0 117490.0 64430.0 118835.0 ;
      RECT  63725.0 120180.0 64430.0 118835.0 ;
      RECT  63725.0 120180.0 64430.0 121525.0 ;
      RECT  63725.0 122870.0 64430.0 121525.0 ;
      RECT  63725.0 122870.0 64430.0 124215.0 ;
      RECT  63725.0 125560.0 64430.0 124215.0 ;
      RECT  63725.0 125560.0 64430.0 126905.0 ;
      RECT  63725.0 128250.0 64430.0 126905.0 ;
      RECT  63725.0 128250.0 64430.0 129595.0 ;
      RECT  63725.0 130940.0 64430.0 129595.0 ;
      RECT  63725.0 130940.0 64430.0 132285.0 ;
      RECT  63725.0 133630.0 64430.0 132285.0 ;
      RECT  63725.0 133630.0 64430.0 134975.0 ;
      RECT  63725.0 136320.0 64430.0 134975.0 ;
      RECT  63725.0 136320.0 64430.0 137665.0 ;
      RECT  63725.0 139010.0 64430.0 137665.0 ;
      RECT  63725.0 139010.0 64430.0 140355.0 ;
      RECT  63725.0 141700.0 64430.0 140355.0 ;
      RECT  63725.0 141700.0 64430.0 143045.0 ;
      RECT  63725.0 144390.0 64430.0 143045.0 ;
      RECT  63725.0 144390.0 64430.0 145735.0 ;
      RECT  63725.0 147080.0 64430.0 145735.0 ;
      RECT  63725.0 147080.0 64430.0 148425.0 ;
      RECT  63725.0 149770.0 64430.0 148425.0 ;
      RECT  63725.0 149770.0 64430.0 151115.0 ;
      RECT  63725.0 152460.0 64430.0 151115.0 ;
      RECT  63725.0 152460.0 64430.0 153805.0 ;
      RECT  63725.0 155150.0 64430.0 153805.0 ;
      RECT  63725.0 155150.0 64430.0 156495.0 ;
      RECT  63725.0 157840.0 64430.0 156495.0 ;
      RECT  63725.0 157840.0 64430.0 159185.0 ;
      RECT  63725.0 160530.0 64430.0 159185.0 ;
      RECT  63725.0 160530.0 64430.0 161875.0 ;
      RECT  63725.0 163220.0 64430.0 161875.0 ;
      RECT  63725.0 163220.0 64430.0 164565.0 ;
      RECT  63725.0 165910.0 64430.0 164565.0 ;
      RECT  63725.0 165910.0 64430.0 167255.0 ;
      RECT  63725.0 168600.0 64430.0 167255.0 ;
      RECT  63725.0 168600.0 64430.0 169945.0 ;
      RECT  63725.0 171290.0 64430.0 169945.0 ;
      RECT  63725.0 171290.0 64430.0 172635.0 ;
      RECT  63725.0 173980.0 64430.0 172635.0 ;
      RECT  63725.0 173980.0 64430.0 175325.0 ;
      RECT  63725.0 176670.0 64430.0 175325.0 ;
      RECT  63725.0 176670.0 64430.0 178015.0 ;
      RECT  63725.0 179360.0 64430.0 178015.0 ;
      RECT  63725.0 179360.0 64430.0 180705.0 ;
      RECT  63725.0 182050.0 64430.0 180705.0 ;
      RECT  63725.0 182050.0 64430.0 183395.0 ;
      RECT  63725.0 184740.0 64430.0 183395.0 ;
      RECT  63725.0 184740.0 64430.0 186085.0 ;
      RECT  63725.0 187430.0 64430.0 186085.0 ;
      RECT  63725.0 187430.0 64430.0 188775.0 ;
      RECT  63725.0 190120.0 64430.0 188775.0 ;
      RECT  63725.0 190120.0 64430.0 191465.0 ;
      RECT  63725.0 192810.0 64430.0 191465.0 ;
      RECT  63725.0 192810.0 64430.0 194155.0 ;
      RECT  63725.0 195500.0 64430.0 194155.0 ;
      RECT  63725.0 195500.0 64430.0 196845.0 ;
      RECT  63725.0 198190.0 64430.0 196845.0 ;
      RECT  63725.0 198190.0 64430.0 199535.0 ;
      RECT  63725.0 200880.0 64430.0 199535.0 ;
      RECT  63725.0 200880.0 64430.0 202225.0 ;
      RECT  63725.0 203570.0 64430.0 202225.0 ;
      RECT  63725.0 203570.0 64430.0 204915.0 ;
      RECT  63725.0 206260.0 64430.0 204915.0 ;
      RECT  64430.0 34100.0 65135.0 35445.0 ;
      RECT  64430.0 36790.0 65135.0 35445.0 ;
      RECT  64430.0 36790.0 65135.0 38135.0 ;
      RECT  64430.0 39480.0 65135.0 38135.0 ;
      RECT  64430.0 39480.0 65135.0 40825.0 ;
      RECT  64430.0 42170.0 65135.0 40825.0 ;
      RECT  64430.0 42170.0 65135.0 43515.0 ;
      RECT  64430.0 44860.0 65135.0 43515.0 ;
      RECT  64430.0 44860.0 65135.0 46205.0 ;
      RECT  64430.0 47550.0 65135.0 46205.0 ;
      RECT  64430.0 47550.0 65135.0 48895.0 ;
      RECT  64430.0 50240.0 65135.0 48895.0 ;
      RECT  64430.0 50240.0 65135.0 51585.0 ;
      RECT  64430.0 52930.0 65135.0 51585.0 ;
      RECT  64430.0 52930.0 65135.0 54275.0 ;
      RECT  64430.0 55620.0 65135.0 54275.0 ;
      RECT  64430.0 55620.0 65135.0 56965.0 ;
      RECT  64430.0 58310.0 65135.0 56965.0 ;
      RECT  64430.0 58310.0 65135.0 59655.0 ;
      RECT  64430.0 61000.0 65135.0 59655.0 ;
      RECT  64430.0 61000.0 65135.0 62345.0 ;
      RECT  64430.0 63690.0 65135.0 62345.0 ;
      RECT  64430.0 63690.0 65135.0 65035.0 ;
      RECT  64430.0 66380.0 65135.0 65035.0 ;
      RECT  64430.0 66380.0 65135.0 67725.0 ;
      RECT  64430.0 69070.0 65135.0 67725.0 ;
      RECT  64430.0 69070.0 65135.0 70415.0 ;
      RECT  64430.0 71760.0 65135.0 70415.0 ;
      RECT  64430.0 71760.0 65135.0 73105.0 ;
      RECT  64430.0 74450.0 65135.0 73105.0 ;
      RECT  64430.0 74450.0 65135.0 75795.0 ;
      RECT  64430.0 77140.0 65135.0 75795.0 ;
      RECT  64430.0 77140.0 65135.0 78485.0 ;
      RECT  64430.0 79830.0 65135.0 78485.0 ;
      RECT  64430.0 79830.0 65135.0 81175.0 ;
      RECT  64430.0 82520.0 65135.0 81175.0 ;
      RECT  64430.0 82520.0 65135.0 83865.0 ;
      RECT  64430.0 85210.0 65135.0 83865.0 ;
      RECT  64430.0 85210.0 65135.0 86555.0 ;
      RECT  64430.0 87900.0 65135.0 86555.0 ;
      RECT  64430.0 87900.0 65135.0 89245.0 ;
      RECT  64430.0 90590.0 65135.0 89245.0 ;
      RECT  64430.0 90590.0 65135.0 91935.0 ;
      RECT  64430.0 93280.0 65135.0 91935.0 ;
      RECT  64430.0 93280.0 65135.0 94625.0 ;
      RECT  64430.0 95970.0 65135.0 94625.0 ;
      RECT  64430.0 95970.0 65135.0 97315.0 ;
      RECT  64430.0 98660.0 65135.0 97315.0 ;
      RECT  64430.0 98660.0 65135.0 100005.0 ;
      RECT  64430.0 101350.0 65135.0 100005.0 ;
      RECT  64430.0 101350.0 65135.0 102695.0 ;
      RECT  64430.0 104040.0 65135.0 102695.0 ;
      RECT  64430.0 104040.0 65135.0 105385.0 ;
      RECT  64430.0 106730.0 65135.0 105385.0 ;
      RECT  64430.0 106730.0 65135.0 108075.0 ;
      RECT  64430.0 109420.0 65135.0 108075.0 ;
      RECT  64430.0 109420.0 65135.0 110765.0 ;
      RECT  64430.0 112110.0 65135.0 110765.0 ;
      RECT  64430.0 112110.0 65135.0 113455.0 ;
      RECT  64430.0 114800.0 65135.0 113455.0 ;
      RECT  64430.0 114800.0 65135.0 116145.0 ;
      RECT  64430.0 117490.0 65135.0 116145.0 ;
      RECT  64430.0 117490.0 65135.0 118835.0 ;
      RECT  64430.0 120180.0 65135.0 118835.0 ;
      RECT  64430.0 120180.0 65135.0 121525.0 ;
      RECT  64430.0 122870.0 65135.0 121525.0 ;
      RECT  64430.0 122870.0 65135.0 124215.0 ;
      RECT  64430.0 125560.0 65135.0 124215.0 ;
      RECT  64430.0 125560.0 65135.0 126905.0 ;
      RECT  64430.0 128250.0 65135.0 126905.0 ;
      RECT  64430.0 128250.0 65135.0 129595.0 ;
      RECT  64430.0 130940.0 65135.0 129595.0 ;
      RECT  64430.0 130940.0 65135.0 132285.0 ;
      RECT  64430.0 133630.0 65135.0 132285.0 ;
      RECT  64430.0 133630.0 65135.0 134975.0 ;
      RECT  64430.0 136320.0 65135.0 134975.0 ;
      RECT  64430.0 136320.0 65135.0 137665.0 ;
      RECT  64430.0 139010.0 65135.0 137665.0 ;
      RECT  64430.0 139010.0 65135.0 140355.0 ;
      RECT  64430.0 141700.0 65135.0 140355.0 ;
      RECT  64430.0 141700.0 65135.0 143045.0 ;
      RECT  64430.0 144390.0 65135.0 143045.0 ;
      RECT  64430.0 144390.0 65135.0 145735.0 ;
      RECT  64430.0 147080.0 65135.0 145735.0 ;
      RECT  64430.0 147080.0 65135.0 148425.0 ;
      RECT  64430.0 149770.0 65135.0 148425.0 ;
      RECT  64430.0 149770.0 65135.0 151115.0 ;
      RECT  64430.0 152460.0 65135.0 151115.0 ;
      RECT  64430.0 152460.0 65135.0 153805.0 ;
      RECT  64430.0 155150.0 65135.0 153805.0 ;
      RECT  64430.0 155150.0 65135.0 156495.0 ;
      RECT  64430.0 157840.0 65135.0 156495.0 ;
      RECT  64430.0 157840.0 65135.0 159185.0 ;
      RECT  64430.0 160530.0 65135.0 159185.0 ;
      RECT  64430.0 160530.0 65135.0 161875.0 ;
      RECT  64430.0 163220.0 65135.0 161875.0 ;
      RECT  64430.0 163220.0 65135.0 164565.0 ;
      RECT  64430.0 165910.0 65135.0 164565.0 ;
      RECT  64430.0 165910.0 65135.0 167255.0 ;
      RECT  64430.0 168600.0 65135.0 167255.0 ;
      RECT  64430.0 168600.0 65135.0 169945.0 ;
      RECT  64430.0 171290.0 65135.0 169945.0 ;
      RECT  64430.0 171290.0 65135.0 172635.0 ;
      RECT  64430.0 173980.0 65135.0 172635.0 ;
      RECT  64430.0 173980.0 65135.0 175325.0 ;
      RECT  64430.0 176670.0 65135.0 175325.0 ;
      RECT  64430.0 176670.0 65135.0 178015.0 ;
      RECT  64430.0 179360.0 65135.0 178015.0 ;
      RECT  64430.0 179360.0 65135.0 180705.0 ;
      RECT  64430.0 182050.0 65135.0 180705.0 ;
      RECT  64430.0 182050.0 65135.0 183395.0 ;
      RECT  64430.0 184740.0 65135.0 183395.0 ;
      RECT  64430.0 184740.0 65135.0 186085.0 ;
      RECT  64430.0 187430.0 65135.0 186085.0 ;
      RECT  64430.0 187430.0 65135.0 188775.0 ;
      RECT  64430.0 190120.0 65135.0 188775.0 ;
      RECT  64430.0 190120.0 65135.0 191465.0 ;
      RECT  64430.0 192810.0 65135.0 191465.0 ;
      RECT  64430.0 192810.0 65135.0 194155.0 ;
      RECT  64430.0 195500.0 65135.0 194155.0 ;
      RECT  64430.0 195500.0 65135.0 196845.0 ;
      RECT  64430.0 198190.0 65135.0 196845.0 ;
      RECT  64430.0 198190.0 65135.0 199535.0 ;
      RECT  64430.0 200880.0 65135.0 199535.0 ;
      RECT  64430.0 200880.0 65135.0 202225.0 ;
      RECT  64430.0 203570.0 65135.0 202225.0 ;
      RECT  64430.0 203570.0 65135.0 204915.0 ;
      RECT  64430.0 206260.0 65135.0 204915.0 ;
      RECT  65135.0 34100.0 65840.0 35445.0 ;
      RECT  65135.0 36790.0 65840.0 35445.0 ;
      RECT  65135.0 36790.0 65840.0 38135.0 ;
      RECT  65135.0 39480.0 65840.0 38135.0 ;
      RECT  65135.0 39480.0 65840.0 40825.0 ;
      RECT  65135.0 42170.0 65840.0 40825.0 ;
      RECT  65135.0 42170.0 65840.0 43515.0 ;
      RECT  65135.0 44860.0 65840.0 43515.0 ;
      RECT  65135.0 44860.0 65840.0 46205.0 ;
      RECT  65135.0 47550.0 65840.0 46205.0 ;
      RECT  65135.0 47550.0 65840.0 48895.0 ;
      RECT  65135.0 50240.0 65840.0 48895.0 ;
      RECT  65135.0 50240.0 65840.0 51585.0 ;
      RECT  65135.0 52930.0 65840.0 51585.0 ;
      RECT  65135.0 52930.0 65840.0 54275.0 ;
      RECT  65135.0 55620.0 65840.0 54275.0 ;
      RECT  65135.0 55620.0 65840.0 56965.0 ;
      RECT  65135.0 58310.0 65840.0 56965.0 ;
      RECT  65135.0 58310.0 65840.0 59655.0 ;
      RECT  65135.0 61000.0 65840.0 59655.0 ;
      RECT  65135.0 61000.0 65840.0 62345.0 ;
      RECT  65135.0 63690.0 65840.0 62345.0 ;
      RECT  65135.0 63690.0 65840.0 65035.0 ;
      RECT  65135.0 66380.0 65840.0 65035.0 ;
      RECT  65135.0 66380.0 65840.0 67725.0 ;
      RECT  65135.0 69070.0 65840.0 67725.0 ;
      RECT  65135.0 69070.0 65840.0 70415.0 ;
      RECT  65135.0 71760.0 65840.0 70415.0 ;
      RECT  65135.0 71760.0 65840.0 73105.0 ;
      RECT  65135.0 74450.0 65840.0 73105.0 ;
      RECT  65135.0 74450.0 65840.0 75795.0 ;
      RECT  65135.0 77140.0 65840.0 75795.0 ;
      RECT  65135.0 77140.0 65840.0 78485.0 ;
      RECT  65135.0 79830.0 65840.0 78485.0 ;
      RECT  65135.0 79830.0 65840.0 81175.0 ;
      RECT  65135.0 82520.0 65840.0 81175.0 ;
      RECT  65135.0 82520.0 65840.0 83865.0 ;
      RECT  65135.0 85210.0 65840.0 83865.0 ;
      RECT  65135.0 85210.0 65840.0 86555.0 ;
      RECT  65135.0 87900.0 65840.0 86555.0 ;
      RECT  65135.0 87900.0 65840.0 89245.0 ;
      RECT  65135.0 90590.0 65840.0 89245.0 ;
      RECT  65135.0 90590.0 65840.0 91935.0 ;
      RECT  65135.0 93280.0 65840.0 91935.0 ;
      RECT  65135.0 93280.0 65840.0 94625.0 ;
      RECT  65135.0 95970.0 65840.0 94625.0 ;
      RECT  65135.0 95970.0 65840.0 97315.0 ;
      RECT  65135.0 98660.0 65840.0 97315.0 ;
      RECT  65135.0 98660.0 65840.0 100005.0 ;
      RECT  65135.0 101350.0 65840.0 100005.0 ;
      RECT  65135.0 101350.0 65840.0 102695.0 ;
      RECT  65135.0 104040.0 65840.0 102695.0 ;
      RECT  65135.0 104040.0 65840.0 105385.0 ;
      RECT  65135.0 106730.0 65840.0 105385.0 ;
      RECT  65135.0 106730.0 65840.0 108075.0 ;
      RECT  65135.0 109420.0 65840.0 108075.0 ;
      RECT  65135.0 109420.0 65840.0 110765.0 ;
      RECT  65135.0 112110.0 65840.0 110765.0 ;
      RECT  65135.0 112110.0 65840.0 113455.0 ;
      RECT  65135.0 114800.0 65840.0 113455.0 ;
      RECT  65135.0 114800.0 65840.0 116145.0 ;
      RECT  65135.0 117490.0 65840.0 116145.0 ;
      RECT  65135.0 117490.0 65840.0 118835.0 ;
      RECT  65135.0 120180.0 65840.0 118835.0 ;
      RECT  65135.0 120180.0 65840.0 121525.0 ;
      RECT  65135.0 122870.0 65840.0 121525.0 ;
      RECT  65135.0 122870.0 65840.0 124215.0 ;
      RECT  65135.0 125560.0 65840.0 124215.0 ;
      RECT  65135.0 125560.0 65840.0 126905.0 ;
      RECT  65135.0 128250.0 65840.0 126905.0 ;
      RECT  65135.0 128250.0 65840.0 129595.0 ;
      RECT  65135.0 130940.0 65840.0 129595.0 ;
      RECT  65135.0 130940.0 65840.0 132285.0 ;
      RECT  65135.0 133630.0 65840.0 132285.0 ;
      RECT  65135.0 133630.0 65840.0 134975.0 ;
      RECT  65135.0 136320.0 65840.0 134975.0 ;
      RECT  65135.0 136320.0 65840.0 137665.0 ;
      RECT  65135.0 139010.0 65840.0 137665.0 ;
      RECT  65135.0 139010.0 65840.0 140355.0 ;
      RECT  65135.0 141700.0 65840.0 140355.0 ;
      RECT  65135.0 141700.0 65840.0 143045.0 ;
      RECT  65135.0 144390.0 65840.0 143045.0 ;
      RECT  65135.0 144390.0 65840.0 145735.0 ;
      RECT  65135.0 147080.0 65840.0 145735.0 ;
      RECT  65135.0 147080.0 65840.0 148425.0 ;
      RECT  65135.0 149770.0 65840.0 148425.0 ;
      RECT  65135.0 149770.0 65840.0 151115.0 ;
      RECT  65135.0 152460.0 65840.0 151115.0 ;
      RECT  65135.0 152460.0 65840.0 153805.0 ;
      RECT  65135.0 155150.0 65840.0 153805.0 ;
      RECT  65135.0 155150.0 65840.0 156495.0 ;
      RECT  65135.0 157840.0 65840.0 156495.0 ;
      RECT  65135.0 157840.0 65840.0 159185.0 ;
      RECT  65135.0 160530.0 65840.0 159185.0 ;
      RECT  65135.0 160530.0 65840.0 161875.0 ;
      RECT  65135.0 163220.0 65840.0 161875.0 ;
      RECT  65135.0 163220.0 65840.0 164565.0 ;
      RECT  65135.0 165910.0 65840.0 164565.0 ;
      RECT  65135.0 165910.0 65840.0 167255.0 ;
      RECT  65135.0 168600.0 65840.0 167255.0 ;
      RECT  65135.0 168600.0 65840.0 169945.0 ;
      RECT  65135.0 171290.0 65840.0 169945.0 ;
      RECT  65135.0 171290.0 65840.0 172635.0 ;
      RECT  65135.0 173980.0 65840.0 172635.0 ;
      RECT  65135.0 173980.0 65840.0 175325.0 ;
      RECT  65135.0 176670.0 65840.0 175325.0 ;
      RECT  65135.0 176670.0 65840.0 178015.0 ;
      RECT  65135.0 179360.0 65840.0 178015.0 ;
      RECT  65135.0 179360.0 65840.0 180705.0 ;
      RECT  65135.0 182050.0 65840.0 180705.0 ;
      RECT  65135.0 182050.0 65840.0 183395.0 ;
      RECT  65135.0 184740.0 65840.0 183395.0 ;
      RECT  65135.0 184740.0 65840.0 186085.0 ;
      RECT  65135.0 187430.0 65840.0 186085.0 ;
      RECT  65135.0 187430.0 65840.0 188775.0 ;
      RECT  65135.0 190120.0 65840.0 188775.0 ;
      RECT  65135.0 190120.0 65840.0 191465.0 ;
      RECT  65135.0 192810.0 65840.0 191465.0 ;
      RECT  65135.0 192810.0 65840.0 194155.0 ;
      RECT  65135.0 195500.0 65840.0 194155.0 ;
      RECT  65135.0 195500.0 65840.0 196845.0 ;
      RECT  65135.0 198190.0 65840.0 196845.0 ;
      RECT  65135.0 198190.0 65840.0 199535.0 ;
      RECT  65135.0 200880.0 65840.0 199535.0 ;
      RECT  65135.0 200880.0 65840.0 202225.0 ;
      RECT  65135.0 203570.0 65840.0 202225.0 ;
      RECT  65135.0 203570.0 65840.0 204915.0 ;
      RECT  65135.0 206260.0 65840.0 204915.0 ;
      RECT  65840.0 34100.0 66545.0 35445.0 ;
      RECT  65840.0 36790.0 66545.0 35445.0 ;
      RECT  65840.0 36790.0 66545.0 38135.0 ;
      RECT  65840.0 39480.0 66545.0 38135.0 ;
      RECT  65840.0 39480.0 66545.0 40825.0 ;
      RECT  65840.0 42170.0 66545.0 40825.0 ;
      RECT  65840.0 42170.0 66545.0 43515.0 ;
      RECT  65840.0 44860.0 66545.0 43515.0 ;
      RECT  65840.0 44860.0 66545.0 46205.0 ;
      RECT  65840.0 47550.0 66545.0 46205.0 ;
      RECT  65840.0 47550.0 66545.0 48895.0 ;
      RECT  65840.0 50240.0 66545.0 48895.0 ;
      RECT  65840.0 50240.0 66545.0 51585.0 ;
      RECT  65840.0 52930.0 66545.0 51585.0 ;
      RECT  65840.0 52930.0 66545.0 54275.0 ;
      RECT  65840.0 55620.0 66545.0 54275.0 ;
      RECT  65840.0 55620.0 66545.0 56965.0 ;
      RECT  65840.0 58310.0 66545.0 56965.0 ;
      RECT  65840.0 58310.0 66545.0 59655.0 ;
      RECT  65840.0 61000.0 66545.0 59655.0 ;
      RECT  65840.0 61000.0 66545.0 62345.0 ;
      RECT  65840.0 63690.0 66545.0 62345.0 ;
      RECT  65840.0 63690.0 66545.0 65035.0 ;
      RECT  65840.0 66380.0 66545.0 65035.0 ;
      RECT  65840.0 66380.0 66545.0 67725.0 ;
      RECT  65840.0 69070.0 66545.0 67725.0 ;
      RECT  65840.0 69070.0 66545.0 70415.0 ;
      RECT  65840.0 71760.0 66545.0 70415.0 ;
      RECT  65840.0 71760.0 66545.0 73105.0 ;
      RECT  65840.0 74450.0 66545.0 73105.0 ;
      RECT  65840.0 74450.0 66545.0 75795.0 ;
      RECT  65840.0 77140.0 66545.0 75795.0 ;
      RECT  65840.0 77140.0 66545.0 78485.0 ;
      RECT  65840.0 79830.0 66545.0 78485.0 ;
      RECT  65840.0 79830.0 66545.0 81175.0 ;
      RECT  65840.0 82520.0 66545.0 81175.0 ;
      RECT  65840.0 82520.0 66545.0 83865.0 ;
      RECT  65840.0 85210.0 66545.0 83865.0 ;
      RECT  65840.0 85210.0 66545.0 86555.0 ;
      RECT  65840.0 87900.0 66545.0 86555.0 ;
      RECT  65840.0 87900.0 66545.0 89245.0 ;
      RECT  65840.0 90590.0 66545.0 89245.0 ;
      RECT  65840.0 90590.0 66545.0 91935.0 ;
      RECT  65840.0 93280.0 66545.0 91935.0 ;
      RECT  65840.0 93280.0 66545.0 94625.0 ;
      RECT  65840.0 95970.0 66545.0 94625.0 ;
      RECT  65840.0 95970.0 66545.0 97315.0 ;
      RECT  65840.0 98660.0 66545.0 97315.0 ;
      RECT  65840.0 98660.0 66545.0 100005.0 ;
      RECT  65840.0 101350.0 66545.0 100005.0 ;
      RECT  65840.0 101350.0 66545.0 102695.0 ;
      RECT  65840.0 104040.0 66545.0 102695.0 ;
      RECT  65840.0 104040.0 66545.0 105385.0 ;
      RECT  65840.0 106730.0 66545.0 105385.0 ;
      RECT  65840.0 106730.0 66545.0 108075.0 ;
      RECT  65840.0 109420.0 66545.0 108075.0 ;
      RECT  65840.0 109420.0 66545.0 110765.0 ;
      RECT  65840.0 112110.0 66545.0 110765.0 ;
      RECT  65840.0 112110.0 66545.0 113455.0 ;
      RECT  65840.0 114800.0 66545.0 113455.0 ;
      RECT  65840.0 114800.0 66545.0 116145.0 ;
      RECT  65840.0 117490.0 66545.0 116145.0 ;
      RECT  65840.0 117490.0 66545.0 118835.0 ;
      RECT  65840.0 120180.0 66545.0 118835.0 ;
      RECT  65840.0 120180.0 66545.0 121525.0 ;
      RECT  65840.0 122870.0 66545.0 121525.0 ;
      RECT  65840.0 122870.0 66545.0 124215.0 ;
      RECT  65840.0 125560.0 66545.0 124215.0 ;
      RECT  65840.0 125560.0 66545.0 126905.0 ;
      RECT  65840.0 128250.0 66545.0 126905.0 ;
      RECT  65840.0 128250.0 66545.0 129595.0 ;
      RECT  65840.0 130940.0 66545.0 129595.0 ;
      RECT  65840.0 130940.0 66545.0 132285.0 ;
      RECT  65840.0 133630.0 66545.0 132285.0 ;
      RECT  65840.0 133630.0 66545.0 134975.0 ;
      RECT  65840.0 136320.0 66545.0 134975.0 ;
      RECT  65840.0 136320.0 66545.0 137665.0 ;
      RECT  65840.0 139010.0 66545.0 137665.0 ;
      RECT  65840.0 139010.0 66545.0 140355.0 ;
      RECT  65840.0 141700.0 66545.0 140355.0 ;
      RECT  65840.0 141700.0 66545.0 143045.0 ;
      RECT  65840.0 144390.0 66545.0 143045.0 ;
      RECT  65840.0 144390.0 66545.0 145735.0 ;
      RECT  65840.0 147080.0 66545.0 145735.0 ;
      RECT  65840.0 147080.0 66545.0 148425.0 ;
      RECT  65840.0 149770.0 66545.0 148425.0 ;
      RECT  65840.0 149770.0 66545.0 151115.0 ;
      RECT  65840.0 152460.0 66545.0 151115.0 ;
      RECT  65840.0 152460.0 66545.0 153805.0 ;
      RECT  65840.0 155150.0 66545.0 153805.0 ;
      RECT  65840.0 155150.0 66545.0 156495.0 ;
      RECT  65840.0 157840.0 66545.0 156495.0 ;
      RECT  65840.0 157840.0 66545.0 159185.0 ;
      RECT  65840.0 160530.0 66545.0 159185.0 ;
      RECT  65840.0 160530.0 66545.0 161875.0 ;
      RECT  65840.0 163220.0 66545.0 161875.0 ;
      RECT  65840.0 163220.0 66545.0 164565.0 ;
      RECT  65840.0 165910.0 66545.0 164565.0 ;
      RECT  65840.0 165910.0 66545.0 167255.0 ;
      RECT  65840.0 168600.0 66545.0 167255.0 ;
      RECT  65840.0 168600.0 66545.0 169945.0 ;
      RECT  65840.0 171290.0 66545.0 169945.0 ;
      RECT  65840.0 171290.0 66545.0 172635.0 ;
      RECT  65840.0 173980.0 66545.0 172635.0 ;
      RECT  65840.0 173980.0 66545.0 175325.0 ;
      RECT  65840.0 176670.0 66545.0 175325.0 ;
      RECT  65840.0 176670.0 66545.0 178015.0 ;
      RECT  65840.0 179360.0 66545.0 178015.0 ;
      RECT  65840.0 179360.0 66545.0 180705.0 ;
      RECT  65840.0 182050.0 66545.0 180705.0 ;
      RECT  65840.0 182050.0 66545.0 183395.0 ;
      RECT  65840.0 184740.0 66545.0 183395.0 ;
      RECT  65840.0 184740.0 66545.0 186085.0 ;
      RECT  65840.0 187430.0 66545.0 186085.0 ;
      RECT  65840.0 187430.0 66545.0 188775.0 ;
      RECT  65840.0 190120.0 66545.0 188775.0 ;
      RECT  65840.0 190120.0 66545.0 191465.0 ;
      RECT  65840.0 192810.0 66545.0 191465.0 ;
      RECT  65840.0 192810.0 66545.0 194155.0 ;
      RECT  65840.0 195500.0 66545.0 194155.0 ;
      RECT  65840.0 195500.0 66545.0 196845.0 ;
      RECT  65840.0 198190.0 66545.0 196845.0 ;
      RECT  65840.0 198190.0 66545.0 199535.0 ;
      RECT  65840.0 200880.0 66545.0 199535.0 ;
      RECT  65840.0 200880.0 66545.0 202225.0 ;
      RECT  65840.0 203570.0 66545.0 202225.0 ;
      RECT  65840.0 203570.0 66545.0 204915.0 ;
      RECT  65840.0 206260.0 66545.0 204915.0 ;
      RECT  66545.0 34100.0 67250.0 35445.0 ;
      RECT  66545.0 36790.0 67250.0 35445.0 ;
      RECT  66545.0 36790.0 67250.0 38135.0 ;
      RECT  66545.0 39480.0 67250.0 38135.0 ;
      RECT  66545.0 39480.0 67250.0 40825.0 ;
      RECT  66545.0 42170.0 67250.0 40825.0 ;
      RECT  66545.0 42170.0 67250.0 43515.0 ;
      RECT  66545.0 44860.0 67250.0 43515.0 ;
      RECT  66545.0 44860.0 67250.0 46205.0 ;
      RECT  66545.0 47550.0 67250.0 46205.0 ;
      RECT  66545.0 47550.0 67250.0 48895.0 ;
      RECT  66545.0 50240.0 67250.0 48895.0 ;
      RECT  66545.0 50240.0 67250.0 51585.0 ;
      RECT  66545.0 52930.0 67250.0 51585.0 ;
      RECT  66545.0 52930.0 67250.0 54275.0 ;
      RECT  66545.0 55620.0 67250.0 54275.0 ;
      RECT  66545.0 55620.0 67250.0 56965.0 ;
      RECT  66545.0 58310.0 67250.0 56965.0 ;
      RECT  66545.0 58310.0 67250.0 59655.0 ;
      RECT  66545.0 61000.0 67250.0 59655.0 ;
      RECT  66545.0 61000.0 67250.0 62345.0 ;
      RECT  66545.0 63690.0 67250.0 62345.0 ;
      RECT  66545.0 63690.0 67250.0 65035.0 ;
      RECT  66545.0 66380.0 67250.0 65035.0 ;
      RECT  66545.0 66380.0 67250.0 67725.0 ;
      RECT  66545.0 69070.0 67250.0 67725.0 ;
      RECT  66545.0 69070.0 67250.0 70415.0 ;
      RECT  66545.0 71760.0 67250.0 70415.0 ;
      RECT  66545.0 71760.0 67250.0 73105.0 ;
      RECT  66545.0 74450.0 67250.0 73105.0 ;
      RECT  66545.0 74450.0 67250.0 75795.0 ;
      RECT  66545.0 77140.0 67250.0 75795.0 ;
      RECT  66545.0 77140.0 67250.0 78485.0 ;
      RECT  66545.0 79830.0 67250.0 78485.0 ;
      RECT  66545.0 79830.0 67250.0 81175.0 ;
      RECT  66545.0 82520.0 67250.0 81175.0 ;
      RECT  66545.0 82520.0 67250.0 83865.0 ;
      RECT  66545.0 85210.0 67250.0 83865.0 ;
      RECT  66545.0 85210.0 67250.0 86555.0 ;
      RECT  66545.0 87900.0 67250.0 86555.0 ;
      RECT  66545.0 87900.0 67250.0 89245.0 ;
      RECT  66545.0 90590.0 67250.0 89245.0 ;
      RECT  66545.0 90590.0 67250.0 91935.0 ;
      RECT  66545.0 93280.0 67250.0 91935.0 ;
      RECT  66545.0 93280.0 67250.0 94625.0 ;
      RECT  66545.0 95970.0 67250.0 94625.0 ;
      RECT  66545.0 95970.0 67250.0 97315.0 ;
      RECT  66545.0 98660.0 67250.0 97315.0 ;
      RECT  66545.0 98660.0 67250.0 100005.0 ;
      RECT  66545.0 101350.0 67250.0 100005.0 ;
      RECT  66545.0 101350.0 67250.0 102695.0 ;
      RECT  66545.0 104040.0 67250.0 102695.0 ;
      RECT  66545.0 104040.0 67250.0 105385.0 ;
      RECT  66545.0 106730.0 67250.0 105385.0 ;
      RECT  66545.0 106730.0 67250.0 108075.0 ;
      RECT  66545.0 109420.0 67250.0 108075.0 ;
      RECT  66545.0 109420.0 67250.0 110765.0 ;
      RECT  66545.0 112110.0 67250.0 110765.0 ;
      RECT  66545.0 112110.0 67250.0 113455.0 ;
      RECT  66545.0 114800.0 67250.0 113455.0 ;
      RECT  66545.0 114800.0 67250.0 116145.0 ;
      RECT  66545.0 117490.0 67250.0 116145.0 ;
      RECT  66545.0 117490.0 67250.0 118835.0 ;
      RECT  66545.0 120180.0 67250.0 118835.0 ;
      RECT  66545.0 120180.0 67250.0 121525.0 ;
      RECT  66545.0 122870.0 67250.0 121525.0 ;
      RECT  66545.0 122870.0 67250.0 124215.0 ;
      RECT  66545.0 125560.0 67250.0 124215.0 ;
      RECT  66545.0 125560.0 67250.0 126905.0 ;
      RECT  66545.0 128250.0 67250.0 126905.0 ;
      RECT  66545.0 128250.0 67250.0 129595.0 ;
      RECT  66545.0 130940.0 67250.0 129595.0 ;
      RECT  66545.0 130940.0 67250.0 132285.0 ;
      RECT  66545.0 133630.0 67250.0 132285.0 ;
      RECT  66545.0 133630.0 67250.0 134975.0 ;
      RECT  66545.0 136320.0 67250.0 134975.0 ;
      RECT  66545.0 136320.0 67250.0 137665.0 ;
      RECT  66545.0 139010.0 67250.0 137665.0 ;
      RECT  66545.0 139010.0 67250.0 140355.0 ;
      RECT  66545.0 141700.0 67250.0 140355.0 ;
      RECT  66545.0 141700.0 67250.0 143045.0 ;
      RECT  66545.0 144390.0 67250.0 143045.0 ;
      RECT  66545.0 144390.0 67250.0 145735.0 ;
      RECT  66545.0 147080.0 67250.0 145735.0 ;
      RECT  66545.0 147080.0 67250.0 148425.0 ;
      RECT  66545.0 149770.0 67250.0 148425.0 ;
      RECT  66545.0 149770.0 67250.0 151115.0 ;
      RECT  66545.0 152460.0 67250.0 151115.0 ;
      RECT  66545.0 152460.0 67250.0 153805.0 ;
      RECT  66545.0 155150.0 67250.0 153805.0 ;
      RECT  66545.0 155150.0 67250.0 156495.0 ;
      RECT  66545.0 157840.0 67250.0 156495.0 ;
      RECT  66545.0 157840.0 67250.0 159185.0 ;
      RECT  66545.0 160530.0 67250.0 159185.0 ;
      RECT  66545.0 160530.0 67250.0 161875.0 ;
      RECT  66545.0 163220.0 67250.0 161875.0 ;
      RECT  66545.0 163220.0 67250.0 164565.0 ;
      RECT  66545.0 165910.0 67250.0 164565.0 ;
      RECT  66545.0 165910.0 67250.0 167255.0 ;
      RECT  66545.0 168600.0 67250.0 167255.0 ;
      RECT  66545.0 168600.0 67250.0 169945.0 ;
      RECT  66545.0 171290.0 67250.0 169945.0 ;
      RECT  66545.0 171290.0 67250.0 172635.0 ;
      RECT  66545.0 173980.0 67250.0 172635.0 ;
      RECT  66545.0 173980.0 67250.0 175325.0 ;
      RECT  66545.0 176670.0 67250.0 175325.0 ;
      RECT  66545.0 176670.0 67250.0 178015.0 ;
      RECT  66545.0 179360.0 67250.0 178015.0 ;
      RECT  66545.0 179360.0 67250.0 180705.0 ;
      RECT  66545.0 182050.0 67250.0 180705.0 ;
      RECT  66545.0 182050.0 67250.0 183395.0 ;
      RECT  66545.0 184740.0 67250.0 183395.0 ;
      RECT  66545.0 184740.0 67250.0 186085.0 ;
      RECT  66545.0 187430.0 67250.0 186085.0 ;
      RECT  66545.0 187430.0 67250.0 188775.0 ;
      RECT  66545.0 190120.0 67250.0 188775.0 ;
      RECT  66545.0 190120.0 67250.0 191465.0 ;
      RECT  66545.0 192810.0 67250.0 191465.0 ;
      RECT  66545.0 192810.0 67250.0 194155.0 ;
      RECT  66545.0 195500.0 67250.0 194155.0 ;
      RECT  66545.0 195500.0 67250.0 196845.0 ;
      RECT  66545.0 198190.0 67250.0 196845.0 ;
      RECT  66545.0 198190.0 67250.0 199535.0 ;
      RECT  66545.0 200880.0 67250.0 199535.0 ;
      RECT  66545.0 200880.0 67250.0 202225.0 ;
      RECT  66545.0 203570.0 67250.0 202225.0 ;
      RECT  66545.0 203570.0 67250.0 204915.0 ;
      RECT  66545.0 206260.0 67250.0 204915.0 ;
      RECT  67250.0 34100.0 67955.0 35445.0 ;
      RECT  67250.0 36790.0 67955.0 35445.0 ;
      RECT  67250.0 36790.0 67955.0 38135.0 ;
      RECT  67250.0 39480.0 67955.0 38135.0 ;
      RECT  67250.0 39480.0 67955.0 40825.0 ;
      RECT  67250.0 42170.0 67955.0 40825.0 ;
      RECT  67250.0 42170.0 67955.0 43515.0 ;
      RECT  67250.0 44860.0 67955.0 43515.0 ;
      RECT  67250.0 44860.0 67955.0 46205.0 ;
      RECT  67250.0 47550.0 67955.0 46205.0 ;
      RECT  67250.0 47550.0 67955.0 48895.0 ;
      RECT  67250.0 50240.0 67955.0 48895.0 ;
      RECT  67250.0 50240.0 67955.0 51585.0 ;
      RECT  67250.0 52930.0 67955.0 51585.0 ;
      RECT  67250.0 52930.0 67955.0 54275.0 ;
      RECT  67250.0 55620.0 67955.0 54275.0 ;
      RECT  67250.0 55620.0 67955.0 56965.0 ;
      RECT  67250.0 58310.0 67955.0 56965.0 ;
      RECT  67250.0 58310.0 67955.0 59655.0 ;
      RECT  67250.0 61000.0 67955.0 59655.0 ;
      RECT  67250.0 61000.0 67955.0 62345.0 ;
      RECT  67250.0 63690.0 67955.0 62345.0 ;
      RECT  67250.0 63690.0 67955.0 65035.0 ;
      RECT  67250.0 66380.0 67955.0 65035.0 ;
      RECT  67250.0 66380.0 67955.0 67725.0 ;
      RECT  67250.0 69070.0 67955.0 67725.0 ;
      RECT  67250.0 69070.0 67955.0 70415.0 ;
      RECT  67250.0 71760.0 67955.0 70415.0 ;
      RECT  67250.0 71760.0 67955.0 73105.0 ;
      RECT  67250.0 74450.0 67955.0 73105.0 ;
      RECT  67250.0 74450.0 67955.0 75795.0 ;
      RECT  67250.0 77140.0 67955.0 75795.0 ;
      RECT  67250.0 77140.0 67955.0 78485.0 ;
      RECT  67250.0 79830.0 67955.0 78485.0 ;
      RECT  67250.0 79830.0 67955.0 81175.0 ;
      RECT  67250.0 82520.0 67955.0 81175.0 ;
      RECT  67250.0 82520.0 67955.0 83865.0 ;
      RECT  67250.0 85210.0 67955.0 83865.0 ;
      RECT  67250.0 85210.0 67955.0 86555.0 ;
      RECT  67250.0 87900.0 67955.0 86555.0 ;
      RECT  67250.0 87900.0 67955.0 89245.0 ;
      RECT  67250.0 90590.0 67955.0 89245.0 ;
      RECT  67250.0 90590.0 67955.0 91935.0 ;
      RECT  67250.0 93280.0 67955.0 91935.0 ;
      RECT  67250.0 93280.0 67955.0 94625.0 ;
      RECT  67250.0 95970.0 67955.0 94625.0 ;
      RECT  67250.0 95970.0 67955.0 97315.0 ;
      RECT  67250.0 98660.0 67955.0 97315.0 ;
      RECT  67250.0 98660.0 67955.0 100005.0 ;
      RECT  67250.0 101350.0 67955.0 100005.0 ;
      RECT  67250.0 101350.0 67955.0 102695.0 ;
      RECT  67250.0 104040.0 67955.0 102695.0 ;
      RECT  67250.0 104040.0 67955.0 105385.0 ;
      RECT  67250.0 106730.0 67955.0 105385.0 ;
      RECT  67250.0 106730.0 67955.0 108075.0 ;
      RECT  67250.0 109420.0 67955.0 108075.0 ;
      RECT  67250.0 109420.0 67955.0 110765.0 ;
      RECT  67250.0 112110.0 67955.0 110765.0 ;
      RECT  67250.0 112110.0 67955.0 113455.0 ;
      RECT  67250.0 114800.0 67955.0 113455.0 ;
      RECT  67250.0 114800.0 67955.0 116145.0 ;
      RECT  67250.0 117490.0 67955.0 116145.0 ;
      RECT  67250.0 117490.0 67955.0 118835.0 ;
      RECT  67250.0 120180.0 67955.0 118835.0 ;
      RECT  67250.0 120180.0 67955.0 121525.0 ;
      RECT  67250.0 122870.0 67955.0 121525.0 ;
      RECT  67250.0 122870.0 67955.0 124215.0 ;
      RECT  67250.0 125560.0 67955.0 124215.0 ;
      RECT  67250.0 125560.0 67955.0 126905.0 ;
      RECT  67250.0 128250.0 67955.0 126905.0 ;
      RECT  67250.0 128250.0 67955.0 129595.0 ;
      RECT  67250.0 130940.0 67955.0 129595.0 ;
      RECT  67250.0 130940.0 67955.0 132285.0 ;
      RECT  67250.0 133630.0 67955.0 132285.0 ;
      RECT  67250.0 133630.0 67955.0 134975.0 ;
      RECT  67250.0 136320.0 67955.0 134975.0 ;
      RECT  67250.0 136320.0 67955.0 137665.0 ;
      RECT  67250.0 139010.0 67955.0 137665.0 ;
      RECT  67250.0 139010.0 67955.0 140355.0 ;
      RECT  67250.0 141700.0 67955.0 140355.0 ;
      RECT  67250.0 141700.0 67955.0 143045.0 ;
      RECT  67250.0 144390.0 67955.0 143045.0 ;
      RECT  67250.0 144390.0 67955.0 145735.0 ;
      RECT  67250.0 147080.0 67955.0 145735.0 ;
      RECT  67250.0 147080.0 67955.0 148425.0 ;
      RECT  67250.0 149770.0 67955.0 148425.0 ;
      RECT  67250.0 149770.0 67955.0 151115.0 ;
      RECT  67250.0 152460.0 67955.0 151115.0 ;
      RECT  67250.0 152460.0 67955.0 153805.0 ;
      RECT  67250.0 155150.0 67955.0 153805.0 ;
      RECT  67250.0 155150.0 67955.0 156495.0 ;
      RECT  67250.0 157840.0 67955.0 156495.0 ;
      RECT  67250.0 157840.0 67955.0 159185.0 ;
      RECT  67250.0 160530.0 67955.0 159185.0 ;
      RECT  67250.0 160530.0 67955.0 161875.0 ;
      RECT  67250.0 163220.0 67955.0 161875.0 ;
      RECT  67250.0 163220.0 67955.0 164565.0 ;
      RECT  67250.0 165910.0 67955.0 164565.0 ;
      RECT  67250.0 165910.0 67955.0 167255.0 ;
      RECT  67250.0 168600.0 67955.0 167255.0 ;
      RECT  67250.0 168600.0 67955.0 169945.0 ;
      RECT  67250.0 171290.0 67955.0 169945.0 ;
      RECT  67250.0 171290.0 67955.0 172635.0 ;
      RECT  67250.0 173980.0 67955.0 172635.0 ;
      RECT  67250.0 173980.0 67955.0 175325.0 ;
      RECT  67250.0 176670.0 67955.0 175325.0 ;
      RECT  67250.0 176670.0 67955.0 178015.0 ;
      RECT  67250.0 179360.0 67955.0 178015.0 ;
      RECT  67250.0 179360.0 67955.0 180705.0 ;
      RECT  67250.0 182050.0 67955.0 180705.0 ;
      RECT  67250.0 182050.0 67955.0 183395.0 ;
      RECT  67250.0 184740.0 67955.0 183395.0 ;
      RECT  67250.0 184740.0 67955.0 186085.0 ;
      RECT  67250.0 187430.0 67955.0 186085.0 ;
      RECT  67250.0 187430.0 67955.0 188775.0 ;
      RECT  67250.0 190120.0 67955.0 188775.0 ;
      RECT  67250.0 190120.0 67955.0 191465.0 ;
      RECT  67250.0 192810.0 67955.0 191465.0 ;
      RECT  67250.0 192810.0 67955.0 194155.0 ;
      RECT  67250.0 195500.0 67955.0 194155.0 ;
      RECT  67250.0 195500.0 67955.0 196845.0 ;
      RECT  67250.0 198190.0 67955.0 196845.0 ;
      RECT  67250.0 198190.0 67955.0 199535.0 ;
      RECT  67250.0 200880.0 67955.0 199535.0 ;
      RECT  67250.0 200880.0 67955.0 202225.0 ;
      RECT  67250.0 203570.0 67955.0 202225.0 ;
      RECT  67250.0 203570.0 67955.0 204915.0 ;
      RECT  67250.0 206260.0 67955.0 204915.0 ;
      RECT  67955.0 34100.0 68660.0 35445.0 ;
      RECT  67955.0 36790.0 68660.0 35445.0 ;
      RECT  67955.0 36790.0 68660.0 38135.0 ;
      RECT  67955.0 39480.0 68660.0 38135.0 ;
      RECT  67955.0 39480.0 68660.0 40825.0 ;
      RECT  67955.0 42170.0 68660.0 40825.0 ;
      RECT  67955.0 42170.0 68660.0 43515.0 ;
      RECT  67955.0 44860.0 68660.0 43515.0 ;
      RECT  67955.0 44860.0 68660.0 46205.0 ;
      RECT  67955.0 47550.0 68660.0 46205.0 ;
      RECT  67955.0 47550.0 68660.0 48895.0 ;
      RECT  67955.0 50240.0 68660.0 48895.0 ;
      RECT  67955.0 50240.0 68660.0 51585.0 ;
      RECT  67955.0 52930.0 68660.0 51585.0 ;
      RECT  67955.0 52930.0 68660.0 54275.0 ;
      RECT  67955.0 55620.0 68660.0 54275.0 ;
      RECT  67955.0 55620.0 68660.0 56965.0 ;
      RECT  67955.0 58310.0 68660.0 56965.0 ;
      RECT  67955.0 58310.0 68660.0 59655.0 ;
      RECT  67955.0 61000.0 68660.0 59655.0 ;
      RECT  67955.0 61000.0 68660.0 62345.0 ;
      RECT  67955.0 63690.0 68660.0 62345.0 ;
      RECT  67955.0 63690.0 68660.0 65035.0 ;
      RECT  67955.0 66380.0 68660.0 65035.0 ;
      RECT  67955.0 66380.0 68660.0 67725.0 ;
      RECT  67955.0 69070.0 68660.0 67725.0 ;
      RECT  67955.0 69070.0 68660.0 70415.0 ;
      RECT  67955.0 71760.0 68660.0 70415.0 ;
      RECT  67955.0 71760.0 68660.0 73105.0 ;
      RECT  67955.0 74450.0 68660.0 73105.0 ;
      RECT  67955.0 74450.0 68660.0 75795.0 ;
      RECT  67955.0 77140.0 68660.0 75795.0 ;
      RECT  67955.0 77140.0 68660.0 78485.0 ;
      RECT  67955.0 79830.0 68660.0 78485.0 ;
      RECT  67955.0 79830.0 68660.0 81175.0 ;
      RECT  67955.0 82520.0 68660.0 81175.0 ;
      RECT  67955.0 82520.0 68660.0 83865.0 ;
      RECT  67955.0 85210.0 68660.0 83865.0 ;
      RECT  67955.0 85210.0 68660.0 86555.0 ;
      RECT  67955.0 87900.0 68660.0 86555.0 ;
      RECT  67955.0 87900.0 68660.0 89245.0 ;
      RECT  67955.0 90590.0 68660.0 89245.0 ;
      RECT  67955.0 90590.0 68660.0 91935.0 ;
      RECT  67955.0 93280.0 68660.0 91935.0 ;
      RECT  67955.0 93280.0 68660.0 94625.0 ;
      RECT  67955.0 95970.0 68660.0 94625.0 ;
      RECT  67955.0 95970.0 68660.0 97315.0 ;
      RECT  67955.0 98660.0 68660.0 97315.0 ;
      RECT  67955.0 98660.0 68660.0 100005.0 ;
      RECT  67955.0 101350.0 68660.0 100005.0 ;
      RECT  67955.0 101350.0 68660.0 102695.0 ;
      RECT  67955.0 104040.0 68660.0 102695.0 ;
      RECT  67955.0 104040.0 68660.0 105385.0 ;
      RECT  67955.0 106730.0 68660.0 105385.0 ;
      RECT  67955.0 106730.0 68660.0 108075.0 ;
      RECT  67955.0 109420.0 68660.0 108075.0 ;
      RECT  67955.0 109420.0 68660.0 110765.0 ;
      RECT  67955.0 112110.0 68660.0 110765.0 ;
      RECT  67955.0 112110.0 68660.0 113455.0 ;
      RECT  67955.0 114800.0 68660.0 113455.0 ;
      RECT  67955.0 114800.0 68660.0 116145.0 ;
      RECT  67955.0 117490.0 68660.0 116145.0 ;
      RECT  67955.0 117490.0 68660.0 118835.0 ;
      RECT  67955.0 120180.0 68660.0 118835.0 ;
      RECT  67955.0 120180.0 68660.0 121525.0 ;
      RECT  67955.0 122870.0 68660.0 121525.0 ;
      RECT  67955.0 122870.0 68660.0 124215.0 ;
      RECT  67955.0 125560.0 68660.0 124215.0 ;
      RECT  67955.0 125560.0 68660.0 126905.0 ;
      RECT  67955.0 128250.0 68660.0 126905.0 ;
      RECT  67955.0 128250.0 68660.0 129595.0 ;
      RECT  67955.0 130940.0 68660.0 129595.0 ;
      RECT  67955.0 130940.0 68660.0 132285.0 ;
      RECT  67955.0 133630.0 68660.0 132285.0 ;
      RECT  67955.0 133630.0 68660.0 134975.0 ;
      RECT  67955.0 136320.0 68660.0 134975.0 ;
      RECT  67955.0 136320.0 68660.0 137665.0 ;
      RECT  67955.0 139010.0 68660.0 137665.0 ;
      RECT  67955.0 139010.0 68660.0 140355.0 ;
      RECT  67955.0 141700.0 68660.0 140355.0 ;
      RECT  67955.0 141700.0 68660.0 143045.0 ;
      RECT  67955.0 144390.0 68660.0 143045.0 ;
      RECT  67955.0 144390.0 68660.0 145735.0 ;
      RECT  67955.0 147080.0 68660.0 145735.0 ;
      RECT  67955.0 147080.0 68660.0 148425.0 ;
      RECT  67955.0 149770.0 68660.0 148425.0 ;
      RECT  67955.0 149770.0 68660.0 151115.0 ;
      RECT  67955.0 152460.0 68660.0 151115.0 ;
      RECT  67955.0 152460.0 68660.0 153805.0 ;
      RECT  67955.0 155150.0 68660.0 153805.0 ;
      RECT  67955.0 155150.0 68660.0 156495.0 ;
      RECT  67955.0 157840.0 68660.0 156495.0 ;
      RECT  67955.0 157840.0 68660.0 159185.0 ;
      RECT  67955.0 160530.0 68660.0 159185.0 ;
      RECT  67955.0 160530.0 68660.0 161875.0 ;
      RECT  67955.0 163220.0 68660.0 161875.0 ;
      RECT  67955.0 163220.0 68660.0 164565.0 ;
      RECT  67955.0 165910.0 68660.0 164565.0 ;
      RECT  67955.0 165910.0 68660.0 167255.0 ;
      RECT  67955.0 168600.0 68660.0 167255.0 ;
      RECT  67955.0 168600.0 68660.0 169945.0 ;
      RECT  67955.0 171290.0 68660.0 169945.0 ;
      RECT  67955.0 171290.0 68660.0 172635.0 ;
      RECT  67955.0 173980.0 68660.0 172635.0 ;
      RECT  67955.0 173980.0 68660.0 175325.0 ;
      RECT  67955.0 176670.0 68660.0 175325.0 ;
      RECT  67955.0 176670.0 68660.0 178015.0 ;
      RECT  67955.0 179360.0 68660.0 178015.0 ;
      RECT  67955.0 179360.0 68660.0 180705.0 ;
      RECT  67955.0 182050.0 68660.0 180705.0 ;
      RECT  67955.0 182050.0 68660.0 183395.0 ;
      RECT  67955.0 184740.0 68660.0 183395.0 ;
      RECT  67955.0 184740.0 68660.0 186085.0 ;
      RECT  67955.0 187430.0 68660.0 186085.0 ;
      RECT  67955.0 187430.0 68660.0 188775.0 ;
      RECT  67955.0 190120.0 68660.0 188775.0 ;
      RECT  67955.0 190120.0 68660.0 191465.0 ;
      RECT  67955.0 192810.0 68660.0 191465.0 ;
      RECT  67955.0 192810.0 68660.0 194155.0 ;
      RECT  67955.0 195500.0 68660.0 194155.0 ;
      RECT  67955.0 195500.0 68660.0 196845.0 ;
      RECT  67955.0 198190.0 68660.0 196845.0 ;
      RECT  67955.0 198190.0 68660.0 199535.0 ;
      RECT  67955.0 200880.0 68660.0 199535.0 ;
      RECT  67955.0 200880.0 68660.0 202225.0 ;
      RECT  67955.0 203570.0 68660.0 202225.0 ;
      RECT  67955.0 203570.0 68660.0 204915.0 ;
      RECT  67955.0 206260.0 68660.0 204915.0 ;
      RECT  68660.0 34100.0 69365.0 35445.0 ;
      RECT  68660.0 36790.0 69365.0 35445.0 ;
      RECT  68660.0 36790.0 69365.0 38135.0 ;
      RECT  68660.0 39480.0 69365.0 38135.0 ;
      RECT  68660.0 39480.0 69365.0 40825.0 ;
      RECT  68660.0 42170.0 69365.0 40825.0 ;
      RECT  68660.0 42170.0 69365.0 43515.0 ;
      RECT  68660.0 44860.0 69365.0 43515.0 ;
      RECT  68660.0 44860.0 69365.0 46205.0 ;
      RECT  68660.0 47550.0 69365.0 46205.0 ;
      RECT  68660.0 47550.0 69365.0 48895.0 ;
      RECT  68660.0 50240.0 69365.0 48895.0 ;
      RECT  68660.0 50240.0 69365.0 51585.0 ;
      RECT  68660.0 52930.0 69365.0 51585.0 ;
      RECT  68660.0 52930.0 69365.0 54275.0 ;
      RECT  68660.0 55620.0 69365.0 54275.0 ;
      RECT  68660.0 55620.0 69365.0 56965.0 ;
      RECT  68660.0 58310.0 69365.0 56965.0 ;
      RECT  68660.0 58310.0 69365.0 59655.0 ;
      RECT  68660.0 61000.0 69365.0 59655.0 ;
      RECT  68660.0 61000.0 69365.0 62345.0 ;
      RECT  68660.0 63690.0 69365.0 62345.0 ;
      RECT  68660.0 63690.0 69365.0 65035.0 ;
      RECT  68660.0 66380.0 69365.0 65035.0 ;
      RECT  68660.0 66380.0 69365.0 67725.0 ;
      RECT  68660.0 69070.0 69365.0 67725.0 ;
      RECT  68660.0 69070.0 69365.0 70415.0 ;
      RECT  68660.0 71760.0 69365.0 70415.0 ;
      RECT  68660.0 71760.0 69365.0 73105.0 ;
      RECT  68660.0 74450.0 69365.0 73105.0 ;
      RECT  68660.0 74450.0 69365.0 75795.0 ;
      RECT  68660.0 77140.0 69365.0 75795.0 ;
      RECT  68660.0 77140.0 69365.0 78485.0 ;
      RECT  68660.0 79830.0 69365.0 78485.0 ;
      RECT  68660.0 79830.0 69365.0 81175.0 ;
      RECT  68660.0 82520.0 69365.0 81175.0 ;
      RECT  68660.0 82520.0 69365.0 83865.0 ;
      RECT  68660.0 85210.0 69365.0 83865.0 ;
      RECT  68660.0 85210.0 69365.0 86555.0 ;
      RECT  68660.0 87900.0 69365.0 86555.0 ;
      RECT  68660.0 87900.0 69365.0 89245.0 ;
      RECT  68660.0 90590.0 69365.0 89245.0 ;
      RECT  68660.0 90590.0 69365.0 91935.0 ;
      RECT  68660.0 93280.0 69365.0 91935.0 ;
      RECT  68660.0 93280.0 69365.0 94625.0 ;
      RECT  68660.0 95970.0 69365.0 94625.0 ;
      RECT  68660.0 95970.0 69365.0 97315.0 ;
      RECT  68660.0 98660.0 69365.0 97315.0 ;
      RECT  68660.0 98660.0 69365.0 100005.0 ;
      RECT  68660.0 101350.0 69365.0 100005.0 ;
      RECT  68660.0 101350.0 69365.0 102695.0 ;
      RECT  68660.0 104040.0 69365.0 102695.0 ;
      RECT  68660.0 104040.0 69365.0 105385.0 ;
      RECT  68660.0 106730.0 69365.0 105385.0 ;
      RECT  68660.0 106730.0 69365.0 108075.0 ;
      RECT  68660.0 109420.0 69365.0 108075.0 ;
      RECT  68660.0 109420.0 69365.0 110765.0 ;
      RECT  68660.0 112110.0 69365.0 110765.0 ;
      RECT  68660.0 112110.0 69365.0 113455.0 ;
      RECT  68660.0 114800.0 69365.0 113455.0 ;
      RECT  68660.0 114800.0 69365.0 116145.0 ;
      RECT  68660.0 117490.0 69365.0 116145.0 ;
      RECT  68660.0 117490.0 69365.0 118835.0 ;
      RECT  68660.0 120180.0 69365.0 118835.0 ;
      RECT  68660.0 120180.0 69365.0 121525.0 ;
      RECT  68660.0 122870.0 69365.0 121525.0 ;
      RECT  68660.0 122870.0 69365.0 124215.0 ;
      RECT  68660.0 125560.0 69365.0 124215.0 ;
      RECT  68660.0 125560.0 69365.0 126905.0 ;
      RECT  68660.0 128250.0 69365.0 126905.0 ;
      RECT  68660.0 128250.0 69365.0 129595.0 ;
      RECT  68660.0 130940.0 69365.0 129595.0 ;
      RECT  68660.0 130940.0 69365.0 132285.0 ;
      RECT  68660.0 133630.0 69365.0 132285.0 ;
      RECT  68660.0 133630.0 69365.0 134975.0 ;
      RECT  68660.0 136320.0 69365.0 134975.0 ;
      RECT  68660.0 136320.0 69365.0 137665.0 ;
      RECT  68660.0 139010.0 69365.0 137665.0 ;
      RECT  68660.0 139010.0 69365.0 140355.0 ;
      RECT  68660.0 141700.0 69365.0 140355.0 ;
      RECT  68660.0 141700.0 69365.0 143045.0 ;
      RECT  68660.0 144390.0 69365.0 143045.0 ;
      RECT  68660.0 144390.0 69365.0 145735.0 ;
      RECT  68660.0 147080.0 69365.0 145735.0 ;
      RECT  68660.0 147080.0 69365.0 148425.0 ;
      RECT  68660.0 149770.0 69365.0 148425.0 ;
      RECT  68660.0 149770.0 69365.0 151115.0 ;
      RECT  68660.0 152460.0 69365.0 151115.0 ;
      RECT  68660.0 152460.0 69365.0 153805.0 ;
      RECT  68660.0 155150.0 69365.0 153805.0 ;
      RECT  68660.0 155150.0 69365.0 156495.0 ;
      RECT  68660.0 157840.0 69365.0 156495.0 ;
      RECT  68660.0 157840.0 69365.0 159185.0 ;
      RECT  68660.0 160530.0 69365.0 159185.0 ;
      RECT  68660.0 160530.0 69365.0 161875.0 ;
      RECT  68660.0 163220.0 69365.0 161875.0 ;
      RECT  68660.0 163220.0 69365.0 164565.0 ;
      RECT  68660.0 165910.0 69365.0 164565.0 ;
      RECT  68660.0 165910.0 69365.0 167255.0 ;
      RECT  68660.0 168600.0 69365.0 167255.0 ;
      RECT  68660.0 168600.0 69365.0 169945.0 ;
      RECT  68660.0 171290.0 69365.0 169945.0 ;
      RECT  68660.0 171290.0 69365.0 172635.0 ;
      RECT  68660.0 173980.0 69365.0 172635.0 ;
      RECT  68660.0 173980.0 69365.0 175325.0 ;
      RECT  68660.0 176670.0 69365.0 175325.0 ;
      RECT  68660.0 176670.0 69365.0 178015.0 ;
      RECT  68660.0 179360.0 69365.0 178015.0 ;
      RECT  68660.0 179360.0 69365.0 180705.0 ;
      RECT  68660.0 182050.0 69365.0 180705.0 ;
      RECT  68660.0 182050.0 69365.0 183395.0 ;
      RECT  68660.0 184740.0 69365.0 183395.0 ;
      RECT  68660.0 184740.0 69365.0 186085.0 ;
      RECT  68660.0 187430.0 69365.0 186085.0 ;
      RECT  68660.0 187430.0 69365.0 188775.0 ;
      RECT  68660.0 190120.0 69365.0 188775.0 ;
      RECT  68660.0 190120.0 69365.0 191465.0 ;
      RECT  68660.0 192810.0 69365.0 191465.0 ;
      RECT  68660.0 192810.0 69365.0 194155.0 ;
      RECT  68660.0 195500.0 69365.0 194155.0 ;
      RECT  68660.0 195500.0 69365.0 196845.0 ;
      RECT  68660.0 198190.0 69365.0 196845.0 ;
      RECT  68660.0 198190.0 69365.0 199535.0 ;
      RECT  68660.0 200880.0 69365.0 199535.0 ;
      RECT  68660.0 200880.0 69365.0 202225.0 ;
      RECT  68660.0 203570.0 69365.0 202225.0 ;
      RECT  68660.0 203570.0 69365.0 204915.0 ;
      RECT  68660.0 206260.0 69365.0 204915.0 ;
      RECT  69365.0 34100.0 70070.0 35445.0 ;
      RECT  69365.0 36790.0 70070.0 35445.0 ;
      RECT  69365.0 36790.0 70070.0 38135.0 ;
      RECT  69365.0 39480.0 70070.0 38135.0 ;
      RECT  69365.0 39480.0 70070.0 40825.0 ;
      RECT  69365.0 42170.0 70070.0 40825.0 ;
      RECT  69365.0 42170.0 70070.0 43515.0 ;
      RECT  69365.0 44860.0 70070.0 43515.0 ;
      RECT  69365.0 44860.0 70070.0 46205.0 ;
      RECT  69365.0 47550.0 70070.0 46205.0 ;
      RECT  69365.0 47550.0 70070.0 48895.0 ;
      RECT  69365.0 50240.0 70070.0 48895.0 ;
      RECT  69365.0 50240.0 70070.0 51585.0 ;
      RECT  69365.0 52930.0 70070.0 51585.0 ;
      RECT  69365.0 52930.0 70070.0 54275.0 ;
      RECT  69365.0 55620.0 70070.0 54275.0 ;
      RECT  69365.0 55620.0 70070.0 56965.0 ;
      RECT  69365.0 58310.0 70070.0 56965.0 ;
      RECT  69365.0 58310.0 70070.0 59655.0 ;
      RECT  69365.0 61000.0 70070.0 59655.0 ;
      RECT  69365.0 61000.0 70070.0 62345.0 ;
      RECT  69365.0 63690.0 70070.0 62345.0 ;
      RECT  69365.0 63690.0 70070.0 65035.0 ;
      RECT  69365.0 66380.0 70070.0 65035.0 ;
      RECT  69365.0 66380.0 70070.0 67725.0 ;
      RECT  69365.0 69070.0 70070.0 67725.0 ;
      RECT  69365.0 69070.0 70070.0 70415.0 ;
      RECT  69365.0 71760.0 70070.0 70415.0 ;
      RECT  69365.0 71760.0 70070.0 73105.0 ;
      RECT  69365.0 74450.0 70070.0 73105.0 ;
      RECT  69365.0 74450.0 70070.0 75795.0 ;
      RECT  69365.0 77140.0 70070.0 75795.0 ;
      RECT  69365.0 77140.0 70070.0 78485.0 ;
      RECT  69365.0 79830.0 70070.0 78485.0 ;
      RECT  69365.0 79830.0 70070.0 81175.0 ;
      RECT  69365.0 82520.0 70070.0 81175.0 ;
      RECT  69365.0 82520.0 70070.0 83865.0 ;
      RECT  69365.0 85210.0 70070.0 83865.0 ;
      RECT  69365.0 85210.0 70070.0 86555.0 ;
      RECT  69365.0 87900.0 70070.0 86555.0 ;
      RECT  69365.0 87900.0 70070.0 89245.0 ;
      RECT  69365.0 90590.0 70070.0 89245.0 ;
      RECT  69365.0 90590.0 70070.0 91935.0 ;
      RECT  69365.0 93280.0 70070.0 91935.0 ;
      RECT  69365.0 93280.0 70070.0 94625.0 ;
      RECT  69365.0 95970.0 70070.0 94625.0 ;
      RECT  69365.0 95970.0 70070.0 97315.0 ;
      RECT  69365.0 98660.0 70070.0 97315.0 ;
      RECT  69365.0 98660.0 70070.0 100005.0 ;
      RECT  69365.0 101350.0 70070.0 100005.0 ;
      RECT  69365.0 101350.0 70070.0 102695.0 ;
      RECT  69365.0 104040.0 70070.0 102695.0 ;
      RECT  69365.0 104040.0 70070.0 105385.0 ;
      RECT  69365.0 106730.0 70070.0 105385.0 ;
      RECT  69365.0 106730.0 70070.0 108075.0 ;
      RECT  69365.0 109420.0 70070.0 108075.0 ;
      RECT  69365.0 109420.0 70070.0 110765.0 ;
      RECT  69365.0 112110.0 70070.0 110765.0 ;
      RECT  69365.0 112110.0 70070.0 113455.0 ;
      RECT  69365.0 114800.0 70070.0 113455.0 ;
      RECT  69365.0 114800.0 70070.0 116145.0 ;
      RECT  69365.0 117490.0 70070.0 116145.0 ;
      RECT  69365.0 117490.0 70070.0 118835.0 ;
      RECT  69365.0 120180.0 70070.0 118835.0 ;
      RECT  69365.0 120180.0 70070.0 121525.0 ;
      RECT  69365.0 122870.0 70070.0 121525.0 ;
      RECT  69365.0 122870.0 70070.0 124215.0 ;
      RECT  69365.0 125560.0 70070.0 124215.0 ;
      RECT  69365.0 125560.0 70070.0 126905.0 ;
      RECT  69365.0 128250.0 70070.0 126905.0 ;
      RECT  69365.0 128250.0 70070.0 129595.0 ;
      RECT  69365.0 130940.0 70070.0 129595.0 ;
      RECT  69365.0 130940.0 70070.0 132285.0 ;
      RECT  69365.0 133630.0 70070.0 132285.0 ;
      RECT  69365.0 133630.0 70070.0 134975.0 ;
      RECT  69365.0 136320.0 70070.0 134975.0 ;
      RECT  69365.0 136320.0 70070.0 137665.0 ;
      RECT  69365.0 139010.0 70070.0 137665.0 ;
      RECT  69365.0 139010.0 70070.0 140355.0 ;
      RECT  69365.0 141700.0 70070.0 140355.0 ;
      RECT  69365.0 141700.0 70070.0 143045.0 ;
      RECT  69365.0 144390.0 70070.0 143045.0 ;
      RECT  69365.0 144390.0 70070.0 145735.0 ;
      RECT  69365.0 147080.0 70070.0 145735.0 ;
      RECT  69365.0 147080.0 70070.0 148425.0 ;
      RECT  69365.0 149770.0 70070.0 148425.0 ;
      RECT  69365.0 149770.0 70070.0 151115.0 ;
      RECT  69365.0 152460.0 70070.0 151115.0 ;
      RECT  69365.0 152460.0 70070.0 153805.0 ;
      RECT  69365.0 155150.0 70070.0 153805.0 ;
      RECT  69365.0 155150.0 70070.0 156495.0 ;
      RECT  69365.0 157840.0 70070.0 156495.0 ;
      RECT  69365.0 157840.0 70070.0 159185.0 ;
      RECT  69365.0 160530.0 70070.0 159185.0 ;
      RECT  69365.0 160530.0 70070.0 161875.0 ;
      RECT  69365.0 163220.0 70070.0 161875.0 ;
      RECT  69365.0 163220.0 70070.0 164565.0 ;
      RECT  69365.0 165910.0 70070.0 164565.0 ;
      RECT  69365.0 165910.0 70070.0 167255.0 ;
      RECT  69365.0 168600.0 70070.0 167255.0 ;
      RECT  69365.0 168600.0 70070.0 169945.0 ;
      RECT  69365.0 171290.0 70070.0 169945.0 ;
      RECT  69365.0 171290.0 70070.0 172635.0 ;
      RECT  69365.0 173980.0 70070.0 172635.0 ;
      RECT  69365.0 173980.0 70070.0 175325.0 ;
      RECT  69365.0 176670.0 70070.0 175325.0 ;
      RECT  69365.0 176670.0 70070.0 178015.0 ;
      RECT  69365.0 179360.0 70070.0 178015.0 ;
      RECT  69365.0 179360.0 70070.0 180705.0 ;
      RECT  69365.0 182050.0 70070.0 180705.0 ;
      RECT  69365.0 182050.0 70070.0 183395.0 ;
      RECT  69365.0 184740.0 70070.0 183395.0 ;
      RECT  69365.0 184740.0 70070.0 186085.0 ;
      RECT  69365.0 187430.0 70070.0 186085.0 ;
      RECT  69365.0 187430.0 70070.0 188775.0 ;
      RECT  69365.0 190120.0 70070.0 188775.0 ;
      RECT  69365.0 190120.0 70070.0 191465.0 ;
      RECT  69365.0 192810.0 70070.0 191465.0 ;
      RECT  69365.0 192810.0 70070.0 194155.0 ;
      RECT  69365.0 195500.0 70070.0 194155.0 ;
      RECT  69365.0 195500.0 70070.0 196845.0 ;
      RECT  69365.0 198190.0 70070.0 196845.0 ;
      RECT  69365.0 198190.0 70070.0 199535.0 ;
      RECT  69365.0 200880.0 70070.0 199535.0 ;
      RECT  69365.0 200880.0 70070.0 202225.0 ;
      RECT  69365.0 203570.0 70070.0 202225.0 ;
      RECT  69365.0 203570.0 70070.0 204915.0 ;
      RECT  69365.0 206260.0 70070.0 204915.0 ;
      RECT  70070.0 34100.0 70775.0 35445.0 ;
      RECT  70070.0 36790.0 70775.0 35445.0 ;
      RECT  70070.0 36790.0 70775.0 38135.0 ;
      RECT  70070.0 39480.0 70775.0 38135.0 ;
      RECT  70070.0 39480.0 70775.0 40825.0 ;
      RECT  70070.0 42170.0 70775.0 40825.0 ;
      RECT  70070.0 42170.0 70775.0 43515.0 ;
      RECT  70070.0 44860.0 70775.0 43515.0 ;
      RECT  70070.0 44860.0 70775.0 46205.0 ;
      RECT  70070.0 47550.0 70775.0 46205.0 ;
      RECT  70070.0 47550.0 70775.0 48895.0 ;
      RECT  70070.0 50240.0 70775.0 48895.0 ;
      RECT  70070.0 50240.0 70775.0 51585.0 ;
      RECT  70070.0 52930.0 70775.0 51585.0 ;
      RECT  70070.0 52930.0 70775.0 54275.0 ;
      RECT  70070.0 55620.0 70775.0 54275.0 ;
      RECT  70070.0 55620.0 70775.0 56965.0 ;
      RECT  70070.0 58310.0 70775.0 56965.0 ;
      RECT  70070.0 58310.0 70775.0 59655.0 ;
      RECT  70070.0 61000.0 70775.0 59655.0 ;
      RECT  70070.0 61000.0 70775.0 62345.0 ;
      RECT  70070.0 63690.0 70775.0 62345.0 ;
      RECT  70070.0 63690.0 70775.0 65035.0 ;
      RECT  70070.0 66380.0 70775.0 65035.0 ;
      RECT  70070.0 66380.0 70775.0 67725.0 ;
      RECT  70070.0 69070.0 70775.0 67725.0 ;
      RECT  70070.0 69070.0 70775.0 70415.0 ;
      RECT  70070.0 71760.0 70775.0 70415.0 ;
      RECT  70070.0 71760.0 70775.0 73105.0 ;
      RECT  70070.0 74450.0 70775.0 73105.0 ;
      RECT  70070.0 74450.0 70775.0 75795.0 ;
      RECT  70070.0 77140.0 70775.0 75795.0 ;
      RECT  70070.0 77140.0 70775.0 78485.0 ;
      RECT  70070.0 79830.0 70775.0 78485.0 ;
      RECT  70070.0 79830.0 70775.0 81175.0 ;
      RECT  70070.0 82520.0 70775.0 81175.0 ;
      RECT  70070.0 82520.0 70775.0 83865.0 ;
      RECT  70070.0 85210.0 70775.0 83865.0 ;
      RECT  70070.0 85210.0 70775.0 86555.0 ;
      RECT  70070.0 87900.0 70775.0 86555.0 ;
      RECT  70070.0 87900.0 70775.0 89245.0 ;
      RECT  70070.0 90590.0 70775.0 89245.0 ;
      RECT  70070.0 90590.0 70775.0 91935.0 ;
      RECT  70070.0 93280.0 70775.0 91935.0 ;
      RECT  70070.0 93280.0 70775.0 94625.0 ;
      RECT  70070.0 95970.0 70775.0 94625.0 ;
      RECT  70070.0 95970.0 70775.0 97315.0 ;
      RECT  70070.0 98660.0 70775.0 97315.0 ;
      RECT  70070.0 98660.0 70775.0 100005.0 ;
      RECT  70070.0 101350.0 70775.0 100005.0 ;
      RECT  70070.0 101350.0 70775.0 102695.0 ;
      RECT  70070.0 104040.0 70775.0 102695.0 ;
      RECT  70070.0 104040.0 70775.0 105385.0 ;
      RECT  70070.0 106730.0 70775.0 105385.0 ;
      RECT  70070.0 106730.0 70775.0 108075.0 ;
      RECT  70070.0 109420.0 70775.0 108075.0 ;
      RECT  70070.0 109420.0 70775.0 110765.0 ;
      RECT  70070.0 112110.0 70775.0 110765.0 ;
      RECT  70070.0 112110.0 70775.0 113455.0 ;
      RECT  70070.0 114800.0 70775.0 113455.0 ;
      RECT  70070.0 114800.0 70775.0 116145.0 ;
      RECT  70070.0 117490.0 70775.0 116145.0 ;
      RECT  70070.0 117490.0 70775.0 118835.0 ;
      RECT  70070.0 120180.0 70775.0 118835.0 ;
      RECT  70070.0 120180.0 70775.0 121525.0 ;
      RECT  70070.0 122870.0 70775.0 121525.0 ;
      RECT  70070.0 122870.0 70775.0 124215.0 ;
      RECT  70070.0 125560.0 70775.0 124215.0 ;
      RECT  70070.0 125560.0 70775.0 126905.0 ;
      RECT  70070.0 128250.0 70775.0 126905.0 ;
      RECT  70070.0 128250.0 70775.0 129595.0 ;
      RECT  70070.0 130940.0 70775.0 129595.0 ;
      RECT  70070.0 130940.0 70775.0 132285.0 ;
      RECT  70070.0 133630.0 70775.0 132285.0 ;
      RECT  70070.0 133630.0 70775.0 134975.0 ;
      RECT  70070.0 136320.0 70775.0 134975.0 ;
      RECT  70070.0 136320.0 70775.0 137665.0 ;
      RECT  70070.0 139010.0 70775.0 137665.0 ;
      RECT  70070.0 139010.0 70775.0 140355.0 ;
      RECT  70070.0 141700.0 70775.0 140355.0 ;
      RECT  70070.0 141700.0 70775.0 143045.0 ;
      RECT  70070.0 144390.0 70775.0 143045.0 ;
      RECT  70070.0 144390.0 70775.0 145735.0 ;
      RECT  70070.0 147080.0 70775.0 145735.0 ;
      RECT  70070.0 147080.0 70775.0 148425.0 ;
      RECT  70070.0 149770.0 70775.0 148425.0 ;
      RECT  70070.0 149770.0 70775.0 151115.0 ;
      RECT  70070.0 152460.0 70775.0 151115.0 ;
      RECT  70070.0 152460.0 70775.0 153805.0 ;
      RECT  70070.0 155150.0 70775.0 153805.0 ;
      RECT  70070.0 155150.0 70775.0 156495.0 ;
      RECT  70070.0 157840.0 70775.0 156495.0 ;
      RECT  70070.0 157840.0 70775.0 159185.0 ;
      RECT  70070.0 160530.0 70775.0 159185.0 ;
      RECT  70070.0 160530.0 70775.0 161875.0 ;
      RECT  70070.0 163220.0 70775.0 161875.0 ;
      RECT  70070.0 163220.0 70775.0 164565.0 ;
      RECT  70070.0 165910.0 70775.0 164565.0 ;
      RECT  70070.0 165910.0 70775.0 167255.0 ;
      RECT  70070.0 168600.0 70775.0 167255.0 ;
      RECT  70070.0 168600.0 70775.0 169945.0 ;
      RECT  70070.0 171290.0 70775.0 169945.0 ;
      RECT  70070.0 171290.0 70775.0 172635.0 ;
      RECT  70070.0 173980.0 70775.0 172635.0 ;
      RECT  70070.0 173980.0 70775.0 175325.0 ;
      RECT  70070.0 176670.0 70775.0 175325.0 ;
      RECT  70070.0 176670.0 70775.0 178015.0 ;
      RECT  70070.0 179360.0 70775.0 178015.0 ;
      RECT  70070.0 179360.0 70775.0 180705.0 ;
      RECT  70070.0 182050.0 70775.0 180705.0 ;
      RECT  70070.0 182050.0 70775.0 183395.0 ;
      RECT  70070.0 184740.0 70775.0 183395.0 ;
      RECT  70070.0 184740.0 70775.0 186085.0 ;
      RECT  70070.0 187430.0 70775.0 186085.0 ;
      RECT  70070.0 187430.0 70775.0 188775.0 ;
      RECT  70070.0 190120.0 70775.0 188775.0 ;
      RECT  70070.0 190120.0 70775.0 191465.0 ;
      RECT  70070.0 192810.0 70775.0 191465.0 ;
      RECT  70070.0 192810.0 70775.0 194155.0 ;
      RECT  70070.0 195500.0 70775.0 194155.0 ;
      RECT  70070.0 195500.0 70775.0 196845.0 ;
      RECT  70070.0 198190.0 70775.0 196845.0 ;
      RECT  70070.0 198190.0 70775.0 199535.0 ;
      RECT  70070.0 200880.0 70775.0 199535.0 ;
      RECT  70070.0 200880.0 70775.0 202225.0 ;
      RECT  70070.0 203570.0 70775.0 202225.0 ;
      RECT  70070.0 203570.0 70775.0 204915.0 ;
      RECT  70070.0 206260.0 70775.0 204915.0 ;
      RECT  70775.0 34100.0 71480.0 35445.0 ;
      RECT  70775.0 36790.0 71480.0 35445.0 ;
      RECT  70775.0 36790.0 71480.0 38135.0 ;
      RECT  70775.0 39480.0 71480.0 38135.0 ;
      RECT  70775.0 39480.0 71480.0 40825.0 ;
      RECT  70775.0 42170.0 71480.0 40825.0 ;
      RECT  70775.0 42170.0 71480.0 43515.0 ;
      RECT  70775.0 44860.0 71480.0 43515.0 ;
      RECT  70775.0 44860.0 71480.0 46205.0 ;
      RECT  70775.0 47550.0 71480.0 46205.0 ;
      RECT  70775.0 47550.0 71480.0 48895.0 ;
      RECT  70775.0 50240.0 71480.0 48895.0 ;
      RECT  70775.0 50240.0 71480.0 51585.0 ;
      RECT  70775.0 52930.0 71480.0 51585.0 ;
      RECT  70775.0 52930.0 71480.0 54275.0 ;
      RECT  70775.0 55620.0 71480.0 54275.0 ;
      RECT  70775.0 55620.0 71480.0 56965.0 ;
      RECT  70775.0 58310.0 71480.0 56965.0 ;
      RECT  70775.0 58310.0 71480.0 59655.0 ;
      RECT  70775.0 61000.0 71480.0 59655.0 ;
      RECT  70775.0 61000.0 71480.0 62345.0 ;
      RECT  70775.0 63690.0 71480.0 62345.0 ;
      RECT  70775.0 63690.0 71480.0 65035.0 ;
      RECT  70775.0 66380.0 71480.0 65035.0 ;
      RECT  70775.0 66380.0 71480.0 67725.0 ;
      RECT  70775.0 69070.0 71480.0 67725.0 ;
      RECT  70775.0 69070.0 71480.0 70415.0 ;
      RECT  70775.0 71760.0 71480.0 70415.0 ;
      RECT  70775.0 71760.0 71480.0 73105.0 ;
      RECT  70775.0 74450.0 71480.0 73105.0 ;
      RECT  70775.0 74450.0 71480.0 75795.0 ;
      RECT  70775.0 77140.0 71480.0 75795.0 ;
      RECT  70775.0 77140.0 71480.0 78485.0 ;
      RECT  70775.0 79830.0 71480.0 78485.0 ;
      RECT  70775.0 79830.0 71480.0 81175.0 ;
      RECT  70775.0 82520.0 71480.0 81175.0 ;
      RECT  70775.0 82520.0 71480.0 83865.0 ;
      RECT  70775.0 85210.0 71480.0 83865.0 ;
      RECT  70775.0 85210.0 71480.0 86555.0 ;
      RECT  70775.0 87900.0 71480.0 86555.0 ;
      RECT  70775.0 87900.0 71480.0 89245.0 ;
      RECT  70775.0 90590.0 71480.0 89245.0 ;
      RECT  70775.0 90590.0 71480.0 91935.0 ;
      RECT  70775.0 93280.0 71480.0 91935.0 ;
      RECT  70775.0 93280.0 71480.0 94625.0 ;
      RECT  70775.0 95970.0 71480.0 94625.0 ;
      RECT  70775.0 95970.0 71480.0 97315.0 ;
      RECT  70775.0 98660.0 71480.0 97315.0 ;
      RECT  70775.0 98660.0 71480.0 100005.0 ;
      RECT  70775.0 101350.0 71480.0 100005.0 ;
      RECT  70775.0 101350.0 71480.0 102695.0 ;
      RECT  70775.0 104040.0 71480.0 102695.0 ;
      RECT  70775.0 104040.0 71480.0 105385.0 ;
      RECT  70775.0 106730.0 71480.0 105385.0 ;
      RECT  70775.0 106730.0 71480.0 108075.0 ;
      RECT  70775.0 109420.0 71480.0 108075.0 ;
      RECT  70775.0 109420.0 71480.0 110765.0 ;
      RECT  70775.0 112110.0 71480.0 110765.0 ;
      RECT  70775.0 112110.0 71480.0 113455.0 ;
      RECT  70775.0 114800.0 71480.0 113455.0 ;
      RECT  70775.0 114800.0 71480.0 116145.0 ;
      RECT  70775.0 117490.0 71480.0 116145.0 ;
      RECT  70775.0 117490.0 71480.0 118835.0 ;
      RECT  70775.0 120180.0 71480.0 118835.0 ;
      RECT  70775.0 120180.0 71480.0 121525.0 ;
      RECT  70775.0 122870.0 71480.0 121525.0 ;
      RECT  70775.0 122870.0 71480.0 124215.0 ;
      RECT  70775.0 125560.0 71480.0 124215.0 ;
      RECT  70775.0 125560.0 71480.0 126905.0 ;
      RECT  70775.0 128250.0 71480.0 126905.0 ;
      RECT  70775.0 128250.0 71480.0 129595.0 ;
      RECT  70775.0 130940.0 71480.0 129595.0 ;
      RECT  70775.0 130940.0 71480.0 132285.0 ;
      RECT  70775.0 133630.0 71480.0 132285.0 ;
      RECT  70775.0 133630.0 71480.0 134975.0 ;
      RECT  70775.0 136320.0 71480.0 134975.0 ;
      RECT  70775.0 136320.0 71480.0 137665.0 ;
      RECT  70775.0 139010.0 71480.0 137665.0 ;
      RECT  70775.0 139010.0 71480.0 140355.0 ;
      RECT  70775.0 141700.0 71480.0 140355.0 ;
      RECT  70775.0 141700.0 71480.0 143045.0 ;
      RECT  70775.0 144390.0 71480.0 143045.0 ;
      RECT  70775.0 144390.0 71480.0 145735.0 ;
      RECT  70775.0 147080.0 71480.0 145735.0 ;
      RECT  70775.0 147080.0 71480.0 148425.0 ;
      RECT  70775.0 149770.0 71480.0 148425.0 ;
      RECT  70775.0 149770.0 71480.0 151115.0 ;
      RECT  70775.0 152460.0 71480.0 151115.0 ;
      RECT  70775.0 152460.0 71480.0 153805.0 ;
      RECT  70775.0 155150.0 71480.0 153805.0 ;
      RECT  70775.0 155150.0 71480.0 156495.0 ;
      RECT  70775.0 157840.0 71480.0 156495.0 ;
      RECT  70775.0 157840.0 71480.0 159185.0 ;
      RECT  70775.0 160530.0 71480.0 159185.0 ;
      RECT  70775.0 160530.0 71480.0 161875.0 ;
      RECT  70775.0 163220.0 71480.0 161875.0 ;
      RECT  70775.0 163220.0 71480.0 164565.0 ;
      RECT  70775.0 165910.0 71480.0 164565.0 ;
      RECT  70775.0 165910.0 71480.0 167255.0 ;
      RECT  70775.0 168600.0 71480.0 167255.0 ;
      RECT  70775.0 168600.0 71480.0 169945.0 ;
      RECT  70775.0 171290.0 71480.0 169945.0 ;
      RECT  70775.0 171290.0 71480.0 172635.0 ;
      RECT  70775.0 173980.0 71480.0 172635.0 ;
      RECT  70775.0 173980.0 71480.0 175325.0 ;
      RECT  70775.0 176670.0 71480.0 175325.0 ;
      RECT  70775.0 176670.0 71480.0 178015.0 ;
      RECT  70775.0 179360.0 71480.0 178015.0 ;
      RECT  70775.0 179360.0 71480.0 180705.0 ;
      RECT  70775.0 182050.0 71480.0 180705.0 ;
      RECT  70775.0 182050.0 71480.0 183395.0 ;
      RECT  70775.0 184740.0 71480.0 183395.0 ;
      RECT  70775.0 184740.0 71480.0 186085.0 ;
      RECT  70775.0 187430.0 71480.0 186085.0 ;
      RECT  70775.0 187430.0 71480.0 188775.0 ;
      RECT  70775.0 190120.0 71480.0 188775.0 ;
      RECT  70775.0 190120.0 71480.0 191465.0 ;
      RECT  70775.0 192810.0 71480.0 191465.0 ;
      RECT  70775.0 192810.0 71480.0 194155.0 ;
      RECT  70775.0 195500.0 71480.0 194155.0 ;
      RECT  70775.0 195500.0 71480.0 196845.0 ;
      RECT  70775.0 198190.0 71480.0 196845.0 ;
      RECT  70775.0 198190.0 71480.0 199535.0 ;
      RECT  70775.0 200880.0 71480.0 199535.0 ;
      RECT  70775.0 200880.0 71480.0 202225.0 ;
      RECT  70775.0 203570.0 71480.0 202225.0 ;
      RECT  70775.0 203570.0 71480.0 204915.0 ;
      RECT  70775.0 206260.0 71480.0 204915.0 ;
      RECT  71480.0 34100.0 72185.0 35445.0 ;
      RECT  71480.0 36790.0 72185.0 35445.0 ;
      RECT  71480.0 36790.0 72185.0 38135.0 ;
      RECT  71480.0 39480.0 72185.0 38135.0 ;
      RECT  71480.0 39480.0 72185.0 40825.0 ;
      RECT  71480.0 42170.0 72185.0 40825.0 ;
      RECT  71480.0 42170.0 72185.0 43515.0 ;
      RECT  71480.0 44860.0 72185.0 43515.0 ;
      RECT  71480.0 44860.0 72185.0 46205.0 ;
      RECT  71480.0 47550.0 72185.0 46205.0 ;
      RECT  71480.0 47550.0 72185.0 48895.0 ;
      RECT  71480.0 50240.0 72185.0 48895.0 ;
      RECT  71480.0 50240.0 72185.0 51585.0 ;
      RECT  71480.0 52930.0 72185.0 51585.0 ;
      RECT  71480.0 52930.0 72185.0 54275.0 ;
      RECT  71480.0 55620.0 72185.0 54275.0 ;
      RECT  71480.0 55620.0 72185.0 56965.0 ;
      RECT  71480.0 58310.0 72185.0 56965.0 ;
      RECT  71480.0 58310.0 72185.0 59655.0 ;
      RECT  71480.0 61000.0 72185.0 59655.0 ;
      RECT  71480.0 61000.0 72185.0 62345.0 ;
      RECT  71480.0 63690.0 72185.0 62345.0 ;
      RECT  71480.0 63690.0 72185.0 65035.0 ;
      RECT  71480.0 66380.0 72185.0 65035.0 ;
      RECT  71480.0 66380.0 72185.0 67725.0 ;
      RECT  71480.0 69070.0 72185.0 67725.0 ;
      RECT  71480.0 69070.0 72185.0 70415.0 ;
      RECT  71480.0 71760.0 72185.0 70415.0 ;
      RECT  71480.0 71760.0 72185.0 73105.0 ;
      RECT  71480.0 74450.0 72185.0 73105.0 ;
      RECT  71480.0 74450.0 72185.0 75795.0 ;
      RECT  71480.0 77140.0 72185.0 75795.0 ;
      RECT  71480.0 77140.0 72185.0 78485.0 ;
      RECT  71480.0 79830.0 72185.0 78485.0 ;
      RECT  71480.0 79830.0 72185.0 81175.0 ;
      RECT  71480.0 82520.0 72185.0 81175.0 ;
      RECT  71480.0 82520.0 72185.0 83865.0 ;
      RECT  71480.0 85210.0 72185.0 83865.0 ;
      RECT  71480.0 85210.0 72185.0 86555.0 ;
      RECT  71480.0 87900.0 72185.0 86555.0 ;
      RECT  71480.0 87900.0 72185.0 89245.0 ;
      RECT  71480.0 90590.0 72185.0 89245.0 ;
      RECT  71480.0 90590.0 72185.0 91935.0 ;
      RECT  71480.0 93280.0 72185.0 91935.0 ;
      RECT  71480.0 93280.0 72185.0 94625.0 ;
      RECT  71480.0 95970.0 72185.0 94625.0 ;
      RECT  71480.0 95970.0 72185.0 97315.0 ;
      RECT  71480.0 98660.0 72185.0 97315.0 ;
      RECT  71480.0 98660.0 72185.0 100005.0 ;
      RECT  71480.0 101350.0 72185.0 100005.0 ;
      RECT  71480.0 101350.0 72185.0 102695.0 ;
      RECT  71480.0 104040.0 72185.0 102695.0 ;
      RECT  71480.0 104040.0 72185.0 105385.0 ;
      RECT  71480.0 106730.0 72185.0 105385.0 ;
      RECT  71480.0 106730.0 72185.0 108075.0 ;
      RECT  71480.0 109420.0 72185.0 108075.0 ;
      RECT  71480.0 109420.0 72185.0 110765.0 ;
      RECT  71480.0 112110.0 72185.0 110765.0 ;
      RECT  71480.0 112110.0 72185.0 113455.0 ;
      RECT  71480.0 114800.0 72185.0 113455.0 ;
      RECT  71480.0 114800.0 72185.0 116145.0 ;
      RECT  71480.0 117490.0 72185.0 116145.0 ;
      RECT  71480.0 117490.0 72185.0 118835.0 ;
      RECT  71480.0 120180.0 72185.0 118835.0 ;
      RECT  71480.0 120180.0 72185.0 121525.0 ;
      RECT  71480.0 122870.0 72185.0 121525.0 ;
      RECT  71480.0 122870.0 72185.0 124215.0 ;
      RECT  71480.0 125560.0 72185.0 124215.0 ;
      RECT  71480.0 125560.0 72185.0 126905.0 ;
      RECT  71480.0 128250.0 72185.0 126905.0 ;
      RECT  71480.0 128250.0 72185.0 129595.0 ;
      RECT  71480.0 130940.0 72185.0 129595.0 ;
      RECT  71480.0 130940.0 72185.0 132285.0 ;
      RECT  71480.0 133630.0 72185.0 132285.0 ;
      RECT  71480.0 133630.0 72185.0 134975.0 ;
      RECT  71480.0 136320.0 72185.0 134975.0 ;
      RECT  71480.0 136320.0 72185.0 137665.0 ;
      RECT  71480.0 139010.0 72185.0 137665.0 ;
      RECT  71480.0 139010.0 72185.0 140355.0 ;
      RECT  71480.0 141700.0 72185.0 140355.0 ;
      RECT  71480.0 141700.0 72185.0 143045.0 ;
      RECT  71480.0 144390.0 72185.0 143045.0 ;
      RECT  71480.0 144390.0 72185.0 145735.0 ;
      RECT  71480.0 147080.0 72185.0 145735.0 ;
      RECT  71480.0 147080.0 72185.0 148425.0 ;
      RECT  71480.0 149770.0 72185.0 148425.0 ;
      RECT  71480.0 149770.0 72185.0 151115.0 ;
      RECT  71480.0 152460.0 72185.0 151115.0 ;
      RECT  71480.0 152460.0 72185.0 153805.0 ;
      RECT  71480.0 155150.0 72185.0 153805.0 ;
      RECT  71480.0 155150.0 72185.0 156495.0 ;
      RECT  71480.0 157840.0 72185.0 156495.0 ;
      RECT  71480.0 157840.0 72185.0 159185.0 ;
      RECT  71480.0 160530.0 72185.0 159185.0 ;
      RECT  71480.0 160530.0 72185.0 161875.0 ;
      RECT  71480.0 163220.0 72185.0 161875.0 ;
      RECT  71480.0 163220.0 72185.0 164565.0 ;
      RECT  71480.0 165910.0 72185.0 164565.0 ;
      RECT  71480.0 165910.0 72185.0 167255.0 ;
      RECT  71480.0 168600.0 72185.0 167255.0 ;
      RECT  71480.0 168600.0 72185.0 169945.0 ;
      RECT  71480.0 171290.0 72185.0 169945.0 ;
      RECT  71480.0 171290.0 72185.0 172635.0 ;
      RECT  71480.0 173980.0 72185.0 172635.0 ;
      RECT  71480.0 173980.0 72185.0 175325.0 ;
      RECT  71480.0 176670.0 72185.0 175325.0 ;
      RECT  71480.0 176670.0 72185.0 178015.0 ;
      RECT  71480.0 179360.0 72185.0 178015.0 ;
      RECT  71480.0 179360.0 72185.0 180705.0 ;
      RECT  71480.0 182050.0 72185.0 180705.0 ;
      RECT  71480.0 182050.0 72185.0 183395.0 ;
      RECT  71480.0 184740.0 72185.0 183395.0 ;
      RECT  71480.0 184740.0 72185.0 186085.0 ;
      RECT  71480.0 187430.0 72185.0 186085.0 ;
      RECT  71480.0 187430.0 72185.0 188775.0 ;
      RECT  71480.0 190120.0 72185.0 188775.0 ;
      RECT  71480.0 190120.0 72185.0 191465.0 ;
      RECT  71480.0 192810.0 72185.0 191465.0 ;
      RECT  71480.0 192810.0 72185.0 194155.0 ;
      RECT  71480.0 195500.0 72185.0 194155.0 ;
      RECT  71480.0 195500.0 72185.0 196845.0 ;
      RECT  71480.0 198190.0 72185.0 196845.0 ;
      RECT  71480.0 198190.0 72185.0 199535.0 ;
      RECT  71480.0 200880.0 72185.0 199535.0 ;
      RECT  71480.0 200880.0 72185.0 202225.0 ;
      RECT  71480.0 203570.0 72185.0 202225.0 ;
      RECT  71480.0 203570.0 72185.0 204915.0 ;
      RECT  71480.0 206260.0 72185.0 204915.0 ;
      RECT  72185.0 34100.0 72890.0 35445.0 ;
      RECT  72185.0 36790.0 72890.0 35445.0 ;
      RECT  72185.0 36790.0 72890.0 38135.0 ;
      RECT  72185.0 39480.0 72890.0 38135.0 ;
      RECT  72185.0 39480.0 72890.0 40825.0 ;
      RECT  72185.0 42170.0 72890.0 40825.0 ;
      RECT  72185.0 42170.0 72890.0 43515.0 ;
      RECT  72185.0 44860.0 72890.0 43515.0 ;
      RECT  72185.0 44860.0 72890.0 46205.0 ;
      RECT  72185.0 47550.0 72890.0 46205.0 ;
      RECT  72185.0 47550.0 72890.0 48895.0 ;
      RECT  72185.0 50240.0 72890.0 48895.0 ;
      RECT  72185.0 50240.0 72890.0 51585.0 ;
      RECT  72185.0 52930.0 72890.0 51585.0 ;
      RECT  72185.0 52930.0 72890.0 54275.0 ;
      RECT  72185.0 55620.0 72890.0 54275.0 ;
      RECT  72185.0 55620.0 72890.0 56965.0 ;
      RECT  72185.0 58310.0 72890.0 56965.0 ;
      RECT  72185.0 58310.0 72890.0 59655.0 ;
      RECT  72185.0 61000.0 72890.0 59655.0 ;
      RECT  72185.0 61000.0 72890.0 62345.0 ;
      RECT  72185.0 63690.0 72890.0 62345.0 ;
      RECT  72185.0 63690.0 72890.0 65035.0 ;
      RECT  72185.0 66380.0 72890.0 65035.0 ;
      RECT  72185.0 66380.0 72890.0 67725.0 ;
      RECT  72185.0 69070.0 72890.0 67725.0 ;
      RECT  72185.0 69070.0 72890.0 70415.0 ;
      RECT  72185.0 71760.0 72890.0 70415.0 ;
      RECT  72185.0 71760.0 72890.0 73105.0 ;
      RECT  72185.0 74450.0 72890.0 73105.0 ;
      RECT  72185.0 74450.0 72890.0 75795.0 ;
      RECT  72185.0 77140.0 72890.0 75795.0 ;
      RECT  72185.0 77140.0 72890.0 78485.0 ;
      RECT  72185.0 79830.0 72890.0 78485.0 ;
      RECT  72185.0 79830.0 72890.0 81175.0 ;
      RECT  72185.0 82520.0 72890.0 81175.0 ;
      RECT  72185.0 82520.0 72890.0 83865.0 ;
      RECT  72185.0 85210.0 72890.0 83865.0 ;
      RECT  72185.0 85210.0 72890.0 86555.0 ;
      RECT  72185.0 87900.0 72890.0 86555.0 ;
      RECT  72185.0 87900.0 72890.0 89245.0 ;
      RECT  72185.0 90590.0 72890.0 89245.0 ;
      RECT  72185.0 90590.0 72890.0 91935.0 ;
      RECT  72185.0 93280.0 72890.0 91935.0 ;
      RECT  72185.0 93280.0 72890.0 94625.0 ;
      RECT  72185.0 95970.0 72890.0 94625.0 ;
      RECT  72185.0 95970.0 72890.0 97315.0 ;
      RECT  72185.0 98660.0 72890.0 97315.0 ;
      RECT  72185.0 98660.0 72890.0 100005.0 ;
      RECT  72185.0 101350.0 72890.0 100005.0 ;
      RECT  72185.0 101350.0 72890.0 102695.0 ;
      RECT  72185.0 104040.0 72890.0 102695.0 ;
      RECT  72185.0 104040.0 72890.0 105385.0 ;
      RECT  72185.0 106730.0 72890.0 105385.0 ;
      RECT  72185.0 106730.0 72890.0 108075.0 ;
      RECT  72185.0 109420.0 72890.0 108075.0 ;
      RECT  72185.0 109420.0 72890.0 110765.0 ;
      RECT  72185.0 112110.0 72890.0 110765.0 ;
      RECT  72185.0 112110.0 72890.0 113455.0 ;
      RECT  72185.0 114800.0 72890.0 113455.0 ;
      RECT  72185.0 114800.0 72890.0 116145.0 ;
      RECT  72185.0 117490.0 72890.0 116145.0 ;
      RECT  72185.0 117490.0 72890.0 118835.0 ;
      RECT  72185.0 120180.0 72890.0 118835.0 ;
      RECT  72185.0 120180.0 72890.0 121525.0 ;
      RECT  72185.0 122870.0 72890.0 121525.0 ;
      RECT  72185.0 122870.0 72890.0 124215.0 ;
      RECT  72185.0 125560.0 72890.0 124215.0 ;
      RECT  72185.0 125560.0 72890.0 126905.0 ;
      RECT  72185.0 128250.0 72890.0 126905.0 ;
      RECT  72185.0 128250.0 72890.0 129595.0 ;
      RECT  72185.0 130940.0 72890.0 129595.0 ;
      RECT  72185.0 130940.0 72890.0 132285.0 ;
      RECT  72185.0 133630.0 72890.0 132285.0 ;
      RECT  72185.0 133630.0 72890.0 134975.0 ;
      RECT  72185.0 136320.0 72890.0 134975.0 ;
      RECT  72185.0 136320.0 72890.0 137665.0 ;
      RECT  72185.0 139010.0 72890.0 137665.0 ;
      RECT  72185.0 139010.0 72890.0 140355.0 ;
      RECT  72185.0 141700.0 72890.0 140355.0 ;
      RECT  72185.0 141700.0 72890.0 143045.0 ;
      RECT  72185.0 144390.0 72890.0 143045.0 ;
      RECT  72185.0 144390.0 72890.0 145735.0 ;
      RECT  72185.0 147080.0 72890.0 145735.0 ;
      RECT  72185.0 147080.0 72890.0 148425.0 ;
      RECT  72185.0 149770.0 72890.0 148425.0 ;
      RECT  72185.0 149770.0 72890.0 151115.0 ;
      RECT  72185.0 152460.0 72890.0 151115.0 ;
      RECT  72185.0 152460.0 72890.0 153805.0 ;
      RECT  72185.0 155150.0 72890.0 153805.0 ;
      RECT  72185.0 155150.0 72890.0 156495.0 ;
      RECT  72185.0 157840.0 72890.0 156495.0 ;
      RECT  72185.0 157840.0 72890.0 159185.0 ;
      RECT  72185.0 160530.0 72890.0 159185.0 ;
      RECT  72185.0 160530.0 72890.0 161875.0 ;
      RECT  72185.0 163220.0 72890.0 161875.0 ;
      RECT  72185.0 163220.0 72890.0 164565.0 ;
      RECT  72185.0 165910.0 72890.0 164565.0 ;
      RECT  72185.0 165910.0 72890.0 167255.0 ;
      RECT  72185.0 168600.0 72890.0 167255.0 ;
      RECT  72185.0 168600.0 72890.0 169945.0 ;
      RECT  72185.0 171290.0 72890.0 169945.0 ;
      RECT  72185.0 171290.0 72890.0 172635.0 ;
      RECT  72185.0 173980.0 72890.0 172635.0 ;
      RECT  72185.0 173980.0 72890.0 175325.0 ;
      RECT  72185.0 176670.0 72890.0 175325.0 ;
      RECT  72185.0 176670.0 72890.0 178015.0 ;
      RECT  72185.0 179360.0 72890.0 178015.0 ;
      RECT  72185.0 179360.0 72890.0 180705.0 ;
      RECT  72185.0 182050.0 72890.0 180705.0 ;
      RECT  72185.0 182050.0 72890.0 183395.0 ;
      RECT  72185.0 184740.0 72890.0 183395.0 ;
      RECT  72185.0 184740.0 72890.0 186085.0 ;
      RECT  72185.0 187430.0 72890.0 186085.0 ;
      RECT  72185.0 187430.0 72890.0 188775.0 ;
      RECT  72185.0 190120.0 72890.0 188775.0 ;
      RECT  72185.0 190120.0 72890.0 191465.0 ;
      RECT  72185.0 192810.0 72890.0 191465.0 ;
      RECT  72185.0 192810.0 72890.0 194155.0 ;
      RECT  72185.0 195500.0 72890.0 194155.0 ;
      RECT  72185.0 195500.0 72890.0 196845.0 ;
      RECT  72185.0 198190.0 72890.0 196845.0 ;
      RECT  72185.0 198190.0 72890.0 199535.0 ;
      RECT  72185.0 200880.0 72890.0 199535.0 ;
      RECT  72185.0 200880.0 72890.0 202225.0 ;
      RECT  72185.0 203570.0 72890.0 202225.0 ;
      RECT  72185.0 203570.0 72890.0 204915.0 ;
      RECT  72185.0 206260.0 72890.0 204915.0 ;
      RECT  72890.0 34100.0 73595.0 35445.0 ;
      RECT  72890.0 36790.0 73595.0 35445.0 ;
      RECT  72890.0 36790.0 73595.0 38135.0 ;
      RECT  72890.0 39480.0 73595.0 38135.0 ;
      RECT  72890.0 39480.0 73595.0 40825.0 ;
      RECT  72890.0 42170.0 73595.0 40825.0 ;
      RECT  72890.0 42170.0 73595.0 43515.0 ;
      RECT  72890.0 44860.0 73595.0 43515.0 ;
      RECT  72890.0 44860.0 73595.0 46205.0 ;
      RECT  72890.0 47550.0 73595.0 46205.0 ;
      RECT  72890.0 47550.0 73595.0 48895.0 ;
      RECT  72890.0 50240.0 73595.0 48895.0 ;
      RECT  72890.0 50240.0 73595.0 51585.0 ;
      RECT  72890.0 52930.0 73595.0 51585.0 ;
      RECT  72890.0 52930.0 73595.0 54275.0 ;
      RECT  72890.0 55620.0 73595.0 54275.0 ;
      RECT  72890.0 55620.0 73595.0 56965.0 ;
      RECT  72890.0 58310.0 73595.0 56965.0 ;
      RECT  72890.0 58310.0 73595.0 59655.0 ;
      RECT  72890.0 61000.0 73595.0 59655.0 ;
      RECT  72890.0 61000.0 73595.0 62345.0 ;
      RECT  72890.0 63690.0 73595.0 62345.0 ;
      RECT  72890.0 63690.0 73595.0 65035.0 ;
      RECT  72890.0 66380.0 73595.0 65035.0 ;
      RECT  72890.0 66380.0 73595.0 67725.0 ;
      RECT  72890.0 69070.0 73595.0 67725.0 ;
      RECT  72890.0 69070.0 73595.0 70415.0 ;
      RECT  72890.0 71760.0 73595.0 70415.0 ;
      RECT  72890.0 71760.0 73595.0 73105.0 ;
      RECT  72890.0 74450.0 73595.0 73105.0 ;
      RECT  72890.0 74450.0 73595.0 75795.0 ;
      RECT  72890.0 77140.0 73595.0 75795.0 ;
      RECT  72890.0 77140.0 73595.0 78485.0 ;
      RECT  72890.0 79830.0 73595.0 78485.0 ;
      RECT  72890.0 79830.0 73595.0 81175.0 ;
      RECT  72890.0 82520.0 73595.0 81175.0 ;
      RECT  72890.0 82520.0 73595.0 83865.0 ;
      RECT  72890.0 85210.0 73595.0 83865.0 ;
      RECT  72890.0 85210.0 73595.0 86555.0 ;
      RECT  72890.0 87900.0 73595.0 86555.0 ;
      RECT  72890.0 87900.0 73595.0 89245.0 ;
      RECT  72890.0 90590.0 73595.0 89245.0 ;
      RECT  72890.0 90590.0 73595.0 91935.0 ;
      RECT  72890.0 93280.0 73595.0 91935.0 ;
      RECT  72890.0 93280.0 73595.0 94625.0 ;
      RECT  72890.0 95970.0 73595.0 94625.0 ;
      RECT  72890.0 95970.0 73595.0 97315.0 ;
      RECT  72890.0 98660.0 73595.0 97315.0 ;
      RECT  72890.0 98660.0 73595.0 100005.0 ;
      RECT  72890.0 101350.0 73595.0 100005.0 ;
      RECT  72890.0 101350.0 73595.0 102695.0 ;
      RECT  72890.0 104040.0 73595.0 102695.0 ;
      RECT  72890.0 104040.0 73595.0 105385.0 ;
      RECT  72890.0 106730.0 73595.0 105385.0 ;
      RECT  72890.0 106730.0 73595.0 108075.0 ;
      RECT  72890.0 109420.0 73595.0 108075.0 ;
      RECT  72890.0 109420.0 73595.0 110765.0 ;
      RECT  72890.0 112110.0 73595.0 110765.0 ;
      RECT  72890.0 112110.0 73595.0 113455.0 ;
      RECT  72890.0 114800.0 73595.0 113455.0 ;
      RECT  72890.0 114800.0 73595.0 116145.0 ;
      RECT  72890.0 117490.0 73595.0 116145.0 ;
      RECT  72890.0 117490.0 73595.0 118835.0 ;
      RECT  72890.0 120180.0 73595.0 118835.0 ;
      RECT  72890.0 120180.0 73595.0 121525.0 ;
      RECT  72890.0 122870.0 73595.0 121525.0 ;
      RECT  72890.0 122870.0 73595.0 124215.0 ;
      RECT  72890.0 125560.0 73595.0 124215.0 ;
      RECT  72890.0 125560.0 73595.0 126905.0 ;
      RECT  72890.0 128250.0 73595.0 126905.0 ;
      RECT  72890.0 128250.0 73595.0 129595.0 ;
      RECT  72890.0 130940.0 73595.0 129595.0 ;
      RECT  72890.0 130940.0 73595.0 132285.0 ;
      RECT  72890.0 133630.0 73595.0 132285.0 ;
      RECT  72890.0 133630.0 73595.0 134975.0 ;
      RECT  72890.0 136320.0 73595.0 134975.0 ;
      RECT  72890.0 136320.0 73595.0 137665.0 ;
      RECT  72890.0 139010.0 73595.0 137665.0 ;
      RECT  72890.0 139010.0 73595.0 140355.0 ;
      RECT  72890.0 141700.0 73595.0 140355.0 ;
      RECT  72890.0 141700.0 73595.0 143045.0 ;
      RECT  72890.0 144390.0 73595.0 143045.0 ;
      RECT  72890.0 144390.0 73595.0 145735.0 ;
      RECT  72890.0 147080.0 73595.0 145735.0 ;
      RECT  72890.0 147080.0 73595.0 148425.0 ;
      RECT  72890.0 149770.0 73595.0 148425.0 ;
      RECT  72890.0 149770.0 73595.0 151115.0 ;
      RECT  72890.0 152460.0 73595.0 151115.0 ;
      RECT  72890.0 152460.0 73595.0 153805.0 ;
      RECT  72890.0 155150.0 73595.0 153805.0 ;
      RECT  72890.0 155150.0 73595.0 156495.0 ;
      RECT  72890.0 157840.0 73595.0 156495.0 ;
      RECT  72890.0 157840.0 73595.0 159185.0 ;
      RECT  72890.0 160530.0 73595.0 159185.0 ;
      RECT  72890.0 160530.0 73595.0 161875.0 ;
      RECT  72890.0 163220.0 73595.0 161875.0 ;
      RECT  72890.0 163220.0 73595.0 164565.0 ;
      RECT  72890.0 165910.0 73595.0 164565.0 ;
      RECT  72890.0 165910.0 73595.0 167255.0 ;
      RECT  72890.0 168600.0 73595.0 167255.0 ;
      RECT  72890.0 168600.0 73595.0 169945.0 ;
      RECT  72890.0 171290.0 73595.0 169945.0 ;
      RECT  72890.0 171290.0 73595.0 172635.0 ;
      RECT  72890.0 173980.0 73595.0 172635.0 ;
      RECT  72890.0 173980.0 73595.0 175325.0 ;
      RECT  72890.0 176670.0 73595.0 175325.0 ;
      RECT  72890.0 176670.0 73595.0 178015.0 ;
      RECT  72890.0 179360.0 73595.0 178015.0 ;
      RECT  72890.0 179360.0 73595.0 180705.0 ;
      RECT  72890.0 182050.0 73595.0 180705.0 ;
      RECT  72890.0 182050.0 73595.0 183395.0 ;
      RECT  72890.0 184740.0 73595.0 183395.0 ;
      RECT  72890.0 184740.0 73595.0 186085.0 ;
      RECT  72890.0 187430.0 73595.0 186085.0 ;
      RECT  72890.0 187430.0 73595.0 188775.0 ;
      RECT  72890.0 190120.0 73595.0 188775.0 ;
      RECT  72890.0 190120.0 73595.0 191465.0 ;
      RECT  72890.0 192810.0 73595.0 191465.0 ;
      RECT  72890.0 192810.0 73595.0 194155.0 ;
      RECT  72890.0 195500.0 73595.0 194155.0 ;
      RECT  72890.0 195500.0 73595.0 196845.0 ;
      RECT  72890.0 198190.0 73595.0 196845.0 ;
      RECT  72890.0 198190.0 73595.0 199535.0 ;
      RECT  72890.0 200880.0 73595.0 199535.0 ;
      RECT  72890.0 200880.0 73595.0 202225.0 ;
      RECT  72890.0 203570.0 73595.0 202225.0 ;
      RECT  72890.0 203570.0 73595.0 204915.0 ;
      RECT  72890.0 206260.0 73595.0 204915.0 ;
      RECT  73595.0 34100.0 74300.0 35445.0 ;
      RECT  73595.0 36790.0 74300.0 35445.0 ;
      RECT  73595.0 36790.0 74300.0 38135.0 ;
      RECT  73595.0 39480.0 74300.0 38135.0 ;
      RECT  73595.0 39480.0 74300.0 40825.0 ;
      RECT  73595.0 42170.0 74300.0 40825.0 ;
      RECT  73595.0 42170.0 74300.0 43515.0 ;
      RECT  73595.0 44860.0 74300.0 43515.0 ;
      RECT  73595.0 44860.0 74300.0 46205.0 ;
      RECT  73595.0 47550.0 74300.0 46205.0 ;
      RECT  73595.0 47550.0 74300.0 48895.0 ;
      RECT  73595.0 50240.0 74300.0 48895.0 ;
      RECT  73595.0 50240.0 74300.0 51585.0 ;
      RECT  73595.0 52930.0 74300.0 51585.0 ;
      RECT  73595.0 52930.0 74300.0 54275.0 ;
      RECT  73595.0 55620.0 74300.0 54275.0 ;
      RECT  73595.0 55620.0 74300.0 56965.0 ;
      RECT  73595.0 58310.0 74300.0 56965.0 ;
      RECT  73595.0 58310.0 74300.0 59655.0 ;
      RECT  73595.0 61000.0 74300.0 59655.0 ;
      RECT  73595.0 61000.0 74300.0 62345.0 ;
      RECT  73595.0 63690.0 74300.0 62345.0 ;
      RECT  73595.0 63690.0 74300.0 65035.0 ;
      RECT  73595.0 66380.0 74300.0 65035.0 ;
      RECT  73595.0 66380.0 74300.0 67725.0 ;
      RECT  73595.0 69070.0 74300.0 67725.0 ;
      RECT  73595.0 69070.0 74300.0 70415.0 ;
      RECT  73595.0 71760.0 74300.0 70415.0 ;
      RECT  73595.0 71760.0 74300.0 73105.0 ;
      RECT  73595.0 74450.0 74300.0 73105.0 ;
      RECT  73595.0 74450.0 74300.0 75795.0 ;
      RECT  73595.0 77140.0 74300.0 75795.0 ;
      RECT  73595.0 77140.0 74300.0 78485.0 ;
      RECT  73595.0 79830.0 74300.0 78485.0 ;
      RECT  73595.0 79830.0 74300.0 81175.0 ;
      RECT  73595.0 82520.0 74300.0 81175.0 ;
      RECT  73595.0 82520.0 74300.0 83865.0 ;
      RECT  73595.0 85210.0 74300.0 83865.0 ;
      RECT  73595.0 85210.0 74300.0 86555.0 ;
      RECT  73595.0 87900.0 74300.0 86555.0 ;
      RECT  73595.0 87900.0 74300.0 89245.0 ;
      RECT  73595.0 90590.0 74300.0 89245.0 ;
      RECT  73595.0 90590.0 74300.0 91935.0 ;
      RECT  73595.0 93280.0 74300.0 91935.0 ;
      RECT  73595.0 93280.0 74300.0 94625.0 ;
      RECT  73595.0 95970.0 74300.0 94625.0 ;
      RECT  73595.0 95970.0 74300.0 97315.0 ;
      RECT  73595.0 98660.0 74300.0 97315.0 ;
      RECT  73595.0 98660.0 74300.0 100005.0 ;
      RECT  73595.0 101350.0 74300.0 100005.0 ;
      RECT  73595.0 101350.0 74300.0 102695.0 ;
      RECT  73595.0 104040.0 74300.0 102695.0 ;
      RECT  73595.0 104040.0 74300.0 105385.0 ;
      RECT  73595.0 106730.0 74300.0 105385.0 ;
      RECT  73595.0 106730.0 74300.0 108075.0 ;
      RECT  73595.0 109420.0 74300.0 108075.0 ;
      RECT  73595.0 109420.0 74300.0 110765.0 ;
      RECT  73595.0 112110.0 74300.0 110765.0 ;
      RECT  73595.0 112110.0 74300.0 113455.0 ;
      RECT  73595.0 114800.0 74300.0 113455.0 ;
      RECT  73595.0 114800.0 74300.0 116145.0 ;
      RECT  73595.0 117490.0 74300.0 116145.0 ;
      RECT  73595.0 117490.0 74300.0 118835.0 ;
      RECT  73595.0 120180.0 74300.0 118835.0 ;
      RECT  73595.0 120180.0 74300.0 121525.0 ;
      RECT  73595.0 122870.0 74300.0 121525.0 ;
      RECT  73595.0 122870.0 74300.0 124215.0 ;
      RECT  73595.0 125560.0 74300.0 124215.0 ;
      RECT  73595.0 125560.0 74300.0 126905.0 ;
      RECT  73595.0 128250.0 74300.0 126905.0 ;
      RECT  73595.0 128250.0 74300.0 129595.0 ;
      RECT  73595.0 130940.0 74300.0 129595.0 ;
      RECT  73595.0 130940.0 74300.0 132285.0 ;
      RECT  73595.0 133630.0 74300.0 132285.0 ;
      RECT  73595.0 133630.0 74300.0 134975.0 ;
      RECT  73595.0 136320.0 74300.0 134975.0 ;
      RECT  73595.0 136320.0 74300.0 137665.0 ;
      RECT  73595.0 139010.0 74300.0 137665.0 ;
      RECT  73595.0 139010.0 74300.0 140355.0 ;
      RECT  73595.0 141700.0 74300.0 140355.0 ;
      RECT  73595.0 141700.0 74300.0 143045.0 ;
      RECT  73595.0 144390.0 74300.0 143045.0 ;
      RECT  73595.0 144390.0 74300.0 145735.0 ;
      RECT  73595.0 147080.0 74300.0 145735.0 ;
      RECT  73595.0 147080.0 74300.0 148425.0 ;
      RECT  73595.0 149770.0 74300.0 148425.0 ;
      RECT  73595.0 149770.0 74300.0 151115.0 ;
      RECT  73595.0 152460.0 74300.0 151115.0 ;
      RECT  73595.0 152460.0 74300.0 153805.0 ;
      RECT  73595.0 155150.0 74300.0 153805.0 ;
      RECT  73595.0 155150.0 74300.0 156495.0 ;
      RECT  73595.0 157840.0 74300.0 156495.0 ;
      RECT  73595.0 157840.0 74300.0 159185.0 ;
      RECT  73595.0 160530.0 74300.0 159185.0 ;
      RECT  73595.0 160530.0 74300.0 161875.0 ;
      RECT  73595.0 163220.0 74300.0 161875.0 ;
      RECT  73595.0 163220.0 74300.0 164565.0 ;
      RECT  73595.0 165910.0 74300.0 164565.0 ;
      RECT  73595.0 165910.0 74300.0 167255.0 ;
      RECT  73595.0 168600.0 74300.0 167255.0 ;
      RECT  73595.0 168600.0 74300.0 169945.0 ;
      RECT  73595.0 171290.0 74300.0 169945.0 ;
      RECT  73595.0 171290.0 74300.0 172635.0 ;
      RECT  73595.0 173980.0 74300.0 172635.0 ;
      RECT  73595.0 173980.0 74300.0 175325.0 ;
      RECT  73595.0 176670.0 74300.0 175325.0 ;
      RECT  73595.0 176670.0 74300.0 178015.0 ;
      RECT  73595.0 179360.0 74300.0 178015.0 ;
      RECT  73595.0 179360.0 74300.0 180705.0 ;
      RECT  73595.0 182050.0 74300.0 180705.0 ;
      RECT  73595.0 182050.0 74300.0 183395.0 ;
      RECT  73595.0 184740.0 74300.0 183395.0 ;
      RECT  73595.0 184740.0 74300.0 186085.0 ;
      RECT  73595.0 187430.0 74300.0 186085.0 ;
      RECT  73595.0 187430.0 74300.0 188775.0 ;
      RECT  73595.0 190120.0 74300.0 188775.0 ;
      RECT  73595.0 190120.0 74300.0 191465.0 ;
      RECT  73595.0 192810.0 74300.0 191465.0 ;
      RECT  73595.0 192810.0 74300.0 194155.0 ;
      RECT  73595.0 195500.0 74300.0 194155.0 ;
      RECT  73595.0 195500.0 74300.0 196845.0 ;
      RECT  73595.0 198190.0 74300.0 196845.0 ;
      RECT  73595.0 198190.0 74300.0 199535.0 ;
      RECT  73595.0 200880.0 74300.0 199535.0 ;
      RECT  73595.0 200880.0 74300.0 202225.0 ;
      RECT  73595.0 203570.0 74300.0 202225.0 ;
      RECT  73595.0 203570.0 74300.0 204915.0 ;
      RECT  73595.0 206260.0 74300.0 204915.0 ;
      RECT  74300.0 34100.0 75005.0 35445.0 ;
      RECT  74300.0 36790.0 75005.0 35445.0 ;
      RECT  74300.0 36790.0 75005.0 38135.0 ;
      RECT  74300.0 39480.0 75005.0 38135.0 ;
      RECT  74300.0 39480.0 75005.0 40825.0 ;
      RECT  74300.0 42170.0 75005.0 40825.0 ;
      RECT  74300.0 42170.0 75005.0 43515.0 ;
      RECT  74300.0 44860.0 75005.0 43515.0 ;
      RECT  74300.0 44860.0 75005.0 46205.0 ;
      RECT  74300.0 47550.0 75005.0 46205.0 ;
      RECT  74300.0 47550.0 75005.0 48895.0 ;
      RECT  74300.0 50240.0 75005.0 48895.0 ;
      RECT  74300.0 50240.0 75005.0 51585.0 ;
      RECT  74300.0 52930.0 75005.0 51585.0 ;
      RECT  74300.0 52930.0 75005.0 54275.0 ;
      RECT  74300.0 55620.0 75005.0 54275.0 ;
      RECT  74300.0 55620.0 75005.0 56965.0 ;
      RECT  74300.0 58310.0 75005.0 56965.0 ;
      RECT  74300.0 58310.0 75005.0 59655.0 ;
      RECT  74300.0 61000.0 75005.0 59655.0 ;
      RECT  74300.0 61000.0 75005.0 62345.0 ;
      RECT  74300.0 63690.0 75005.0 62345.0 ;
      RECT  74300.0 63690.0 75005.0 65035.0 ;
      RECT  74300.0 66380.0 75005.0 65035.0 ;
      RECT  74300.0 66380.0 75005.0 67725.0 ;
      RECT  74300.0 69070.0 75005.0 67725.0 ;
      RECT  74300.0 69070.0 75005.0 70415.0 ;
      RECT  74300.0 71760.0 75005.0 70415.0 ;
      RECT  74300.0 71760.0 75005.0 73105.0 ;
      RECT  74300.0 74450.0 75005.0 73105.0 ;
      RECT  74300.0 74450.0 75005.0 75795.0 ;
      RECT  74300.0 77140.0 75005.0 75795.0 ;
      RECT  74300.0 77140.0 75005.0 78485.0 ;
      RECT  74300.0 79830.0 75005.0 78485.0 ;
      RECT  74300.0 79830.0 75005.0 81175.0 ;
      RECT  74300.0 82520.0 75005.0 81175.0 ;
      RECT  74300.0 82520.0 75005.0 83865.0 ;
      RECT  74300.0 85210.0 75005.0 83865.0 ;
      RECT  74300.0 85210.0 75005.0 86555.0 ;
      RECT  74300.0 87900.0 75005.0 86555.0 ;
      RECT  74300.0 87900.0 75005.0 89245.0 ;
      RECT  74300.0 90590.0 75005.0 89245.0 ;
      RECT  74300.0 90590.0 75005.0 91935.0 ;
      RECT  74300.0 93280.0 75005.0 91935.0 ;
      RECT  74300.0 93280.0 75005.0 94625.0 ;
      RECT  74300.0 95970.0 75005.0 94625.0 ;
      RECT  74300.0 95970.0 75005.0 97315.0 ;
      RECT  74300.0 98660.0 75005.0 97315.0 ;
      RECT  74300.0 98660.0 75005.0 100005.0 ;
      RECT  74300.0 101350.0 75005.0 100005.0 ;
      RECT  74300.0 101350.0 75005.0 102695.0 ;
      RECT  74300.0 104040.0 75005.0 102695.0 ;
      RECT  74300.0 104040.0 75005.0 105385.0 ;
      RECT  74300.0 106730.0 75005.0 105385.0 ;
      RECT  74300.0 106730.0 75005.0 108075.0 ;
      RECT  74300.0 109420.0 75005.0 108075.0 ;
      RECT  74300.0 109420.0 75005.0 110765.0 ;
      RECT  74300.0 112110.0 75005.0 110765.0 ;
      RECT  74300.0 112110.0 75005.0 113455.0 ;
      RECT  74300.0 114800.0 75005.0 113455.0 ;
      RECT  74300.0 114800.0 75005.0 116145.0 ;
      RECT  74300.0 117490.0 75005.0 116145.0 ;
      RECT  74300.0 117490.0 75005.0 118835.0 ;
      RECT  74300.0 120180.0 75005.0 118835.0 ;
      RECT  74300.0 120180.0 75005.0 121525.0 ;
      RECT  74300.0 122870.0 75005.0 121525.0 ;
      RECT  74300.0 122870.0 75005.0 124215.0 ;
      RECT  74300.0 125560.0 75005.0 124215.0 ;
      RECT  74300.0 125560.0 75005.0 126905.0 ;
      RECT  74300.0 128250.0 75005.0 126905.0 ;
      RECT  74300.0 128250.0 75005.0 129595.0 ;
      RECT  74300.0 130940.0 75005.0 129595.0 ;
      RECT  74300.0 130940.0 75005.0 132285.0 ;
      RECT  74300.0 133630.0 75005.0 132285.0 ;
      RECT  74300.0 133630.0 75005.0 134975.0 ;
      RECT  74300.0 136320.0 75005.0 134975.0 ;
      RECT  74300.0 136320.0 75005.0 137665.0 ;
      RECT  74300.0 139010.0 75005.0 137665.0 ;
      RECT  74300.0 139010.0 75005.0 140355.0 ;
      RECT  74300.0 141700.0 75005.0 140355.0 ;
      RECT  74300.0 141700.0 75005.0 143045.0 ;
      RECT  74300.0 144390.0 75005.0 143045.0 ;
      RECT  74300.0 144390.0 75005.0 145735.0 ;
      RECT  74300.0 147080.0 75005.0 145735.0 ;
      RECT  74300.0 147080.0 75005.0 148425.0 ;
      RECT  74300.0 149770.0 75005.0 148425.0 ;
      RECT  74300.0 149770.0 75005.0 151115.0 ;
      RECT  74300.0 152460.0 75005.0 151115.0 ;
      RECT  74300.0 152460.0 75005.0 153805.0 ;
      RECT  74300.0 155150.0 75005.0 153805.0 ;
      RECT  74300.0 155150.0 75005.0 156495.0 ;
      RECT  74300.0 157840.0 75005.0 156495.0 ;
      RECT  74300.0 157840.0 75005.0 159185.0 ;
      RECT  74300.0 160530.0 75005.0 159185.0 ;
      RECT  74300.0 160530.0 75005.0 161875.0 ;
      RECT  74300.0 163220.0 75005.0 161875.0 ;
      RECT  74300.0 163220.0 75005.0 164565.0 ;
      RECT  74300.0 165910.0 75005.0 164565.0 ;
      RECT  74300.0 165910.0 75005.0 167255.0 ;
      RECT  74300.0 168600.0 75005.0 167255.0 ;
      RECT  74300.0 168600.0 75005.0 169945.0 ;
      RECT  74300.0 171290.0 75005.0 169945.0 ;
      RECT  74300.0 171290.0 75005.0 172635.0 ;
      RECT  74300.0 173980.0 75005.0 172635.0 ;
      RECT  74300.0 173980.0 75005.0 175325.0 ;
      RECT  74300.0 176670.0 75005.0 175325.0 ;
      RECT  74300.0 176670.0 75005.0 178015.0 ;
      RECT  74300.0 179360.0 75005.0 178015.0 ;
      RECT  74300.0 179360.0 75005.0 180705.0 ;
      RECT  74300.0 182050.0 75005.0 180705.0 ;
      RECT  74300.0 182050.0 75005.0 183395.0 ;
      RECT  74300.0 184740.0 75005.0 183395.0 ;
      RECT  74300.0 184740.0 75005.0 186085.0 ;
      RECT  74300.0 187430.0 75005.0 186085.0 ;
      RECT  74300.0 187430.0 75005.0 188775.0 ;
      RECT  74300.0 190120.0 75005.0 188775.0 ;
      RECT  74300.0 190120.0 75005.0 191465.0 ;
      RECT  74300.0 192810.0 75005.0 191465.0 ;
      RECT  74300.0 192810.0 75005.0 194155.0 ;
      RECT  74300.0 195500.0 75005.0 194155.0 ;
      RECT  74300.0 195500.0 75005.0 196845.0 ;
      RECT  74300.0 198190.0 75005.0 196845.0 ;
      RECT  74300.0 198190.0 75005.0 199535.0 ;
      RECT  74300.0 200880.0 75005.0 199535.0 ;
      RECT  74300.0 200880.0 75005.0 202225.0 ;
      RECT  74300.0 203570.0 75005.0 202225.0 ;
      RECT  74300.0 203570.0 75005.0 204915.0 ;
      RECT  74300.0 206260.0 75005.0 204915.0 ;
      RECT  75005.0 34100.0 75710.0 35445.0 ;
      RECT  75005.0 36790.0 75710.0 35445.0 ;
      RECT  75005.0 36790.0 75710.0 38135.0 ;
      RECT  75005.0 39480.0 75710.0 38135.0 ;
      RECT  75005.0 39480.0 75710.0 40825.0 ;
      RECT  75005.0 42170.0 75710.0 40825.0 ;
      RECT  75005.0 42170.0 75710.0 43515.0 ;
      RECT  75005.0 44860.0 75710.0 43515.0 ;
      RECT  75005.0 44860.0 75710.0 46205.0 ;
      RECT  75005.0 47550.0 75710.0 46205.0 ;
      RECT  75005.0 47550.0 75710.0 48895.0 ;
      RECT  75005.0 50240.0 75710.0 48895.0 ;
      RECT  75005.0 50240.0 75710.0 51585.0 ;
      RECT  75005.0 52930.0 75710.0 51585.0 ;
      RECT  75005.0 52930.0 75710.0 54275.0 ;
      RECT  75005.0 55620.0 75710.0 54275.0 ;
      RECT  75005.0 55620.0 75710.0 56965.0 ;
      RECT  75005.0 58310.0 75710.0 56965.0 ;
      RECT  75005.0 58310.0 75710.0 59655.0 ;
      RECT  75005.0 61000.0 75710.0 59655.0 ;
      RECT  75005.0 61000.0 75710.0 62345.0 ;
      RECT  75005.0 63690.0 75710.0 62345.0 ;
      RECT  75005.0 63690.0 75710.0 65035.0 ;
      RECT  75005.0 66380.0 75710.0 65035.0 ;
      RECT  75005.0 66380.0 75710.0 67725.0 ;
      RECT  75005.0 69070.0 75710.0 67725.0 ;
      RECT  75005.0 69070.0 75710.0 70415.0 ;
      RECT  75005.0 71760.0 75710.0 70415.0 ;
      RECT  75005.0 71760.0 75710.0 73105.0 ;
      RECT  75005.0 74450.0 75710.0 73105.0 ;
      RECT  75005.0 74450.0 75710.0 75795.0 ;
      RECT  75005.0 77140.0 75710.0 75795.0 ;
      RECT  75005.0 77140.0 75710.0 78485.0 ;
      RECT  75005.0 79830.0 75710.0 78485.0 ;
      RECT  75005.0 79830.0 75710.0 81175.0 ;
      RECT  75005.0 82520.0 75710.0 81175.0 ;
      RECT  75005.0 82520.0 75710.0 83865.0 ;
      RECT  75005.0 85210.0 75710.0 83865.0 ;
      RECT  75005.0 85210.0 75710.0 86555.0 ;
      RECT  75005.0 87900.0 75710.0 86555.0 ;
      RECT  75005.0 87900.0 75710.0 89245.0 ;
      RECT  75005.0 90590.0 75710.0 89245.0 ;
      RECT  75005.0 90590.0 75710.0 91935.0 ;
      RECT  75005.0 93280.0 75710.0 91935.0 ;
      RECT  75005.0 93280.0 75710.0 94625.0 ;
      RECT  75005.0 95970.0 75710.0 94625.0 ;
      RECT  75005.0 95970.0 75710.0 97315.0 ;
      RECT  75005.0 98660.0 75710.0 97315.0 ;
      RECT  75005.0 98660.0 75710.0 100005.0 ;
      RECT  75005.0 101350.0 75710.0 100005.0 ;
      RECT  75005.0 101350.0 75710.0 102695.0 ;
      RECT  75005.0 104040.0 75710.0 102695.0 ;
      RECT  75005.0 104040.0 75710.0 105385.0 ;
      RECT  75005.0 106730.0 75710.0 105385.0 ;
      RECT  75005.0 106730.0 75710.0 108075.0 ;
      RECT  75005.0 109420.0 75710.0 108075.0 ;
      RECT  75005.0 109420.0 75710.0 110765.0 ;
      RECT  75005.0 112110.0 75710.0 110765.0 ;
      RECT  75005.0 112110.0 75710.0 113455.0 ;
      RECT  75005.0 114800.0 75710.0 113455.0 ;
      RECT  75005.0 114800.0 75710.0 116145.0 ;
      RECT  75005.0 117490.0 75710.0 116145.0 ;
      RECT  75005.0 117490.0 75710.0 118835.0 ;
      RECT  75005.0 120180.0 75710.0 118835.0 ;
      RECT  75005.0 120180.0 75710.0 121525.0 ;
      RECT  75005.0 122870.0 75710.0 121525.0 ;
      RECT  75005.0 122870.0 75710.0 124215.0 ;
      RECT  75005.0 125560.0 75710.0 124215.0 ;
      RECT  75005.0 125560.0 75710.0 126905.0 ;
      RECT  75005.0 128250.0 75710.0 126905.0 ;
      RECT  75005.0 128250.0 75710.0 129595.0 ;
      RECT  75005.0 130940.0 75710.0 129595.0 ;
      RECT  75005.0 130940.0 75710.0 132285.0 ;
      RECT  75005.0 133630.0 75710.0 132285.0 ;
      RECT  75005.0 133630.0 75710.0 134975.0 ;
      RECT  75005.0 136320.0 75710.0 134975.0 ;
      RECT  75005.0 136320.0 75710.0 137665.0 ;
      RECT  75005.0 139010.0 75710.0 137665.0 ;
      RECT  75005.0 139010.0 75710.0 140355.0 ;
      RECT  75005.0 141700.0 75710.0 140355.0 ;
      RECT  75005.0 141700.0 75710.0 143045.0 ;
      RECT  75005.0 144390.0 75710.0 143045.0 ;
      RECT  75005.0 144390.0 75710.0 145735.0 ;
      RECT  75005.0 147080.0 75710.0 145735.0 ;
      RECT  75005.0 147080.0 75710.0 148425.0 ;
      RECT  75005.0 149770.0 75710.0 148425.0 ;
      RECT  75005.0 149770.0 75710.0 151115.0 ;
      RECT  75005.0 152460.0 75710.0 151115.0 ;
      RECT  75005.0 152460.0 75710.0 153805.0 ;
      RECT  75005.0 155150.0 75710.0 153805.0 ;
      RECT  75005.0 155150.0 75710.0 156495.0 ;
      RECT  75005.0 157840.0 75710.0 156495.0 ;
      RECT  75005.0 157840.0 75710.0 159185.0 ;
      RECT  75005.0 160530.0 75710.0 159185.0 ;
      RECT  75005.0 160530.0 75710.0 161875.0 ;
      RECT  75005.0 163220.0 75710.0 161875.0 ;
      RECT  75005.0 163220.0 75710.0 164565.0 ;
      RECT  75005.0 165910.0 75710.0 164565.0 ;
      RECT  75005.0 165910.0 75710.0 167255.0 ;
      RECT  75005.0 168600.0 75710.0 167255.0 ;
      RECT  75005.0 168600.0 75710.0 169945.0 ;
      RECT  75005.0 171290.0 75710.0 169945.0 ;
      RECT  75005.0 171290.0 75710.0 172635.0 ;
      RECT  75005.0 173980.0 75710.0 172635.0 ;
      RECT  75005.0 173980.0 75710.0 175325.0 ;
      RECT  75005.0 176670.0 75710.0 175325.0 ;
      RECT  75005.0 176670.0 75710.0 178015.0 ;
      RECT  75005.0 179360.0 75710.0 178015.0 ;
      RECT  75005.0 179360.0 75710.0 180705.0 ;
      RECT  75005.0 182050.0 75710.0 180705.0 ;
      RECT  75005.0 182050.0 75710.0 183395.0 ;
      RECT  75005.0 184740.0 75710.0 183395.0 ;
      RECT  75005.0 184740.0 75710.0 186085.0 ;
      RECT  75005.0 187430.0 75710.0 186085.0 ;
      RECT  75005.0 187430.0 75710.0 188775.0 ;
      RECT  75005.0 190120.0 75710.0 188775.0 ;
      RECT  75005.0 190120.0 75710.0 191465.0 ;
      RECT  75005.0 192810.0 75710.0 191465.0 ;
      RECT  75005.0 192810.0 75710.0 194155.0 ;
      RECT  75005.0 195500.0 75710.0 194155.0 ;
      RECT  75005.0 195500.0 75710.0 196845.0 ;
      RECT  75005.0 198190.0 75710.0 196845.0 ;
      RECT  75005.0 198190.0 75710.0 199535.0 ;
      RECT  75005.0 200880.0 75710.0 199535.0 ;
      RECT  75005.0 200880.0 75710.0 202225.0 ;
      RECT  75005.0 203570.0 75710.0 202225.0 ;
      RECT  75005.0 203570.0 75710.0 204915.0 ;
      RECT  75005.0 206260.0 75710.0 204915.0 ;
      RECT  75710.0 34100.0 76415.0 35445.0 ;
      RECT  75710.0 36790.0 76415.0 35445.0 ;
      RECT  75710.0 36790.0 76415.0 38135.0 ;
      RECT  75710.0 39480.0 76415.0 38135.0 ;
      RECT  75710.0 39480.0 76415.0 40825.0 ;
      RECT  75710.0 42170.0 76415.0 40825.0 ;
      RECT  75710.0 42170.0 76415.0 43515.0 ;
      RECT  75710.0 44860.0 76415.0 43515.0 ;
      RECT  75710.0 44860.0 76415.0 46205.0 ;
      RECT  75710.0 47550.0 76415.0 46205.0 ;
      RECT  75710.0 47550.0 76415.0 48895.0 ;
      RECT  75710.0 50240.0 76415.0 48895.0 ;
      RECT  75710.0 50240.0 76415.0 51585.0 ;
      RECT  75710.0 52930.0 76415.0 51585.0 ;
      RECT  75710.0 52930.0 76415.0 54275.0 ;
      RECT  75710.0 55620.0 76415.0 54275.0 ;
      RECT  75710.0 55620.0 76415.0 56965.0 ;
      RECT  75710.0 58310.0 76415.0 56965.0 ;
      RECT  75710.0 58310.0 76415.0 59655.0 ;
      RECT  75710.0 61000.0 76415.0 59655.0 ;
      RECT  75710.0 61000.0 76415.0 62345.0 ;
      RECT  75710.0 63690.0 76415.0 62345.0 ;
      RECT  75710.0 63690.0 76415.0 65035.0 ;
      RECT  75710.0 66380.0 76415.0 65035.0 ;
      RECT  75710.0 66380.0 76415.0 67725.0 ;
      RECT  75710.0 69070.0 76415.0 67725.0 ;
      RECT  75710.0 69070.0 76415.0 70415.0 ;
      RECT  75710.0 71760.0 76415.0 70415.0 ;
      RECT  75710.0 71760.0 76415.0 73105.0 ;
      RECT  75710.0 74450.0 76415.0 73105.0 ;
      RECT  75710.0 74450.0 76415.0 75795.0 ;
      RECT  75710.0 77140.0 76415.0 75795.0 ;
      RECT  75710.0 77140.0 76415.0 78485.0 ;
      RECT  75710.0 79830.0 76415.0 78485.0 ;
      RECT  75710.0 79830.0 76415.0 81175.0 ;
      RECT  75710.0 82520.0 76415.0 81175.0 ;
      RECT  75710.0 82520.0 76415.0 83865.0 ;
      RECT  75710.0 85210.0 76415.0 83865.0 ;
      RECT  75710.0 85210.0 76415.0 86555.0 ;
      RECT  75710.0 87900.0 76415.0 86555.0 ;
      RECT  75710.0 87900.0 76415.0 89245.0 ;
      RECT  75710.0 90590.0 76415.0 89245.0 ;
      RECT  75710.0 90590.0 76415.0 91935.0 ;
      RECT  75710.0 93280.0 76415.0 91935.0 ;
      RECT  75710.0 93280.0 76415.0 94625.0 ;
      RECT  75710.0 95970.0 76415.0 94625.0 ;
      RECT  75710.0 95970.0 76415.0 97315.0 ;
      RECT  75710.0 98660.0 76415.0 97315.0 ;
      RECT  75710.0 98660.0 76415.0 100005.0 ;
      RECT  75710.0 101350.0 76415.0 100005.0 ;
      RECT  75710.0 101350.0 76415.0 102695.0 ;
      RECT  75710.0 104040.0 76415.0 102695.0 ;
      RECT  75710.0 104040.0 76415.0 105385.0 ;
      RECT  75710.0 106730.0 76415.0 105385.0 ;
      RECT  75710.0 106730.0 76415.0 108075.0 ;
      RECT  75710.0 109420.0 76415.0 108075.0 ;
      RECT  75710.0 109420.0 76415.0 110765.0 ;
      RECT  75710.0 112110.0 76415.0 110765.0 ;
      RECT  75710.0 112110.0 76415.0 113455.0 ;
      RECT  75710.0 114800.0 76415.0 113455.0 ;
      RECT  75710.0 114800.0 76415.0 116145.0 ;
      RECT  75710.0 117490.0 76415.0 116145.0 ;
      RECT  75710.0 117490.0 76415.0 118835.0 ;
      RECT  75710.0 120180.0 76415.0 118835.0 ;
      RECT  75710.0 120180.0 76415.0 121525.0 ;
      RECT  75710.0 122870.0 76415.0 121525.0 ;
      RECT  75710.0 122870.0 76415.0 124215.0 ;
      RECT  75710.0 125560.0 76415.0 124215.0 ;
      RECT  75710.0 125560.0 76415.0 126905.0 ;
      RECT  75710.0 128250.0 76415.0 126905.0 ;
      RECT  75710.0 128250.0 76415.0 129595.0 ;
      RECT  75710.0 130940.0 76415.0 129595.0 ;
      RECT  75710.0 130940.0 76415.0 132285.0 ;
      RECT  75710.0 133630.0 76415.0 132285.0 ;
      RECT  75710.0 133630.0 76415.0 134975.0 ;
      RECT  75710.0 136320.0 76415.0 134975.0 ;
      RECT  75710.0 136320.0 76415.0 137665.0 ;
      RECT  75710.0 139010.0 76415.0 137665.0 ;
      RECT  75710.0 139010.0 76415.0 140355.0 ;
      RECT  75710.0 141700.0 76415.0 140355.0 ;
      RECT  75710.0 141700.0 76415.0 143045.0 ;
      RECT  75710.0 144390.0 76415.0 143045.0 ;
      RECT  75710.0 144390.0 76415.0 145735.0 ;
      RECT  75710.0 147080.0 76415.0 145735.0 ;
      RECT  75710.0 147080.0 76415.0 148425.0 ;
      RECT  75710.0 149770.0 76415.0 148425.0 ;
      RECT  75710.0 149770.0 76415.0 151115.0 ;
      RECT  75710.0 152460.0 76415.0 151115.0 ;
      RECT  75710.0 152460.0 76415.0 153805.0 ;
      RECT  75710.0 155150.0 76415.0 153805.0 ;
      RECT  75710.0 155150.0 76415.0 156495.0 ;
      RECT  75710.0 157840.0 76415.0 156495.0 ;
      RECT  75710.0 157840.0 76415.0 159185.0 ;
      RECT  75710.0 160530.0 76415.0 159185.0 ;
      RECT  75710.0 160530.0 76415.0 161875.0 ;
      RECT  75710.0 163220.0 76415.0 161875.0 ;
      RECT  75710.0 163220.0 76415.0 164565.0 ;
      RECT  75710.0 165910.0 76415.0 164565.0 ;
      RECT  75710.0 165910.0 76415.0 167255.0 ;
      RECT  75710.0 168600.0 76415.0 167255.0 ;
      RECT  75710.0 168600.0 76415.0 169945.0 ;
      RECT  75710.0 171290.0 76415.0 169945.0 ;
      RECT  75710.0 171290.0 76415.0 172635.0 ;
      RECT  75710.0 173980.0 76415.0 172635.0 ;
      RECT  75710.0 173980.0 76415.0 175325.0 ;
      RECT  75710.0 176670.0 76415.0 175325.0 ;
      RECT  75710.0 176670.0 76415.0 178015.0 ;
      RECT  75710.0 179360.0 76415.0 178015.0 ;
      RECT  75710.0 179360.0 76415.0 180705.0 ;
      RECT  75710.0 182050.0 76415.0 180705.0 ;
      RECT  75710.0 182050.0 76415.0 183395.0 ;
      RECT  75710.0 184740.0 76415.0 183395.0 ;
      RECT  75710.0 184740.0 76415.0 186085.0 ;
      RECT  75710.0 187430.0 76415.0 186085.0 ;
      RECT  75710.0 187430.0 76415.0 188775.0 ;
      RECT  75710.0 190120.0 76415.0 188775.0 ;
      RECT  75710.0 190120.0 76415.0 191465.0 ;
      RECT  75710.0 192810.0 76415.0 191465.0 ;
      RECT  75710.0 192810.0 76415.0 194155.0 ;
      RECT  75710.0 195500.0 76415.0 194155.0 ;
      RECT  75710.0 195500.0 76415.0 196845.0 ;
      RECT  75710.0 198190.0 76415.0 196845.0 ;
      RECT  75710.0 198190.0 76415.0 199535.0 ;
      RECT  75710.0 200880.0 76415.0 199535.0 ;
      RECT  75710.0 200880.0 76415.0 202225.0 ;
      RECT  75710.0 203570.0 76415.0 202225.0 ;
      RECT  75710.0 203570.0 76415.0 204915.0 ;
      RECT  75710.0 206260.0 76415.0 204915.0 ;
      RECT  76415.0 34100.0 77120.0 35445.0 ;
      RECT  76415.0 36790.0 77120.0 35445.0 ;
      RECT  76415.0 36790.0 77120.0 38135.0 ;
      RECT  76415.0 39480.0 77120.0 38135.0 ;
      RECT  76415.0 39480.0 77120.0 40825.0 ;
      RECT  76415.0 42170.0 77120.0 40825.0 ;
      RECT  76415.0 42170.0 77120.0 43515.0 ;
      RECT  76415.0 44860.0 77120.0 43515.0 ;
      RECT  76415.0 44860.0 77120.0 46205.0 ;
      RECT  76415.0 47550.0 77120.0 46205.0 ;
      RECT  76415.0 47550.0 77120.0 48895.0 ;
      RECT  76415.0 50240.0 77120.0 48895.0 ;
      RECT  76415.0 50240.0 77120.0 51585.0 ;
      RECT  76415.0 52930.0 77120.0 51585.0 ;
      RECT  76415.0 52930.0 77120.0 54275.0 ;
      RECT  76415.0 55620.0 77120.0 54275.0 ;
      RECT  76415.0 55620.0 77120.0 56965.0 ;
      RECT  76415.0 58310.0 77120.0 56965.0 ;
      RECT  76415.0 58310.0 77120.0 59655.0 ;
      RECT  76415.0 61000.0 77120.0 59655.0 ;
      RECT  76415.0 61000.0 77120.0 62345.0 ;
      RECT  76415.0 63690.0 77120.0 62345.0 ;
      RECT  76415.0 63690.0 77120.0 65035.0 ;
      RECT  76415.0 66380.0 77120.0 65035.0 ;
      RECT  76415.0 66380.0 77120.0 67725.0 ;
      RECT  76415.0 69070.0 77120.0 67725.0 ;
      RECT  76415.0 69070.0 77120.0 70415.0 ;
      RECT  76415.0 71760.0 77120.0 70415.0 ;
      RECT  76415.0 71760.0 77120.0 73105.0 ;
      RECT  76415.0 74450.0 77120.0 73105.0 ;
      RECT  76415.0 74450.0 77120.0 75795.0 ;
      RECT  76415.0 77140.0 77120.0 75795.0 ;
      RECT  76415.0 77140.0 77120.0 78485.0 ;
      RECT  76415.0 79830.0 77120.0 78485.0 ;
      RECT  76415.0 79830.0 77120.0 81175.0 ;
      RECT  76415.0 82520.0 77120.0 81175.0 ;
      RECT  76415.0 82520.0 77120.0 83865.0 ;
      RECT  76415.0 85210.0 77120.0 83865.0 ;
      RECT  76415.0 85210.0 77120.0 86555.0 ;
      RECT  76415.0 87900.0 77120.0 86555.0 ;
      RECT  76415.0 87900.0 77120.0 89245.0 ;
      RECT  76415.0 90590.0 77120.0 89245.0 ;
      RECT  76415.0 90590.0 77120.0 91935.0 ;
      RECT  76415.0 93280.0 77120.0 91935.0 ;
      RECT  76415.0 93280.0 77120.0 94625.0 ;
      RECT  76415.0 95970.0 77120.0 94625.0 ;
      RECT  76415.0 95970.0 77120.0 97315.0 ;
      RECT  76415.0 98660.0 77120.0 97315.0 ;
      RECT  76415.0 98660.0 77120.0 100005.0 ;
      RECT  76415.0 101350.0 77120.0 100005.0 ;
      RECT  76415.0 101350.0 77120.0 102695.0 ;
      RECT  76415.0 104040.0 77120.0 102695.0 ;
      RECT  76415.0 104040.0 77120.0 105385.0 ;
      RECT  76415.0 106730.0 77120.0 105385.0 ;
      RECT  76415.0 106730.0 77120.0 108075.0 ;
      RECT  76415.0 109420.0 77120.0 108075.0 ;
      RECT  76415.0 109420.0 77120.0 110765.0 ;
      RECT  76415.0 112110.0 77120.0 110765.0 ;
      RECT  76415.0 112110.0 77120.0 113455.0 ;
      RECT  76415.0 114800.0 77120.0 113455.0 ;
      RECT  76415.0 114800.0 77120.0 116145.0 ;
      RECT  76415.0 117490.0 77120.0 116145.0 ;
      RECT  76415.0 117490.0 77120.0 118835.0 ;
      RECT  76415.0 120180.0 77120.0 118835.0 ;
      RECT  76415.0 120180.0 77120.0 121525.0 ;
      RECT  76415.0 122870.0 77120.0 121525.0 ;
      RECT  76415.0 122870.0 77120.0 124215.0 ;
      RECT  76415.0 125560.0 77120.0 124215.0 ;
      RECT  76415.0 125560.0 77120.0 126905.0 ;
      RECT  76415.0 128250.0 77120.0 126905.0 ;
      RECT  76415.0 128250.0 77120.0 129595.0 ;
      RECT  76415.0 130940.0 77120.0 129595.0 ;
      RECT  76415.0 130940.0 77120.0 132285.0 ;
      RECT  76415.0 133630.0 77120.0 132285.0 ;
      RECT  76415.0 133630.0 77120.0 134975.0 ;
      RECT  76415.0 136320.0 77120.0 134975.0 ;
      RECT  76415.0 136320.0 77120.0 137665.0 ;
      RECT  76415.0 139010.0 77120.0 137665.0 ;
      RECT  76415.0 139010.0 77120.0 140355.0 ;
      RECT  76415.0 141700.0 77120.0 140355.0 ;
      RECT  76415.0 141700.0 77120.0 143045.0 ;
      RECT  76415.0 144390.0 77120.0 143045.0 ;
      RECT  76415.0 144390.0 77120.0 145735.0 ;
      RECT  76415.0 147080.0 77120.0 145735.0 ;
      RECT  76415.0 147080.0 77120.0 148425.0 ;
      RECT  76415.0 149770.0 77120.0 148425.0 ;
      RECT  76415.0 149770.0 77120.0 151115.0 ;
      RECT  76415.0 152460.0 77120.0 151115.0 ;
      RECT  76415.0 152460.0 77120.0 153805.0 ;
      RECT  76415.0 155150.0 77120.0 153805.0 ;
      RECT  76415.0 155150.0 77120.0 156495.0 ;
      RECT  76415.0 157840.0 77120.0 156495.0 ;
      RECT  76415.0 157840.0 77120.0 159185.0 ;
      RECT  76415.0 160530.0 77120.0 159185.0 ;
      RECT  76415.0 160530.0 77120.0 161875.0 ;
      RECT  76415.0 163220.0 77120.0 161875.0 ;
      RECT  76415.0 163220.0 77120.0 164565.0 ;
      RECT  76415.0 165910.0 77120.0 164565.0 ;
      RECT  76415.0 165910.0 77120.0 167255.0 ;
      RECT  76415.0 168600.0 77120.0 167255.0 ;
      RECT  76415.0 168600.0 77120.0 169945.0 ;
      RECT  76415.0 171290.0 77120.0 169945.0 ;
      RECT  76415.0 171290.0 77120.0 172635.0 ;
      RECT  76415.0 173980.0 77120.0 172635.0 ;
      RECT  76415.0 173980.0 77120.0 175325.0 ;
      RECT  76415.0 176670.0 77120.0 175325.0 ;
      RECT  76415.0 176670.0 77120.0 178015.0 ;
      RECT  76415.0 179360.0 77120.0 178015.0 ;
      RECT  76415.0 179360.0 77120.0 180705.0 ;
      RECT  76415.0 182050.0 77120.0 180705.0 ;
      RECT  76415.0 182050.0 77120.0 183395.0 ;
      RECT  76415.0 184740.0 77120.0 183395.0 ;
      RECT  76415.0 184740.0 77120.0 186085.0 ;
      RECT  76415.0 187430.0 77120.0 186085.0 ;
      RECT  76415.0 187430.0 77120.0 188775.0 ;
      RECT  76415.0 190120.0 77120.0 188775.0 ;
      RECT  76415.0 190120.0 77120.0 191465.0 ;
      RECT  76415.0 192810.0 77120.0 191465.0 ;
      RECT  76415.0 192810.0 77120.0 194155.0 ;
      RECT  76415.0 195500.0 77120.0 194155.0 ;
      RECT  76415.0 195500.0 77120.0 196845.0 ;
      RECT  76415.0 198190.0 77120.0 196845.0 ;
      RECT  76415.0 198190.0 77120.0 199535.0 ;
      RECT  76415.0 200880.0 77120.0 199535.0 ;
      RECT  76415.0 200880.0 77120.0 202225.0 ;
      RECT  76415.0 203570.0 77120.0 202225.0 ;
      RECT  76415.0 203570.0 77120.0 204915.0 ;
      RECT  76415.0 206260.0 77120.0 204915.0 ;
      RECT  77120.0 34100.0 77825.0 35445.0 ;
      RECT  77120.0 36790.0 77825.0 35445.0 ;
      RECT  77120.0 36790.0 77825.0 38135.0 ;
      RECT  77120.0 39480.0 77825.0 38135.0 ;
      RECT  77120.0 39480.0 77825.0 40825.0 ;
      RECT  77120.0 42170.0 77825.0 40825.0 ;
      RECT  77120.0 42170.0 77825.0 43515.0 ;
      RECT  77120.0 44860.0 77825.0 43515.0 ;
      RECT  77120.0 44860.0 77825.0 46205.0 ;
      RECT  77120.0 47550.0 77825.0 46205.0 ;
      RECT  77120.0 47550.0 77825.0 48895.0 ;
      RECT  77120.0 50240.0 77825.0 48895.0 ;
      RECT  77120.0 50240.0 77825.0 51585.0 ;
      RECT  77120.0 52930.0 77825.0 51585.0 ;
      RECT  77120.0 52930.0 77825.0 54275.0 ;
      RECT  77120.0 55620.0 77825.0 54275.0 ;
      RECT  77120.0 55620.0 77825.0 56965.0 ;
      RECT  77120.0 58310.0 77825.0 56965.0 ;
      RECT  77120.0 58310.0 77825.0 59655.0 ;
      RECT  77120.0 61000.0 77825.0 59655.0 ;
      RECT  77120.0 61000.0 77825.0 62345.0 ;
      RECT  77120.0 63690.0 77825.0 62345.0 ;
      RECT  77120.0 63690.0 77825.0 65035.0 ;
      RECT  77120.0 66380.0 77825.0 65035.0 ;
      RECT  77120.0 66380.0 77825.0 67725.0 ;
      RECT  77120.0 69070.0 77825.0 67725.0 ;
      RECT  77120.0 69070.0 77825.0 70415.0 ;
      RECT  77120.0 71760.0 77825.0 70415.0 ;
      RECT  77120.0 71760.0 77825.0 73105.0 ;
      RECT  77120.0 74450.0 77825.0 73105.0 ;
      RECT  77120.0 74450.0 77825.0 75795.0 ;
      RECT  77120.0 77140.0 77825.0 75795.0 ;
      RECT  77120.0 77140.0 77825.0 78485.0 ;
      RECT  77120.0 79830.0 77825.0 78485.0 ;
      RECT  77120.0 79830.0 77825.0 81175.0 ;
      RECT  77120.0 82520.0 77825.0 81175.0 ;
      RECT  77120.0 82520.0 77825.0 83865.0 ;
      RECT  77120.0 85210.0 77825.0 83865.0 ;
      RECT  77120.0 85210.0 77825.0 86555.0 ;
      RECT  77120.0 87900.0 77825.0 86555.0 ;
      RECT  77120.0 87900.0 77825.0 89245.0 ;
      RECT  77120.0 90590.0 77825.0 89245.0 ;
      RECT  77120.0 90590.0 77825.0 91935.0 ;
      RECT  77120.0 93280.0 77825.0 91935.0 ;
      RECT  77120.0 93280.0 77825.0 94625.0 ;
      RECT  77120.0 95970.0 77825.0 94625.0 ;
      RECT  77120.0 95970.0 77825.0 97315.0 ;
      RECT  77120.0 98660.0 77825.0 97315.0 ;
      RECT  77120.0 98660.0 77825.0 100005.0 ;
      RECT  77120.0 101350.0 77825.0 100005.0 ;
      RECT  77120.0 101350.0 77825.0 102695.0 ;
      RECT  77120.0 104040.0 77825.0 102695.0 ;
      RECT  77120.0 104040.0 77825.0 105385.0 ;
      RECT  77120.0 106730.0 77825.0 105385.0 ;
      RECT  77120.0 106730.0 77825.0 108075.0 ;
      RECT  77120.0 109420.0 77825.0 108075.0 ;
      RECT  77120.0 109420.0 77825.0 110765.0 ;
      RECT  77120.0 112110.0 77825.0 110765.0 ;
      RECT  77120.0 112110.0 77825.0 113455.0 ;
      RECT  77120.0 114800.0 77825.0 113455.0 ;
      RECT  77120.0 114800.0 77825.0 116145.0 ;
      RECT  77120.0 117490.0 77825.0 116145.0 ;
      RECT  77120.0 117490.0 77825.0 118835.0 ;
      RECT  77120.0 120180.0 77825.0 118835.0 ;
      RECT  77120.0 120180.0 77825.0 121525.0 ;
      RECT  77120.0 122870.0 77825.0 121525.0 ;
      RECT  77120.0 122870.0 77825.0 124215.0 ;
      RECT  77120.0 125560.0 77825.0 124215.0 ;
      RECT  77120.0 125560.0 77825.0 126905.0 ;
      RECT  77120.0 128250.0 77825.0 126905.0 ;
      RECT  77120.0 128250.0 77825.0 129595.0 ;
      RECT  77120.0 130940.0 77825.0 129595.0 ;
      RECT  77120.0 130940.0 77825.0 132285.0 ;
      RECT  77120.0 133630.0 77825.0 132285.0 ;
      RECT  77120.0 133630.0 77825.0 134975.0 ;
      RECT  77120.0 136320.0 77825.0 134975.0 ;
      RECT  77120.0 136320.0 77825.0 137665.0 ;
      RECT  77120.0 139010.0 77825.0 137665.0 ;
      RECT  77120.0 139010.0 77825.0 140355.0 ;
      RECT  77120.0 141700.0 77825.0 140355.0 ;
      RECT  77120.0 141700.0 77825.0 143045.0 ;
      RECT  77120.0 144390.0 77825.0 143045.0 ;
      RECT  77120.0 144390.0 77825.0 145735.0 ;
      RECT  77120.0 147080.0 77825.0 145735.0 ;
      RECT  77120.0 147080.0 77825.0 148425.0 ;
      RECT  77120.0 149770.0 77825.0 148425.0 ;
      RECT  77120.0 149770.0 77825.0 151115.0 ;
      RECT  77120.0 152460.0 77825.0 151115.0 ;
      RECT  77120.0 152460.0 77825.0 153805.0 ;
      RECT  77120.0 155150.0 77825.0 153805.0 ;
      RECT  77120.0 155150.0 77825.0 156495.0 ;
      RECT  77120.0 157840.0 77825.0 156495.0 ;
      RECT  77120.0 157840.0 77825.0 159185.0 ;
      RECT  77120.0 160530.0 77825.0 159185.0 ;
      RECT  77120.0 160530.0 77825.0 161875.0 ;
      RECT  77120.0 163220.0 77825.0 161875.0 ;
      RECT  77120.0 163220.0 77825.0 164565.0 ;
      RECT  77120.0 165910.0 77825.0 164565.0 ;
      RECT  77120.0 165910.0 77825.0 167255.0 ;
      RECT  77120.0 168600.0 77825.0 167255.0 ;
      RECT  77120.0 168600.0 77825.0 169945.0 ;
      RECT  77120.0 171290.0 77825.0 169945.0 ;
      RECT  77120.0 171290.0 77825.0 172635.0 ;
      RECT  77120.0 173980.0 77825.0 172635.0 ;
      RECT  77120.0 173980.0 77825.0 175325.0 ;
      RECT  77120.0 176670.0 77825.0 175325.0 ;
      RECT  77120.0 176670.0 77825.0 178015.0 ;
      RECT  77120.0 179360.0 77825.0 178015.0 ;
      RECT  77120.0 179360.0 77825.0 180705.0 ;
      RECT  77120.0 182050.0 77825.0 180705.0 ;
      RECT  77120.0 182050.0 77825.0 183395.0 ;
      RECT  77120.0 184740.0 77825.0 183395.0 ;
      RECT  77120.0 184740.0 77825.0 186085.0 ;
      RECT  77120.0 187430.0 77825.0 186085.0 ;
      RECT  77120.0 187430.0 77825.0 188775.0 ;
      RECT  77120.0 190120.0 77825.0 188775.0 ;
      RECT  77120.0 190120.0 77825.0 191465.0 ;
      RECT  77120.0 192810.0 77825.0 191465.0 ;
      RECT  77120.0 192810.0 77825.0 194155.0 ;
      RECT  77120.0 195500.0 77825.0 194155.0 ;
      RECT  77120.0 195500.0 77825.0 196845.0 ;
      RECT  77120.0 198190.0 77825.0 196845.0 ;
      RECT  77120.0 198190.0 77825.0 199535.0 ;
      RECT  77120.0 200880.0 77825.0 199535.0 ;
      RECT  77120.0 200880.0 77825.0 202225.0 ;
      RECT  77120.0 203570.0 77825.0 202225.0 ;
      RECT  77120.0 203570.0 77825.0 204915.0 ;
      RECT  77120.0 206260.0 77825.0 204915.0 ;
      RECT  77825.0 34100.0 78530.0 35445.0 ;
      RECT  77825.0 36790.0 78530.0 35445.0 ;
      RECT  77825.0 36790.0 78530.0 38135.0 ;
      RECT  77825.0 39480.0 78530.0 38135.0 ;
      RECT  77825.0 39480.0 78530.0 40825.0 ;
      RECT  77825.0 42170.0 78530.0 40825.0 ;
      RECT  77825.0 42170.0 78530.0 43515.0 ;
      RECT  77825.0 44860.0 78530.0 43515.0 ;
      RECT  77825.0 44860.0 78530.0 46205.0 ;
      RECT  77825.0 47550.0 78530.0 46205.0 ;
      RECT  77825.0 47550.0 78530.0 48895.0 ;
      RECT  77825.0 50240.0 78530.0 48895.0 ;
      RECT  77825.0 50240.0 78530.0 51585.0 ;
      RECT  77825.0 52930.0 78530.0 51585.0 ;
      RECT  77825.0 52930.0 78530.0 54275.0 ;
      RECT  77825.0 55620.0 78530.0 54275.0 ;
      RECT  77825.0 55620.0 78530.0 56965.0 ;
      RECT  77825.0 58310.0 78530.0 56965.0 ;
      RECT  77825.0 58310.0 78530.0 59655.0 ;
      RECT  77825.0 61000.0 78530.0 59655.0 ;
      RECT  77825.0 61000.0 78530.0 62345.0 ;
      RECT  77825.0 63690.0 78530.0 62345.0 ;
      RECT  77825.0 63690.0 78530.0 65035.0 ;
      RECT  77825.0 66380.0 78530.0 65035.0 ;
      RECT  77825.0 66380.0 78530.0 67725.0 ;
      RECT  77825.0 69070.0 78530.0 67725.0 ;
      RECT  77825.0 69070.0 78530.0 70415.0 ;
      RECT  77825.0 71760.0 78530.0 70415.0 ;
      RECT  77825.0 71760.0 78530.0 73105.0 ;
      RECT  77825.0 74450.0 78530.0 73105.0 ;
      RECT  77825.0 74450.0 78530.0 75795.0 ;
      RECT  77825.0 77140.0 78530.0 75795.0 ;
      RECT  77825.0 77140.0 78530.0 78485.0 ;
      RECT  77825.0 79830.0 78530.0 78485.0 ;
      RECT  77825.0 79830.0 78530.0 81175.0 ;
      RECT  77825.0 82520.0 78530.0 81175.0 ;
      RECT  77825.0 82520.0 78530.0 83865.0 ;
      RECT  77825.0 85210.0 78530.0 83865.0 ;
      RECT  77825.0 85210.0 78530.0 86555.0 ;
      RECT  77825.0 87900.0 78530.0 86555.0 ;
      RECT  77825.0 87900.0 78530.0 89245.0 ;
      RECT  77825.0 90590.0 78530.0 89245.0 ;
      RECT  77825.0 90590.0 78530.0 91935.0 ;
      RECT  77825.0 93280.0 78530.0 91935.0 ;
      RECT  77825.0 93280.0 78530.0 94625.0 ;
      RECT  77825.0 95970.0 78530.0 94625.0 ;
      RECT  77825.0 95970.0 78530.0 97315.0 ;
      RECT  77825.0 98660.0 78530.0 97315.0 ;
      RECT  77825.0 98660.0 78530.0 100005.0 ;
      RECT  77825.0 101350.0 78530.0 100005.0 ;
      RECT  77825.0 101350.0 78530.0 102695.0 ;
      RECT  77825.0 104040.0 78530.0 102695.0 ;
      RECT  77825.0 104040.0 78530.0 105385.0 ;
      RECT  77825.0 106730.0 78530.0 105385.0 ;
      RECT  77825.0 106730.0 78530.0 108075.0 ;
      RECT  77825.0 109420.0 78530.0 108075.0 ;
      RECT  77825.0 109420.0 78530.0 110765.0 ;
      RECT  77825.0 112110.0 78530.0 110765.0 ;
      RECT  77825.0 112110.0 78530.0 113455.0 ;
      RECT  77825.0 114800.0 78530.0 113455.0 ;
      RECT  77825.0 114800.0 78530.0 116145.0 ;
      RECT  77825.0 117490.0 78530.0 116145.0 ;
      RECT  77825.0 117490.0 78530.0 118835.0 ;
      RECT  77825.0 120180.0 78530.0 118835.0 ;
      RECT  77825.0 120180.0 78530.0 121525.0 ;
      RECT  77825.0 122870.0 78530.0 121525.0 ;
      RECT  77825.0 122870.0 78530.0 124215.0 ;
      RECT  77825.0 125560.0 78530.0 124215.0 ;
      RECT  77825.0 125560.0 78530.0 126905.0 ;
      RECT  77825.0 128250.0 78530.0 126905.0 ;
      RECT  77825.0 128250.0 78530.0 129595.0 ;
      RECT  77825.0 130940.0 78530.0 129595.0 ;
      RECT  77825.0 130940.0 78530.0 132285.0 ;
      RECT  77825.0 133630.0 78530.0 132285.0 ;
      RECT  77825.0 133630.0 78530.0 134975.0 ;
      RECT  77825.0 136320.0 78530.0 134975.0 ;
      RECT  77825.0 136320.0 78530.0 137665.0 ;
      RECT  77825.0 139010.0 78530.0 137665.0 ;
      RECT  77825.0 139010.0 78530.0 140355.0 ;
      RECT  77825.0 141700.0 78530.0 140355.0 ;
      RECT  77825.0 141700.0 78530.0 143045.0 ;
      RECT  77825.0 144390.0 78530.0 143045.0 ;
      RECT  77825.0 144390.0 78530.0 145735.0 ;
      RECT  77825.0 147080.0 78530.0 145735.0 ;
      RECT  77825.0 147080.0 78530.0 148425.0 ;
      RECT  77825.0 149770.0 78530.0 148425.0 ;
      RECT  77825.0 149770.0 78530.0 151115.0 ;
      RECT  77825.0 152460.0 78530.0 151115.0 ;
      RECT  77825.0 152460.0 78530.0 153805.0 ;
      RECT  77825.0 155150.0 78530.0 153805.0 ;
      RECT  77825.0 155150.0 78530.0 156495.0 ;
      RECT  77825.0 157840.0 78530.0 156495.0 ;
      RECT  77825.0 157840.0 78530.0 159185.0 ;
      RECT  77825.0 160530.0 78530.0 159185.0 ;
      RECT  77825.0 160530.0 78530.0 161875.0 ;
      RECT  77825.0 163220.0 78530.0 161875.0 ;
      RECT  77825.0 163220.0 78530.0 164565.0 ;
      RECT  77825.0 165910.0 78530.0 164565.0 ;
      RECT  77825.0 165910.0 78530.0 167255.0 ;
      RECT  77825.0 168600.0 78530.0 167255.0 ;
      RECT  77825.0 168600.0 78530.0 169945.0 ;
      RECT  77825.0 171290.0 78530.0 169945.0 ;
      RECT  77825.0 171290.0 78530.0 172635.0 ;
      RECT  77825.0 173980.0 78530.0 172635.0 ;
      RECT  77825.0 173980.0 78530.0 175325.0 ;
      RECT  77825.0 176670.0 78530.0 175325.0 ;
      RECT  77825.0 176670.0 78530.0 178015.0 ;
      RECT  77825.0 179360.0 78530.0 178015.0 ;
      RECT  77825.0 179360.0 78530.0 180705.0 ;
      RECT  77825.0 182050.0 78530.0 180705.0 ;
      RECT  77825.0 182050.0 78530.0 183395.0 ;
      RECT  77825.0 184740.0 78530.0 183395.0 ;
      RECT  77825.0 184740.0 78530.0 186085.0 ;
      RECT  77825.0 187430.0 78530.0 186085.0 ;
      RECT  77825.0 187430.0 78530.0 188775.0 ;
      RECT  77825.0 190120.0 78530.0 188775.0 ;
      RECT  77825.0 190120.0 78530.0 191465.0 ;
      RECT  77825.0 192810.0 78530.0 191465.0 ;
      RECT  77825.0 192810.0 78530.0 194155.0 ;
      RECT  77825.0 195500.0 78530.0 194155.0 ;
      RECT  77825.0 195500.0 78530.0 196845.0 ;
      RECT  77825.0 198190.0 78530.0 196845.0 ;
      RECT  77825.0 198190.0 78530.0 199535.0 ;
      RECT  77825.0 200880.0 78530.0 199535.0 ;
      RECT  77825.0 200880.0 78530.0 202225.0 ;
      RECT  77825.0 203570.0 78530.0 202225.0 ;
      RECT  77825.0 203570.0 78530.0 204915.0 ;
      RECT  77825.0 206260.0 78530.0 204915.0 ;
      RECT  78530.0 34100.0 79235.0 35445.0 ;
      RECT  78530.0 36790.0 79235.0 35445.0 ;
      RECT  78530.0 36790.0 79235.0 38135.0 ;
      RECT  78530.0 39480.0 79235.0 38135.0 ;
      RECT  78530.0 39480.0 79235.0 40825.0 ;
      RECT  78530.0 42170.0 79235.0 40825.0 ;
      RECT  78530.0 42170.0 79235.0 43515.0 ;
      RECT  78530.0 44860.0 79235.0 43515.0 ;
      RECT  78530.0 44860.0 79235.0 46205.0 ;
      RECT  78530.0 47550.0 79235.0 46205.0 ;
      RECT  78530.0 47550.0 79235.0 48895.0 ;
      RECT  78530.0 50240.0 79235.0 48895.0 ;
      RECT  78530.0 50240.0 79235.0 51585.0 ;
      RECT  78530.0 52930.0 79235.0 51585.0 ;
      RECT  78530.0 52930.0 79235.0 54275.0 ;
      RECT  78530.0 55620.0 79235.0 54275.0 ;
      RECT  78530.0 55620.0 79235.0 56965.0 ;
      RECT  78530.0 58310.0 79235.0 56965.0 ;
      RECT  78530.0 58310.0 79235.0 59655.0 ;
      RECT  78530.0 61000.0 79235.0 59655.0 ;
      RECT  78530.0 61000.0 79235.0 62345.0 ;
      RECT  78530.0 63690.0 79235.0 62345.0 ;
      RECT  78530.0 63690.0 79235.0 65035.0 ;
      RECT  78530.0 66380.0 79235.0 65035.0 ;
      RECT  78530.0 66380.0 79235.0 67725.0 ;
      RECT  78530.0 69070.0 79235.0 67725.0 ;
      RECT  78530.0 69070.0 79235.0 70415.0 ;
      RECT  78530.0 71760.0 79235.0 70415.0 ;
      RECT  78530.0 71760.0 79235.0 73105.0 ;
      RECT  78530.0 74450.0 79235.0 73105.0 ;
      RECT  78530.0 74450.0 79235.0 75795.0 ;
      RECT  78530.0 77140.0 79235.0 75795.0 ;
      RECT  78530.0 77140.0 79235.0 78485.0 ;
      RECT  78530.0 79830.0 79235.0 78485.0 ;
      RECT  78530.0 79830.0 79235.0 81175.0 ;
      RECT  78530.0 82520.0 79235.0 81175.0 ;
      RECT  78530.0 82520.0 79235.0 83865.0 ;
      RECT  78530.0 85210.0 79235.0 83865.0 ;
      RECT  78530.0 85210.0 79235.0 86555.0 ;
      RECT  78530.0 87900.0 79235.0 86555.0 ;
      RECT  78530.0 87900.0 79235.0 89245.0 ;
      RECT  78530.0 90590.0 79235.0 89245.0 ;
      RECT  78530.0 90590.0 79235.0 91935.0 ;
      RECT  78530.0 93280.0 79235.0 91935.0 ;
      RECT  78530.0 93280.0 79235.0 94625.0 ;
      RECT  78530.0 95970.0 79235.0 94625.0 ;
      RECT  78530.0 95970.0 79235.0 97315.0 ;
      RECT  78530.0 98660.0 79235.0 97315.0 ;
      RECT  78530.0 98660.0 79235.0 100005.0 ;
      RECT  78530.0 101350.0 79235.0 100005.0 ;
      RECT  78530.0 101350.0 79235.0 102695.0 ;
      RECT  78530.0 104040.0 79235.0 102695.0 ;
      RECT  78530.0 104040.0 79235.0 105385.0 ;
      RECT  78530.0 106730.0 79235.0 105385.0 ;
      RECT  78530.0 106730.0 79235.0 108075.0 ;
      RECT  78530.0 109420.0 79235.0 108075.0 ;
      RECT  78530.0 109420.0 79235.0 110765.0 ;
      RECT  78530.0 112110.0 79235.0 110765.0 ;
      RECT  78530.0 112110.0 79235.0 113455.0 ;
      RECT  78530.0 114800.0 79235.0 113455.0 ;
      RECT  78530.0 114800.0 79235.0 116145.0 ;
      RECT  78530.0 117490.0 79235.0 116145.0 ;
      RECT  78530.0 117490.0 79235.0 118835.0 ;
      RECT  78530.0 120180.0 79235.0 118835.0 ;
      RECT  78530.0 120180.0 79235.0 121525.0 ;
      RECT  78530.0 122870.0 79235.0 121525.0 ;
      RECT  78530.0 122870.0 79235.0 124215.0 ;
      RECT  78530.0 125560.0 79235.0 124215.0 ;
      RECT  78530.0 125560.0 79235.0 126905.0 ;
      RECT  78530.0 128250.0 79235.0 126905.0 ;
      RECT  78530.0 128250.0 79235.0 129595.0 ;
      RECT  78530.0 130940.0 79235.0 129595.0 ;
      RECT  78530.0 130940.0 79235.0 132285.0 ;
      RECT  78530.0 133630.0 79235.0 132285.0 ;
      RECT  78530.0 133630.0 79235.0 134975.0 ;
      RECT  78530.0 136320.0 79235.0 134975.0 ;
      RECT  78530.0 136320.0 79235.0 137665.0 ;
      RECT  78530.0 139010.0 79235.0 137665.0 ;
      RECT  78530.0 139010.0 79235.0 140355.0 ;
      RECT  78530.0 141700.0 79235.0 140355.0 ;
      RECT  78530.0 141700.0 79235.0 143045.0 ;
      RECT  78530.0 144390.0 79235.0 143045.0 ;
      RECT  78530.0 144390.0 79235.0 145735.0 ;
      RECT  78530.0 147080.0 79235.0 145735.0 ;
      RECT  78530.0 147080.0 79235.0 148425.0 ;
      RECT  78530.0 149770.0 79235.0 148425.0 ;
      RECT  78530.0 149770.0 79235.0 151115.0 ;
      RECT  78530.0 152460.0 79235.0 151115.0 ;
      RECT  78530.0 152460.0 79235.0 153805.0 ;
      RECT  78530.0 155150.0 79235.0 153805.0 ;
      RECT  78530.0 155150.0 79235.0 156495.0 ;
      RECT  78530.0 157840.0 79235.0 156495.0 ;
      RECT  78530.0 157840.0 79235.0 159185.0 ;
      RECT  78530.0 160530.0 79235.0 159185.0 ;
      RECT  78530.0 160530.0 79235.0 161875.0 ;
      RECT  78530.0 163220.0 79235.0 161875.0 ;
      RECT  78530.0 163220.0 79235.0 164565.0 ;
      RECT  78530.0 165910.0 79235.0 164565.0 ;
      RECT  78530.0 165910.0 79235.0 167255.0 ;
      RECT  78530.0 168600.0 79235.0 167255.0 ;
      RECT  78530.0 168600.0 79235.0 169945.0 ;
      RECT  78530.0 171290.0 79235.0 169945.0 ;
      RECT  78530.0 171290.0 79235.0 172635.0 ;
      RECT  78530.0 173980.0 79235.0 172635.0 ;
      RECT  78530.0 173980.0 79235.0 175325.0 ;
      RECT  78530.0 176670.0 79235.0 175325.0 ;
      RECT  78530.0 176670.0 79235.0 178015.0 ;
      RECT  78530.0 179360.0 79235.0 178015.0 ;
      RECT  78530.0 179360.0 79235.0 180705.0 ;
      RECT  78530.0 182050.0 79235.0 180705.0 ;
      RECT  78530.0 182050.0 79235.0 183395.0 ;
      RECT  78530.0 184740.0 79235.0 183395.0 ;
      RECT  78530.0 184740.0 79235.0 186085.0 ;
      RECT  78530.0 187430.0 79235.0 186085.0 ;
      RECT  78530.0 187430.0 79235.0 188775.0 ;
      RECT  78530.0 190120.0 79235.0 188775.0 ;
      RECT  78530.0 190120.0 79235.0 191465.0 ;
      RECT  78530.0 192810.0 79235.0 191465.0 ;
      RECT  78530.0 192810.0 79235.0 194155.0 ;
      RECT  78530.0 195500.0 79235.0 194155.0 ;
      RECT  78530.0 195500.0 79235.0 196845.0 ;
      RECT  78530.0 198190.0 79235.0 196845.0 ;
      RECT  78530.0 198190.0 79235.0 199535.0 ;
      RECT  78530.0 200880.0 79235.0 199535.0 ;
      RECT  78530.0 200880.0 79235.0 202225.0 ;
      RECT  78530.0 203570.0 79235.0 202225.0 ;
      RECT  78530.0 203570.0 79235.0 204915.0 ;
      RECT  78530.0 206260.0 79235.0 204915.0 ;
      RECT  79235.0 34100.0 79940.0 35445.0 ;
      RECT  79235.0 36790.0 79940.0 35445.0 ;
      RECT  79235.0 36790.0 79940.0 38135.0 ;
      RECT  79235.0 39480.0 79940.0 38135.0 ;
      RECT  79235.0 39480.0 79940.0 40825.0 ;
      RECT  79235.0 42170.0 79940.0 40825.0 ;
      RECT  79235.0 42170.0 79940.0 43515.0 ;
      RECT  79235.0 44860.0 79940.0 43515.0 ;
      RECT  79235.0 44860.0 79940.0 46205.0 ;
      RECT  79235.0 47550.0 79940.0 46205.0 ;
      RECT  79235.0 47550.0 79940.0 48895.0 ;
      RECT  79235.0 50240.0 79940.0 48895.0 ;
      RECT  79235.0 50240.0 79940.0 51585.0 ;
      RECT  79235.0 52930.0 79940.0 51585.0 ;
      RECT  79235.0 52930.0 79940.0 54275.0 ;
      RECT  79235.0 55620.0 79940.0 54275.0 ;
      RECT  79235.0 55620.0 79940.0 56965.0 ;
      RECT  79235.0 58310.0 79940.0 56965.0 ;
      RECT  79235.0 58310.0 79940.0 59655.0 ;
      RECT  79235.0 61000.0 79940.0 59655.0 ;
      RECT  79235.0 61000.0 79940.0 62345.0 ;
      RECT  79235.0 63690.0 79940.0 62345.0 ;
      RECT  79235.0 63690.0 79940.0 65035.0 ;
      RECT  79235.0 66380.0 79940.0 65035.0 ;
      RECT  79235.0 66380.0 79940.0 67725.0 ;
      RECT  79235.0 69070.0 79940.0 67725.0 ;
      RECT  79235.0 69070.0 79940.0 70415.0 ;
      RECT  79235.0 71760.0 79940.0 70415.0 ;
      RECT  79235.0 71760.0 79940.0 73105.0 ;
      RECT  79235.0 74450.0 79940.0 73105.0 ;
      RECT  79235.0 74450.0 79940.0 75795.0 ;
      RECT  79235.0 77140.0 79940.0 75795.0 ;
      RECT  79235.0 77140.0 79940.0 78485.0 ;
      RECT  79235.0 79830.0 79940.0 78485.0 ;
      RECT  79235.0 79830.0 79940.0 81175.0 ;
      RECT  79235.0 82520.0 79940.0 81175.0 ;
      RECT  79235.0 82520.0 79940.0 83865.0 ;
      RECT  79235.0 85210.0 79940.0 83865.0 ;
      RECT  79235.0 85210.0 79940.0 86555.0 ;
      RECT  79235.0 87900.0 79940.0 86555.0 ;
      RECT  79235.0 87900.0 79940.0 89245.0 ;
      RECT  79235.0 90590.0 79940.0 89245.0 ;
      RECT  79235.0 90590.0 79940.0 91935.0 ;
      RECT  79235.0 93280.0 79940.0 91935.0 ;
      RECT  79235.0 93280.0 79940.0 94625.0 ;
      RECT  79235.0 95970.0 79940.0 94625.0 ;
      RECT  79235.0 95970.0 79940.0 97315.0 ;
      RECT  79235.0 98660.0 79940.0 97315.0 ;
      RECT  79235.0 98660.0 79940.0 100005.0 ;
      RECT  79235.0 101350.0 79940.0 100005.0 ;
      RECT  79235.0 101350.0 79940.0 102695.0 ;
      RECT  79235.0 104040.0 79940.0 102695.0 ;
      RECT  79235.0 104040.0 79940.0 105385.0 ;
      RECT  79235.0 106730.0 79940.0 105385.0 ;
      RECT  79235.0 106730.0 79940.0 108075.0 ;
      RECT  79235.0 109420.0 79940.0 108075.0 ;
      RECT  79235.0 109420.0 79940.0 110765.0 ;
      RECT  79235.0 112110.0 79940.0 110765.0 ;
      RECT  79235.0 112110.0 79940.0 113455.0 ;
      RECT  79235.0 114800.0 79940.0 113455.0 ;
      RECT  79235.0 114800.0 79940.0 116145.0 ;
      RECT  79235.0 117490.0 79940.0 116145.0 ;
      RECT  79235.0 117490.0 79940.0 118835.0 ;
      RECT  79235.0 120180.0 79940.0 118835.0 ;
      RECT  79235.0 120180.0 79940.0 121525.0 ;
      RECT  79235.0 122870.0 79940.0 121525.0 ;
      RECT  79235.0 122870.0 79940.0 124215.0 ;
      RECT  79235.0 125560.0 79940.0 124215.0 ;
      RECT  79235.0 125560.0 79940.0 126905.0 ;
      RECT  79235.0 128250.0 79940.0 126905.0 ;
      RECT  79235.0 128250.0 79940.0 129595.0 ;
      RECT  79235.0 130940.0 79940.0 129595.0 ;
      RECT  79235.0 130940.0 79940.0 132285.0 ;
      RECT  79235.0 133630.0 79940.0 132285.0 ;
      RECT  79235.0 133630.0 79940.0 134975.0 ;
      RECT  79235.0 136320.0 79940.0 134975.0 ;
      RECT  79235.0 136320.0 79940.0 137665.0 ;
      RECT  79235.0 139010.0 79940.0 137665.0 ;
      RECT  79235.0 139010.0 79940.0 140355.0 ;
      RECT  79235.0 141700.0 79940.0 140355.0 ;
      RECT  79235.0 141700.0 79940.0 143045.0 ;
      RECT  79235.0 144390.0 79940.0 143045.0 ;
      RECT  79235.0 144390.0 79940.0 145735.0 ;
      RECT  79235.0 147080.0 79940.0 145735.0 ;
      RECT  79235.0 147080.0 79940.0 148425.0 ;
      RECT  79235.0 149770.0 79940.0 148425.0 ;
      RECT  79235.0 149770.0 79940.0 151115.0 ;
      RECT  79235.0 152460.0 79940.0 151115.0 ;
      RECT  79235.0 152460.0 79940.0 153805.0 ;
      RECT  79235.0 155150.0 79940.0 153805.0 ;
      RECT  79235.0 155150.0 79940.0 156495.0 ;
      RECT  79235.0 157840.0 79940.0 156495.0 ;
      RECT  79235.0 157840.0 79940.0 159185.0 ;
      RECT  79235.0 160530.0 79940.0 159185.0 ;
      RECT  79235.0 160530.0 79940.0 161875.0 ;
      RECT  79235.0 163220.0 79940.0 161875.0 ;
      RECT  79235.0 163220.0 79940.0 164565.0 ;
      RECT  79235.0 165910.0 79940.0 164565.0 ;
      RECT  79235.0 165910.0 79940.0 167255.0 ;
      RECT  79235.0 168600.0 79940.0 167255.0 ;
      RECT  79235.0 168600.0 79940.0 169945.0 ;
      RECT  79235.0 171290.0 79940.0 169945.0 ;
      RECT  79235.0 171290.0 79940.0 172635.0 ;
      RECT  79235.0 173980.0 79940.0 172635.0 ;
      RECT  79235.0 173980.0 79940.0 175325.0 ;
      RECT  79235.0 176670.0 79940.0 175325.0 ;
      RECT  79235.0 176670.0 79940.0 178015.0 ;
      RECT  79235.0 179360.0 79940.0 178015.0 ;
      RECT  79235.0 179360.0 79940.0 180705.0 ;
      RECT  79235.0 182050.0 79940.0 180705.0 ;
      RECT  79235.0 182050.0 79940.0 183395.0 ;
      RECT  79235.0 184740.0 79940.0 183395.0 ;
      RECT  79235.0 184740.0 79940.0 186085.0 ;
      RECT  79235.0 187430.0 79940.0 186085.0 ;
      RECT  79235.0 187430.0 79940.0 188775.0 ;
      RECT  79235.0 190120.0 79940.0 188775.0 ;
      RECT  79235.0 190120.0 79940.0 191465.0 ;
      RECT  79235.0 192810.0 79940.0 191465.0 ;
      RECT  79235.0 192810.0 79940.0 194155.0 ;
      RECT  79235.0 195500.0 79940.0 194155.0 ;
      RECT  79235.0 195500.0 79940.0 196845.0 ;
      RECT  79235.0 198190.0 79940.0 196845.0 ;
      RECT  79235.0 198190.0 79940.0 199535.0 ;
      RECT  79235.0 200880.0 79940.0 199535.0 ;
      RECT  79235.0 200880.0 79940.0 202225.0 ;
      RECT  79235.0 203570.0 79940.0 202225.0 ;
      RECT  79235.0 203570.0 79940.0 204915.0 ;
      RECT  79235.0 206260.0 79940.0 204915.0 ;
      RECT  79940.0 34100.0 80645.0 35445.0 ;
      RECT  79940.0 36790.0 80645.0 35445.0 ;
      RECT  79940.0 36790.0 80645.0 38135.0 ;
      RECT  79940.0 39480.0 80645.0 38135.0 ;
      RECT  79940.0 39480.0 80645.0 40825.0 ;
      RECT  79940.0 42170.0 80645.0 40825.0 ;
      RECT  79940.0 42170.0 80645.0 43515.0 ;
      RECT  79940.0 44860.0 80645.0 43515.0 ;
      RECT  79940.0 44860.0 80645.0 46205.0 ;
      RECT  79940.0 47550.0 80645.0 46205.0 ;
      RECT  79940.0 47550.0 80645.0 48895.0 ;
      RECT  79940.0 50240.0 80645.0 48895.0 ;
      RECT  79940.0 50240.0 80645.0 51585.0 ;
      RECT  79940.0 52930.0 80645.0 51585.0 ;
      RECT  79940.0 52930.0 80645.0 54275.0 ;
      RECT  79940.0 55620.0 80645.0 54275.0 ;
      RECT  79940.0 55620.0 80645.0 56965.0 ;
      RECT  79940.0 58310.0 80645.0 56965.0 ;
      RECT  79940.0 58310.0 80645.0 59655.0 ;
      RECT  79940.0 61000.0 80645.0 59655.0 ;
      RECT  79940.0 61000.0 80645.0 62345.0 ;
      RECT  79940.0 63690.0 80645.0 62345.0 ;
      RECT  79940.0 63690.0 80645.0 65035.0 ;
      RECT  79940.0 66380.0 80645.0 65035.0 ;
      RECT  79940.0 66380.0 80645.0 67725.0 ;
      RECT  79940.0 69070.0 80645.0 67725.0 ;
      RECT  79940.0 69070.0 80645.0 70415.0 ;
      RECT  79940.0 71760.0 80645.0 70415.0 ;
      RECT  79940.0 71760.0 80645.0 73105.0 ;
      RECT  79940.0 74450.0 80645.0 73105.0 ;
      RECT  79940.0 74450.0 80645.0 75795.0 ;
      RECT  79940.0 77140.0 80645.0 75795.0 ;
      RECT  79940.0 77140.0 80645.0 78485.0 ;
      RECT  79940.0 79830.0 80645.0 78485.0 ;
      RECT  79940.0 79830.0 80645.0 81175.0 ;
      RECT  79940.0 82520.0 80645.0 81175.0 ;
      RECT  79940.0 82520.0 80645.0 83865.0 ;
      RECT  79940.0 85210.0 80645.0 83865.0 ;
      RECT  79940.0 85210.0 80645.0 86555.0 ;
      RECT  79940.0 87900.0 80645.0 86555.0 ;
      RECT  79940.0 87900.0 80645.0 89245.0 ;
      RECT  79940.0 90590.0 80645.0 89245.0 ;
      RECT  79940.0 90590.0 80645.0 91935.0 ;
      RECT  79940.0 93280.0 80645.0 91935.0 ;
      RECT  79940.0 93280.0 80645.0 94625.0 ;
      RECT  79940.0 95970.0 80645.0 94625.0 ;
      RECT  79940.0 95970.0 80645.0 97315.0 ;
      RECT  79940.0 98660.0 80645.0 97315.0 ;
      RECT  79940.0 98660.0 80645.0 100005.0 ;
      RECT  79940.0 101350.0 80645.0 100005.0 ;
      RECT  79940.0 101350.0 80645.0 102695.0 ;
      RECT  79940.0 104040.0 80645.0 102695.0 ;
      RECT  79940.0 104040.0 80645.0 105385.0 ;
      RECT  79940.0 106730.0 80645.0 105385.0 ;
      RECT  79940.0 106730.0 80645.0 108075.0 ;
      RECT  79940.0 109420.0 80645.0 108075.0 ;
      RECT  79940.0 109420.0 80645.0 110765.0 ;
      RECT  79940.0 112110.0 80645.0 110765.0 ;
      RECT  79940.0 112110.0 80645.0 113455.0 ;
      RECT  79940.0 114800.0 80645.0 113455.0 ;
      RECT  79940.0 114800.0 80645.0 116145.0 ;
      RECT  79940.0 117490.0 80645.0 116145.0 ;
      RECT  79940.0 117490.0 80645.0 118835.0 ;
      RECT  79940.0 120180.0 80645.0 118835.0 ;
      RECT  79940.0 120180.0 80645.0 121525.0 ;
      RECT  79940.0 122870.0 80645.0 121525.0 ;
      RECT  79940.0 122870.0 80645.0 124215.0 ;
      RECT  79940.0 125560.0 80645.0 124215.0 ;
      RECT  79940.0 125560.0 80645.0 126905.0 ;
      RECT  79940.0 128250.0 80645.0 126905.0 ;
      RECT  79940.0 128250.0 80645.0 129595.0 ;
      RECT  79940.0 130940.0 80645.0 129595.0 ;
      RECT  79940.0 130940.0 80645.0 132285.0 ;
      RECT  79940.0 133630.0 80645.0 132285.0 ;
      RECT  79940.0 133630.0 80645.0 134975.0 ;
      RECT  79940.0 136320.0 80645.0 134975.0 ;
      RECT  79940.0 136320.0 80645.0 137665.0 ;
      RECT  79940.0 139010.0 80645.0 137665.0 ;
      RECT  79940.0 139010.0 80645.0 140355.0 ;
      RECT  79940.0 141700.0 80645.0 140355.0 ;
      RECT  79940.0 141700.0 80645.0 143045.0 ;
      RECT  79940.0 144390.0 80645.0 143045.0 ;
      RECT  79940.0 144390.0 80645.0 145735.0 ;
      RECT  79940.0 147080.0 80645.0 145735.0 ;
      RECT  79940.0 147080.0 80645.0 148425.0 ;
      RECT  79940.0 149770.0 80645.0 148425.0 ;
      RECT  79940.0 149770.0 80645.0 151115.0 ;
      RECT  79940.0 152460.0 80645.0 151115.0 ;
      RECT  79940.0 152460.0 80645.0 153805.0 ;
      RECT  79940.0 155150.0 80645.0 153805.0 ;
      RECT  79940.0 155150.0 80645.0 156495.0 ;
      RECT  79940.0 157840.0 80645.0 156495.0 ;
      RECT  79940.0 157840.0 80645.0 159185.0 ;
      RECT  79940.0 160530.0 80645.0 159185.0 ;
      RECT  79940.0 160530.0 80645.0 161875.0 ;
      RECT  79940.0 163220.0 80645.0 161875.0 ;
      RECT  79940.0 163220.0 80645.0 164565.0 ;
      RECT  79940.0 165910.0 80645.0 164565.0 ;
      RECT  79940.0 165910.0 80645.0 167255.0 ;
      RECT  79940.0 168600.0 80645.0 167255.0 ;
      RECT  79940.0 168600.0 80645.0 169945.0 ;
      RECT  79940.0 171290.0 80645.0 169945.0 ;
      RECT  79940.0 171290.0 80645.0 172635.0 ;
      RECT  79940.0 173980.0 80645.0 172635.0 ;
      RECT  79940.0 173980.0 80645.0 175325.0 ;
      RECT  79940.0 176670.0 80645.0 175325.0 ;
      RECT  79940.0 176670.0 80645.0 178015.0 ;
      RECT  79940.0 179360.0 80645.0 178015.0 ;
      RECT  79940.0 179360.0 80645.0 180705.0 ;
      RECT  79940.0 182050.0 80645.0 180705.0 ;
      RECT  79940.0 182050.0 80645.0 183395.0 ;
      RECT  79940.0 184740.0 80645.0 183395.0 ;
      RECT  79940.0 184740.0 80645.0 186085.0 ;
      RECT  79940.0 187430.0 80645.0 186085.0 ;
      RECT  79940.0 187430.0 80645.0 188775.0 ;
      RECT  79940.0 190120.0 80645.0 188775.0 ;
      RECT  79940.0 190120.0 80645.0 191465.0 ;
      RECT  79940.0 192810.0 80645.0 191465.0 ;
      RECT  79940.0 192810.0 80645.0 194155.0 ;
      RECT  79940.0 195500.0 80645.0 194155.0 ;
      RECT  79940.0 195500.0 80645.0 196845.0 ;
      RECT  79940.0 198190.0 80645.0 196845.0 ;
      RECT  79940.0 198190.0 80645.0 199535.0 ;
      RECT  79940.0 200880.0 80645.0 199535.0 ;
      RECT  79940.0 200880.0 80645.0 202225.0 ;
      RECT  79940.0 203570.0 80645.0 202225.0 ;
      RECT  79940.0 203570.0 80645.0 204915.0 ;
      RECT  79940.0 206260.0 80645.0 204915.0 ;
      RECT  80645.0 34100.0 81350.0 35445.0 ;
      RECT  80645.0 36790.0 81350.0 35445.0 ;
      RECT  80645.0 36790.0 81350.0 38135.0 ;
      RECT  80645.0 39480.0 81350.0 38135.0 ;
      RECT  80645.0 39480.0 81350.0 40825.0 ;
      RECT  80645.0 42170.0 81350.0 40825.0 ;
      RECT  80645.0 42170.0 81350.0 43515.0 ;
      RECT  80645.0 44860.0 81350.0 43515.0 ;
      RECT  80645.0 44860.0 81350.0 46205.0 ;
      RECT  80645.0 47550.0 81350.0 46205.0 ;
      RECT  80645.0 47550.0 81350.0 48895.0 ;
      RECT  80645.0 50240.0 81350.0 48895.0 ;
      RECT  80645.0 50240.0 81350.0 51585.0 ;
      RECT  80645.0 52930.0 81350.0 51585.0 ;
      RECT  80645.0 52930.0 81350.0 54275.0 ;
      RECT  80645.0 55620.0 81350.0 54275.0 ;
      RECT  80645.0 55620.0 81350.0 56965.0 ;
      RECT  80645.0 58310.0 81350.0 56965.0 ;
      RECT  80645.0 58310.0 81350.0 59655.0 ;
      RECT  80645.0 61000.0 81350.0 59655.0 ;
      RECT  80645.0 61000.0 81350.0 62345.0 ;
      RECT  80645.0 63690.0 81350.0 62345.0 ;
      RECT  80645.0 63690.0 81350.0 65035.0 ;
      RECT  80645.0 66380.0 81350.0 65035.0 ;
      RECT  80645.0 66380.0 81350.0 67725.0 ;
      RECT  80645.0 69070.0 81350.0 67725.0 ;
      RECT  80645.0 69070.0 81350.0 70415.0 ;
      RECT  80645.0 71760.0 81350.0 70415.0 ;
      RECT  80645.0 71760.0 81350.0 73105.0 ;
      RECT  80645.0 74450.0 81350.0 73105.0 ;
      RECT  80645.0 74450.0 81350.0 75795.0 ;
      RECT  80645.0 77140.0 81350.0 75795.0 ;
      RECT  80645.0 77140.0 81350.0 78485.0 ;
      RECT  80645.0 79830.0 81350.0 78485.0 ;
      RECT  80645.0 79830.0 81350.0 81175.0 ;
      RECT  80645.0 82520.0 81350.0 81175.0 ;
      RECT  80645.0 82520.0 81350.0 83865.0 ;
      RECT  80645.0 85210.0 81350.0 83865.0 ;
      RECT  80645.0 85210.0 81350.0 86555.0 ;
      RECT  80645.0 87900.0 81350.0 86555.0 ;
      RECT  80645.0 87900.0 81350.0 89245.0 ;
      RECT  80645.0 90590.0 81350.0 89245.0 ;
      RECT  80645.0 90590.0 81350.0 91935.0 ;
      RECT  80645.0 93280.0 81350.0 91935.0 ;
      RECT  80645.0 93280.0 81350.0 94625.0 ;
      RECT  80645.0 95970.0 81350.0 94625.0 ;
      RECT  80645.0 95970.0 81350.0 97315.0 ;
      RECT  80645.0 98660.0 81350.0 97315.0 ;
      RECT  80645.0 98660.0 81350.0 100005.0 ;
      RECT  80645.0 101350.0 81350.0 100005.0 ;
      RECT  80645.0 101350.0 81350.0 102695.0 ;
      RECT  80645.0 104040.0 81350.0 102695.0 ;
      RECT  80645.0 104040.0 81350.0 105385.0 ;
      RECT  80645.0 106730.0 81350.0 105385.0 ;
      RECT  80645.0 106730.0 81350.0 108075.0 ;
      RECT  80645.0 109420.0 81350.0 108075.0 ;
      RECT  80645.0 109420.0 81350.0 110765.0 ;
      RECT  80645.0 112110.0 81350.0 110765.0 ;
      RECT  80645.0 112110.0 81350.0 113455.0 ;
      RECT  80645.0 114800.0 81350.0 113455.0 ;
      RECT  80645.0 114800.0 81350.0 116145.0 ;
      RECT  80645.0 117490.0 81350.0 116145.0 ;
      RECT  80645.0 117490.0 81350.0 118835.0 ;
      RECT  80645.0 120180.0 81350.0 118835.0 ;
      RECT  80645.0 120180.0 81350.0 121525.0 ;
      RECT  80645.0 122870.0 81350.0 121525.0 ;
      RECT  80645.0 122870.0 81350.0 124215.0 ;
      RECT  80645.0 125560.0 81350.0 124215.0 ;
      RECT  80645.0 125560.0 81350.0 126905.0 ;
      RECT  80645.0 128250.0 81350.0 126905.0 ;
      RECT  80645.0 128250.0 81350.0 129595.0 ;
      RECT  80645.0 130940.0 81350.0 129595.0 ;
      RECT  80645.0 130940.0 81350.0 132285.0 ;
      RECT  80645.0 133630.0 81350.0 132285.0 ;
      RECT  80645.0 133630.0 81350.0 134975.0 ;
      RECT  80645.0 136320.0 81350.0 134975.0 ;
      RECT  80645.0 136320.0 81350.0 137665.0 ;
      RECT  80645.0 139010.0 81350.0 137665.0 ;
      RECT  80645.0 139010.0 81350.0 140355.0 ;
      RECT  80645.0 141700.0 81350.0 140355.0 ;
      RECT  80645.0 141700.0 81350.0 143045.0 ;
      RECT  80645.0 144390.0 81350.0 143045.0 ;
      RECT  80645.0 144390.0 81350.0 145735.0 ;
      RECT  80645.0 147080.0 81350.0 145735.0 ;
      RECT  80645.0 147080.0 81350.0 148425.0 ;
      RECT  80645.0 149770.0 81350.0 148425.0 ;
      RECT  80645.0 149770.0 81350.0 151115.0 ;
      RECT  80645.0 152460.0 81350.0 151115.0 ;
      RECT  80645.0 152460.0 81350.0 153805.0 ;
      RECT  80645.0 155150.0 81350.0 153805.0 ;
      RECT  80645.0 155150.0 81350.0 156495.0 ;
      RECT  80645.0 157840.0 81350.0 156495.0 ;
      RECT  80645.0 157840.0 81350.0 159185.0 ;
      RECT  80645.0 160530.0 81350.0 159185.0 ;
      RECT  80645.0 160530.0 81350.0 161875.0 ;
      RECT  80645.0 163220.0 81350.0 161875.0 ;
      RECT  80645.0 163220.0 81350.0 164565.0 ;
      RECT  80645.0 165910.0 81350.0 164565.0 ;
      RECT  80645.0 165910.0 81350.0 167255.0 ;
      RECT  80645.0 168600.0 81350.0 167255.0 ;
      RECT  80645.0 168600.0 81350.0 169945.0 ;
      RECT  80645.0 171290.0 81350.0 169945.0 ;
      RECT  80645.0 171290.0 81350.0 172635.0 ;
      RECT  80645.0 173980.0 81350.0 172635.0 ;
      RECT  80645.0 173980.0 81350.0 175325.0 ;
      RECT  80645.0 176670.0 81350.0 175325.0 ;
      RECT  80645.0 176670.0 81350.0 178015.0 ;
      RECT  80645.0 179360.0 81350.0 178015.0 ;
      RECT  80645.0 179360.0 81350.0 180705.0 ;
      RECT  80645.0 182050.0 81350.0 180705.0 ;
      RECT  80645.0 182050.0 81350.0 183395.0 ;
      RECT  80645.0 184740.0 81350.0 183395.0 ;
      RECT  80645.0 184740.0 81350.0 186085.0 ;
      RECT  80645.0 187430.0 81350.0 186085.0 ;
      RECT  80645.0 187430.0 81350.0 188775.0 ;
      RECT  80645.0 190120.0 81350.0 188775.0 ;
      RECT  80645.0 190120.0 81350.0 191465.0 ;
      RECT  80645.0 192810.0 81350.0 191465.0 ;
      RECT  80645.0 192810.0 81350.0 194155.0 ;
      RECT  80645.0 195500.0 81350.0 194155.0 ;
      RECT  80645.0 195500.0 81350.0 196845.0 ;
      RECT  80645.0 198190.0 81350.0 196845.0 ;
      RECT  80645.0 198190.0 81350.0 199535.0 ;
      RECT  80645.0 200880.0 81350.0 199535.0 ;
      RECT  80645.0 200880.0 81350.0 202225.0 ;
      RECT  80645.0 203570.0 81350.0 202225.0 ;
      RECT  80645.0 203570.0 81350.0 204915.0 ;
      RECT  80645.0 206260.0 81350.0 204915.0 ;
      RECT  81350.0 34100.0 82055.0 35445.0 ;
      RECT  81350.0 36790.0 82055.0 35445.0 ;
      RECT  81350.0 36790.0 82055.0 38135.0 ;
      RECT  81350.0 39480.0 82055.0 38135.0 ;
      RECT  81350.0 39480.0 82055.0 40825.0 ;
      RECT  81350.0 42170.0 82055.0 40825.0 ;
      RECT  81350.0 42170.0 82055.0 43515.0 ;
      RECT  81350.0 44860.0 82055.0 43515.0 ;
      RECT  81350.0 44860.0 82055.0 46205.0 ;
      RECT  81350.0 47550.0 82055.0 46205.0 ;
      RECT  81350.0 47550.0 82055.0 48895.0 ;
      RECT  81350.0 50240.0 82055.0 48895.0 ;
      RECT  81350.0 50240.0 82055.0 51585.0 ;
      RECT  81350.0 52930.0 82055.0 51585.0 ;
      RECT  81350.0 52930.0 82055.0 54275.0 ;
      RECT  81350.0 55620.0 82055.0 54275.0 ;
      RECT  81350.0 55620.0 82055.0 56965.0 ;
      RECT  81350.0 58310.0 82055.0 56965.0 ;
      RECT  81350.0 58310.0 82055.0 59655.0 ;
      RECT  81350.0 61000.0 82055.0 59655.0 ;
      RECT  81350.0 61000.0 82055.0 62345.0 ;
      RECT  81350.0 63690.0 82055.0 62345.0 ;
      RECT  81350.0 63690.0 82055.0 65035.0 ;
      RECT  81350.0 66380.0 82055.0 65035.0 ;
      RECT  81350.0 66380.0 82055.0 67725.0 ;
      RECT  81350.0 69070.0 82055.0 67725.0 ;
      RECT  81350.0 69070.0 82055.0 70415.0 ;
      RECT  81350.0 71760.0 82055.0 70415.0 ;
      RECT  81350.0 71760.0 82055.0 73105.0 ;
      RECT  81350.0 74450.0 82055.0 73105.0 ;
      RECT  81350.0 74450.0 82055.0 75795.0 ;
      RECT  81350.0 77140.0 82055.0 75795.0 ;
      RECT  81350.0 77140.0 82055.0 78485.0 ;
      RECT  81350.0 79830.0 82055.0 78485.0 ;
      RECT  81350.0 79830.0 82055.0 81175.0 ;
      RECT  81350.0 82520.0 82055.0 81175.0 ;
      RECT  81350.0 82520.0 82055.0 83865.0 ;
      RECT  81350.0 85210.0 82055.0 83865.0 ;
      RECT  81350.0 85210.0 82055.0 86555.0 ;
      RECT  81350.0 87900.0 82055.0 86555.0 ;
      RECT  81350.0 87900.0 82055.0 89245.0 ;
      RECT  81350.0 90590.0 82055.0 89245.0 ;
      RECT  81350.0 90590.0 82055.0 91935.0 ;
      RECT  81350.0 93280.0 82055.0 91935.0 ;
      RECT  81350.0 93280.0 82055.0 94625.0 ;
      RECT  81350.0 95970.0 82055.0 94625.0 ;
      RECT  81350.0 95970.0 82055.0 97315.0 ;
      RECT  81350.0 98660.0 82055.0 97315.0 ;
      RECT  81350.0 98660.0 82055.0 100005.0 ;
      RECT  81350.0 101350.0 82055.0 100005.0 ;
      RECT  81350.0 101350.0 82055.0 102695.0 ;
      RECT  81350.0 104040.0 82055.0 102695.0 ;
      RECT  81350.0 104040.0 82055.0 105385.0 ;
      RECT  81350.0 106730.0 82055.0 105385.0 ;
      RECT  81350.0 106730.0 82055.0 108075.0 ;
      RECT  81350.0 109420.0 82055.0 108075.0 ;
      RECT  81350.0 109420.0 82055.0 110765.0 ;
      RECT  81350.0 112110.0 82055.0 110765.0 ;
      RECT  81350.0 112110.0 82055.0 113455.0 ;
      RECT  81350.0 114800.0 82055.0 113455.0 ;
      RECT  81350.0 114800.0 82055.0 116145.0 ;
      RECT  81350.0 117490.0 82055.0 116145.0 ;
      RECT  81350.0 117490.0 82055.0 118835.0 ;
      RECT  81350.0 120180.0 82055.0 118835.0 ;
      RECT  81350.0 120180.0 82055.0 121525.0 ;
      RECT  81350.0 122870.0 82055.0 121525.0 ;
      RECT  81350.0 122870.0 82055.0 124215.0 ;
      RECT  81350.0 125560.0 82055.0 124215.0 ;
      RECT  81350.0 125560.0 82055.0 126905.0 ;
      RECT  81350.0 128250.0 82055.0 126905.0 ;
      RECT  81350.0 128250.0 82055.0 129595.0 ;
      RECT  81350.0 130940.0 82055.0 129595.0 ;
      RECT  81350.0 130940.0 82055.0 132285.0 ;
      RECT  81350.0 133630.0 82055.0 132285.0 ;
      RECT  81350.0 133630.0 82055.0 134975.0 ;
      RECT  81350.0 136320.0 82055.0 134975.0 ;
      RECT  81350.0 136320.0 82055.0 137665.0 ;
      RECT  81350.0 139010.0 82055.0 137665.0 ;
      RECT  81350.0 139010.0 82055.0 140355.0 ;
      RECT  81350.0 141700.0 82055.0 140355.0 ;
      RECT  81350.0 141700.0 82055.0 143045.0 ;
      RECT  81350.0 144390.0 82055.0 143045.0 ;
      RECT  81350.0 144390.0 82055.0 145735.0 ;
      RECT  81350.0 147080.0 82055.0 145735.0 ;
      RECT  81350.0 147080.0 82055.0 148425.0 ;
      RECT  81350.0 149770.0 82055.0 148425.0 ;
      RECT  81350.0 149770.0 82055.0 151115.0 ;
      RECT  81350.0 152460.0 82055.0 151115.0 ;
      RECT  81350.0 152460.0 82055.0 153805.0 ;
      RECT  81350.0 155150.0 82055.0 153805.0 ;
      RECT  81350.0 155150.0 82055.0 156495.0 ;
      RECT  81350.0 157840.0 82055.0 156495.0 ;
      RECT  81350.0 157840.0 82055.0 159185.0 ;
      RECT  81350.0 160530.0 82055.0 159185.0 ;
      RECT  81350.0 160530.0 82055.0 161875.0 ;
      RECT  81350.0 163220.0 82055.0 161875.0 ;
      RECT  81350.0 163220.0 82055.0 164565.0 ;
      RECT  81350.0 165910.0 82055.0 164565.0 ;
      RECT  81350.0 165910.0 82055.0 167255.0 ;
      RECT  81350.0 168600.0 82055.0 167255.0 ;
      RECT  81350.0 168600.0 82055.0 169945.0 ;
      RECT  81350.0 171290.0 82055.0 169945.0 ;
      RECT  81350.0 171290.0 82055.0 172635.0 ;
      RECT  81350.0 173980.0 82055.0 172635.0 ;
      RECT  81350.0 173980.0 82055.0 175325.0 ;
      RECT  81350.0 176670.0 82055.0 175325.0 ;
      RECT  81350.0 176670.0 82055.0 178015.0 ;
      RECT  81350.0 179360.0 82055.0 178015.0 ;
      RECT  81350.0 179360.0 82055.0 180705.0 ;
      RECT  81350.0 182050.0 82055.0 180705.0 ;
      RECT  81350.0 182050.0 82055.0 183395.0 ;
      RECT  81350.0 184740.0 82055.0 183395.0 ;
      RECT  81350.0 184740.0 82055.0 186085.0 ;
      RECT  81350.0 187430.0 82055.0 186085.0 ;
      RECT  81350.0 187430.0 82055.0 188775.0 ;
      RECT  81350.0 190120.0 82055.0 188775.0 ;
      RECT  81350.0 190120.0 82055.0 191465.0 ;
      RECT  81350.0 192810.0 82055.0 191465.0 ;
      RECT  81350.0 192810.0 82055.0 194155.0 ;
      RECT  81350.0 195500.0 82055.0 194155.0 ;
      RECT  81350.0 195500.0 82055.0 196845.0 ;
      RECT  81350.0 198190.0 82055.0 196845.0 ;
      RECT  81350.0 198190.0 82055.0 199535.0 ;
      RECT  81350.0 200880.0 82055.0 199535.0 ;
      RECT  81350.0 200880.0 82055.0 202225.0 ;
      RECT  81350.0 203570.0 82055.0 202225.0 ;
      RECT  81350.0 203570.0 82055.0 204915.0 ;
      RECT  81350.0 206260.0 82055.0 204915.0 ;
      RECT  82055.0 34100.0 82760.0 35445.0 ;
      RECT  82055.0 36790.0 82760.0 35445.0 ;
      RECT  82055.0 36790.0 82760.0 38135.0 ;
      RECT  82055.0 39480.0 82760.0 38135.0 ;
      RECT  82055.0 39480.0 82760.0 40825.0 ;
      RECT  82055.0 42170.0 82760.0 40825.0 ;
      RECT  82055.0 42170.0 82760.0 43515.0 ;
      RECT  82055.0 44860.0 82760.0 43515.0 ;
      RECT  82055.0 44860.0 82760.0 46205.0 ;
      RECT  82055.0 47550.0 82760.0 46205.0 ;
      RECT  82055.0 47550.0 82760.0 48895.0 ;
      RECT  82055.0 50240.0 82760.0 48895.0 ;
      RECT  82055.0 50240.0 82760.0 51585.0 ;
      RECT  82055.0 52930.0 82760.0 51585.0 ;
      RECT  82055.0 52930.0 82760.0 54275.0 ;
      RECT  82055.0 55620.0 82760.0 54275.0 ;
      RECT  82055.0 55620.0 82760.0 56965.0 ;
      RECT  82055.0 58310.0 82760.0 56965.0 ;
      RECT  82055.0 58310.0 82760.0 59655.0 ;
      RECT  82055.0 61000.0 82760.0 59655.0 ;
      RECT  82055.0 61000.0 82760.0 62345.0 ;
      RECT  82055.0 63690.0 82760.0 62345.0 ;
      RECT  82055.0 63690.0 82760.0 65035.0 ;
      RECT  82055.0 66380.0 82760.0 65035.0 ;
      RECT  82055.0 66380.0 82760.0 67725.0 ;
      RECT  82055.0 69070.0 82760.0 67725.0 ;
      RECT  82055.0 69070.0 82760.0 70415.0 ;
      RECT  82055.0 71760.0 82760.0 70415.0 ;
      RECT  82055.0 71760.0 82760.0 73105.0 ;
      RECT  82055.0 74450.0 82760.0 73105.0 ;
      RECT  82055.0 74450.0 82760.0 75795.0 ;
      RECT  82055.0 77140.0 82760.0 75795.0 ;
      RECT  82055.0 77140.0 82760.0 78485.0 ;
      RECT  82055.0 79830.0 82760.0 78485.0 ;
      RECT  82055.0 79830.0 82760.0 81175.0 ;
      RECT  82055.0 82520.0 82760.0 81175.0 ;
      RECT  82055.0 82520.0 82760.0 83865.0 ;
      RECT  82055.0 85210.0 82760.0 83865.0 ;
      RECT  82055.0 85210.0 82760.0 86555.0 ;
      RECT  82055.0 87900.0 82760.0 86555.0 ;
      RECT  82055.0 87900.0 82760.0 89245.0 ;
      RECT  82055.0 90590.0 82760.0 89245.0 ;
      RECT  82055.0 90590.0 82760.0 91935.0 ;
      RECT  82055.0 93280.0 82760.0 91935.0 ;
      RECT  82055.0 93280.0 82760.0 94625.0 ;
      RECT  82055.0 95970.0 82760.0 94625.0 ;
      RECT  82055.0 95970.0 82760.0 97315.0 ;
      RECT  82055.0 98660.0 82760.0 97315.0 ;
      RECT  82055.0 98660.0 82760.0 100005.0 ;
      RECT  82055.0 101350.0 82760.0 100005.0 ;
      RECT  82055.0 101350.0 82760.0 102695.0 ;
      RECT  82055.0 104040.0 82760.0 102695.0 ;
      RECT  82055.0 104040.0 82760.0 105385.0 ;
      RECT  82055.0 106730.0 82760.0 105385.0 ;
      RECT  82055.0 106730.0 82760.0 108075.0 ;
      RECT  82055.0 109420.0 82760.0 108075.0 ;
      RECT  82055.0 109420.0 82760.0 110765.0 ;
      RECT  82055.0 112110.0 82760.0 110765.0 ;
      RECT  82055.0 112110.0 82760.0 113455.0 ;
      RECT  82055.0 114800.0 82760.0 113455.0 ;
      RECT  82055.0 114800.0 82760.0 116145.0 ;
      RECT  82055.0 117490.0 82760.0 116145.0 ;
      RECT  82055.0 117490.0 82760.0 118835.0 ;
      RECT  82055.0 120180.0 82760.0 118835.0 ;
      RECT  82055.0 120180.0 82760.0 121525.0 ;
      RECT  82055.0 122870.0 82760.0 121525.0 ;
      RECT  82055.0 122870.0 82760.0 124215.0 ;
      RECT  82055.0 125560.0 82760.0 124215.0 ;
      RECT  82055.0 125560.0 82760.0 126905.0 ;
      RECT  82055.0 128250.0 82760.0 126905.0 ;
      RECT  82055.0 128250.0 82760.0 129595.0 ;
      RECT  82055.0 130940.0 82760.0 129595.0 ;
      RECT  82055.0 130940.0 82760.0 132285.0 ;
      RECT  82055.0 133630.0 82760.0 132285.0 ;
      RECT  82055.0 133630.0 82760.0 134975.0 ;
      RECT  82055.0 136320.0 82760.0 134975.0 ;
      RECT  82055.0 136320.0 82760.0 137665.0 ;
      RECT  82055.0 139010.0 82760.0 137665.0 ;
      RECT  82055.0 139010.0 82760.0 140355.0 ;
      RECT  82055.0 141700.0 82760.0 140355.0 ;
      RECT  82055.0 141700.0 82760.0 143045.0 ;
      RECT  82055.0 144390.0 82760.0 143045.0 ;
      RECT  82055.0 144390.0 82760.0 145735.0 ;
      RECT  82055.0 147080.0 82760.0 145735.0 ;
      RECT  82055.0 147080.0 82760.0 148425.0 ;
      RECT  82055.0 149770.0 82760.0 148425.0 ;
      RECT  82055.0 149770.0 82760.0 151115.0 ;
      RECT  82055.0 152460.0 82760.0 151115.0 ;
      RECT  82055.0 152460.0 82760.0 153805.0 ;
      RECT  82055.0 155150.0 82760.0 153805.0 ;
      RECT  82055.0 155150.0 82760.0 156495.0 ;
      RECT  82055.0 157840.0 82760.0 156495.0 ;
      RECT  82055.0 157840.0 82760.0 159185.0 ;
      RECT  82055.0 160530.0 82760.0 159185.0 ;
      RECT  82055.0 160530.0 82760.0 161875.0 ;
      RECT  82055.0 163220.0 82760.0 161875.0 ;
      RECT  82055.0 163220.0 82760.0 164565.0 ;
      RECT  82055.0 165910.0 82760.0 164565.0 ;
      RECT  82055.0 165910.0 82760.0 167255.0 ;
      RECT  82055.0 168600.0 82760.0 167255.0 ;
      RECT  82055.0 168600.0 82760.0 169945.0 ;
      RECT  82055.0 171290.0 82760.0 169945.0 ;
      RECT  82055.0 171290.0 82760.0 172635.0 ;
      RECT  82055.0 173980.0 82760.0 172635.0 ;
      RECT  82055.0 173980.0 82760.0 175325.0 ;
      RECT  82055.0 176670.0 82760.0 175325.0 ;
      RECT  82055.0 176670.0 82760.0 178015.0 ;
      RECT  82055.0 179360.0 82760.0 178015.0 ;
      RECT  82055.0 179360.0 82760.0 180705.0 ;
      RECT  82055.0 182050.0 82760.0 180705.0 ;
      RECT  82055.0 182050.0 82760.0 183395.0 ;
      RECT  82055.0 184740.0 82760.0 183395.0 ;
      RECT  82055.0 184740.0 82760.0 186085.0 ;
      RECT  82055.0 187430.0 82760.0 186085.0 ;
      RECT  82055.0 187430.0 82760.0 188775.0 ;
      RECT  82055.0 190120.0 82760.0 188775.0 ;
      RECT  82055.0 190120.0 82760.0 191465.0 ;
      RECT  82055.0 192810.0 82760.0 191465.0 ;
      RECT  82055.0 192810.0 82760.0 194155.0 ;
      RECT  82055.0 195500.0 82760.0 194155.0 ;
      RECT  82055.0 195500.0 82760.0 196845.0 ;
      RECT  82055.0 198190.0 82760.0 196845.0 ;
      RECT  82055.0 198190.0 82760.0 199535.0 ;
      RECT  82055.0 200880.0 82760.0 199535.0 ;
      RECT  82055.0 200880.0 82760.0 202225.0 ;
      RECT  82055.0 203570.0 82760.0 202225.0 ;
      RECT  82055.0 203570.0 82760.0 204915.0 ;
      RECT  82055.0 206260.0 82760.0 204915.0 ;
      RECT  82760.0 34100.0 83465.0 35445.0 ;
      RECT  82760.0 36790.0 83465.0 35445.0 ;
      RECT  82760.0 36790.0 83465.0 38135.0 ;
      RECT  82760.0 39480.0 83465.0 38135.0 ;
      RECT  82760.0 39480.0 83465.0 40825.0 ;
      RECT  82760.0 42170.0 83465.0 40825.0 ;
      RECT  82760.0 42170.0 83465.0 43515.0 ;
      RECT  82760.0 44860.0 83465.0 43515.0 ;
      RECT  82760.0 44860.0 83465.0 46205.0 ;
      RECT  82760.0 47550.0 83465.0 46205.0 ;
      RECT  82760.0 47550.0 83465.0 48895.0 ;
      RECT  82760.0 50240.0 83465.0 48895.0 ;
      RECT  82760.0 50240.0 83465.0 51585.0 ;
      RECT  82760.0 52930.0 83465.0 51585.0 ;
      RECT  82760.0 52930.0 83465.0 54275.0 ;
      RECT  82760.0 55620.0 83465.0 54275.0 ;
      RECT  82760.0 55620.0 83465.0 56965.0 ;
      RECT  82760.0 58310.0 83465.0 56965.0 ;
      RECT  82760.0 58310.0 83465.0 59655.0 ;
      RECT  82760.0 61000.0 83465.0 59655.0 ;
      RECT  82760.0 61000.0 83465.0 62345.0 ;
      RECT  82760.0 63690.0 83465.0 62345.0 ;
      RECT  82760.0 63690.0 83465.0 65035.0 ;
      RECT  82760.0 66380.0 83465.0 65035.0 ;
      RECT  82760.0 66380.0 83465.0 67725.0 ;
      RECT  82760.0 69070.0 83465.0 67725.0 ;
      RECT  82760.0 69070.0 83465.0 70415.0 ;
      RECT  82760.0 71760.0 83465.0 70415.0 ;
      RECT  82760.0 71760.0 83465.0 73105.0 ;
      RECT  82760.0 74450.0 83465.0 73105.0 ;
      RECT  82760.0 74450.0 83465.0 75795.0 ;
      RECT  82760.0 77140.0 83465.0 75795.0 ;
      RECT  82760.0 77140.0 83465.0 78485.0 ;
      RECT  82760.0 79830.0 83465.0 78485.0 ;
      RECT  82760.0 79830.0 83465.0 81175.0 ;
      RECT  82760.0 82520.0 83465.0 81175.0 ;
      RECT  82760.0 82520.0 83465.0 83865.0 ;
      RECT  82760.0 85210.0 83465.0 83865.0 ;
      RECT  82760.0 85210.0 83465.0 86555.0 ;
      RECT  82760.0 87900.0 83465.0 86555.0 ;
      RECT  82760.0 87900.0 83465.0 89245.0 ;
      RECT  82760.0 90590.0 83465.0 89245.0 ;
      RECT  82760.0 90590.0 83465.0 91935.0 ;
      RECT  82760.0 93280.0 83465.0 91935.0 ;
      RECT  82760.0 93280.0 83465.0 94625.0 ;
      RECT  82760.0 95970.0 83465.0 94625.0 ;
      RECT  82760.0 95970.0 83465.0 97315.0 ;
      RECT  82760.0 98660.0 83465.0 97315.0 ;
      RECT  82760.0 98660.0 83465.0 100005.0 ;
      RECT  82760.0 101350.0 83465.0 100005.0 ;
      RECT  82760.0 101350.0 83465.0 102695.0 ;
      RECT  82760.0 104040.0 83465.0 102695.0 ;
      RECT  82760.0 104040.0 83465.0 105385.0 ;
      RECT  82760.0 106730.0 83465.0 105385.0 ;
      RECT  82760.0 106730.0 83465.0 108075.0 ;
      RECT  82760.0 109420.0 83465.0 108075.0 ;
      RECT  82760.0 109420.0 83465.0 110765.0 ;
      RECT  82760.0 112110.0 83465.0 110765.0 ;
      RECT  82760.0 112110.0 83465.0 113455.0 ;
      RECT  82760.0 114800.0 83465.0 113455.0 ;
      RECT  82760.0 114800.0 83465.0 116145.0 ;
      RECT  82760.0 117490.0 83465.0 116145.0 ;
      RECT  82760.0 117490.0 83465.0 118835.0 ;
      RECT  82760.0 120180.0 83465.0 118835.0 ;
      RECT  82760.0 120180.0 83465.0 121525.0 ;
      RECT  82760.0 122870.0 83465.0 121525.0 ;
      RECT  82760.0 122870.0 83465.0 124215.0 ;
      RECT  82760.0 125560.0 83465.0 124215.0 ;
      RECT  82760.0 125560.0 83465.0 126905.0 ;
      RECT  82760.0 128250.0 83465.0 126905.0 ;
      RECT  82760.0 128250.0 83465.0 129595.0 ;
      RECT  82760.0 130940.0 83465.0 129595.0 ;
      RECT  82760.0 130940.0 83465.0 132285.0 ;
      RECT  82760.0 133630.0 83465.0 132285.0 ;
      RECT  82760.0 133630.0 83465.0 134975.0 ;
      RECT  82760.0 136320.0 83465.0 134975.0 ;
      RECT  82760.0 136320.0 83465.0 137665.0 ;
      RECT  82760.0 139010.0 83465.0 137665.0 ;
      RECT  82760.0 139010.0 83465.0 140355.0 ;
      RECT  82760.0 141700.0 83465.0 140355.0 ;
      RECT  82760.0 141700.0 83465.0 143045.0 ;
      RECT  82760.0 144390.0 83465.0 143045.0 ;
      RECT  82760.0 144390.0 83465.0 145735.0 ;
      RECT  82760.0 147080.0 83465.0 145735.0 ;
      RECT  82760.0 147080.0 83465.0 148425.0 ;
      RECT  82760.0 149770.0 83465.0 148425.0 ;
      RECT  82760.0 149770.0 83465.0 151115.0 ;
      RECT  82760.0 152460.0 83465.0 151115.0 ;
      RECT  82760.0 152460.0 83465.0 153805.0 ;
      RECT  82760.0 155150.0 83465.0 153805.0 ;
      RECT  82760.0 155150.0 83465.0 156495.0 ;
      RECT  82760.0 157840.0 83465.0 156495.0 ;
      RECT  82760.0 157840.0 83465.0 159185.0 ;
      RECT  82760.0 160530.0 83465.0 159185.0 ;
      RECT  82760.0 160530.0 83465.0 161875.0 ;
      RECT  82760.0 163220.0 83465.0 161875.0 ;
      RECT  82760.0 163220.0 83465.0 164565.0 ;
      RECT  82760.0 165910.0 83465.0 164565.0 ;
      RECT  82760.0 165910.0 83465.0 167255.0 ;
      RECT  82760.0 168600.0 83465.0 167255.0 ;
      RECT  82760.0 168600.0 83465.0 169945.0 ;
      RECT  82760.0 171290.0 83465.0 169945.0 ;
      RECT  82760.0 171290.0 83465.0 172635.0 ;
      RECT  82760.0 173980.0 83465.0 172635.0 ;
      RECT  82760.0 173980.0 83465.0 175325.0 ;
      RECT  82760.0 176670.0 83465.0 175325.0 ;
      RECT  82760.0 176670.0 83465.0 178015.0 ;
      RECT  82760.0 179360.0 83465.0 178015.0 ;
      RECT  82760.0 179360.0 83465.0 180705.0 ;
      RECT  82760.0 182050.0 83465.0 180705.0 ;
      RECT  82760.0 182050.0 83465.0 183395.0 ;
      RECT  82760.0 184740.0 83465.0 183395.0 ;
      RECT  82760.0 184740.0 83465.0 186085.0 ;
      RECT  82760.0 187430.0 83465.0 186085.0 ;
      RECT  82760.0 187430.0 83465.0 188775.0 ;
      RECT  82760.0 190120.0 83465.0 188775.0 ;
      RECT  82760.0 190120.0 83465.0 191465.0 ;
      RECT  82760.0 192810.0 83465.0 191465.0 ;
      RECT  82760.0 192810.0 83465.0 194155.0 ;
      RECT  82760.0 195500.0 83465.0 194155.0 ;
      RECT  82760.0 195500.0 83465.0 196845.0 ;
      RECT  82760.0 198190.0 83465.0 196845.0 ;
      RECT  82760.0 198190.0 83465.0 199535.0 ;
      RECT  82760.0 200880.0 83465.0 199535.0 ;
      RECT  82760.0 200880.0 83465.0 202225.0 ;
      RECT  82760.0 203570.0 83465.0 202225.0 ;
      RECT  82760.0 203570.0 83465.0 204915.0 ;
      RECT  82760.0 206260.0 83465.0 204915.0 ;
      RECT  83465.0 34100.0 84170.0 35445.0 ;
      RECT  83465.0 36790.0 84170.0 35445.0 ;
      RECT  83465.0 36790.0 84170.0 38135.0 ;
      RECT  83465.0 39480.0 84170.0 38135.0 ;
      RECT  83465.0 39480.0 84170.0 40825.0 ;
      RECT  83465.0 42170.0 84170.0 40825.0 ;
      RECT  83465.0 42170.0 84170.0 43515.0 ;
      RECT  83465.0 44860.0 84170.0 43515.0 ;
      RECT  83465.0 44860.0 84170.0 46205.0 ;
      RECT  83465.0 47550.0 84170.0 46205.0 ;
      RECT  83465.0 47550.0 84170.0 48895.0 ;
      RECT  83465.0 50240.0 84170.0 48895.0 ;
      RECT  83465.0 50240.0 84170.0 51585.0 ;
      RECT  83465.0 52930.0 84170.0 51585.0 ;
      RECT  83465.0 52930.0 84170.0 54275.0 ;
      RECT  83465.0 55620.0 84170.0 54275.0 ;
      RECT  83465.0 55620.0 84170.0 56965.0 ;
      RECT  83465.0 58310.0 84170.0 56965.0 ;
      RECT  83465.0 58310.0 84170.0 59655.0 ;
      RECT  83465.0 61000.0 84170.0 59655.0 ;
      RECT  83465.0 61000.0 84170.0 62345.0 ;
      RECT  83465.0 63690.0 84170.0 62345.0 ;
      RECT  83465.0 63690.0 84170.0 65035.0 ;
      RECT  83465.0 66380.0 84170.0 65035.0 ;
      RECT  83465.0 66380.0 84170.0 67725.0 ;
      RECT  83465.0 69070.0 84170.0 67725.0 ;
      RECT  83465.0 69070.0 84170.0 70415.0 ;
      RECT  83465.0 71760.0 84170.0 70415.0 ;
      RECT  83465.0 71760.0 84170.0 73105.0 ;
      RECT  83465.0 74450.0 84170.0 73105.0 ;
      RECT  83465.0 74450.0 84170.0 75795.0 ;
      RECT  83465.0 77140.0 84170.0 75795.0 ;
      RECT  83465.0 77140.0 84170.0 78485.0 ;
      RECT  83465.0 79830.0 84170.0 78485.0 ;
      RECT  83465.0 79830.0 84170.0 81175.0 ;
      RECT  83465.0 82520.0 84170.0 81175.0 ;
      RECT  83465.0 82520.0 84170.0 83865.0 ;
      RECT  83465.0 85210.0 84170.0 83865.0 ;
      RECT  83465.0 85210.0 84170.0 86555.0 ;
      RECT  83465.0 87900.0 84170.0 86555.0 ;
      RECT  83465.0 87900.0 84170.0 89245.0 ;
      RECT  83465.0 90590.0 84170.0 89245.0 ;
      RECT  83465.0 90590.0 84170.0 91935.0 ;
      RECT  83465.0 93280.0 84170.0 91935.0 ;
      RECT  83465.0 93280.0 84170.0 94625.0 ;
      RECT  83465.0 95970.0 84170.0 94625.0 ;
      RECT  83465.0 95970.0 84170.0 97315.0 ;
      RECT  83465.0 98660.0 84170.0 97315.0 ;
      RECT  83465.0 98660.0 84170.0 100005.0 ;
      RECT  83465.0 101350.0 84170.0 100005.0 ;
      RECT  83465.0 101350.0 84170.0 102695.0 ;
      RECT  83465.0 104040.0 84170.0 102695.0 ;
      RECT  83465.0 104040.0 84170.0 105385.0 ;
      RECT  83465.0 106730.0 84170.0 105385.0 ;
      RECT  83465.0 106730.0 84170.0 108075.0 ;
      RECT  83465.0 109420.0 84170.0 108075.0 ;
      RECT  83465.0 109420.0 84170.0 110765.0 ;
      RECT  83465.0 112110.0 84170.0 110765.0 ;
      RECT  83465.0 112110.0 84170.0 113455.0 ;
      RECT  83465.0 114800.0 84170.0 113455.0 ;
      RECT  83465.0 114800.0 84170.0 116145.0 ;
      RECT  83465.0 117490.0 84170.0 116145.0 ;
      RECT  83465.0 117490.0 84170.0 118835.0 ;
      RECT  83465.0 120180.0 84170.0 118835.0 ;
      RECT  83465.0 120180.0 84170.0 121525.0 ;
      RECT  83465.0 122870.0 84170.0 121525.0 ;
      RECT  83465.0 122870.0 84170.0 124215.0 ;
      RECT  83465.0 125560.0 84170.0 124215.0 ;
      RECT  83465.0 125560.0 84170.0 126905.0 ;
      RECT  83465.0 128250.0 84170.0 126905.0 ;
      RECT  83465.0 128250.0 84170.0 129595.0 ;
      RECT  83465.0 130940.0 84170.0 129595.0 ;
      RECT  83465.0 130940.0 84170.0 132285.0 ;
      RECT  83465.0 133630.0 84170.0 132285.0 ;
      RECT  83465.0 133630.0 84170.0 134975.0 ;
      RECT  83465.0 136320.0 84170.0 134975.0 ;
      RECT  83465.0 136320.0 84170.0 137665.0 ;
      RECT  83465.0 139010.0 84170.0 137665.0 ;
      RECT  83465.0 139010.0 84170.0 140355.0 ;
      RECT  83465.0 141700.0 84170.0 140355.0 ;
      RECT  83465.0 141700.0 84170.0 143045.0 ;
      RECT  83465.0 144390.0 84170.0 143045.0 ;
      RECT  83465.0 144390.0 84170.0 145735.0 ;
      RECT  83465.0 147080.0 84170.0 145735.0 ;
      RECT  83465.0 147080.0 84170.0 148425.0 ;
      RECT  83465.0 149770.0 84170.0 148425.0 ;
      RECT  83465.0 149770.0 84170.0 151115.0 ;
      RECT  83465.0 152460.0 84170.0 151115.0 ;
      RECT  83465.0 152460.0 84170.0 153805.0 ;
      RECT  83465.0 155150.0 84170.0 153805.0 ;
      RECT  83465.0 155150.0 84170.0 156495.0 ;
      RECT  83465.0 157840.0 84170.0 156495.0 ;
      RECT  83465.0 157840.0 84170.0 159185.0 ;
      RECT  83465.0 160530.0 84170.0 159185.0 ;
      RECT  83465.0 160530.0 84170.0 161875.0 ;
      RECT  83465.0 163220.0 84170.0 161875.0 ;
      RECT  83465.0 163220.0 84170.0 164565.0 ;
      RECT  83465.0 165910.0 84170.0 164565.0 ;
      RECT  83465.0 165910.0 84170.0 167255.0 ;
      RECT  83465.0 168600.0 84170.0 167255.0 ;
      RECT  83465.0 168600.0 84170.0 169945.0 ;
      RECT  83465.0 171290.0 84170.0 169945.0 ;
      RECT  83465.0 171290.0 84170.0 172635.0 ;
      RECT  83465.0 173980.0 84170.0 172635.0 ;
      RECT  83465.0 173980.0 84170.0 175325.0 ;
      RECT  83465.0 176670.0 84170.0 175325.0 ;
      RECT  83465.0 176670.0 84170.0 178015.0 ;
      RECT  83465.0 179360.0 84170.0 178015.0 ;
      RECT  83465.0 179360.0 84170.0 180705.0 ;
      RECT  83465.0 182050.0 84170.0 180705.0 ;
      RECT  83465.0 182050.0 84170.0 183395.0 ;
      RECT  83465.0 184740.0 84170.0 183395.0 ;
      RECT  83465.0 184740.0 84170.0 186085.0 ;
      RECT  83465.0 187430.0 84170.0 186085.0 ;
      RECT  83465.0 187430.0 84170.0 188775.0 ;
      RECT  83465.0 190120.0 84170.0 188775.0 ;
      RECT  83465.0 190120.0 84170.0 191465.0 ;
      RECT  83465.0 192810.0 84170.0 191465.0 ;
      RECT  83465.0 192810.0 84170.0 194155.0 ;
      RECT  83465.0 195500.0 84170.0 194155.0 ;
      RECT  83465.0 195500.0 84170.0 196845.0 ;
      RECT  83465.0 198190.0 84170.0 196845.0 ;
      RECT  83465.0 198190.0 84170.0 199535.0 ;
      RECT  83465.0 200880.0 84170.0 199535.0 ;
      RECT  83465.0 200880.0 84170.0 202225.0 ;
      RECT  83465.0 203570.0 84170.0 202225.0 ;
      RECT  83465.0 203570.0 84170.0 204915.0 ;
      RECT  83465.0 206260.0 84170.0 204915.0 ;
      RECT  84170.0 34100.0 84875.0 35445.0 ;
      RECT  84170.0 36790.0 84875.0 35445.0 ;
      RECT  84170.0 36790.0 84875.0 38135.0 ;
      RECT  84170.0 39480.0 84875.0 38135.0 ;
      RECT  84170.0 39480.0 84875.0 40825.0 ;
      RECT  84170.0 42170.0 84875.0 40825.0 ;
      RECT  84170.0 42170.0 84875.0 43515.0 ;
      RECT  84170.0 44860.0 84875.0 43515.0 ;
      RECT  84170.0 44860.0 84875.0 46205.0 ;
      RECT  84170.0 47550.0 84875.0 46205.0 ;
      RECT  84170.0 47550.0 84875.0 48895.0 ;
      RECT  84170.0 50240.0 84875.0 48895.0 ;
      RECT  84170.0 50240.0 84875.0 51585.0 ;
      RECT  84170.0 52930.0 84875.0 51585.0 ;
      RECT  84170.0 52930.0 84875.0 54275.0 ;
      RECT  84170.0 55620.0 84875.0 54275.0 ;
      RECT  84170.0 55620.0 84875.0 56965.0 ;
      RECT  84170.0 58310.0 84875.0 56965.0 ;
      RECT  84170.0 58310.0 84875.0 59655.0 ;
      RECT  84170.0 61000.0 84875.0 59655.0 ;
      RECT  84170.0 61000.0 84875.0 62345.0 ;
      RECT  84170.0 63690.0 84875.0 62345.0 ;
      RECT  84170.0 63690.0 84875.0 65035.0 ;
      RECT  84170.0 66380.0 84875.0 65035.0 ;
      RECT  84170.0 66380.0 84875.0 67725.0 ;
      RECT  84170.0 69070.0 84875.0 67725.0 ;
      RECT  84170.0 69070.0 84875.0 70415.0 ;
      RECT  84170.0 71760.0 84875.0 70415.0 ;
      RECT  84170.0 71760.0 84875.0 73105.0 ;
      RECT  84170.0 74450.0 84875.0 73105.0 ;
      RECT  84170.0 74450.0 84875.0 75795.0 ;
      RECT  84170.0 77140.0 84875.0 75795.0 ;
      RECT  84170.0 77140.0 84875.0 78485.0 ;
      RECT  84170.0 79830.0 84875.0 78485.0 ;
      RECT  84170.0 79830.0 84875.0 81175.0 ;
      RECT  84170.0 82520.0 84875.0 81175.0 ;
      RECT  84170.0 82520.0 84875.0 83865.0 ;
      RECT  84170.0 85210.0 84875.0 83865.0 ;
      RECT  84170.0 85210.0 84875.0 86555.0 ;
      RECT  84170.0 87900.0 84875.0 86555.0 ;
      RECT  84170.0 87900.0 84875.0 89245.0 ;
      RECT  84170.0 90590.0 84875.0 89245.0 ;
      RECT  84170.0 90590.0 84875.0 91935.0 ;
      RECT  84170.0 93280.0 84875.0 91935.0 ;
      RECT  84170.0 93280.0 84875.0 94625.0 ;
      RECT  84170.0 95970.0 84875.0 94625.0 ;
      RECT  84170.0 95970.0 84875.0 97315.0 ;
      RECT  84170.0 98660.0 84875.0 97315.0 ;
      RECT  84170.0 98660.0 84875.0 100005.0 ;
      RECT  84170.0 101350.0 84875.0 100005.0 ;
      RECT  84170.0 101350.0 84875.0 102695.0 ;
      RECT  84170.0 104040.0 84875.0 102695.0 ;
      RECT  84170.0 104040.0 84875.0 105385.0 ;
      RECT  84170.0 106730.0 84875.0 105385.0 ;
      RECT  84170.0 106730.0 84875.0 108075.0 ;
      RECT  84170.0 109420.0 84875.0 108075.0 ;
      RECT  84170.0 109420.0 84875.0 110765.0 ;
      RECT  84170.0 112110.0 84875.0 110765.0 ;
      RECT  84170.0 112110.0 84875.0 113455.0 ;
      RECT  84170.0 114800.0 84875.0 113455.0 ;
      RECT  84170.0 114800.0 84875.0 116145.0 ;
      RECT  84170.0 117490.0 84875.0 116145.0 ;
      RECT  84170.0 117490.0 84875.0 118835.0 ;
      RECT  84170.0 120180.0 84875.0 118835.0 ;
      RECT  84170.0 120180.0 84875.0 121525.0 ;
      RECT  84170.0 122870.0 84875.0 121525.0 ;
      RECT  84170.0 122870.0 84875.0 124215.0 ;
      RECT  84170.0 125560.0 84875.0 124215.0 ;
      RECT  84170.0 125560.0 84875.0 126905.0 ;
      RECT  84170.0 128250.0 84875.0 126905.0 ;
      RECT  84170.0 128250.0 84875.0 129595.0 ;
      RECT  84170.0 130940.0 84875.0 129595.0 ;
      RECT  84170.0 130940.0 84875.0 132285.0 ;
      RECT  84170.0 133630.0 84875.0 132285.0 ;
      RECT  84170.0 133630.0 84875.0 134975.0 ;
      RECT  84170.0 136320.0 84875.0 134975.0 ;
      RECT  84170.0 136320.0 84875.0 137665.0 ;
      RECT  84170.0 139010.0 84875.0 137665.0 ;
      RECT  84170.0 139010.0 84875.0 140355.0 ;
      RECT  84170.0 141700.0 84875.0 140355.0 ;
      RECT  84170.0 141700.0 84875.0 143045.0 ;
      RECT  84170.0 144390.0 84875.0 143045.0 ;
      RECT  84170.0 144390.0 84875.0 145735.0 ;
      RECT  84170.0 147080.0 84875.0 145735.0 ;
      RECT  84170.0 147080.0 84875.0 148425.0 ;
      RECT  84170.0 149770.0 84875.0 148425.0 ;
      RECT  84170.0 149770.0 84875.0 151115.0 ;
      RECT  84170.0 152460.0 84875.0 151115.0 ;
      RECT  84170.0 152460.0 84875.0 153805.0 ;
      RECT  84170.0 155150.0 84875.0 153805.0 ;
      RECT  84170.0 155150.0 84875.0 156495.0 ;
      RECT  84170.0 157840.0 84875.0 156495.0 ;
      RECT  84170.0 157840.0 84875.0 159185.0 ;
      RECT  84170.0 160530.0 84875.0 159185.0 ;
      RECT  84170.0 160530.0 84875.0 161875.0 ;
      RECT  84170.0 163220.0 84875.0 161875.0 ;
      RECT  84170.0 163220.0 84875.0 164565.0 ;
      RECT  84170.0 165910.0 84875.0 164565.0 ;
      RECT  84170.0 165910.0 84875.0 167255.0 ;
      RECT  84170.0 168600.0 84875.0 167255.0 ;
      RECT  84170.0 168600.0 84875.0 169945.0 ;
      RECT  84170.0 171290.0 84875.0 169945.0 ;
      RECT  84170.0 171290.0 84875.0 172635.0 ;
      RECT  84170.0 173980.0 84875.0 172635.0 ;
      RECT  84170.0 173980.0 84875.0 175325.0 ;
      RECT  84170.0 176670.0 84875.0 175325.0 ;
      RECT  84170.0 176670.0 84875.0 178015.0 ;
      RECT  84170.0 179360.0 84875.0 178015.0 ;
      RECT  84170.0 179360.0 84875.0 180705.0 ;
      RECT  84170.0 182050.0 84875.0 180705.0 ;
      RECT  84170.0 182050.0 84875.0 183395.0 ;
      RECT  84170.0 184740.0 84875.0 183395.0 ;
      RECT  84170.0 184740.0 84875.0 186085.0 ;
      RECT  84170.0 187430.0 84875.0 186085.0 ;
      RECT  84170.0 187430.0 84875.0 188775.0 ;
      RECT  84170.0 190120.0 84875.0 188775.0 ;
      RECT  84170.0 190120.0 84875.0 191465.0 ;
      RECT  84170.0 192810.0 84875.0 191465.0 ;
      RECT  84170.0 192810.0 84875.0 194155.0 ;
      RECT  84170.0 195500.0 84875.0 194155.0 ;
      RECT  84170.0 195500.0 84875.0 196845.0 ;
      RECT  84170.0 198190.0 84875.0 196845.0 ;
      RECT  84170.0 198190.0 84875.0 199535.0 ;
      RECT  84170.0 200880.0 84875.0 199535.0 ;
      RECT  84170.0 200880.0 84875.0 202225.0 ;
      RECT  84170.0 203570.0 84875.0 202225.0 ;
      RECT  84170.0 203570.0 84875.0 204915.0 ;
      RECT  84170.0 206260.0 84875.0 204915.0 ;
      RECT  84875.0 34100.0 85580.0 35445.0 ;
      RECT  84875.0 36790.0 85580.0 35445.0 ;
      RECT  84875.0 36790.0 85580.0 38135.0 ;
      RECT  84875.0 39480.0 85580.0 38135.0 ;
      RECT  84875.0 39480.0 85580.0 40825.0 ;
      RECT  84875.0 42170.0 85580.0 40825.0 ;
      RECT  84875.0 42170.0 85580.0 43515.0 ;
      RECT  84875.0 44860.0 85580.0 43515.0 ;
      RECT  84875.0 44860.0 85580.0 46205.0 ;
      RECT  84875.0 47550.0 85580.0 46205.0 ;
      RECT  84875.0 47550.0 85580.0 48895.0 ;
      RECT  84875.0 50240.0 85580.0 48895.0 ;
      RECT  84875.0 50240.0 85580.0 51585.0 ;
      RECT  84875.0 52930.0 85580.0 51585.0 ;
      RECT  84875.0 52930.0 85580.0 54275.0 ;
      RECT  84875.0 55620.0 85580.0 54275.0 ;
      RECT  84875.0 55620.0 85580.0 56965.0 ;
      RECT  84875.0 58310.0 85580.0 56965.0 ;
      RECT  84875.0 58310.0 85580.0 59655.0 ;
      RECT  84875.0 61000.0 85580.0 59655.0 ;
      RECT  84875.0 61000.0 85580.0 62345.0 ;
      RECT  84875.0 63690.0 85580.0 62345.0 ;
      RECT  84875.0 63690.0 85580.0 65035.0 ;
      RECT  84875.0 66380.0 85580.0 65035.0 ;
      RECT  84875.0 66380.0 85580.0 67725.0 ;
      RECT  84875.0 69070.0 85580.0 67725.0 ;
      RECT  84875.0 69070.0 85580.0 70415.0 ;
      RECT  84875.0 71760.0 85580.0 70415.0 ;
      RECT  84875.0 71760.0 85580.0 73105.0 ;
      RECT  84875.0 74450.0 85580.0 73105.0 ;
      RECT  84875.0 74450.0 85580.0 75795.0 ;
      RECT  84875.0 77140.0 85580.0 75795.0 ;
      RECT  84875.0 77140.0 85580.0 78485.0 ;
      RECT  84875.0 79830.0 85580.0 78485.0 ;
      RECT  84875.0 79830.0 85580.0 81175.0 ;
      RECT  84875.0 82520.0 85580.0 81175.0 ;
      RECT  84875.0 82520.0 85580.0 83865.0 ;
      RECT  84875.0 85210.0 85580.0 83865.0 ;
      RECT  84875.0 85210.0 85580.0 86555.0 ;
      RECT  84875.0 87900.0 85580.0 86555.0 ;
      RECT  84875.0 87900.0 85580.0 89245.0 ;
      RECT  84875.0 90590.0 85580.0 89245.0 ;
      RECT  84875.0 90590.0 85580.0 91935.0 ;
      RECT  84875.0 93280.0 85580.0 91935.0 ;
      RECT  84875.0 93280.0 85580.0 94625.0 ;
      RECT  84875.0 95970.0 85580.0 94625.0 ;
      RECT  84875.0 95970.0 85580.0 97315.0 ;
      RECT  84875.0 98660.0 85580.0 97315.0 ;
      RECT  84875.0 98660.0 85580.0 100005.0 ;
      RECT  84875.0 101350.0 85580.0 100005.0 ;
      RECT  84875.0 101350.0 85580.0 102695.0 ;
      RECT  84875.0 104040.0 85580.0 102695.0 ;
      RECT  84875.0 104040.0 85580.0 105385.0 ;
      RECT  84875.0 106730.0 85580.0 105385.0 ;
      RECT  84875.0 106730.0 85580.0 108075.0 ;
      RECT  84875.0 109420.0 85580.0 108075.0 ;
      RECT  84875.0 109420.0 85580.0 110765.0 ;
      RECT  84875.0 112110.0 85580.0 110765.0 ;
      RECT  84875.0 112110.0 85580.0 113455.0 ;
      RECT  84875.0 114800.0 85580.0 113455.0 ;
      RECT  84875.0 114800.0 85580.0 116145.0 ;
      RECT  84875.0 117490.0 85580.0 116145.0 ;
      RECT  84875.0 117490.0 85580.0 118835.0 ;
      RECT  84875.0 120180.0 85580.0 118835.0 ;
      RECT  84875.0 120180.0 85580.0 121525.0 ;
      RECT  84875.0 122870.0 85580.0 121525.0 ;
      RECT  84875.0 122870.0 85580.0 124215.0 ;
      RECT  84875.0 125560.0 85580.0 124215.0 ;
      RECT  84875.0 125560.0 85580.0 126905.0 ;
      RECT  84875.0 128250.0 85580.0 126905.0 ;
      RECT  84875.0 128250.0 85580.0 129595.0 ;
      RECT  84875.0 130940.0 85580.0 129595.0 ;
      RECT  84875.0 130940.0 85580.0 132285.0 ;
      RECT  84875.0 133630.0 85580.0 132285.0 ;
      RECT  84875.0 133630.0 85580.0 134975.0 ;
      RECT  84875.0 136320.0 85580.0 134975.0 ;
      RECT  84875.0 136320.0 85580.0 137665.0 ;
      RECT  84875.0 139010.0 85580.0 137665.0 ;
      RECT  84875.0 139010.0 85580.0 140355.0 ;
      RECT  84875.0 141700.0 85580.0 140355.0 ;
      RECT  84875.0 141700.0 85580.0 143045.0 ;
      RECT  84875.0 144390.0 85580.0 143045.0 ;
      RECT  84875.0 144390.0 85580.0 145735.0 ;
      RECT  84875.0 147080.0 85580.0 145735.0 ;
      RECT  84875.0 147080.0 85580.0 148425.0 ;
      RECT  84875.0 149770.0 85580.0 148425.0 ;
      RECT  84875.0 149770.0 85580.0 151115.0 ;
      RECT  84875.0 152460.0 85580.0 151115.0 ;
      RECT  84875.0 152460.0 85580.0 153805.0 ;
      RECT  84875.0 155150.0 85580.0 153805.0 ;
      RECT  84875.0 155150.0 85580.0 156495.0 ;
      RECT  84875.0 157840.0 85580.0 156495.0 ;
      RECT  84875.0 157840.0 85580.0 159185.0 ;
      RECT  84875.0 160530.0 85580.0 159185.0 ;
      RECT  84875.0 160530.0 85580.0 161875.0 ;
      RECT  84875.0 163220.0 85580.0 161875.0 ;
      RECT  84875.0 163220.0 85580.0 164565.0 ;
      RECT  84875.0 165910.0 85580.0 164565.0 ;
      RECT  84875.0 165910.0 85580.0 167255.0 ;
      RECT  84875.0 168600.0 85580.0 167255.0 ;
      RECT  84875.0 168600.0 85580.0 169945.0 ;
      RECT  84875.0 171290.0 85580.0 169945.0 ;
      RECT  84875.0 171290.0 85580.0 172635.0 ;
      RECT  84875.0 173980.0 85580.0 172635.0 ;
      RECT  84875.0 173980.0 85580.0 175325.0 ;
      RECT  84875.0 176670.0 85580.0 175325.0 ;
      RECT  84875.0 176670.0 85580.0 178015.0 ;
      RECT  84875.0 179360.0 85580.0 178015.0 ;
      RECT  84875.0 179360.0 85580.0 180705.0 ;
      RECT  84875.0 182050.0 85580.0 180705.0 ;
      RECT  84875.0 182050.0 85580.0 183395.0 ;
      RECT  84875.0 184740.0 85580.0 183395.0 ;
      RECT  84875.0 184740.0 85580.0 186085.0 ;
      RECT  84875.0 187430.0 85580.0 186085.0 ;
      RECT  84875.0 187430.0 85580.0 188775.0 ;
      RECT  84875.0 190120.0 85580.0 188775.0 ;
      RECT  84875.0 190120.0 85580.0 191465.0 ;
      RECT  84875.0 192810.0 85580.0 191465.0 ;
      RECT  84875.0 192810.0 85580.0 194155.0 ;
      RECT  84875.0 195500.0 85580.0 194155.0 ;
      RECT  84875.0 195500.0 85580.0 196845.0 ;
      RECT  84875.0 198190.0 85580.0 196845.0 ;
      RECT  84875.0 198190.0 85580.0 199535.0 ;
      RECT  84875.0 200880.0 85580.0 199535.0 ;
      RECT  84875.0 200880.0 85580.0 202225.0 ;
      RECT  84875.0 203570.0 85580.0 202225.0 ;
      RECT  84875.0 203570.0 85580.0 204915.0 ;
      RECT  84875.0 206260.0 85580.0 204915.0 ;
      RECT  85580.0 34100.0 86285.0 35445.0 ;
      RECT  85580.0 36790.0 86285.0 35445.0 ;
      RECT  85580.0 36790.0 86285.0 38135.0 ;
      RECT  85580.0 39480.0 86285.0 38135.0 ;
      RECT  85580.0 39480.0 86285.0 40825.0 ;
      RECT  85580.0 42170.0 86285.0 40825.0 ;
      RECT  85580.0 42170.0 86285.0 43515.0 ;
      RECT  85580.0 44860.0 86285.0 43515.0 ;
      RECT  85580.0 44860.0 86285.0 46205.0 ;
      RECT  85580.0 47550.0 86285.0 46205.0 ;
      RECT  85580.0 47550.0 86285.0 48895.0 ;
      RECT  85580.0 50240.0 86285.0 48895.0 ;
      RECT  85580.0 50240.0 86285.0 51585.0 ;
      RECT  85580.0 52930.0 86285.0 51585.0 ;
      RECT  85580.0 52930.0 86285.0 54275.0 ;
      RECT  85580.0 55620.0 86285.0 54275.0 ;
      RECT  85580.0 55620.0 86285.0 56965.0 ;
      RECT  85580.0 58310.0 86285.0 56965.0 ;
      RECT  85580.0 58310.0 86285.0 59655.0 ;
      RECT  85580.0 61000.0 86285.0 59655.0 ;
      RECT  85580.0 61000.0 86285.0 62345.0 ;
      RECT  85580.0 63690.0 86285.0 62345.0 ;
      RECT  85580.0 63690.0 86285.0 65035.0 ;
      RECT  85580.0 66380.0 86285.0 65035.0 ;
      RECT  85580.0 66380.0 86285.0 67725.0 ;
      RECT  85580.0 69070.0 86285.0 67725.0 ;
      RECT  85580.0 69070.0 86285.0 70415.0 ;
      RECT  85580.0 71760.0 86285.0 70415.0 ;
      RECT  85580.0 71760.0 86285.0 73105.0 ;
      RECT  85580.0 74450.0 86285.0 73105.0 ;
      RECT  85580.0 74450.0 86285.0 75795.0 ;
      RECT  85580.0 77140.0 86285.0 75795.0 ;
      RECT  85580.0 77140.0 86285.0 78485.0 ;
      RECT  85580.0 79830.0 86285.0 78485.0 ;
      RECT  85580.0 79830.0 86285.0 81175.0 ;
      RECT  85580.0 82520.0 86285.0 81175.0 ;
      RECT  85580.0 82520.0 86285.0 83865.0 ;
      RECT  85580.0 85210.0 86285.0 83865.0 ;
      RECT  85580.0 85210.0 86285.0 86555.0 ;
      RECT  85580.0 87900.0 86285.0 86555.0 ;
      RECT  85580.0 87900.0 86285.0 89245.0 ;
      RECT  85580.0 90590.0 86285.0 89245.0 ;
      RECT  85580.0 90590.0 86285.0 91935.0 ;
      RECT  85580.0 93280.0 86285.0 91935.0 ;
      RECT  85580.0 93280.0 86285.0 94625.0 ;
      RECT  85580.0 95970.0 86285.0 94625.0 ;
      RECT  85580.0 95970.0 86285.0 97315.0 ;
      RECT  85580.0 98660.0 86285.0 97315.0 ;
      RECT  85580.0 98660.0 86285.0 100005.0 ;
      RECT  85580.0 101350.0 86285.0 100005.0 ;
      RECT  85580.0 101350.0 86285.0 102695.0 ;
      RECT  85580.0 104040.0 86285.0 102695.0 ;
      RECT  85580.0 104040.0 86285.0 105385.0 ;
      RECT  85580.0 106730.0 86285.0 105385.0 ;
      RECT  85580.0 106730.0 86285.0 108075.0 ;
      RECT  85580.0 109420.0 86285.0 108075.0 ;
      RECT  85580.0 109420.0 86285.0 110765.0 ;
      RECT  85580.0 112110.0 86285.0 110765.0 ;
      RECT  85580.0 112110.0 86285.0 113455.0 ;
      RECT  85580.0 114800.0 86285.0 113455.0 ;
      RECT  85580.0 114800.0 86285.0 116145.0 ;
      RECT  85580.0 117490.0 86285.0 116145.0 ;
      RECT  85580.0 117490.0 86285.0 118835.0 ;
      RECT  85580.0 120180.0 86285.0 118835.0 ;
      RECT  85580.0 120180.0 86285.0 121525.0 ;
      RECT  85580.0 122870.0 86285.0 121525.0 ;
      RECT  85580.0 122870.0 86285.0 124215.0 ;
      RECT  85580.0 125560.0 86285.0 124215.0 ;
      RECT  85580.0 125560.0 86285.0 126905.0 ;
      RECT  85580.0 128250.0 86285.0 126905.0 ;
      RECT  85580.0 128250.0 86285.0 129595.0 ;
      RECT  85580.0 130940.0 86285.0 129595.0 ;
      RECT  85580.0 130940.0 86285.0 132285.0 ;
      RECT  85580.0 133630.0 86285.0 132285.0 ;
      RECT  85580.0 133630.0 86285.0 134975.0 ;
      RECT  85580.0 136320.0 86285.0 134975.0 ;
      RECT  85580.0 136320.0 86285.0 137665.0 ;
      RECT  85580.0 139010.0 86285.0 137665.0 ;
      RECT  85580.0 139010.0 86285.0 140355.0 ;
      RECT  85580.0 141700.0 86285.0 140355.0 ;
      RECT  85580.0 141700.0 86285.0 143045.0 ;
      RECT  85580.0 144390.0 86285.0 143045.0 ;
      RECT  85580.0 144390.0 86285.0 145735.0 ;
      RECT  85580.0 147080.0 86285.0 145735.0 ;
      RECT  85580.0 147080.0 86285.0 148425.0 ;
      RECT  85580.0 149770.0 86285.0 148425.0 ;
      RECT  85580.0 149770.0 86285.0 151115.0 ;
      RECT  85580.0 152460.0 86285.0 151115.0 ;
      RECT  85580.0 152460.0 86285.0 153805.0 ;
      RECT  85580.0 155150.0 86285.0 153805.0 ;
      RECT  85580.0 155150.0 86285.0 156495.0 ;
      RECT  85580.0 157840.0 86285.0 156495.0 ;
      RECT  85580.0 157840.0 86285.0 159185.0 ;
      RECT  85580.0 160530.0 86285.0 159185.0 ;
      RECT  85580.0 160530.0 86285.0 161875.0 ;
      RECT  85580.0 163220.0 86285.0 161875.0 ;
      RECT  85580.0 163220.0 86285.0 164565.0 ;
      RECT  85580.0 165910.0 86285.0 164565.0 ;
      RECT  85580.0 165910.0 86285.0 167255.0 ;
      RECT  85580.0 168600.0 86285.0 167255.0 ;
      RECT  85580.0 168600.0 86285.0 169945.0 ;
      RECT  85580.0 171290.0 86285.0 169945.0 ;
      RECT  85580.0 171290.0 86285.0 172635.0 ;
      RECT  85580.0 173980.0 86285.0 172635.0 ;
      RECT  85580.0 173980.0 86285.0 175325.0 ;
      RECT  85580.0 176670.0 86285.0 175325.0 ;
      RECT  85580.0 176670.0 86285.0 178015.0 ;
      RECT  85580.0 179360.0 86285.0 178015.0 ;
      RECT  85580.0 179360.0 86285.0 180705.0 ;
      RECT  85580.0 182050.0 86285.0 180705.0 ;
      RECT  85580.0 182050.0 86285.0 183395.0 ;
      RECT  85580.0 184740.0 86285.0 183395.0 ;
      RECT  85580.0 184740.0 86285.0 186085.0 ;
      RECT  85580.0 187430.0 86285.0 186085.0 ;
      RECT  85580.0 187430.0 86285.0 188775.0 ;
      RECT  85580.0 190120.0 86285.0 188775.0 ;
      RECT  85580.0 190120.0 86285.0 191465.0 ;
      RECT  85580.0 192810.0 86285.0 191465.0 ;
      RECT  85580.0 192810.0 86285.0 194155.0 ;
      RECT  85580.0 195500.0 86285.0 194155.0 ;
      RECT  85580.0 195500.0 86285.0 196845.0 ;
      RECT  85580.0 198190.0 86285.0 196845.0 ;
      RECT  85580.0 198190.0 86285.0 199535.0 ;
      RECT  85580.0 200880.0 86285.0 199535.0 ;
      RECT  85580.0 200880.0 86285.0 202225.0 ;
      RECT  85580.0 203570.0 86285.0 202225.0 ;
      RECT  85580.0 203570.0 86285.0 204915.0 ;
      RECT  85580.0 206260.0 86285.0 204915.0 ;
      RECT  86285.0 34100.0 86990.0 35445.0 ;
      RECT  86285.0 36790.0 86990.0 35445.0 ;
      RECT  86285.0 36790.0 86990.0 38135.0 ;
      RECT  86285.0 39480.0 86990.0 38135.0 ;
      RECT  86285.0 39480.0 86990.0 40825.0 ;
      RECT  86285.0 42170.0 86990.0 40825.0 ;
      RECT  86285.0 42170.0 86990.0 43515.0 ;
      RECT  86285.0 44860.0 86990.0 43515.0 ;
      RECT  86285.0 44860.0 86990.0 46205.0 ;
      RECT  86285.0 47550.0 86990.0 46205.0 ;
      RECT  86285.0 47550.0 86990.0 48895.0 ;
      RECT  86285.0 50240.0 86990.0 48895.0 ;
      RECT  86285.0 50240.0 86990.0 51585.0 ;
      RECT  86285.0 52930.0 86990.0 51585.0 ;
      RECT  86285.0 52930.0 86990.0 54275.0 ;
      RECT  86285.0 55620.0 86990.0 54275.0 ;
      RECT  86285.0 55620.0 86990.0 56965.0 ;
      RECT  86285.0 58310.0 86990.0 56965.0 ;
      RECT  86285.0 58310.0 86990.0 59655.0 ;
      RECT  86285.0 61000.0 86990.0 59655.0 ;
      RECT  86285.0 61000.0 86990.0 62345.0 ;
      RECT  86285.0 63690.0 86990.0 62345.0 ;
      RECT  86285.0 63690.0 86990.0 65035.0 ;
      RECT  86285.0 66380.0 86990.0 65035.0 ;
      RECT  86285.0 66380.0 86990.0 67725.0 ;
      RECT  86285.0 69070.0 86990.0 67725.0 ;
      RECT  86285.0 69070.0 86990.0 70415.0 ;
      RECT  86285.0 71760.0 86990.0 70415.0 ;
      RECT  86285.0 71760.0 86990.0 73105.0 ;
      RECT  86285.0 74450.0 86990.0 73105.0 ;
      RECT  86285.0 74450.0 86990.0 75795.0 ;
      RECT  86285.0 77140.0 86990.0 75795.0 ;
      RECT  86285.0 77140.0 86990.0 78485.0 ;
      RECT  86285.0 79830.0 86990.0 78485.0 ;
      RECT  86285.0 79830.0 86990.0 81175.0 ;
      RECT  86285.0 82520.0 86990.0 81175.0 ;
      RECT  86285.0 82520.0 86990.0 83865.0 ;
      RECT  86285.0 85210.0 86990.0 83865.0 ;
      RECT  86285.0 85210.0 86990.0 86555.0 ;
      RECT  86285.0 87900.0 86990.0 86555.0 ;
      RECT  86285.0 87900.0 86990.0 89245.0 ;
      RECT  86285.0 90590.0 86990.0 89245.0 ;
      RECT  86285.0 90590.0 86990.0 91935.0 ;
      RECT  86285.0 93280.0 86990.0 91935.0 ;
      RECT  86285.0 93280.0 86990.0 94625.0 ;
      RECT  86285.0 95970.0 86990.0 94625.0 ;
      RECT  86285.0 95970.0 86990.0 97315.0 ;
      RECT  86285.0 98660.0 86990.0 97315.0 ;
      RECT  86285.0 98660.0 86990.0 100005.0 ;
      RECT  86285.0 101350.0 86990.0 100005.0 ;
      RECT  86285.0 101350.0 86990.0 102695.0 ;
      RECT  86285.0 104040.0 86990.0 102695.0 ;
      RECT  86285.0 104040.0 86990.0 105385.0 ;
      RECT  86285.0 106730.0 86990.0 105385.0 ;
      RECT  86285.0 106730.0 86990.0 108075.0 ;
      RECT  86285.0 109420.0 86990.0 108075.0 ;
      RECT  86285.0 109420.0 86990.0 110765.0 ;
      RECT  86285.0 112110.0 86990.0 110765.0 ;
      RECT  86285.0 112110.0 86990.0 113455.0 ;
      RECT  86285.0 114800.0 86990.0 113455.0 ;
      RECT  86285.0 114800.0 86990.0 116145.0 ;
      RECT  86285.0 117490.0 86990.0 116145.0 ;
      RECT  86285.0 117490.0 86990.0 118835.0 ;
      RECT  86285.0 120180.0 86990.0 118835.0 ;
      RECT  86285.0 120180.0 86990.0 121525.0 ;
      RECT  86285.0 122870.0 86990.0 121525.0 ;
      RECT  86285.0 122870.0 86990.0 124215.0 ;
      RECT  86285.0 125560.0 86990.0 124215.0 ;
      RECT  86285.0 125560.0 86990.0 126905.0 ;
      RECT  86285.0 128250.0 86990.0 126905.0 ;
      RECT  86285.0 128250.0 86990.0 129595.0 ;
      RECT  86285.0 130940.0 86990.0 129595.0 ;
      RECT  86285.0 130940.0 86990.0 132285.0 ;
      RECT  86285.0 133630.0 86990.0 132285.0 ;
      RECT  86285.0 133630.0 86990.0 134975.0 ;
      RECT  86285.0 136320.0 86990.0 134975.0 ;
      RECT  86285.0 136320.0 86990.0 137665.0 ;
      RECT  86285.0 139010.0 86990.0 137665.0 ;
      RECT  86285.0 139010.0 86990.0 140355.0 ;
      RECT  86285.0 141700.0 86990.0 140355.0 ;
      RECT  86285.0 141700.0 86990.0 143045.0 ;
      RECT  86285.0 144390.0 86990.0 143045.0 ;
      RECT  86285.0 144390.0 86990.0 145735.0 ;
      RECT  86285.0 147080.0 86990.0 145735.0 ;
      RECT  86285.0 147080.0 86990.0 148425.0 ;
      RECT  86285.0 149770.0 86990.0 148425.0 ;
      RECT  86285.0 149770.0 86990.0 151115.0 ;
      RECT  86285.0 152460.0 86990.0 151115.0 ;
      RECT  86285.0 152460.0 86990.0 153805.0 ;
      RECT  86285.0 155150.0 86990.0 153805.0 ;
      RECT  86285.0 155150.0 86990.0 156495.0 ;
      RECT  86285.0 157840.0 86990.0 156495.0 ;
      RECT  86285.0 157840.0 86990.0 159185.0 ;
      RECT  86285.0 160530.0 86990.0 159185.0 ;
      RECT  86285.0 160530.0 86990.0 161875.0 ;
      RECT  86285.0 163220.0 86990.0 161875.0 ;
      RECT  86285.0 163220.0 86990.0 164565.0 ;
      RECT  86285.0 165910.0 86990.0 164565.0 ;
      RECT  86285.0 165910.0 86990.0 167255.0 ;
      RECT  86285.0 168600.0 86990.0 167255.0 ;
      RECT  86285.0 168600.0 86990.0 169945.0 ;
      RECT  86285.0 171290.0 86990.0 169945.0 ;
      RECT  86285.0 171290.0 86990.0 172635.0 ;
      RECT  86285.0 173980.0 86990.0 172635.0 ;
      RECT  86285.0 173980.0 86990.0 175325.0 ;
      RECT  86285.0 176670.0 86990.0 175325.0 ;
      RECT  86285.0 176670.0 86990.0 178015.0 ;
      RECT  86285.0 179360.0 86990.0 178015.0 ;
      RECT  86285.0 179360.0 86990.0 180705.0 ;
      RECT  86285.0 182050.0 86990.0 180705.0 ;
      RECT  86285.0 182050.0 86990.0 183395.0 ;
      RECT  86285.0 184740.0 86990.0 183395.0 ;
      RECT  86285.0 184740.0 86990.0 186085.0 ;
      RECT  86285.0 187430.0 86990.0 186085.0 ;
      RECT  86285.0 187430.0 86990.0 188775.0 ;
      RECT  86285.0 190120.0 86990.0 188775.0 ;
      RECT  86285.0 190120.0 86990.0 191465.0 ;
      RECT  86285.0 192810.0 86990.0 191465.0 ;
      RECT  86285.0 192810.0 86990.0 194155.0 ;
      RECT  86285.0 195500.0 86990.0 194155.0 ;
      RECT  86285.0 195500.0 86990.0 196845.0 ;
      RECT  86285.0 198190.0 86990.0 196845.0 ;
      RECT  86285.0 198190.0 86990.0 199535.0 ;
      RECT  86285.0 200880.0 86990.0 199535.0 ;
      RECT  86285.0 200880.0 86990.0 202225.0 ;
      RECT  86285.0 203570.0 86990.0 202225.0 ;
      RECT  86285.0 203570.0 86990.0 204915.0 ;
      RECT  86285.0 206260.0 86990.0 204915.0 ;
      RECT  86990.0 34100.0 87695.0 35445.0 ;
      RECT  86990.0 36790.0 87695.0 35445.0 ;
      RECT  86990.0 36790.0 87695.0 38135.0 ;
      RECT  86990.0 39480.0 87695.0 38135.0 ;
      RECT  86990.0 39480.0 87695.0 40825.0 ;
      RECT  86990.0 42170.0 87695.0 40825.0 ;
      RECT  86990.0 42170.0 87695.0 43515.0 ;
      RECT  86990.0 44860.0 87695.0 43515.0 ;
      RECT  86990.0 44860.0 87695.0 46205.0 ;
      RECT  86990.0 47550.0 87695.0 46205.0 ;
      RECT  86990.0 47550.0 87695.0 48895.0 ;
      RECT  86990.0 50240.0 87695.0 48895.0 ;
      RECT  86990.0 50240.0 87695.0 51585.0 ;
      RECT  86990.0 52930.0 87695.0 51585.0 ;
      RECT  86990.0 52930.0 87695.0 54275.0 ;
      RECT  86990.0 55620.0 87695.0 54275.0 ;
      RECT  86990.0 55620.0 87695.0 56965.0 ;
      RECT  86990.0 58310.0 87695.0 56965.0 ;
      RECT  86990.0 58310.0 87695.0 59655.0 ;
      RECT  86990.0 61000.0 87695.0 59655.0 ;
      RECT  86990.0 61000.0 87695.0 62345.0 ;
      RECT  86990.0 63690.0 87695.0 62345.0 ;
      RECT  86990.0 63690.0 87695.0 65035.0 ;
      RECT  86990.0 66380.0 87695.0 65035.0 ;
      RECT  86990.0 66380.0 87695.0 67725.0 ;
      RECT  86990.0 69070.0 87695.0 67725.0 ;
      RECT  86990.0 69070.0 87695.0 70415.0 ;
      RECT  86990.0 71760.0 87695.0 70415.0 ;
      RECT  86990.0 71760.0 87695.0 73105.0 ;
      RECT  86990.0 74450.0 87695.0 73105.0 ;
      RECT  86990.0 74450.0 87695.0 75795.0 ;
      RECT  86990.0 77140.0 87695.0 75795.0 ;
      RECT  86990.0 77140.0 87695.0 78485.0 ;
      RECT  86990.0 79830.0 87695.0 78485.0 ;
      RECT  86990.0 79830.0 87695.0 81175.0 ;
      RECT  86990.0 82520.0 87695.0 81175.0 ;
      RECT  86990.0 82520.0 87695.0 83865.0 ;
      RECT  86990.0 85210.0 87695.0 83865.0 ;
      RECT  86990.0 85210.0 87695.0 86555.0 ;
      RECT  86990.0 87900.0 87695.0 86555.0 ;
      RECT  86990.0 87900.0 87695.0 89245.0 ;
      RECT  86990.0 90590.0 87695.0 89245.0 ;
      RECT  86990.0 90590.0 87695.0 91935.0 ;
      RECT  86990.0 93280.0 87695.0 91935.0 ;
      RECT  86990.0 93280.0 87695.0 94625.0 ;
      RECT  86990.0 95970.0 87695.0 94625.0 ;
      RECT  86990.0 95970.0 87695.0 97315.0 ;
      RECT  86990.0 98660.0 87695.0 97315.0 ;
      RECT  86990.0 98660.0 87695.0 100005.0 ;
      RECT  86990.0 101350.0 87695.0 100005.0 ;
      RECT  86990.0 101350.0 87695.0 102695.0 ;
      RECT  86990.0 104040.0 87695.0 102695.0 ;
      RECT  86990.0 104040.0 87695.0 105385.0 ;
      RECT  86990.0 106730.0 87695.0 105385.0 ;
      RECT  86990.0 106730.0 87695.0 108075.0 ;
      RECT  86990.0 109420.0 87695.0 108075.0 ;
      RECT  86990.0 109420.0 87695.0 110765.0 ;
      RECT  86990.0 112110.0 87695.0 110765.0 ;
      RECT  86990.0 112110.0 87695.0 113455.0 ;
      RECT  86990.0 114800.0 87695.0 113455.0 ;
      RECT  86990.0 114800.0 87695.0 116145.0 ;
      RECT  86990.0 117490.0 87695.0 116145.0 ;
      RECT  86990.0 117490.0 87695.0 118835.0 ;
      RECT  86990.0 120180.0 87695.0 118835.0 ;
      RECT  86990.0 120180.0 87695.0 121525.0 ;
      RECT  86990.0 122870.0 87695.0 121525.0 ;
      RECT  86990.0 122870.0 87695.0 124215.0 ;
      RECT  86990.0 125560.0 87695.0 124215.0 ;
      RECT  86990.0 125560.0 87695.0 126905.0 ;
      RECT  86990.0 128250.0 87695.0 126905.0 ;
      RECT  86990.0 128250.0 87695.0 129595.0 ;
      RECT  86990.0 130940.0 87695.0 129595.0 ;
      RECT  86990.0 130940.0 87695.0 132285.0 ;
      RECT  86990.0 133630.0 87695.0 132285.0 ;
      RECT  86990.0 133630.0 87695.0 134975.0 ;
      RECT  86990.0 136320.0 87695.0 134975.0 ;
      RECT  86990.0 136320.0 87695.0 137665.0 ;
      RECT  86990.0 139010.0 87695.0 137665.0 ;
      RECT  86990.0 139010.0 87695.0 140355.0 ;
      RECT  86990.0 141700.0 87695.0 140355.0 ;
      RECT  86990.0 141700.0 87695.0 143045.0 ;
      RECT  86990.0 144390.0 87695.0 143045.0 ;
      RECT  86990.0 144390.0 87695.0 145735.0 ;
      RECT  86990.0 147080.0 87695.0 145735.0 ;
      RECT  86990.0 147080.0 87695.0 148425.0 ;
      RECT  86990.0 149770.0 87695.0 148425.0 ;
      RECT  86990.0 149770.0 87695.0 151115.0 ;
      RECT  86990.0 152460.0 87695.0 151115.0 ;
      RECT  86990.0 152460.0 87695.0 153805.0 ;
      RECT  86990.0 155150.0 87695.0 153805.0 ;
      RECT  86990.0 155150.0 87695.0 156495.0 ;
      RECT  86990.0 157840.0 87695.0 156495.0 ;
      RECT  86990.0 157840.0 87695.0 159185.0 ;
      RECT  86990.0 160530.0 87695.0 159185.0 ;
      RECT  86990.0 160530.0 87695.0 161875.0 ;
      RECT  86990.0 163220.0 87695.0 161875.0 ;
      RECT  86990.0 163220.0 87695.0 164565.0 ;
      RECT  86990.0 165910.0 87695.0 164565.0 ;
      RECT  86990.0 165910.0 87695.0 167255.0 ;
      RECT  86990.0 168600.0 87695.0 167255.0 ;
      RECT  86990.0 168600.0 87695.0 169945.0 ;
      RECT  86990.0 171290.0 87695.0 169945.0 ;
      RECT  86990.0 171290.0 87695.0 172635.0 ;
      RECT  86990.0 173980.0 87695.0 172635.0 ;
      RECT  86990.0 173980.0 87695.0 175325.0 ;
      RECT  86990.0 176670.0 87695.0 175325.0 ;
      RECT  86990.0 176670.0 87695.0 178015.0 ;
      RECT  86990.0 179360.0 87695.0 178015.0 ;
      RECT  86990.0 179360.0 87695.0 180705.0 ;
      RECT  86990.0 182050.0 87695.0 180705.0 ;
      RECT  86990.0 182050.0 87695.0 183395.0 ;
      RECT  86990.0 184740.0 87695.0 183395.0 ;
      RECT  86990.0 184740.0 87695.0 186085.0 ;
      RECT  86990.0 187430.0 87695.0 186085.0 ;
      RECT  86990.0 187430.0 87695.0 188775.0 ;
      RECT  86990.0 190120.0 87695.0 188775.0 ;
      RECT  86990.0 190120.0 87695.0 191465.0 ;
      RECT  86990.0 192810.0 87695.0 191465.0 ;
      RECT  86990.0 192810.0 87695.0 194155.0 ;
      RECT  86990.0 195500.0 87695.0 194155.0 ;
      RECT  86990.0 195500.0 87695.0 196845.0 ;
      RECT  86990.0 198190.0 87695.0 196845.0 ;
      RECT  86990.0 198190.0 87695.0 199535.0 ;
      RECT  86990.0 200880.0 87695.0 199535.0 ;
      RECT  86990.0 200880.0 87695.0 202225.0 ;
      RECT  86990.0 203570.0 87695.0 202225.0 ;
      RECT  86990.0 203570.0 87695.0 204915.0 ;
      RECT  86990.0 206260.0 87695.0 204915.0 ;
      RECT  87695.0 34100.0 88400.0 35445.0 ;
      RECT  87695.0 36790.0 88400.0 35445.0 ;
      RECT  87695.0 36790.0 88400.0 38135.0 ;
      RECT  87695.0 39480.0 88400.0 38135.0 ;
      RECT  87695.0 39480.0 88400.0 40825.0 ;
      RECT  87695.0 42170.0 88400.0 40825.0 ;
      RECT  87695.0 42170.0 88400.0 43515.0 ;
      RECT  87695.0 44860.0 88400.0 43515.0 ;
      RECT  87695.0 44860.0 88400.0 46205.0 ;
      RECT  87695.0 47550.0 88400.0 46205.0 ;
      RECT  87695.0 47550.0 88400.0 48895.0 ;
      RECT  87695.0 50240.0 88400.0 48895.0 ;
      RECT  87695.0 50240.0 88400.0 51585.0 ;
      RECT  87695.0 52930.0 88400.0 51585.0 ;
      RECT  87695.0 52930.0 88400.0 54275.0 ;
      RECT  87695.0 55620.0 88400.0 54275.0 ;
      RECT  87695.0 55620.0 88400.0 56965.0 ;
      RECT  87695.0 58310.0 88400.0 56965.0 ;
      RECT  87695.0 58310.0 88400.0 59655.0 ;
      RECT  87695.0 61000.0 88400.0 59655.0 ;
      RECT  87695.0 61000.0 88400.0 62345.0 ;
      RECT  87695.0 63690.0 88400.0 62345.0 ;
      RECT  87695.0 63690.0 88400.0 65035.0 ;
      RECT  87695.0 66380.0 88400.0 65035.0 ;
      RECT  87695.0 66380.0 88400.0 67725.0 ;
      RECT  87695.0 69070.0 88400.0 67725.0 ;
      RECT  87695.0 69070.0 88400.0 70415.0 ;
      RECT  87695.0 71760.0 88400.0 70415.0 ;
      RECT  87695.0 71760.0 88400.0 73105.0 ;
      RECT  87695.0 74450.0 88400.0 73105.0 ;
      RECT  87695.0 74450.0 88400.0 75795.0 ;
      RECT  87695.0 77140.0 88400.0 75795.0 ;
      RECT  87695.0 77140.0 88400.0 78485.0 ;
      RECT  87695.0 79830.0 88400.0 78485.0 ;
      RECT  87695.0 79830.0 88400.0 81175.0 ;
      RECT  87695.0 82520.0 88400.0 81175.0 ;
      RECT  87695.0 82520.0 88400.0 83865.0 ;
      RECT  87695.0 85210.0 88400.0 83865.0 ;
      RECT  87695.0 85210.0 88400.0 86555.0 ;
      RECT  87695.0 87900.0 88400.0 86555.0 ;
      RECT  87695.0 87900.0 88400.0 89245.0 ;
      RECT  87695.0 90590.0 88400.0 89245.0 ;
      RECT  87695.0 90590.0 88400.0 91935.0 ;
      RECT  87695.0 93280.0 88400.0 91935.0 ;
      RECT  87695.0 93280.0 88400.0 94625.0 ;
      RECT  87695.0 95970.0 88400.0 94625.0 ;
      RECT  87695.0 95970.0 88400.0 97315.0 ;
      RECT  87695.0 98660.0 88400.0 97315.0 ;
      RECT  87695.0 98660.0 88400.0 100005.0 ;
      RECT  87695.0 101350.0 88400.0 100005.0 ;
      RECT  87695.0 101350.0 88400.0 102695.0 ;
      RECT  87695.0 104040.0 88400.0 102695.0 ;
      RECT  87695.0 104040.0 88400.0 105385.0 ;
      RECT  87695.0 106730.0 88400.0 105385.0 ;
      RECT  87695.0 106730.0 88400.0 108075.0 ;
      RECT  87695.0 109420.0 88400.0 108075.0 ;
      RECT  87695.0 109420.0 88400.0 110765.0 ;
      RECT  87695.0 112110.0 88400.0 110765.0 ;
      RECT  87695.0 112110.0 88400.0 113455.0 ;
      RECT  87695.0 114800.0 88400.0 113455.0 ;
      RECT  87695.0 114800.0 88400.0 116145.0 ;
      RECT  87695.0 117490.0 88400.0 116145.0 ;
      RECT  87695.0 117490.0 88400.0 118835.0 ;
      RECT  87695.0 120180.0 88400.0 118835.0 ;
      RECT  87695.0 120180.0 88400.0 121525.0 ;
      RECT  87695.0 122870.0 88400.0 121525.0 ;
      RECT  87695.0 122870.0 88400.0 124215.0 ;
      RECT  87695.0 125560.0 88400.0 124215.0 ;
      RECT  87695.0 125560.0 88400.0 126905.0 ;
      RECT  87695.0 128250.0 88400.0 126905.0 ;
      RECT  87695.0 128250.0 88400.0 129595.0 ;
      RECT  87695.0 130940.0 88400.0 129595.0 ;
      RECT  87695.0 130940.0 88400.0 132285.0 ;
      RECT  87695.0 133630.0 88400.0 132285.0 ;
      RECT  87695.0 133630.0 88400.0 134975.0 ;
      RECT  87695.0 136320.0 88400.0 134975.0 ;
      RECT  87695.0 136320.0 88400.0 137665.0 ;
      RECT  87695.0 139010.0 88400.0 137665.0 ;
      RECT  87695.0 139010.0 88400.0 140355.0 ;
      RECT  87695.0 141700.0 88400.0 140355.0 ;
      RECT  87695.0 141700.0 88400.0 143045.0 ;
      RECT  87695.0 144390.0 88400.0 143045.0 ;
      RECT  87695.0 144390.0 88400.0 145735.0 ;
      RECT  87695.0 147080.0 88400.0 145735.0 ;
      RECT  87695.0 147080.0 88400.0 148425.0 ;
      RECT  87695.0 149770.0 88400.0 148425.0 ;
      RECT  87695.0 149770.0 88400.0 151115.0 ;
      RECT  87695.0 152460.0 88400.0 151115.0 ;
      RECT  87695.0 152460.0 88400.0 153805.0 ;
      RECT  87695.0 155150.0 88400.0 153805.0 ;
      RECT  87695.0 155150.0 88400.0 156495.0 ;
      RECT  87695.0 157840.0 88400.0 156495.0 ;
      RECT  87695.0 157840.0 88400.0 159185.0 ;
      RECT  87695.0 160530.0 88400.0 159185.0 ;
      RECT  87695.0 160530.0 88400.0 161875.0 ;
      RECT  87695.0 163220.0 88400.0 161875.0 ;
      RECT  87695.0 163220.0 88400.0 164565.0 ;
      RECT  87695.0 165910.0 88400.0 164565.0 ;
      RECT  87695.0 165910.0 88400.0 167255.0 ;
      RECT  87695.0 168600.0 88400.0 167255.0 ;
      RECT  87695.0 168600.0 88400.0 169945.0 ;
      RECT  87695.0 171290.0 88400.0 169945.0 ;
      RECT  87695.0 171290.0 88400.0 172635.0 ;
      RECT  87695.0 173980.0 88400.0 172635.0 ;
      RECT  87695.0 173980.0 88400.0 175325.0 ;
      RECT  87695.0 176670.0 88400.0 175325.0 ;
      RECT  87695.0 176670.0 88400.0 178015.0 ;
      RECT  87695.0 179360.0 88400.0 178015.0 ;
      RECT  87695.0 179360.0 88400.0 180705.0 ;
      RECT  87695.0 182050.0 88400.0 180705.0 ;
      RECT  87695.0 182050.0 88400.0 183395.0 ;
      RECT  87695.0 184740.0 88400.0 183395.0 ;
      RECT  87695.0 184740.0 88400.0 186085.0 ;
      RECT  87695.0 187430.0 88400.0 186085.0 ;
      RECT  87695.0 187430.0 88400.0 188775.0 ;
      RECT  87695.0 190120.0 88400.0 188775.0 ;
      RECT  87695.0 190120.0 88400.0 191465.0 ;
      RECT  87695.0 192810.0 88400.0 191465.0 ;
      RECT  87695.0 192810.0 88400.0 194155.0 ;
      RECT  87695.0 195500.0 88400.0 194155.0 ;
      RECT  87695.0 195500.0 88400.0 196845.0 ;
      RECT  87695.0 198190.0 88400.0 196845.0 ;
      RECT  87695.0 198190.0 88400.0 199535.0 ;
      RECT  87695.0 200880.0 88400.0 199535.0 ;
      RECT  87695.0 200880.0 88400.0 202225.0 ;
      RECT  87695.0 203570.0 88400.0 202225.0 ;
      RECT  87695.0 203570.0 88400.0 204915.0 ;
      RECT  87695.0 206260.0 88400.0 204915.0 ;
      RECT  88400.0 34100.0 89105.0 35445.0 ;
      RECT  88400.0 36790.0 89105.0 35445.0 ;
      RECT  88400.0 36790.0 89105.0 38135.0 ;
      RECT  88400.0 39480.0 89105.0 38135.0 ;
      RECT  88400.0 39480.0 89105.0 40825.0 ;
      RECT  88400.0 42170.0 89105.0 40825.0 ;
      RECT  88400.0 42170.0 89105.0 43515.0 ;
      RECT  88400.0 44860.0 89105.0 43515.0 ;
      RECT  88400.0 44860.0 89105.0 46205.0 ;
      RECT  88400.0 47550.0 89105.0 46205.0 ;
      RECT  88400.0 47550.0 89105.0 48895.0 ;
      RECT  88400.0 50240.0 89105.0 48895.0 ;
      RECT  88400.0 50240.0 89105.0 51585.0 ;
      RECT  88400.0 52930.0 89105.0 51585.0 ;
      RECT  88400.0 52930.0 89105.0 54275.0 ;
      RECT  88400.0 55620.0 89105.0 54275.0 ;
      RECT  88400.0 55620.0 89105.0 56965.0 ;
      RECT  88400.0 58310.0 89105.0 56965.0 ;
      RECT  88400.0 58310.0 89105.0 59655.0 ;
      RECT  88400.0 61000.0 89105.0 59655.0 ;
      RECT  88400.0 61000.0 89105.0 62345.0 ;
      RECT  88400.0 63690.0 89105.0 62345.0 ;
      RECT  88400.0 63690.0 89105.0 65035.0 ;
      RECT  88400.0 66380.0 89105.0 65035.0 ;
      RECT  88400.0 66380.0 89105.0 67725.0 ;
      RECT  88400.0 69070.0 89105.0 67725.0 ;
      RECT  88400.0 69070.0 89105.0 70415.0 ;
      RECT  88400.0 71760.0 89105.0 70415.0 ;
      RECT  88400.0 71760.0 89105.0 73105.0 ;
      RECT  88400.0 74450.0 89105.0 73105.0 ;
      RECT  88400.0 74450.0 89105.0 75795.0 ;
      RECT  88400.0 77140.0 89105.0 75795.0 ;
      RECT  88400.0 77140.0 89105.0 78485.0 ;
      RECT  88400.0 79830.0 89105.0 78485.0 ;
      RECT  88400.0 79830.0 89105.0 81175.0 ;
      RECT  88400.0 82520.0 89105.0 81175.0 ;
      RECT  88400.0 82520.0 89105.0 83865.0 ;
      RECT  88400.0 85210.0 89105.0 83865.0 ;
      RECT  88400.0 85210.0 89105.0 86555.0 ;
      RECT  88400.0 87900.0 89105.0 86555.0 ;
      RECT  88400.0 87900.0 89105.0 89245.0 ;
      RECT  88400.0 90590.0 89105.0 89245.0 ;
      RECT  88400.0 90590.0 89105.0 91935.0 ;
      RECT  88400.0 93280.0 89105.0 91935.0 ;
      RECT  88400.0 93280.0 89105.0 94625.0 ;
      RECT  88400.0 95970.0 89105.0 94625.0 ;
      RECT  88400.0 95970.0 89105.0 97315.0 ;
      RECT  88400.0 98660.0 89105.0 97315.0 ;
      RECT  88400.0 98660.0 89105.0 100005.0 ;
      RECT  88400.0 101350.0 89105.0 100005.0 ;
      RECT  88400.0 101350.0 89105.0 102695.0 ;
      RECT  88400.0 104040.0 89105.0 102695.0 ;
      RECT  88400.0 104040.0 89105.0 105385.0 ;
      RECT  88400.0 106730.0 89105.0 105385.0 ;
      RECT  88400.0 106730.0 89105.0 108075.0 ;
      RECT  88400.0 109420.0 89105.0 108075.0 ;
      RECT  88400.0 109420.0 89105.0 110765.0 ;
      RECT  88400.0 112110.0 89105.0 110765.0 ;
      RECT  88400.0 112110.0 89105.0 113455.0 ;
      RECT  88400.0 114800.0 89105.0 113455.0 ;
      RECT  88400.0 114800.0 89105.0 116145.0 ;
      RECT  88400.0 117490.0 89105.0 116145.0 ;
      RECT  88400.0 117490.0 89105.0 118835.0 ;
      RECT  88400.0 120180.0 89105.0 118835.0 ;
      RECT  88400.0 120180.0 89105.0 121525.0 ;
      RECT  88400.0 122870.0 89105.0 121525.0 ;
      RECT  88400.0 122870.0 89105.0 124215.0 ;
      RECT  88400.0 125560.0 89105.0 124215.0 ;
      RECT  88400.0 125560.0 89105.0 126905.0 ;
      RECT  88400.0 128250.0 89105.0 126905.0 ;
      RECT  88400.0 128250.0 89105.0 129595.0 ;
      RECT  88400.0 130940.0 89105.0 129595.0 ;
      RECT  88400.0 130940.0 89105.0 132285.0 ;
      RECT  88400.0 133630.0 89105.0 132285.0 ;
      RECT  88400.0 133630.0 89105.0 134975.0 ;
      RECT  88400.0 136320.0 89105.0 134975.0 ;
      RECT  88400.0 136320.0 89105.0 137665.0 ;
      RECT  88400.0 139010.0 89105.0 137665.0 ;
      RECT  88400.0 139010.0 89105.0 140355.0 ;
      RECT  88400.0 141700.0 89105.0 140355.0 ;
      RECT  88400.0 141700.0 89105.0 143045.0 ;
      RECT  88400.0 144390.0 89105.0 143045.0 ;
      RECT  88400.0 144390.0 89105.0 145735.0 ;
      RECT  88400.0 147080.0 89105.0 145735.0 ;
      RECT  88400.0 147080.0 89105.0 148425.0 ;
      RECT  88400.0 149770.0 89105.0 148425.0 ;
      RECT  88400.0 149770.0 89105.0 151115.0 ;
      RECT  88400.0 152460.0 89105.0 151115.0 ;
      RECT  88400.0 152460.0 89105.0 153805.0 ;
      RECT  88400.0 155150.0 89105.0 153805.0 ;
      RECT  88400.0 155150.0 89105.0 156495.0 ;
      RECT  88400.0 157840.0 89105.0 156495.0 ;
      RECT  88400.0 157840.0 89105.0 159185.0 ;
      RECT  88400.0 160530.0 89105.0 159185.0 ;
      RECT  88400.0 160530.0 89105.0 161875.0 ;
      RECT  88400.0 163220.0 89105.0 161875.0 ;
      RECT  88400.0 163220.0 89105.0 164565.0 ;
      RECT  88400.0 165910.0 89105.0 164565.0 ;
      RECT  88400.0 165910.0 89105.0 167255.0 ;
      RECT  88400.0 168600.0 89105.0 167255.0 ;
      RECT  88400.0 168600.0 89105.0 169945.0 ;
      RECT  88400.0 171290.0 89105.0 169945.0 ;
      RECT  88400.0 171290.0 89105.0 172635.0 ;
      RECT  88400.0 173980.0 89105.0 172635.0 ;
      RECT  88400.0 173980.0 89105.0 175325.0 ;
      RECT  88400.0 176670.0 89105.0 175325.0 ;
      RECT  88400.0 176670.0 89105.0 178015.0 ;
      RECT  88400.0 179360.0 89105.0 178015.0 ;
      RECT  88400.0 179360.0 89105.0 180705.0 ;
      RECT  88400.0 182050.0 89105.0 180705.0 ;
      RECT  88400.0 182050.0 89105.0 183395.0 ;
      RECT  88400.0 184740.0 89105.0 183395.0 ;
      RECT  88400.0 184740.0 89105.0 186085.0 ;
      RECT  88400.0 187430.0 89105.0 186085.0 ;
      RECT  88400.0 187430.0 89105.0 188775.0 ;
      RECT  88400.0 190120.0 89105.0 188775.0 ;
      RECT  88400.0 190120.0 89105.0 191465.0 ;
      RECT  88400.0 192810.0 89105.0 191465.0 ;
      RECT  88400.0 192810.0 89105.0 194155.0 ;
      RECT  88400.0 195500.0 89105.0 194155.0 ;
      RECT  88400.0 195500.0 89105.0 196845.0 ;
      RECT  88400.0 198190.0 89105.0 196845.0 ;
      RECT  88400.0 198190.0 89105.0 199535.0 ;
      RECT  88400.0 200880.0 89105.0 199535.0 ;
      RECT  88400.0 200880.0 89105.0 202225.0 ;
      RECT  88400.0 203570.0 89105.0 202225.0 ;
      RECT  88400.0 203570.0 89105.0 204915.0 ;
      RECT  88400.0 206260.0 89105.0 204915.0 ;
      RECT  89105.0 34100.0 89810.0 35445.0 ;
      RECT  89105.0 36790.0 89810.0 35445.0 ;
      RECT  89105.0 36790.0 89810.0 38135.0 ;
      RECT  89105.0 39480.0 89810.0 38135.0 ;
      RECT  89105.0 39480.0 89810.0 40825.0 ;
      RECT  89105.0 42170.0 89810.0 40825.0 ;
      RECT  89105.0 42170.0 89810.0 43515.0 ;
      RECT  89105.0 44860.0 89810.0 43515.0 ;
      RECT  89105.0 44860.0 89810.0 46205.0 ;
      RECT  89105.0 47550.0 89810.0 46205.0 ;
      RECT  89105.0 47550.0 89810.0 48895.0 ;
      RECT  89105.0 50240.0 89810.0 48895.0 ;
      RECT  89105.0 50240.0 89810.0 51585.0 ;
      RECT  89105.0 52930.0 89810.0 51585.0 ;
      RECT  89105.0 52930.0 89810.0 54275.0 ;
      RECT  89105.0 55620.0 89810.0 54275.0 ;
      RECT  89105.0 55620.0 89810.0 56965.0 ;
      RECT  89105.0 58310.0 89810.0 56965.0 ;
      RECT  89105.0 58310.0 89810.0 59655.0 ;
      RECT  89105.0 61000.0 89810.0 59655.0 ;
      RECT  89105.0 61000.0 89810.0 62345.0 ;
      RECT  89105.0 63690.0 89810.0 62345.0 ;
      RECT  89105.0 63690.0 89810.0 65035.0 ;
      RECT  89105.0 66380.0 89810.0 65035.0 ;
      RECT  89105.0 66380.0 89810.0 67725.0 ;
      RECT  89105.0 69070.0 89810.0 67725.0 ;
      RECT  89105.0 69070.0 89810.0 70415.0 ;
      RECT  89105.0 71760.0 89810.0 70415.0 ;
      RECT  89105.0 71760.0 89810.0 73105.0 ;
      RECT  89105.0 74450.0 89810.0 73105.0 ;
      RECT  89105.0 74450.0 89810.0 75795.0 ;
      RECT  89105.0 77140.0 89810.0 75795.0 ;
      RECT  89105.0 77140.0 89810.0 78485.0 ;
      RECT  89105.0 79830.0 89810.0 78485.0 ;
      RECT  89105.0 79830.0 89810.0 81175.0 ;
      RECT  89105.0 82520.0 89810.0 81175.0 ;
      RECT  89105.0 82520.0 89810.0 83865.0 ;
      RECT  89105.0 85210.0 89810.0 83865.0 ;
      RECT  89105.0 85210.0 89810.0 86555.0 ;
      RECT  89105.0 87900.0 89810.0 86555.0 ;
      RECT  89105.0 87900.0 89810.0 89245.0 ;
      RECT  89105.0 90590.0 89810.0 89245.0 ;
      RECT  89105.0 90590.0 89810.0 91935.0 ;
      RECT  89105.0 93280.0 89810.0 91935.0 ;
      RECT  89105.0 93280.0 89810.0 94625.0 ;
      RECT  89105.0 95970.0 89810.0 94625.0 ;
      RECT  89105.0 95970.0 89810.0 97315.0 ;
      RECT  89105.0 98660.0 89810.0 97315.0 ;
      RECT  89105.0 98660.0 89810.0 100005.0 ;
      RECT  89105.0 101350.0 89810.0 100005.0 ;
      RECT  89105.0 101350.0 89810.0 102695.0 ;
      RECT  89105.0 104040.0 89810.0 102695.0 ;
      RECT  89105.0 104040.0 89810.0 105385.0 ;
      RECT  89105.0 106730.0 89810.0 105385.0 ;
      RECT  89105.0 106730.0 89810.0 108075.0 ;
      RECT  89105.0 109420.0 89810.0 108075.0 ;
      RECT  89105.0 109420.0 89810.0 110765.0 ;
      RECT  89105.0 112110.0 89810.0 110765.0 ;
      RECT  89105.0 112110.0 89810.0 113455.0 ;
      RECT  89105.0 114800.0 89810.0 113455.0 ;
      RECT  89105.0 114800.0 89810.0 116145.0 ;
      RECT  89105.0 117490.0 89810.0 116145.0 ;
      RECT  89105.0 117490.0 89810.0 118835.0 ;
      RECT  89105.0 120180.0 89810.0 118835.0 ;
      RECT  89105.0 120180.0 89810.0 121525.0 ;
      RECT  89105.0 122870.0 89810.0 121525.0 ;
      RECT  89105.0 122870.0 89810.0 124215.0 ;
      RECT  89105.0 125560.0 89810.0 124215.0 ;
      RECT  89105.0 125560.0 89810.0 126905.0 ;
      RECT  89105.0 128250.0 89810.0 126905.0 ;
      RECT  89105.0 128250.0 89810.0 129595.0 ;
      RECT  89105.0 130940.0 89810.0 129595.0 ;
      RECT  89105.0 130940.0 89810.0 132285.0 ;
      RECT  89105.0 133630.0 89810.0 132285.0 ;
      RECT  89105.0 133630.0 89810.0 134975.0 ;
      RECT  89105.0 136320.0 89810.0 134975.0 ;
      RECT  89105.0 136320.0 89810.0 137665.0 ;
      RECT  89105.0 139010.0 89810.0 137665.0 ;
      RECT  89105.0 139010.0 89810.0 140355.0 ;
      RECT  89105.0 141700.0 89810.0 140355.0 ;
      RECT  89105.0 141700.0 89810.0 143045.0 ;
      RECT  89105.0 144390.0 89810.0 143045.0 ;
      RECT  89105.0 144390.0 89810.0 145735.0 ;
      RECT  89105.0 147080.0 89810.0 145735.0 ;
      RECT  89105.0 147080.0 89810.0 148425.0 ;
      RECT  89105.0 149770.0 89810.0 148425.0 ;
      RECT  89105.0 149770.0 89810.0 151115.0 ;
      RECT  89105.0 152460.0 89810.0 151115.0 ;
      RECT  89105.0 152460.0 89810.0 153805.0 ;
      RECT  89105.0 155150.0 89810.0 153805.0 ;
      RECT  89105.0 155150.0 89810.0 156495.0 ;
      RECT  89105.0 157840.0 89810.0 156495.0 ;
      RECT  89105.0 157840.0 89810.0 159185.0 ;
      RECT  89105.0 160530.0 89810.0 159185.0 ;
      RECT  89105.0 160530.0 89810.0 161875.0 ;
      RECT  89105.0 163220.0 89810.0 161875.0 ;
      RECT  89105.0 163220.0 89810.0 164565.0 ;
      RECT  89105.0 165910.0 89810.0 164565.0 ;
      RECT  89105.0 165910.0 89810.0 167255.0 ;
      RECT  89105.0 168600.0 89810.0 167255.0 ;
      RECT  89105.0 168600.0 89810.0 169945.0 ;
      RECT  89105.0 171290.0 89810.0 169945.0 ;
      RECT  89105.0 171290.0 89810.0 172635.0 ;
      RECT  89105.0 173980.0 89810.0 172635.0 ;
      RECT  89105.0 173980.0 89810.0 175325.0 ;
      RECT  89105.0 176670.0 89810.0 175325.0 ;
      RECT  89105.0 176670.0 89810.0 178015.0 ;
      RECT  89105.0 179360.0 89810.0 178015.0 ;
      RECT  89105.0 179360.0 89810.0 180705.0 ;
      RECT  89105.0 182050.0 89810.0 180705.0 ;
      RECT  89105.0 182050.0 89810.0 183395.0 ;
      RECT  89105.0 184740.0 89810.0 183395.0 ;
      RECT  89105.0 184740.0 89810.0 186085.0 ;
      RECT  89105.0 187430.0 89810.0 186085.0 ;
      RECT  89105.0 187430.0 89810.0 188775.0 ;
      RECT  89105.0 190120.0 89810.0 188775.0 ;
      RECT  89105.0 190120.0 89810.0 191465.0 ;
      RECT  89105.0 192810.0 89810.0 191465.0 ;
      RECT  89105.0 192810.0 89810.0 194155.0 ;
      RECT  89105.0 195500.0 89810.0 194155.0 ;
      RECT  89105.0 195500.0 89810.0 196845.0 ;
      RECT  89105.0 198190.0 89810.0 196845.0 ;
      RECT  89105.0 198190.0 89810.0 199535.0 ;
      RECT  89105.0 200880.0 89810.0 199535.0 ;
      RECT  89105.0 200880.0 89810.0 202225.0 ;
      RECT  89105.0 203570.0 89810.0 202225.0 ;
      RECT  89105.0 203570.0 89810.0 204915.0 ;
      RECT  89105.0 206260.0 89810.0 204915.0 ;
      RECT  89810.0 34100.0 90515.0 35445.0 ;
      RECT  89810.0 36790.0 90515.0 35445.0 ;
      RECT  89810.0 36790.0 90515.0 38135.0 ;
      RECT  89810.0 39480.0 90515.0 38135.0 ;
      RECT  89810.0 39480.0 90515.0 40825.0 ;
      RECT  89810.0 42170.0 90515.0 40825.0 ;
      RECT  89810.0 42170.0 90515.0 43515.0 ;
      RECT  89810.0 44860.0 90515.0 43515.0 ;
      RECT  89810.0 44860.0 90515.0 46205.0 ;
      RECT  89810.0 47550.0 90515.0 46205.0 ;
      RECT  89810.0 47550.0 90515.0 48895.0 ;
      RECT  89810.0 50240.0 90515.0 48895.0 ;
      RECT  89810.0 50240.0 90515.0 51585.0 ;
      RECT  89810.0 52930.0 90515.0 51585.0 ;
      RECT  89810.0 52930.0 90515.0 54275.0 ;
      RECT  89810.0 55620.0 90515.0 54275.0 ;
      RECT  89810.0 55620.0 90515.0 56965.0 ;
      RECT  89810.0 58310.0 90515.0 56965.0 ;
      RECT  89810.0 58310.0 90515.0 59655.0 ;
      RECT  89810.0 61000.0 90515.0 59655.0 ;
      RECT  89810.0 61000.0 90515.0 62345.0 ;
      RECT  89810.0 63690.0 90515.0 62345.0 ;
      RECT  89810.0 63690.0 90515.0 65035.0 ;
      RECT  89810.0 66380.0 90515.0 65035.0 ;
      RECT  89810.0 66380.0 90515.0 67725.0 ;
      RECT  89810.0 69070.0 90515.0 67725.0 ;
      RECT  89810.0 69070.0 90515.0 70415.0 ;
      RECT  89810.0 71760.0 90515.0 70415.0 ;
      RECT  89810.0 71760.0 90515.0 73105.0 ;
      RECT  89810.0 74450.0 90515.0 73105.0 ;
      RECT  89810.0 74450.0 90515.0 75795.0 ;
      RECT  89810.0 77140.0 90515.0 75795.0 ;
      RECT  89810.0 77140.0 90515.0 78485.0 ;
      RECT  89810.0 79830.0 90515.0 78485.0 ;
      RECT  89810.0 79830.0 90515.0 81175.0 ;
      RECT  89810.0 82520.0 90515.0 81175.0 ;
      RECT  89810.0 82520.0 90515.0 83865.0 ;
      RECT  89810.0 85210.0 90515.0 83865.0 ;
      RECT  89810.0 85210.0 90515.0 86555.0 ;
      RECT  89810.0 87900.0 90515.0 86555.0 ;
      RECT  89810.0 87900.0 90515.0 89245.0 ;
      RECT  89810.0 90590.0 90515.0 89245.0 ;
      RECT  89810.0 90590.0 90515.0 91935.0 ;
      RECT  89810.0 93280.0 90515.0 91935.0 ;
      RECT  89810.0 93280.0 90515.0 94625.0 ;
      RECT  89810.0 95970.0 90515.0 94625.0 ;
      RECT  89810.0 95970.0 90515.0 97315.0 ;
      RECT  89810.0 98660.0 90515.0 97315.0 ;
      RECT  89810.0 98660.0 90515.0 100005.0 ;
      RECT  89810.0 101350.0 90515.0 100005.0 ;
      RECT  89810.0 101350.0 90515.0 102695.0 ;
      RECT  89810.0 104040.0 90515.0 102695.0 ;
      RECT  89810.0 104040.0 90515.0 105385.0 ;
      RECT  89810.0 106730.0 90515.0 105385.0 ;
      RECT  89810.0 106730.0 90515.0 108075.0 ;
      RECT  89810.0 109420.0 90515.0 108075.0 ;
      RECT  89810.0 109420.0 90515.0 110765.0 ;
      RECT  89810.0 112110.0 90515.0 110765.0 ;
      RECT  89810.0 112110.0 90515.0 113455.0 ;
      RECT  89810.0 114800.0 90515.0 113455.0 ;
      RECT  89810.0 114800.0 90515.0 116145.0 ;
      RECT  89810.0 117490.0 90515.0 116145.0 ;
      RECT  89810.0 117490.0 90515.0 118835.0 ;
      RECT  89810.0 120180.0 90515.0 118835.0 ;
      RECT  89810.0 120180.0 90515.0 121525.0 ;
      RECT  89810.0 122870.0 90515.0 121525.0 ;
      RECT  89810.0 122870.0 90515.0 124215.0 ;
      RECT  89810.0 125560.0 90515.0 124215.0 ;
      RECT  89810.0 125560.0 90515.0 126905.0 ;
      RECT  89810.0 128250.0 90515.0 126905.0 ;
      RECT  89810.0 128250.0 90515.0 129595.0 ;
      RECT  89810.0 130940.0 90515.0 129595.0 ;
      RECT  89810.0 130940.0 90515.0 132285.0 ;
      RECT  89810.0 133630.0 90515.0 132285.0 ;
      RECT  89810.0 133630.0 90515.0 134975.0 ;
      RECT  89810.0 136320.0 90515.0 134975.0 ;
      RECT  89810.0 136320.0 90515.0 137665.0 ;
      RECT  89810.0 139010.0 90515.0 137665.0 ;
      RECT  89810.0 139010.0 90515.0 140355.0 ;
      RECT  89810.0 141700.0 90515.0 140355.0 ;
      RECT  89810.0 141700.0 90515.0 143045.0 ;
      RECT  89810.0 144390.0 90515.0 143045.0 ;
      RECT  89810.0 144390.0 90515.0 145735.0 ;
      RECT  89810.0 147080.0 90515.0 145735.0 ;
      RECT  89810.0 147080.0 90515.0 148425.0 ;
      RECT  89810.0 149770.0 90515.0 148425.0 ;
      RECT  89810.0 149770.0 90515.0 151115.0 ;
      RECT  89810.0 152460.0 90515.0 151115.0 ;
      RECT  89810.0 152460.0 90515.0 153805.0 ;
      RECT  89810.0 155150.0 90515.0 153805.0 ;
      RECT  89810.0 155150.0 90515.0 156495.0 ;
      RECT  89810.0 157840.0 90515.0 156495.0 ;
      RECT  89810.0 157840.0 90515.0 159185.0 ;
      RECT  89810.0 160530.0 90515.0 159185.0 ;
      RECT  89810.0 160530.0 90515.0 161875.0 ;
      RECT  89810.0 163220.0 90515.0 161875.0 ;
      RECT  89810.0 163220.0 90515.0 164565.0 ;
      RECT  89810.0 165910.0 90515.0 164565.0 ;
      RECT  89810.0 165910.0 90515.0 167255.0 ;
      RECT  89810.0 168600.0 90515.0 167255.0 ;
      RECT  89810.0 168600.0 90515.0 169945.0 ;
      RECT  89810.0 171290.0 90515.0 169945.0 ;
      RECT  89810.0 171290.0 90515.0 172635.0 ;
      RECT  89810.0 173980.0 90515.0 172635.0 ;
      RECT  89810.0 173980.0 90515.0 175325.0 ;
      RECT  89810.0 176670.0 90515.0 175325.0 ;
      RECT  89810.0 176670.0 90515.0 178015.0 ;
      RECT  89810.0 179360.0 90515.0 178015.0 ;
      RECT  89810.0 179360.0 90515.0 180705.0 ;
      RECT  89810.0 182050.0 90515.0 180705.0 ;
      RECT  89810.0 182050.0 90515.0 183395.0 ;
      RECT  89810.0 184740.0 90515.0 183395.0 ;
      RECT  89810.0 184740.0 90515.0 186085.0 ;
      RECT  89810.0 187430.0 90515.0 186085.0 ;
      RECT  89810.0 187430.0 90515.0 188775.0 ;
      RECT  89810.0 190120.0 90515.0 188775.0 ;
      RECT  89810.0 190120.0 90515.0 191465.0 ;
      RECT  89810.0 192810.0 90515.0 191465.0 ;
      RECT  89810.0 192810.0 90515.0 194155.0 ;
      RECT  89810.0 195500.0 90515.0 194155.0 ;
      RECT  89810.0 195500.0 90515.0 196845.0 ;
      RECT  89810.0 198190.0 90515.0 196845.0 ;
      RECT  89810.0 198190.0 90515.0 199535.0 ;
      RECT  89810.0 200880.0 90515.0 199535.0 ;
      RECT  89810.0 200880.0 90515.0 202225.0 ;
      RECT  89810.0 203570.0 90515.0 202225.0 ;
      RECT  89810.0 203570.0 90515.0 204915.0 ;
      RECT  89810.0 206260.0 90515.0 204915.0 ;
      RECT  90515.0 34100.0 91220.0 35445.0 ;
      RECT  90515.0 36790.0 91220.0 35445.0 ;
      RECT  90515.0 36790.0 91220.0 38135.0 ;
      RECT  90515.0 39480.0 91220.0 38135.0 ;
      RECT  90515.0 39480.0 91220.0 40825.0 ;
      RECT  90515.0 42170.0 91220.0 40825.0 ;
      RECT  90515.0 42170.0 91220.0 43515.0 ;
      RECT  90515.0 44860.0 91220.0 43515.0 ;
      RECT  90515.0 44860.0 91220.0 46205.0 ;
      RECT  90515.0 47550.0 91220.0 46205.0 ;
      RECT  90515.0 47550.0 91220.0 48895.0 ;
      RECT  90515.0 50240.0 91220.0 48895.0 ;
      RECT  90515.0 50240.0 91220.0 51585.0 ;
      RECT  90515.0 52930.0 91220.0 51585.0 ;
      RECT  90515.0 52930.0 91220.0 54275.0 ;
      RECT  90515.0 55620.0 91220.0 54275.0 ;
      RECT  90515.0 55620.0 91220.0 56965.0 ;
      RECT  90515.0 58310.0 91220.0 56965.0 ;
      RECT  90515.0 58310.0 91220.0 59655.0 ;
      RECT  90515.0 61000.0 91220.0 59655.0 ;
      RECT  90515.0 61000.0 91220.0 62345.0 ;
      RECT  90515.0 63690.0 91220.0 62345.0 ;
      RECT  90515.0 63690.0 91220.0 65035.0 ;
      RECT  90515.0 66380.0 91220.0 65035.0 ;
      RECT  90515.0 66380.0 91220.0 67725.0 ;
      RECT  90515.0 69070.0 91220.0 67725.0 ;
      RECT  90515.0 69070.0 91220.0 70415.0 ;
      RECT  90515.0 71760.0 91220.0 70415.0 ;
      RECT  90515.0 71760.0 91220.0 73105.0 ;
      RECT  90515.0 74450.0 91220.0 73105.0 ;
      RECT  90515.0 74450.0 91220.0 75795.0 ;
      RECT  90515.0 77140.0 91220.0 75795.0 ;
      RECT  90515.0 77140.0 91220.0 78485.0 ;
      RECT  90515.0 79830.0 91220.0 78485.0 ;
      RECT  90515.0 79830.0 91220.0 81175.0 ;
      RECT  90515.0 82520.0 91220.0 81175.0 ;
      RECT  90515.0 82520.0 91220.0 83865.0 ;
      RECT  90515.0 85210.0 91220.0 83865.0 ;
      RECT  90515.0 85210.0 91220.0 86555.0 ;
      RECT  90515.0 87900.0 91220.0 86555.0 ;
      RECT  90515.0 87900.0 91220.0 89245.0 ;
      RECT  90515.0 90590.0 91220.0 89245.0 ;
      RECT  90515.0 90590.0 91220.0 91935.0 ;
      RECT  90515.0 93280.0 91220.0 91935.0 ;
      RECT  90515.0 93280.0 91220.0 94625.0 ;
      RECT  90515.0 95970.0 91220.0 94625.0 ;
      RECT  90515.0 95970.0 91220.0 97315.0 ;
      RECT  90515.0 98660.0 91220.0 97315.0 ;
      RECT  90515.0 98660.0 91220.0 100005.0 ;
      RECT  90515.0 101350.0 91220.0 100005.0 ;
      RECT  90515.0 101350.0 91220.0 102695.0 ;
      RECT  90515.0 104040.0 91220.0 102695.0 ;
      RECT  90515.0 104040.0 91220.0 105385.0 ;
      RECT  90515.0 106730.0 91220.0 105385.0 ;
      RECT  90515.0 106730.0 91220.0 108075.0 ;
      RECT  90515.0 109420.0 91220.0 108075.0 ;
      RECT  90515.0 109420.0 91220.0 110765.0 ;
      RECT  90515.0 112110.0 91220.0 110765.0 ;
      RECT  90515.0 112110.0 91220.0 113455.0 ;
      RECT  90515.0 114800.0 91220.0 113455.0 ;
      RECT  90515.0 114800.0 91220.0 116145.0 ;
      RECT  90515.0 117490.0 91220.0 116145.0 ;
      RECT  90515.0 117490.0 91220.0 118835.0 ;
      RECT  90515.0 120180.0 91220.0 118835.0 ;
      RECT  90515.0 120180.0 91220.0 121525.0 ;
      RECT  90515.0 122870.0 91220.0 121525.0 ;
      RECT  90515.0 122870.0 91220.0 124215.0 ;
      RECT  90515.0 125560.0 91220.0 124215.0 ;
      RECT  90515.0 125560.0 91220.0 126905.0 ;
      RECT  90515.0 128250.0 91220.0 126905.0 ;
      RECT  90515.0 128250.0 91220.0 129595.0 ;
      RECT  90515.0 130940.0 91220.0 129595.0 ;
      RECT  90515.0 130940.0 91220.0 132285.0 ;
      RECT  90515.0 133630.0 91220.0 132285.0 ;
      RECT  90515.0 133630.0 91220.0 134975.0 ;
      RECT  90515.0 136320.0 91220.0 134975.0 ;
      RECT  90515.0 136320.0 91220.0 137665.0 ;
      RECT  90515.0 139010.0 91220.0 137665.0 ;
      RECT  90515.0 139010.0 91220.0 140355.0 ;
      RECT  90515.0 141700.0 91220.0 140355.0 ;
      RECT  90515.0 141700.0 91220.0 143045.0 ;
      RECT  90515.0 144390.0 91220.0 143045.0 ;
      RECT  90515.0 144390.0 91220.0 145735.0 ;
      RECT  90515.0 147080.0 91220.0 145735.0 ;
      RECT  90515.0 147080.0 91220.0 148425.0 ;
      RECT  90515.0 149770.0 91220.0 148425.0 ;
      RECT  90515.0 149770.0 91220.0 151115.0 ;
      RECT  90515.0 152460.0 91220.0 151115.0 ;
      RECT  90515.0 152460.0 91220.0 153805.0 ;
      RECT  90515.0 155150.0 91220.0 153805.0 ;
      RECT  90515.0 155150.0 91220.0 156495.0 ;
      RECT  90515.0 157840.0 91220.0 156495.0 ;
      RECT  90515.0 157840.0 91220.0 159185.0 ;
      RECT  90515.0 160530.0 91220.0 159185.0 ;
      RECT  90515.0 160530.0 91220.0 161875.0 ;
      RECT  90515.0 163220.0 91220.0 161875.0 ;
      RECT  90515.0 163220.0 91220.0 164565.0 ;
      RECT  90515.0 165910.0 91220.0 164565.0 ;
      RECT  90515.0 165910.0 91220.0 167255.0 ;
      RECT  90515.0 168600.0 91220.0 167255.0 ;
      RECT  90515.0 168600.0 91220.0 169945.0 ;
      RECT  90515.0 171290.0 91220.0 169945.0 ;
      RECT  90515.0 171290.0 91220.0 172635.0 ;
      RECT  90515.0 173980.0 91220.0 172635.0 ;
      RECT  90515.0 173980.0 91220.0 175325.0 ;
      RECT  90515.0 176670.0 91220.0 175325.0 ;
      RECT  90515.0 176670.0 91220.0 178015.0 ;
      RECT  90515.0 179360.0 91220.0 178015.0 ;
      RECT  90515.0 179360.0 91220.0 180705.0 ;
      RECT  90515.0 182050.0 91220.0 180705.0 ;
      RECT  90515.0 182050.0 91220.0 183395.0 ;
      RECT  90515.0 184740.0 91220.0 183395.0 ;
      RECT  90515.0 184740.0 91220.0 186085.0 ;
      RECT  90515.0 187430.0 91220.0 186085.0 ;
      RECT  90515.0 187430.0 91220.0 188775.0 ;
      RECT  90515.0 190120.0 91220.0 188775.0 ;
      RECT  90515.0 190120.0 91220.0 191465.0 ;
      RECT  90515.0 192810.0 91220.0 191465.0 ;
      RECT  90515.0 192810.0 91220.0 194155.0 ;
      RECT  90515.0 195500.0 91220.0 194155.0 ;
      RECT  90515.0 195500.0 91220.0 196845.0 ;
      RECT  90515.0 198190.0 91220.0 196845.0 ;
      RECT  90515.0 198190.0 91220.0 199535.0 ;
      RECT  90515.0 200880.0 91220.0 199535.0 ;
      RECT  90515.0 200880.0 91220.0 202225.0 ;
      RECT  90515.0 203570.0 91220.0 202225.0 ;
      RECT  90515.0 203570.0 91220.0 204915.0 ;
      RECT  90515.0 206260.0 91220.0 204915.0 ;
      RECT  91220.0 34100.0 91925.0 35445.0 ;
      RECT  91220.0 36790.0 91925.0 35445.0 ;
      RECT  91220.0 36790.0 91925.0 38135.0 ;
      RECT  91220.0 39480.0 91925.0 38135.0 ;
      RECT  91220.0 39480.0 91925.0 40825.0 ;
      RECT  91220.0 42170.0 91925.0 40825.0 ;
      RECT  91220.0 42170.0 91925.0 43515.0 ;
      RECT  91220.0 44860.0 91925.0 43515.0 ;
      RECT  91220.0 44860.0 91925.0 46205.0 ;
      RECT  91220.0 47550.0 91925.0 46205.0 ;
      RECT  91220.0 47550.0 91925.0 48895.0 ;
      RECT  91220.0 50240.0 91925.0 48895.0 ;
      RECT  91220.0 50240.0 91925.0 51585.0 ;
      RECT  91220.0 52930.0 91925.0 51585.0 ;
      RECT  91220.0 52930.0 91925.0 54275.0 ;
      RECT  91220.0 55620.0 91925.0 54275.0 ;
      RECT  91220.0 55620.0 91925.0 56965.0 ;
      RECT  91220.0 58310.0 91925.0 56965.0 ;
      RECT  91220.0 58310.0 91925.0 59655.0 ;
      RECT  91220.0 61000.0 91925.0 59655.0 ;
      RECT  91220.0 61000.0 91925.0 62345.0 ;
      RECT  91220.0 63690.0 91925.0 62345.0 ;
      RECT  91220.0 63690.0 91925.0 65035.0 ;
      RECT  91220.0 66380.0 91925.0 65035.0 ;
      RECT  91220.0 66380.0 91925.0 67725.0 ;
      RECT  91220.0 69070.0 91925.0 67725.0 ;
      RECT  91220.0 69070.0 91925.0 70415.0 ;
      RECT  91220.0 71760.0 91925.0 70415.0 ;
      RECT  91220.0 71760.0 91925.0 73105.0 ;
      RECT  91220.0 74450.0 91925.0 73105.0 ;
      RECT  91220.0 74450.0 91925.0 75795.0 ;
      RECT  91220.0 77140.0 91925.0 75795.0 ;
      RECT  91220.0 77140.0 91925.0 78485.0 ;
      RECT  91220.0 79830.0 91925.0 78485.0 ;
      RECT  91220.0 79830.0 91925.0 81175.0 ;
      RECT  91220.0 82520.0 91925.0 81175.0 ;
      RECT  91220.0 82520.0 91925.0 83865.0 ;
      RECT  91220.0 85210.0 91925.0 83865.0 ;
      RECT  91220.0 85210.0 91925.0 86555.0 ;
      RECT  91220.0 87900.0 91925.0 86555.0 ;
      RECT  91220.0 87900.0 91925.0 89245.0 ;
      RECT  91220.0 90590.0 91925.0 89245.0 ;
      RECT  91220.0 90590.0 91925.0 91935.0 ;
      RECT  91220.0 93280.0 91925.0 91935.0 ;
      RECT  91220.0 93280.0 91925.0 94625.0 ;
      RECT  91220.0 95970.0 91925.0 94625.0 ;
      RECT  91220.0 95970.0 91925.0 97315.0 ;
      RECT  91220.0 98660.0 91925.0 97315.0 ;
      RECT  91220.0 98660.0 91925.0 100005.0 ;
      RECT  91220.0 101350.0 91925.0 100005.0 ;
      RECT  91220.0 101350.0 91925.0 102695.0 ;
      RECT  91220.0 104040.0 91925.0 102695.0 ;
      RECT  91220.0 104040.0 91925.0 105385.0 ;
      RECT  91220.0 106730.0 91925.0 105385.0 ;
      RECT  91220.0 106730.0 91925.0 108075.0 ;
      RECT  91220.0 109420.0 91925.0 108075.0 ;
      RECT  91220.0 109420.0 91925.0 110765.0 ;
      RECT  91220.0 112110.0 91925.0 110765.0 ;
      RECT  91220.0 112110.0 91925.0 113455.0 ;
      RECT  91220.0 114800.0 91925.0 113455.0 ;
      RECT  91220.0 114800.0 91925.0 116145.0 ;
      RECT  91220.0 117490.0 91925.0 116145.0 ;
      RECT  91220.0 117490.0 91925.0 118835.0 ;
      RECT  91220.0 120180.0 91925.0 118835.0 ;
      RECT  91220.0 120180.0 91925.0 121525.0 ;
      RECT  91220.0 122870.0 91925.0 121525.0 ;
      RECT  91220.0 122870.0 91925.0 124215.0 ;
      RECT  91220.0 125560.0 91925.0 124215.0 ;
      RECT  91220.0 125560.0 91925.0 126905.0 ;
      RECT  91220.0 128250.0 91925.0 126905.0 ;
      RECT  91220.0 128250.0 91925.0 129595.0 ;
      RECT  91220.0 130940.0 91925.0 129595.0 ;
      RECT  91220.0 130940.0 91925.0 132285.0 ;
      RECT  91220.0 133630.0 91925.0 132285.0 ;
      RECT  91220.0 133630.0 91925.0 134975.0 ;
      RECT  91220.0 136320.0 91925.0 134975.0 ;
      RECT  91220.0 136320.0 91925.0 137665.0 ;
      RECT  91220.0 139010.0 91925.0 137665.0 ;
      RECT  91220.0 139010.0 91925.0 140355.0 ;
      RECT  91220.0 141700.0 91925.0 140355.0 ;
      RECT  91220.0 141700.0 91925.0 143045.0 ;
      RECT  91220.0 144390.0 91925.0 143045.0 ;
      RECT  91220.0 144390.0 91925.0 145735.0 ;
      RECT  91220.0 147080.0 91925.0 145735.0 ;
      RECT  91220.0 147080.0 91925.0 148425.0 ;
      RECT  91220.0 149770.0 91925.0 148425.0 ;
      RECT  91220.0 149770.0 91925.0 151115.0 ;
      RECT  91220.0 152460.0 91925.0 151115.0 ;
      RECT  91220.0 152460.0 91925.0 153805.0 ;
      RECT  91220.0 155150.0 91925.0 153805.0 ;
      RECT  91220.0 155150.0 91925.0 156495.0 ;
      RECT  91220.0 157840.0 91925.0 156495.0 ;
      RECT  91220.0 157840.0 91925.0 159185.0 ;
      RECT  91220.0 160530.0 91925.0 159185.0 ;
      RECT  91220.0 160530.0 91925.0 161875.0 ;
      RECT  91220.0 163220.0 91925.0 161875.0 ;
      RECT  91220.0 163220.0 91925.0 164565.0 ;
      RECT  91220.0 165910.0 91925.0 164565.0 ;
      RECT  91220.0 165910.0 91925.0 167255.0 ;
      RECT  91220.0 168600.0 91925.0 167255.0 ;
      RECT  91220.0 168600.0 91925.0 169945.0 ;
      RECT  91220.0 171290.0 91925.0 169945.0 ;
      RECT  91220.0 171290.0 91925.0 172635.0 ;
      RECT  91220.0 173980.0 91925.0 172635.0 ;
      RECT  91220.0 173980.0 91925.0 175325.0 ;
      RECT  91220.0 176670.0 91925.0 175325.0 ;
      RECT  91220.0 176670.0 91925.0 178015.0 ;
      RECT  91220.0 179360.0 91925.0 178015.0 ;
      RECT  91220.0 179360.0 91925.0 180705.0 ;
      RECT  91220.0 182050.0 91925.0 180705.0 ;
      RECT  91220.0 182050.0 91925.0 183395.0 ;
      RECT  91220.0 184740.0 91925.0 183395.0 ;
      RECT  91220.0 184740.0 91925.0 186085.0 ;
      RECT  91220.0 187430.0 91925.0 186085.0 ;
      RECT  91220.0 187430.0 91925.0 188775.0 ;
      RECT  91220.0 190120.0 91925.0 188775.0 ;
      RECT  91220.0 190120.0 91925.0 191465.0 ;
      RECT  91220.0 192810.0 91925.0 191465.0 ;
      RECT  91220.0 192810.0 91925.0 194155.0 ;
      RECT  91220.0 195500.0 91925.0 194155.0 ;
      RECT  91220.0 195500.0 91925.0 196845.0 ;
      RECT  91220.0 198190.0 91925.0 196845.0 ;
      RECT  91220.0 198190.0 91925.0 199535.0 ;
      RECT  91220.0 200880.0 91925.0 199535.0 ;
      RECT  91220.0 200880.0 91925.0 202225.0 ;
      RECT  91220.0 203570.0 91925.0 202225.0 ;
      RECT  91220.0 203570.0 91925.0 204915.0 ;
      RECT  91220.0 206260.0 91925.0 204915.0 ;
      RECT  91925.0 34100.0 92630.0 35445.0 ;
      RECT  91925.0 36790.0 92630.0 35445.0 ;
      RECT  91925.0 36790.0 92630.0 38135.0 ;
      RECT  91925.0 39480.0 92630.0 38135.0 ;
      RECT  91925.0 39480.0 92630.0 40825.0 ;
      RECT  91925.0 42170.0 92630.0 40825.0 ;
      RECT  91925.0 42170.0 92630.0 43515.0 ;
      RECT  91925.0 44860.0 92630.0 43515.0 ;
      RECT  91925.0 44860.0 92630.0 46205.0 ;
      RECT  91925.0 47550.0 92630.0 46205.0 ;
      RECT  91925.0 47550.0 92630.0 48895.0 ;
      RECT  91925.0 50240.0 92630.0 48895.0 ;
      RECT  91925.0 50240.0 92630.0 51585.0 ;
      RECT  91925.0 52930.0 92630.0 51585.0 ;
      RECT  91925.0 52930.0 92630.0 54275.0 ;
      RECT  91925.0 55620.0 92630.0 54275.0 ;
      RECT  91925.0 55620.0 92630.0 56965.0 ;
      RECT  91925.0 58310.0 92630.0 56965.0 ;
      RECT  91925.0 58310.0 92630.0 59655.0 ;
      RECT  91925.0 61000.0 92630.0 59655.0 ;
      RECT  91925.0 61000.0 92630.0 62345.0 ;
      RECT  91925.0 63690.0 92630.0 62345.0 ;
      RECT  91925.0 63690.0 92630.0 65035.0 ;
      RECT  91925.0 66380.0 92630.0 65035.0 ;
      RECT  91925.0 66380.0 92630.0 67725.0 ;
      RECT  91925.0 69070.0 92630.0 67725.0 ;
      RECT  91925.0 69070.0 92630.0 70415.0 ;
      RECT  91925.0 71760.0 92630.0 70415.0 ;
      RECT  91925.0 71760.0 92630.0 73105.0 ;
      RECT  91925.0 74450.0 92630.0 73105.0 ;
      RECT  91925.0 74450.0 92630.0 75795.0 ;
      RECT  91925.0 77140.0 92630.0 75795.0 ;
      RECT  91925.0 77140.0 92630.0 78485.0 ;
      RECT  91925.0 79830.0 92630.0 78485.0 ;
      RECT  91925.0 79830.0 92630.0 81175.0 ;
      RECT  91925.0 82520.0 92630.0 81175.0 ;
      RECT  91925.0 82520.0 92630.0 83865.0 ;
      RECT  91925.0 85210.0 92630.0 83865.0 ;
      RECT  91925.0 85210.0 92630.0 86555.0 ;
      RECT  91925.0 87900.0 92630.0 86555.0 ;
      RECT  91925.0 87900.0 92630.0 89245.0 ;
      RECT  91925.0 90590.0 92630.0 89245.0 ;
      RECT  91925.0 90590.0 92630.0 91935.0 ;
      RECT  91925.0 93280.0 92630.0 91935.0 ;
      RECT  91925.0 93280.0 92630.0 94625.0 ;
      RECT  91925.0 95970.0 92630.0 94625.0 ;
      RECT  91925.0 95970.0 92630.0 97315.0 ;
      RECT  91925.0 98660.0 92630.0 97315.0 ;
      RECT  91925.0 98660.0 92630.0 100005.0 ;
      RECT  91925.0 101350.0 92630.0 100005.0 ;
      RECT  91925.0 101350.0 92630.0 102695.0 ;
      RECT  91925.0 104040.0 92630.0 102695.0 ;
      RECT  91925.0 104040.0 92630.0 105385.0 ;
      RECT  91925.0 106730.0 92630.0 105385.0 ;
      RECT  91925.0 106730.0 92630.0 108075.0 ;
      RECT  91925.0 109420.0 92630.0 108075.0 ;
      RECT  91925.0 109420.0 92630.0 110765.0 ;
      RECT  91925.0 112110.0 92630.0 110765.0 ;
      RECT  91925.0 112110.0 92630.0 113455.0 ;
      RECT  91925.0 114800.0 92630.0 113455.0 ;
      RECT  91925.0 114800.0 92630.0 116145.0 ;
      RECT  91925.0 117490.0 92630.0 116145.0 ;
      RECT  91925.0 117490.0 92630.0 118835.0 ;
      RECT  91925.0 120180.0 92630.0 118835.0 ;
      RECT  91925.0 120180.0 92630.0 121525.0 ;
      RECT  91925.0 122870.0 92630.0 121525.0 ;
      RECT  91925.0 122870.0 92630.0 124215.0 ;
      RECT  91925.0 125560.0 92630.0 124215.0 ;
      RECT  91925.0 125560.0 92630.0 126905.0 ;
      RECT  91925.0 128250.0 92630.0 126905.0 ;
      RECT  91925.0 128250.0 92630.0 129595.0 ;
      RECT  91925.0 130940.0 92630.0 129595.0 ;
      RECT  91925.0 130940.0 92630.0 132285.0 ;
      RECT  91925.0 133630.0 92630.0 132285.0 ;
      RECT  91925.0 133630.0 92630.0 134975.0 ;
      RECT  91925.0 136320.0 92630.0 134975.0 ;
      RECT  91925.0 136320.0 92630.0 137665.0 ;
      RECT  91925.0 139010.0 92630.0 137665.0 ;
      RECT  91925.0 139010.0 92630.0 140355.0 ;
      RECT  91925.0 141700.0 92630.0 140355.0 ;
      RECT  91925.0 141700.0 92630.0 143045.0 ;
      RECT  91925.0 144390.0 92630.0 143045.0 ;
      RECT  91925.0 144390.0 92630.0 145735.0 ;
      RECT  91925.0 147080.0 92630.0 145735.0 ;
      RECT  91925.0 147080.0 92630.0 148425.0 ;
      RECT  91925.0 149770.0 92630.0 148425.0 ;
      RECT  91925.0 149770.0 92630.0 151115.0 ;
      RECT  91925.0 152460.0 92630.0 151115.0 ;
      RECT  91925.0 152460.0 92630.0 153805.0 ;
      RECT  91925.0 155150.0 92630.0 153805.0 ;
      RECT  91925.0 155150.0 92630.0 156495.0 ;
      RECT  91925.0 157840.0 92630.0 156495.0 ;
      RECT  91925.0 157840.0 92630.0 159185.0 ;
      RECT  91925.0 160530.0 92630.0 159185.0 ;
      RECT  91925.0 160530.0 92630.0 161875.0 ;
      RECT  91925.0 163220.0 92630.0 161875.0 ;
      RECT  91925.0 163220.0 92630.0 164565.0 ;
      RECT  91925.0 165910.0 92630.0 164565.0 ;
      RECT  91925.0 165910.0 92630.0 167255.0 ;
      RECT  91925.0 168600.0 92630.0 167255.0 ;
      RECT  91925.0 168600.0 92630.0 169945.0 ;
      RECT  91925.0 171290.0 92630.0 169945.0 ;
      RECT  91925.0 171290.0 92630.0 172635.0 ;
      RECT  91925.0 173980.0 92630.0 172635.0 ;
      RECT  91925.0 173980.0 92630.0 175325.0 ;
      RECT  91925.0 176670.0 92630.0 175325.0 ;
      RECT  91925.0 176670.0 92630.0 178015.0 ;
      RECT  91925.0 179360.0 92630.0 178015.0 ;
      RECT  91925.0 179360.0 92630.0 180705.0 ;
      RECT  91925.0 182050.0 92630.0 180705.0 ;
      RECT  91925.0 182050.0 92630.0 183395.0 ;
      RECT  91925.0 184740.0 92630.0 183395.0 ;
      RECT  91925.0 184740.0 92630.0 186085.0 ;
      RECT  91925.0 187430.0 92630.0 186085.0 ;
      RECT  91925.0 187430.0 92630.0 188775.0 ;
      RECT  91925.0 190120.0 92630.0 188775.0 ;
      RECT  91925.0 190120.0 92630.0 191465.0 ;
      RECT  91925.0 192810.0 92630.0 191465.0 ;
      RECT  91925.0 192810.0 92630.0 194155.0 ;
      RECT  91925.0 195500.0 92630.0 194155.0 ;
      RECT  91925.0 195500.0 92630.0 196845.0 ;
      RECT  91925.0 198190.0 92630.0 196845.0 ;
      RECT  91925.0 198190.0 92630.0 199535.0 ;
      RECT  91925.0 200880.0 92630.0 199535.0 ;
      RECT  91925.0 200880.0 92630.0 202225.0 ;
      RECT  91925.0 203570.0 92630.0 202225.0 ;
      RECT  91925.0 203570.0 92630.0 204915.0 ;
      RECT  91925.0 206260.0 92630.0 204915.0 ;
      RECT  92630.0 34100.0 93335.0 35445.0 ;
      RECT  92630.0 36790.0 93335.0 35445.0 ;
      RECT  92630.0 36790.0 93335.0 38135.0 ;
      RECT  92630.0 39480.0 93335.0 38135.0 ;
      RECT  92630.0 39480.0 93335.0 40825.0 ;
      RECT  92630.0 42170.0 93335.0 40825.0 ;
      RECT  92630.0 42170.0 93335.0 43515.0 ;
      RECT  92630.0 44860.0 93335.0 43515.0 ;
      RECT  92630.0 44860.0 93335.0 46205.0 ;
      RECT  92630.0 47550.0 93335.0 46205.0 ;
      RECT  92630.0 47550.0 93335.0 48895.0 ;
      RECT  92630.0 50240.0 93335.0 48895.0 ;
      RECT  92630.0 50240.0 93335.0 51585.0 ;
      RECT  92630.0 52930.0 93335.0 51585.0 ;
      RECT  92630.0 52930.0 93335.0 54275.0 ;
      RECT  92630.0 55620.0 93335.0 54275.0 ;
      RECT  92630.0 55620.0 93335.0 56965.0 ;
      RECT  92630.0 58310.0 93335.0 56965.0 ;
      RECT  92630.0 58310.0 93335.0 59655.0 ;
      RECT  92630.0 61000.0 93335.0 59655.0 ;
      RECT  92630.0 61000.0 93335.0 62345.0 ;
      RECT  92630.0 63690.0 93335.0 62345.0 ;
      RECT  92630.0 63690.0 93335.0 65035.0 ;
      RECT  92630.0 66380.0 93335.0 65035.0 ;
      RECT  92630.0 66380.0 93335.0 67725.0 ;
      RECT  92630.0 69070.0 93335.0 67725.0 ;
      RECT  92630.0 69070.0 93335.0 70415.0 ;
      RECT  92630.0 71760.0 93335.0 70415.0 ;
      RECT  92630.0 71760.0 93335.0 73105.0 ;
      RECT  92630.0 74450.0 93335.0 73105.0 ;
      RECT  92630.0 74450.0 93335.0 75795.0 ;
      RECT  92630.0 77140.0 93335.0 75795.0 ;
      RECT  92630.0 77140.0 93335.0 78485.0 ;
      RECT  92630.0 79830.0 93335.0 78485.0 ;
      RECT  92630.0 79830.0 93335.0 81175.0 ;
      RECT  92630.0 82520.0 93335.0 81175.0 ;
      RECT  92630.0 82520.0 93335.0 83865.0 ;
      RECT  92630.0 85210.0 93335.0 83865.0 ;
      RECT  92630.0 85210.0 93335.0 86555.0 ;
      RECT  92630.0 87900.0 93335.0 86555.0 ;
      RECT  92630.0 87900.0 93335.0 89245.0 ;
      RECT  92630.0 90590.0 93335.0 89245.0 ;
      RECT  92630.0 90590.0 93335.0 91935.0 ;
      RECT  92630.0 93280.0 93335.0 91935.0 ;
      RECT  92630.0 93280.0 93335.0 94625.0 ;
      RECT  92630.0 95970.0 93335.0 94625.0 ;
      RECT  92630.0 95970.0 93335.0 97315.0 ;
      RECT  92630.0 98660.0 93335.0 97315.0 ;
      RECT  92630.0 98660.0 93335.0 100005.0 ;
      RECT  92630.0 101350.0 93335.0 100005.0 ;
      RECT  92630.0 101350.0 93335.0 102695.0 ;
      RECT  92630.0 104040.0 93335.0 102695.0 ;
      RECT  92630.0 104040.0 93335.0 105385.0 ;
      RECT  92630.0 106730.0 93335.0 105385.0 ;
      RECT  92630.0 106730.0 93335.0 108075.0 ;
      RECT  92630.0 109420.0 93335.0 108075.0 ;
      RECT  92630.0 109420.0 93335.0 110765.0 ;
      RECT  92630.0 112110.0 93335.0 110765.0 ;
      RECT  92630.0 112110.0 93335.0 113455.0 ;
      RECT  92630.0 114800.0 93335.0 113455.0 ;
      RECT  92630.0 114800.0 93335.0 116145.0 ;
      RECT  92630.0 117490.0 93335.0 116145.0 ;
      RECT  92630.0 117490.0 93335.0 118835.0 ;
      RECT  92630.0 120180.0 93335.0 118835.0 ;
      RECT  92630.0 120180.0 93335.0 121525.0 ;
      RECT  92630.0 122870.0 93335.0 121525.0 ;
      RECT  92630.0 122870.0 93335.0 124215.0 ;
      RECT  92630.0 125560.0 93335.0 124215.0 ;
      RECT  92630.0 125560.0 93335.0 126905.0 ;
      RECT  92630.0 128250.0 93335.0 126905.0 ;
      RECT  92630.0 128250.0 93335.0 129595.0 ;
      RECT  92630.0 130940.0 93335.0 129595.0 ;
      RECT  92630.0 130940.0 93335.0 132285.0 ;
      RECT  92630.0 133630.0 93335.0 132285.0 ;
      RECT  92630.0 133630.0 93335.0 134975.0 ;
      RECT  92630.0 136320.0 93335.0 134975.0 ;
      RECT  92630.0 136320.0 93335.0 137665.0 ;
      RECT  92630.0 139010.0 93335.0 137665.0 ;
      RECT  92630.0 139010.0 93335.0 140355.0 ;
      RECT  92630.0 141700.0 93335.0 140355.0 ;
      RECT  92630.0 141700.0 93335.0 143045.0 ;
      RECT  92630.0 144390.0 93335.0 143045.0 ;
      RECT  92630.0 144390.0 93335.0 145735.0 ;
      RECT  92630.0 147080.0 93335.0 145735.0 ;
      RECT  92630.0 147080.0 93335.0 148425.0 ;
      RECT  92630.0 149770.0 93335.0 148425.0 ;
      RECT  92630.0 149770.0 93335.0 151115.0 ;
      RECT  92630.0 152460.0 93335.0 151115.0 ;
      RECT  92630.0 152460.0 93335.0 153805.0 ;
      RECT  92630.0 155150.0 93335.0 153805.0 ;
      RECT  92630.0 155150.0 93335.0 156495.0 ;
      RECT  92630.0 157840.0 93335.0 156495.0 ;
      RECT  92630.0 157840.0 93335.0 159185.0 ;
      RECT  92630.0 160530.0 93335.0 159185.0 ;
      RECT  92630.0 160530.0 93335.0 161875.0 ;
      RECT  92630.0 163220.0 93335.0 161875.0 ;
      RECT  92630.0 163220.0 93335.0 164565.0 ;
      RECT  92630.0 165910.0 93335.0 164565.0 ;
      RECT  92630.0 165910.0 93335.0 167255.0 ;
      RECT  92630.0 168600.0 93335.0 167255.0 ;
      RECT  92630.0 168600.0 93335.0 169945.0 ;
      RECT  92630.0 171290.0 93335.0 169945.0 ;
      RECT  92630.0 171290.0 93335.0 172635.0 ;
      RECT  92630.0 173980.0 93335.0 172635.0 ;
      RECT  92630.0 173980.0 93335.0 175325.0 ;
      RECT  92630.0 176670.0 93335.0 175325.0 ;
      RECT  92630.0 176670.0 93335.0 178015.0 ;
      RECT  92630.0 179360.0 93335.0 178015.0 ;
      RECT  92630.0 179360.0 93335.0 180705.0 ;
      RECT  92630.0 182050.0 93335.0 180705.0 ;
      RECT  92630.0 182050.0 93335.0 183395.0 ;
      RECT  92630.0 184740.0 93335.0 183395.0 ;
      RECT  92630.0 184740.0 93335.0 186085.0 ;
      RECT  92630.0 187430.0 93335.0 186085.0 ;
      RECT  92630.0 187430.0 93335.0 188775.0 ;
      RECT  92630.0 190120.0 93335.0 188775.0 ;
      RECT  92630.0 190120.0 93335.0 191465.0 ;
      RECT  92630.0 192810.0 93335.0 191465.0 ;
      RECT  92630.0 192810.0 93335.0 194155.0 ;
      RECT  92630.0 195500.0 93335.0 194155.0 ;
      RECT  92630.0 195500.0 93335.0 196845.0 ;
      RECT  92630.0 198190.0 93335.0 196845.0 ;
      RECT  92630.0 198190.0 93335.0 199535.0 ;
      RECT  92630.0 200880.0 93335.0 199535.0 ;
      RECT  92630.0 200880.0 93335.0 202225.0 ;
      RECT  92630.0 203570.0 93335.0 202225.0 ;
      RECT  92630.0 203570.0 93335.0 204915.0 ;
      RECT  92630.0 206260.0 93335.0 204915.0 ;
      RECT  93335.0 34100.0 94040.0 35445.0 ;
      RECT  93335.0 36790.0 94040.0 35445.0 ;
      RECT  93335.0 36790.0 94040.0 38135.0 ;
      RECT  93335.0 39480.0 94040.0 38135.0 ;
      RECT  93335.0 39480.0 94040.0 40825.0 ;
      RECT  93335.0 42170.0 94040.0 40825.0 ;
      RECT  93335.0 42170.0 94040.0 43515.0 ;
      RECT  93335.0 44860.0 94040.0 43515.0 ;
      RECT  93335.0 44860.0 94040.0 46205.0 ;
      RECT  93335.0 47550.0 94040.0 46205.0 ;
      RECT  93335.0 47550.0 94040.0 48895.0 ;
      RECT  93335.0 50240.0 94040.0 48895.0 ;
      RECT  93335.0 50240.0 94040.0 51585.0 ;
      RECT  93335.0 52930.0 94040.0 51585.0 ;
      RECT  93335.0 52930.0 94040.0 54275.0 ;
      RECT  93335.0 55620.0 94040.0 54275.0 ;
      RECT  93335.0 55620.0 94040.0 56965.0 ;
      RECT  93335.0 58310.0 94040.0 56965.0 ;
      RECT  93335.0 58310.0 94040.0 59655.0 ;
      RECT  93335.0 61000.0 94040.0 59655.0 ;
      RECT  93335.0 61000.0 94040.0 62345.0 ;
      RECT  93335.0 63690.0 94040.0 62345.0 ;
      RECT  93335.0 63690.0 94040.0 65035.0 ;
      RECT  93335.0 66380.0 94040.0 65035.0 ;
      RECT  93335.0 66380.0 94040.0 67725.0 ;
      RECT  93335.0 69070.0 94040.0 67725.0 ;
      RECT  93335.0 69070.0 94040.0 70415.0 ;
      RECT  93335.0 71760.0 94040.0 70415.0 ;
      RECT  93335.0 71760.0 94040.0 73105.0 ;
      RECT  93335.0 74450.0 94040.0 73105.0 ;
      RECT  93335.0 74450.0 94040.0 75795.0 ;
      RECT  93335.0 77140.0 94040.0 75795.0 ;
      RECT  93335.0 77140.0 94040.0 78485.0 ;
      RECT  93335.0 79830.0 94040.0 78485.0 ;
      RECT  93335.0 79830.0 94040.0 81175.0 ;
      RECT  93335.0 82520.0 94040.0 81175.0 ;
      RECT  93335.0 82520.0 94040.0 83865.0 ;
      RECT  93335.0 85210.0 94040.0 83865.0 ;
      RECT  93335.0 85210.0 94040.0 86555.0 ;
      RECT  93335.0 87900.0 94040.0 86555.0 ;
      RECT  93335.0 87900.0 94040.0 89245.0 ;
      RECT  93335.0 90590.0 94040.0 89245.0 ;
      RECT  93335.0 90590.0 94040.0 91935.0 ;
      RECT  93335.0 93280.0 94040.0 91935.0 ;
      RECT  93335.0 93280.0 94040.0 94625.0 ;
      RECT  93335.0 95970.0 94040.0 94625.0 ;
      RECT  93335.0 95970.0 94040.0 97315.0 ;
      RECT  93335.0 98660.0 94040.0 97315.0 ;
      RECT  93335.0 98660.0 94040.0 100005.0 ;
      RECT  93335.0 101350.0 94040.0 100005.0 ;
      RECT  93335.0 101350.0 94040.0 102695.0 ;
      RECT  93335.0 104040.0 94040.0 102695.0 ;
      RECT  93335.0 104040.0 94040.0 105385.0 ;
      RECT  93335.0 106730.0 94040.0 105385.0 ;
      RECT  93335.0 106730.0 94040.0 108075.0 ;
      RECT  93335.0 109420.0 94040.0 108075.0 ;
      RECT  93335.0 109420.0 94040.0 110765.0 ;
      RECT  93335.0 112110.0 94040.0 110765.0 ;
      RECT  93335.0 112110.0 94040.0 113455.0 ;
      RECT  93335.0 114800.0 94040.0 113455.0 ;
      RECT  93335.0 114800.0 94040.0 116145.0 ;
      RECT  93335.0 117490.0 94040.0 116145.0 ;
      RECT  93335.0 117490.0 94040.0 118835.0 ;
      RECT  93335.0 120180.0 94040.0 118835.0 ;
      RECT  93335.0 120180.0 94040.0 121525.0 ;
      RECT  93335.0 122870.0 94040.0 121525.0 ;
      RECT  93335.0 122870.0 94040.0 124215.0 ;
      RECT  93335.0 125560.0 94040.0 124215.0 ;
      RECT  93335.0 125560.0 94040.0 126905.0 ;
      RECT  93335.0 128250.0 94040.0 126905.0 ;
      RECT  93335.0 128250.0 94040.0 129595.0 ;
      RECT  93335.0 130940.0 94040.0 129595.0 ;
      RECT  93335.0 130940.0 94040.0 132285.0 ;
      RECT  93335.0 133630.0 94040.0 132285.0 ;
      RECT  93335.0 133630.0 94040.0 134975.0 ;
      RECT  93335.0 136320.0 94040.0 134975.0 ;
      RECT  93335.0 136320.0 94040.0 137665.0 ;
      RECT  93335.0 139010.0 94040.0 137665.0 ;
      RECT  93335.0 139010.0 94040.0 140355.0 ;
      RECT  93335.0 141700.0 94040.0 140355.0 ;
      RECT  93335.0 141700.0 94040.0 143045.0 ;
      RECT  93335.0 144390.0 94040.0 143045.0 ;
      RECT  93335.0 144390.0 94040.0 145735.0 ;
      RECT  93335.0 147080.0 94040.0 145735.0 ;
      RECT  93335.0 147080.0 94040.0 148425.0 ;
      RECT  93335.0 149770.0 94040.0 148425.0 ;
      RECT  93335.0 149770.0 94040.0 151115.0 ;
      RECT  93335.0 152460.0 94040.0 151115.0 ;
      RECT  93335.0 152460.0 94040.0 153805.0 ;
      RECT  93335.0 155150.0 94040.0 153805.0 ;
      RECT  93335.0 155150.0 94040.0 156495.0 ;
      RECT  93335.0 157840.0 94040.0 156495.0 ;
      RECT  93335.0 157840.0 94040.0 159185.0 ;
      RECT  93335.0 160530.0 94040.0 159185.0 ;
      RECT  93335.0 160530.0 94040.0 161875.0 ;
      RECT  93335.0 163220.0 94040.0 161875.0 ;
      RECT  93335.0 163220.0 94040.0 164565.0 ;
      RECT  93335.0 165910.0 94040.0 164565.0 ;
      RECT  93335.0 165910.0 94040.0 167255.0 ;
      RECT  93335.0 168600.0 94040.0 167255.0 ;
      RECT  93335.0 168600.0 94040.0 169945.0 ;
      RECT  93335.0 171290.0 94040.0 169945.0 ;
      RECT  93335.0 171290.0 94040.0 172635.0 ;
      RECT  93335.0 173980.0 94040.0 172635.0 ;
      RECT  93335.0 173980.0 94040.0 175325.0 ;
      RECT  93335.0 176670.0 94040.0 175325.0 ;
      RECT  93335.0 176670.0 94040.0 178015.0 ;
      RECT  93335.0 179360.0 94040.0 178015.0 ;
      RECT  93335.0 179360.0 94040.0 180705.0 ;
      RECT  93335.0 182050.0 94040.0 180705.0 ;
      RECT  93335.0 182050.0 94040.0 183395.0 ;
      RECT  93335.0 184740.0 94040.0 183395.0 ;
      RECT  93335.0 184740.0 94040.0 186085.0 ;
      RECT  93335.0 187430.0 94040.0 186085.0 ;
      RECT  93335.0 187430.0 94040.0 188775.0 ;
      RECT  93335.0 190120.0 94040.0 188775.0 ;
      RECT  93335.0 190120.0 94040.0 191465.0 ;
      RECT  93335.0 192810.0 94040.0 191465.0 ;
      RECT  93335.0 192810.0 94040.0 194155.0 ;
      RECT  93335.0 195500.0 94040.0 194155.0 ;
      RECT  93335.0 195500.0 94040.0 196845.0 ;
      RECT  93335.0 198190.0 94040.0 196845.0 ;
      RECT  93335.0 198190.0 94040.0 199535.0 ;
      RECT  93335.0 200880.0 94040.0 199535.0 ;
      RECT  93335.0 200880.0 94040.0 202225.0 ;
      RECT  93335.0 203570.0 94040.0 202225.0 ;
      RECT  93335.0 203570.0 94040.0 204915.0 ;
      RECT  93335.0 206260.0 94040.0 204915.0 ;
      RECT  94040.0 34100.0 94745.0 35445.0 ;
      RECT  94040.0 36790.0 94745.0 35445.0 ;
      RECT  94040.0 36790.0 94745.0 38135.0 ;
      RECT  94040.0 39480.0 94745.0 38135.0 ;
      RECT  94040.0 39480.0 94745.0 40825.0 ;
      RECT  94040.0 42170.0 94745.0 40825.0 ;
      RECT  94040.0 42170.0 94745.0 43515.0 ;
      RECT  94040.0 44860.0 94745.0 43515.0 ;
      RECT  94040.0 44860.0 94745.0 46205.0 ;
      RECT  94040.0 47550.0 94745.0 46205.0 ;
      RECT  94040.0 47550.0 94745.0 48895.0 ;
      RECT  94040.0 50240.0 94745.0 48895.0 ;
      RECT  94040.0 50240.0 94745.0 51585.0 ;
      RECT  94040.0 52930.0 94745.0 51585.0 ;
      RECT  94040.0 52930.0 94745.0 54275.0 ;
      RECT  94040.0 55620.0 94745.0 54275.0 ;
      RECT  94040.0 55620.0 94745.0 56965.0 ;
      RECT  94040.0 58310.0 94745.0 56965.0 ;
      RECT  94040.0 58310.0 94745.0 59655.0 ;
      RECT  94040.0 61000.0 94745.0 59655.0 ;
      RECT  94040.0 61000.0 94745.0 62345.0 ;
      RECT  94040.0 63690.0 94745.0 62345.0 ;
      RECT  94040.0 63690.0 94745.0 65035.0 ;
      RECT  94040.0 66380.0 94745.0 65035.0 ;
      RECT  94040.0 66380.0 94745.0 67725.0 ;
      RECT  94040.0 69070.0 94745.0 67725.0 ;
      RECT  94040.0 69070.0 94745.0 70415.0 ;
      RECT  94040.0 71760.0 94745.0 70415.0 ;
      RECT  94040.0 71760.0 94745.0 73105.0 ;
      RECT  94040.0 74450.0 94745.0 73105.0 ;
      RECT  94040.0 74450.0 94745.0 75795.0 ;
      RECT  94040.0 77140.0 94745.0 75795.0 ;
      RECT  94040.0 77140.0 94745.0 78485.0 ;
      RECT  94040.0 79830.0 94745.0 78485.0 ;
      RECT  94040.0 79830.0 94745.0 81175.0 ;
      RECT  94040.0 82520.0 94745.0 81175.0 ;
      RECT  94040.0 82520.0 94745.0 83865.0 ;
      RECT  94040.0 85210.0 94745.0 83865.0 ;
      RECT  94040.0 85210.0 94745.0 86555.0 ;
      RECT  94040.0 87900.0 94745.0 86555.0 ;
      RECT  94040.0 87900.0 94745.0 89245.0 ;
      RECT  94040.0 90590.0 94745.0 89245.0 ;
      RECT  94040.0 90590.0 94745.0 91935.0 ;
      RECT  94040.0 93280.0 94745.0 91935.0 ;
      RECT  94040.0 93280.0 94745.0 94625.0 ;
      RECT  94040.0 95970.0 94745.0 94625.0 ;
      RECT  94040.0 95970.0 94745.0 97315.0 ;
      RECT  94040.0 98660.0 94745.0 97315.0 ;
      RECT  94040.0 98660.0 94745.0 100005.0 ;
      RECT  94040.0 101350.0 94745.0 100005.0 ;
      RECT  94040.0 101350.0 94745.0 102695.0 ;
      RECT  94040.0 104040.0 94745.0 102695.0 ;
      RECT  94040.0 104040.0 94745.0 105385.0 ;
      RECT  94040.0 106730.0 94745.0 105385.0 ;
      RECT  94040.0 106730.0 94745.0 108075.0 ;
      RECT  94040.0 109420.0 94745.0 108075.0 ;
      RECT  94040.0 109420.0 94745.0 110765.0 ;
      RECT  94040.0 112110.0 94745.0 110765.0 ;
      RECT  94040.0 112110.0 94745.0 113455.0 ;
      RECT  94040.0 114800.0 94745.0 113455.0 ;
      RECT  94040.0 114800.0 94745.0 116145.0 ;
      RECT  94040.0 117490.0 94745.0 116145.0 ;
      RECT  94040.0 117490.0 94745.0 118835.0 ;
      RECT  94040.0 120180.0 94745.0 118835.0 ;
      RECT  94040.0 120180.0 94745.0 121525.0 ;
      RECT  94040.0 122870.0 94745.0 121525.0 ;
      RECT  94040.0 122870.0 94745.0 124215.0 ;
      RECT  94040.0 125560.0 94745.0 124215.0 ;
      RECT  94040.0 125560.0 94745.0 126905.0 ;
      RECT  94040.0 128250.0 94745.0 126905.0 ;
      RECT  94040.0 128250.0 94745.0 129595.0 ;
      RECT  94040.0 130940.0 94745.0 129595.0 ;
      RECT  94040.0 130940.0 94745.0 132285.0 ;
      RECT  94040.0 133630.0 94745.0 132285.0 ;
      RECT  94040.0 133630.0 94745.0 134975.0 ;
      RECT  94040.0 136320.0 94745.0 134975.0 ;
      RECT  94040.0 136320.0 94745.0 137665.0 ;
      RECT  94040.0 139010.0 94745.0 137665.0 ;
      RECT  94040.0 139010.0 94745.0 140355.0 ;
      RECT  94040.0 141700.0 94745.0 140355.0 ;
      RECT  94040.0 141700.0 94745.0 143045.0 ;
      RECT  94040.0 144390.0 94745.0 143045.0 ;
      RECT  94040.0 144390.0 94745.0 145735.0 ;
      RECT  94040.0 147080.0 94745.0 145735.0 ;
      RECT  94040.0 147080.0 94745.0 148425.0 ;
      RECT  94040.0 149770.0 94745.0 148425.0 ;
      RECT  94040.0 149770.0 94745.0 151115.0 ;
      RECT  94040.0 152460.0 94745.0 151115.0 ;
      RECT  94040.0 152460.0 94745.0 153805.0 ;
      RECT  94040.0 155150.0 94745.0 153805.0 ;
      RECT  94040.0 155150.0 94745.0 156495.0 ;
      RECT  94040.0 157840.0 94745.0 156495.0 ;
      RECT  94040.0 157840.0 94745.0 159185.0 ;
      RECT  94040.0 160530.0 94745.0 159185.0 ;
      RECT  94040.0 160530.0 94745.0 161875.0 ;
      RECT  94040.0 163220.0 94745.0 161875.0 ;
      RECT  94040.0 163220.0 94745.0 164565.0 ;
      RECT  94040.0 165910.0 94745.0 164565.0 ;
      RECT  94040.0 165910.0 94745.0 167255.0 ;
      RECT  94040.0 168600.0 94745.0 167255.0 ;
      RECT  94040.0 168600.0 94745.0 169945.0 ;
      RECT  94040.0 171290.0 94745.0 169945.0 ;
      RECT  94040.0 171290.0 94745.0 172635.0 ;
      RECT  94040.0 173980.0 94745.0 172635.0 ;
      RECT  94040.0 173980.0 94745.0 175325.0 ;
      RECT  94040.0 176670.0 94745.0 175325.0 ;
      RECT  94040.0 176670.0 94745.0 178015.0 ;
      RECT  94040.0 179360.0 94745.0 178015.0 ;
      RECT  94040.0 179360.0 94745.0 180705.0 ;
      RECT  94040.0 182050.0 94745.0 180705.0 ;
      RECT  94040.0 182050.0 94745.0 183395.0 ;
      RECT  94040.0 184740.0 94745.0 183395.0 ;
      RECT  94040.0 184740.0 94745.0 186085.0 ;
      RECT  94040.0 187430.0 94745.0 186085.0 ;
      RECT  94040.0 187430.0 94745.0 188775.0 ;
      RECT  94040.0 190120.0 94745.0 188775.0 ;
      RECT  94040.0 190120.0 94745.0 191465.0 ;
      RECT  94040.0 192810.0 94745.0 191465.0 ;
      RECT  94040.0 192810.0 94745.0 194155.0 ;
      RECT  94040.0 195500.0 94745.0 194155.0 ;
      RECT  94040.0 195500.0 94745.0 196845.0 ;
      RECT  94040.0 198190.0 94745.0 196845.0 ;
      RECT  94040.0 198190.0 94745.0 199535.0 ;
      RECT  94040.0 200880.0 94745.0 199535.0 ;
      RECT  94040.0 200880.0 94745.0 202225.0 ;
      RECT  94040.0 203570.0 94745.0 202225.0 ;
      RECT  94040.0 203570.0 94745.0 204915.0 ;
      RECT  94040.0 206260.0 94745.0 204915.0 ;
      RECT  94745.0 34100.0 95450.0 35445.0 ;
      RECT  94745.0 36790.0 95450.0 35445.0 ;
      RECT  94745.0 36790.0 95450.0 38135.0 ;
      RECT  94745.0 39480.0 95450.0 38135.0 ;
      RECT  94745.0 39480.0 95450.0 40825.0 ;
      RECT  94745.0 42170.0 95450.0 40825.0 ;
      RECT  94745.0 42170.0 95450.0 43515.0 ;
      RECT  94745.0 44860.0 95450.0 43515.0 ;
      RECT  94745.0 44860.0 95450.0 46205.0 ;
      RECT  94745.0 47550.0 95450.0 46205.0 ;
      RECT  94745.0 47550.0 95450.0 48895.0 ;
      RECT  94745.0 50240.0 95450.0 48895.0 ;
      RECT  94745.0 50240.0 95450.0 51585.0 ;
      RECT  94745.0 52930.0 95450.0 51585.0 ;
      RECT  94745.0 52930.0 95450.0 54275.0 ;
      RECT  94745.0 55620.0 95450.0 54275.0 ;
      RECT  94745.0 55620.0 95450.0 56965.0 ;
      RECT  94745.0 58310.0 95450.0 56965.0 ;
      RECT  94745.0 58310.0 95450.0 59655.0 ;
      RECT  94745.0 61000.0 95450.0 59655.0 ;
      RECT  94745.0 61000.0 95450.0 62345.0 ;
      RECT  94745.0 63690.0 95450.0 62345.0 ;
      RECT  94745.0 63690.0 95450.0 65035.0 ;
      RECT  94745.0 66380.0 95450.0 65035.0 ;
      RECT  94745.0 66380.0 95450.0 67725.0 ;
      RECT  94745.0 69070.0 95450.0 67725.0 ;
      RECT  94745.0 69070.0 95450.0 70415.0 ;
      RECT  94745.0 71760.0 95450.0 70415.0 ;
      RECT  94745.0 71760.0 95450.0 73105.0 ;
      RECT  94745.0 74450.0 95450.0 73105.0 ;
      RECT  94745.0 74450.0 95450.0 75795.0 ;
      RECT  94745.0 77140.0 95450.0 75795.0 ;
      RECT  94745.0 77140.0 95450.0 78485.0 ;
      RECT  94745.0 79830.0 95450.0 78485.0 ;
      RECT  94745.0 79830.0 95450.0 81175.0 ;
      RECT  94745.0 82520.0 95450.0 81175.0 ;
      RECT  94745.0 82520.0 95450.0 83865.0 ;
      RECT  94745.0 85210.0 95450.0 83865.0 ;
      RECT  94745.0 85210.0 95450.0 86555.0 ;
      RECT  94745.0 87900.0 95450.0 86555.0 ;
      RECT  94745.0 87900.0 95450.0 89245.0 ;
      RECT  94745.0 90590.0 95450.0 89245.0 ;
      RECT  94745.0 90590.0 95450.0 91935.0 ;
      RECT  94745.0 93280.0 95450.0 91935.0 ;
      RECT  94745.0 93280.0 95450.0 94625.0 ;
      RECT  94745.0 95970.0 95450.0 94625.0 ;
      RECT  94745.0 95970.0 95450.0 97315.0 ;
      RECT  94745.0 98660.0 95450.0 97315.0 ;
      RECT  94745.0 98660.0 95450.0 100005.0 ;
      RECT  94745.0 101350.0 95450.0 100005.0 ;
      RECT  94745.0 101350.0 95450.0 102695.0 ;
      RECT  94745.0 104040.0 95450.0 102695.0 ;
      RECT  94745.0 104040.0 95450.0 105385.0 ;
      RECT  94745.0 106730.0 95450.0 105385.0 ;
      RECT  94745.0 106730.0 95450.0 108075.0 ;
      RECT  94745.0 109420.0 95450.0 108075.0 ;
      RECT  94745.0 109420.0 95450.0 110765.0 ;
      RECT  94745.0 112110.0 95450.0 110765.0 ;
      RECT  94745.0 112110.0 95450.0 113455.0 ;
      RECT  94745.0 114800.0 95450.0 113455.0 ;
      RECT  94745.0 114800.0 95450.0 116145.0 ;
      RECT  94745.0 117490.0 95450.0 116145.0 ;
      RECT  94745.0 117490.0 95450.0 118835.0 ;
      RECT  94745.0 120180.0 95450.0 118835.0 ;
      RECT  94745.0 120180.0 95450.0 121525.0 ;
      RECT  94745.0 122870.0 95450.0 121525.0 ;
      RECT  94745.0 122870.0 95450.0 124215.0 ;
      RECT  94745.0 125560.0 95450.0 124215.0 ;
      RECT  94745.0 125560.0 95450.0 126905.0 ;
      RECT  94745.0 128250.0 95450.0 126905.0 ;
      RECT  94745.0 128250.0 95450.0 129595.0 ;
      RECT  94745.0 130940.0 95450.0 129595.0 ;
      RECT  94745.0 130940.0 95450.0 132285.0 ;
      RECT  94745.0 133630.0 95450.0 132285.0 ;
      RECT  94745.0 133630.0 95450.0 134975.0 ;
      RECT  94745.0 136320.0 95450.0 134975.0 ;
      RECT  94745.0 136320.0 95450.0 137665.0 ;
      RECT  94745.0 139010.0 95450.0 137665.0 ;
      RECT  94745.0 139010.0 95450.0 140355.0 ;
      RECT  94745.0 141700.0 95450.0 140355.0 ;
      RECT  94745.0 141700.0 95450.0 143045.0 ;
      RECT  94745.0 144390.0 95450.0 143045.0 ;
      RECT  94745.0 144390.0 95450.0 145735.0 ;
      RECT  94745.0 147080.0 95450.0 145735.0 ;
      RECT  94745.0 147080.0 95450.0 148425.0 ;
      RECT  94745.0 149770.0 95450.0 148425.0 ;
      RECT  94745.0 149770.0 95450.0 151115.0 ;
      RECT  94745.0 152460.0 95450.0 151115.0 ;
      RECT  94745.0 152460.0 95450.0 153805.0 ;
      RECT  94745.0 155150.0 95450.0 153805.0 ;
      RECT  94745.0 155150.0 95450.0 156495.0 ;
      RECT  94745.0 157840.0 95450.0 156495.0 ;
      RECT  94745.0 157840.0 95450.0 159185.0 ;
      RECT  94745.0 160530.0 95450.0 159185.0 ;
      RECT  94745.0 160530.0 95450.0 161875.0 ;
      RECT  94745.0 163220.0 95450.0 161875.0 ;
      RECT  94745.0 163220.0 95450.0 164565.0 ;
      RECT  94745.0 165910.0 95450.0 164565.0 ;
      RECT  94745.0 165910.0 95450.0 167255.0 ;
      RECT  94745.0 168600.0 95450.0 167255.0 ;
      RECT  94745.0 168600.0 95450.0 169945.0 ;
      RECT  94745.0 171290.0 95450.0 169945.0 ;
      RECT  94745.0 171290.0 95450.0 172635.0 ;
      RECT  94745.0 173980.0 95450.0 172635.0 ;
      RECT  94745.0 173980.0 95450.0 175325.0 ;
      RECT  94745.0 176670.0 95450.0 175325.0 ;
      RECT  94745.0 176670.0 95450.0 178015.0 ;
      RECT  94745.0 179360.0 95450.0 178015.0 ;
      RECT  94745.0 179360.0 95450.0 180705.0 ;
      RECT  94745.0 182050.0 95450.0 180705.0 ;
      RECT  94745.0 182050.0 95450.0 183395.0 ;
      RECT  94745.0 184740.0 95450.0 183395.0 ;
      RECT  94745.0 184740.0 95450.0 186085.0 ;
      RECT  94745.0 187430.0 95450.0 186085.0 ;
      RECT  94745.0 187430.0 95450.0 188775.0 ;
      RECT  94745.0 190120.0 95450.0 188775.0 ;
      RECT  94745.0 190120.0 95450.0 191465.0 ;
      RECT  94745.0 192810.0 95450.0 191465.0 ;
      RECT  94745.0 192810.0 95450.0 194155.0 ;
      RECT  94745.0 195500.0 95450.0 194155.0 ;
      RECT  94745.0 195500.0 95450.0 196845.0 ;
      RECT  94745.0 198190.0 95450.0 196845.0 ;
      RECT  94745.0 198190.0 95450.0 199535.0 ;
      RECT  94745.0 200880.0 95450.0 199535.0 ;
      RECT  94745.0 200880.0 95450.0 202225.0 ;
      RECT  94745.0 203570.0 95450.0 202225.0 ;
      RECT  94745.0 203570.0 95450.0 204915.0 ;
      RECT  94745.0 206260.0 95450.0 204915.0 ;
      RECT  95450.0 34100.0 96155.0 35445.0 ;
      RECT  95450.0 36790.0 96155.0 35445.0 ;
      RECT  95450.0 36790.0 96155.0 38135.0 ;
      RECT  95450.0 39480.0 96155.0 38135.0 ;
      RECT  95450.0 39480.0 96155.0 40825.0 ;
      RECT  95450.0 42170.0 96155.0 40825.0 ;
      RECT  95450.0 42170.0 96155.0 43515.0 ;
      RECT  95450.0 44860.0 96155.0 43515.0 ;
      RECT  95450.0 44860.0 96155.0 46205.0 ;
      RECT  95450.0 47550.0 96155.0 46205.0 ;
      RECT  95450.0 47550.0 96155.0 48895.0 ;
      RECT  95450.0 50240.0 96155.0 48895.0 ;
      RECT  95450.0 50240.0 96155.0 51585.0 ;
      RECT  95450.0 52930.0 96155.0 51585.0 ;
      RECT  95450.0 52930.0 96155.0 54275.0 ;
      RECT  95450.0 55620.0 96155.0 54275.0 ;
      RECT  95450.0 55620.0 96155.0 56965.0 ;
      RECT  95450.0 58310.0 96155.0 56965.0 ;
      RECT  95450.0 58310.0 96155.0 59655.0 ;
      RECT  95450.0 61000.0 96155.0 59655.0 ;
      RECT  95450.0 61000.0 96155.0 62345.0 ;
      RECT  95450.0 63690.0 96155.0 62345.0 ;
      RECT  95450.0 63690.0 96155.0 65035.0 ;
      RECT  95450.0 66380.0 96155.0 65035.0 ;
      RECT  95450.0 66380.0 96155.0 67725.0 ;
      RECT  95450.0 69070.0 96155.0 67725.0 ;
      RECT  95450.0 69070.0 96155.0 70415.0 ;
      RECT  95450.0 71760.0 96155.0 70415.0 ;
      RECT  95450.0 71760.0 96155.0 73105.0 ;
      RECT  95450.0 74450.0 96155.0 73105.0 ;
      RECT  95450.0 74450.0 96155.0 75795.0 ;
      RECT  95450.0 77140.0 96155.0 75795.0 ;
      RECT  95450.0 77140.0 96155.0 78485.0 ;
      RECT  95450.0 79830.0 96155.0 78485.0 ;
      RECT  95450.0 79830.0 96155.0 81175.0 ;
      RECT  95450.0 82520.0 96155.0 81175.0 ;
      RECT  95450.0 82520.0 96155.0 83865.0 ;
      RECT  95450.0 85210.0 96155.0 83865.0 ;
      RECT  95450.0 85210.0 96155.0 86555.0 ;
      RECT  95450.0 87900.0 96155.0 86555.0 ;
      RECT  95450.0 87900.0 96155.0 89245.0 ;
      RECT  95450.0 90590.0 96155.0 89245.0 ;
      RECT  95450.0 90590.0 96155.0 91935.0 ;
      RECT  95450.0 93280.0 96155.0 91935.0 ;
      RECT  95450.0 93280.0 96155.0 94625.0 ;
      RECT  95450.0 95970.0 96155.0 94625.0 ;
      RECT  95450.0 95970.0 96155.0 97315.0 ;
      RECT  95450.0 98660.0 96155.0 97315.0 ;
      RECT  95450.0 98660.0 96155.0 100005.0 ;
      RECT  95450.0 101350.0 96155.0 100005.0 ;
      RECT  95450.0 101350.0 96155.0 102695.0 ;
      RECT  95450.0 104040.0 96155.0 102695.0 ;
      RECT  95450.0 104040.0 96155.0 105385.0 ;
      RECT  95450.0 106730.0 96155.0 105385.0 ;
      RECT  95450.0 106730.0 96155.0 108075.0 ;
      RECT  95450.0 109420.0 96155.0 108075.0 ;
      RECT  95450.0 109420.0 96155.0 110765.0 ;
      RECT  95450.0 112110.0 96155.0 110765.0 ;
      RECT  95450.0 112110.0 96155.0 113455.0 ;
      RECT  95450.0 114800.0 96155.0 113455.0 ;
      RECT  95450.0 114800.0 96155.0 116145.0 ;
      RECT  95450.0 117490.0 96155.0 116145.0 ;
      RECT  95450.0 117490.0 96155.0 118835.0 ;
      RECT  95450.0 120180.0 96155.0 118835.0 ;
      RECT  95450.0 120180.0 96155.0 121525.0 ;
      RECT  95450.0 122870.0 96155.0 121525.0 ;
      RECT  95450.0 122870.0 96155.0 124215.0 ;
      RECT  95450.0 125560.0 96155.0 124215.0 ;
      RECT  95450.0 125560.0 96155.0 126905.0 ;
      RECT  95450.0 128250.0 96155.0 126905.0 ;
      RECT  95450.0 128250.0 96155.0 129595.0 ;
      RECT  95450.0 130940.0 96155.0 129595.0 ;
      RECT  95450.0 130940.0 96155.0 132285.0 ;
      RECT  95450.0 133630.0 96155.0 132285.0 ;
      RECT  95450.0 133630.0 96155.0 134975.0 ;
      RECT  95450.0 136320.0 96155.0 134975.0 ;
      RECT  95450.0 136320.0 96155.0 137665.0 ;
      RECT  95450.0 139010.0 96155.0 137665.0 ;
      RECT  95450.0 139010.0 96155.0 140355.0 ;
      RECT  95450.0 141700.0 96155.0 140355.0 ;
      RECT  95450.0 141700.0 96155.0 143045.0 ;
      RECT  95450.0 144390.0 96155.0 143045.0 ;
      RECT  95450.0 144390.0 96155.0 145735.0 ;
      RECT  95450.0 147080.0 96155.0 145735.0 ;
      RECT  95450.0 147080.0 96155.0 148425.0 ;
      RECT  95450.0 149770.0 96155.0 148425.0 ;
      RECT  95450.0 149770.0 96155.0 151115.0 ;
      RECT  95450.0 152460.0 96155.0 151115.0 ;
      RECT  95450.0 152460.0 96155.0 153805.0 ;
      RECT  95450.0 155150.0 96155.0 153805.0 ;
      RECT  95450.0 155150.0 96155.0 156495.0 ;
      RECT  95450.0 157840.0 96155.0 156495.0 ;
      RECT  95450.0 157840.0 96155.0 159185.0 ;
      RECT  95450.0 160530.0 96155.0 159185.0 ;
      RECT  95450.0 160530.0 96155.0 161875.0 ;
      RECT  95450.0 163220.0 96155.0 161875.0 ;
      RECT  95450.0 163220.0 96155.0 164565.0 ;
      RECT  95450.0 165910.0 96155.0 164565.0 ;
      RECT  95450.0 165910.0 96155.0 167255.0 ;
      RECT  95450.0 168600.0 96155.0 167255.0 ;
      RECT  95450.0 168600.0 96155.0 169945.0 ;
      RECT  95450.0 171290.0 96155.0 169945.0 ;
      RECT  95450.0 171290.0 96155.0 172635.0 ;
      RECT  95450.0 173980.0 96155.0 172635.0 ;
      RECT  95450.0 173980.0 96155.0 175325.0 ;
      RECT  95450.0 176670.0 96155.0 175325.0 ;
      RECT  95450.0 176670.0 96155.0 178015.0 ;
      RECT  95450.0 179360.0 96155.0 178015.0 ;
      RECT  95450.0 179360.0 96155.0 180705.0 ;
      RECT  95450.0 182050.0 96155.0 180705.0 ;
      RECT  95450.0 182050.0 96155.0 183395.0 ;
      RECT  95450.0 184740.0 96155.0 183395.0 ;
      RECT  95450.0 184740.0 96155.0 186085.0 ;
      RECT  95450.0 187430.0 96155.0 186085.0 ;
      RECT  95450.0 187430.0 96155.0 188775.0 ;
      RECT  95450.0 190120.0 96155.0 188775.0 ;
      RECT  95450.0 190120.0 96155.0 191465.0 ;
      RECT  95450.0 192810.0 96155.0 191465.0 ;
      RECT  95450.0 192810.0 96155.0 194155.0 ;
      RECT  95450.0 195500.0 96155.0 194155.0 ;
      RECT  95450.0 195500.0 96155.0 196845.0 ;
      RECT  95450.0 198190.0 96155.0 196845.0 ;
      RECT  95450.0 198190.0 96155.0 199535.0 ;
      RECT  95450.0 200880.0 96155.0 199535.0 ;
      RECT  95450.0 200880.0 96155.0 202225.0 ;
      RECT  95450.0 203570.0 96155.0 202225.0 ;
      RECT  95450.0 203570.0 96155.0 204915.0 ;
      RECT  95450.0 206260.0 96155.0 204915.0 ;
      RECT  96155.0 34100.0 96860.0 35445.0 ;
      RECT  96155.0 36790.0 96860.0 35445.0 ;
      RECT  96155.0 36790.0 96860.0 38135.0 ;
      RECT  96155.0 39480.0 96860.0 38135.0 ;
      RECT  96155.0 39480.0 96860.0 40825.0 ;
      RECT  96155.0 42170.0 96860.0 40825.0 ;
      RECT  96155.0 42170.0 96860.0 43515.0 ;
      RECT  96155.0 44860.0 96860.0 43515.0 ;
      RECT  96155.0 44860.0 96860.0 46205.0 ;
      RECT  96155.0 47550.0 96860.0 46205.0 ;
      RECT  96155.0 47550.0 96860.0 48895.0 ;
      RECT  96155.0 50240.0 96860.0 48895.0 ;
      RECT  96155.0 50240.0 96860.0 51585.0 ;
      RECT  96155.0 52930.0 96860.0 51585.0 ;
      RECT  96155.0 52930.0 96860.0 54275.0 ;
      RECT  96155.0 55620.0 96860.0 54275.0 ;
      RECT  96155.0 55620.0 96860.0 56965.0 ;
      RECT  96155.0 58310.0 96860.0 56965.0 ;
      RECT  96155.0 58310.0 96860.0 59655.0 ;
      RECT  96155.0 61000.0 96860.0 59655.0 ;
      RECT  96155.0 61000.0 96860.0 62345.0 ;
      RECT  96155.0 63690.0 96860.0 62345.0 ;
      RECT  96155.0 63690.0 96860.0 65035.0 ;
      RECT  96155.0 66380.0 96860.0 65035.0 ;
      RECT  96155.0 66380.0 96860.0 67725.0 ;
      RECT  96155.0 69070.0 96860.0 67725.0 ;
      RECT  96155.0 69070.0 96860.0 70415.0 ;
      RECT  96155.0 71760.0 96860.0 70415.0 ;
      RECT  96155.0 71760.0 96860.0 73105.0 ;
      RECT  96155.0 74450.0 96860.0 73105.0 ;
      RECT  96155.0 74450.0 96860.0 75795.0 ;
      RECT  96155.0 77140.0 96860.0 75795.0 ;
      RECT  96155.0 77140.0 96860.0 78485.0 ;
      RECT  96155.0 79830.0 96860.0 78485.0 ;
      RECT  96155.0 79830.0 96860.0 81175.0 ;
      RECT  96155.0 82520.0 96860.0 81175.0 ;
      RECT  96155.0 82520.0 96860.0 83865.0 ;
      RECT  96155.0 85210.0 96860.0 83865.0 ;
      RECT  96155.0 85210.0 96860.0 86555.0 ;
      RECT  96155.0 87900.0 96860.0 86555.0 ;
      RECT  96155.0 87900.0 96860.0 89245.0 ;
      RECT  96155.0 90590.0 96860.0 89245.0 ;
      RECT  96155.0 90590.0 96860.0 91935.0 ;
      RECT  96155.0 93280.0 96860.0 91935.0 ;
      RECT  96155.0 93280.0 96860.0 94625.0 ;
      RECT  96155.0 95970.0 96860.0 94625.0 ;
      RECT  96155.0 95970.0 96860.0 97315.0 ;
      RECT  96155.0 98660.0 96860.0 97315.0 ;
      RECT  96155.0 98660.0 96860.0 100005.0 ;
      RECT  96155.0 101350.0 96860.0 100005.0 ;
      RECT  96155.0 101350.0 96860.0 102695.0 ;
      RECT  96155.0 104040.0 96860.0 102695.0 ;
      RECT  96155.0 104040.0 96860.0 105385.0 ;
      RECT  96155.0 106730.0 96860.0 105385.0 ;
      RECT  96155.0 106730.0 96860.0 108075.0 ;
      RECT  96155.0 109420.0 96860.0 108075.0 ;
      RECT  96155.0 109420.0 96860.0 110765.0 ;
      RECT  96155.0 112110.0 96860.0 110765.0 ;
      RECT  96155.0 112110.0 96860.0 113455.0 ;
      RECT  96155.0 114800.0 96860.0 113455.0 ;
      RECT  96155.0 114800.0 96860.0 116145.0 ;
      RECT  96155.0 117490.0 96860.0 116145.0 ;
      RECT  96155.0 117490.0 96860.0 118835.0 ;
      RECT  96155.0 120180.0 96860.0 118835.0 ;
      RECT  96155.0 120180.0 96860.0 121525.0 ;
      RECT  96155.0 122870.0 96860.0 121525.0 ;
      RECT  96155.0 122870.0 96860.0 124215.0 ;
      RECT  96155.0 125560.0 96860.0 124215.0 ;
      RECT  96155.0 125560.0 96860.0 126905.0 ;
      RECT  96155.0 128250.0 96860.0 126905.0 ;
      RECT  96155.0 128250.0 96860.0 129595.0 ;
      RECT  96155.0 130940.0 96860.0 129595.0 ;
      RECT  96155.0 130940.0 96860.0 132285.0 ;
      RECT  96155.0 133630.0 96860.0 132285.0 ;
      RECT  96155.0 133630.0 96860.0 134975.0 ;
      RECT  96155.0 136320.0 96860.0 134975.0 ;
      RECT  96155.0 136320.0 96860.0 137665.0 ;
      RECT  96155.0 139010.0 96860.0 137665.0 ;
      RECT  96155.0 139010.0 96860.0 140355.0 ;
      RECT  96155.0 141700.0 96860.0 140355.0 ;
      RECT  96155.0 141700.0 96860.0 143045.0 ;
      RECT  96155.0 144390.0 96860.0 143045.0 ;
      RECT  96155.0 144390.0 96860.0 145735.0 ;
      RECT  96155.0 147080.0 96860.0 145735.0 ;
      RECT  96155.0 147080.0 96860.0 148425.0 ;
      RECT  96155.0 149770.0 96860.0 148425.0 ;
      RECT  96155.0 149770.0 96860.0 151115.0 ;
      RECT  96155.0 152460.0 96860.0 151115.0 ;
      RECT  96155.0 152460.0 96860.0 153805.0 ;
      RECT  96155.0 155150.0 96860.0 153805.0 ;
      RECT  96155.0 155150.0 96860.0 156495.0 ;
      RECT  96155.0 157840.0 96860.0 156495.0 ;
      RECT  96155.0 157840.0 96860.0 159185.0 ;
      RECT  96155.0 160530.0 96860.0 159185.0 ;
      RECT  96155.0 160530.0 96860.0 161875.0 ;
      RECT  96155.0 163220.0 96860.0 161875.0 ;
      RECT  96155.0 163220.0 96860.0 164565.0 ;
      RECT  96155.0 165910.0 96860.0 164565.0 ;
      RECT  96155.0 165910.0 96860.0 167255.0 ;
      RECT  96155.0 168600.0 96860.0 167255.0 ;
      RECT  96155.0 168600.0 96860.0 169945.0 ;
      RECT  96155.0 171290.0 96860.0 169945.0 ;
      RECT  96155.0 171290.0 96860.0 172635.0 ;
      RECT  96155.0 173980.0 96860.0 172635.0 ;
      RECT  96155.0 173980.0 96860.0 175325.0 ;
      RECT  96155.0 176670.0 96860.0 175325.0 ;
      RECT  96155.0 176670.0 96860.0 178015.0 ;
      RECT  96155.0 179360.0 96860.0 178015.0 ;
      RECT  96155.0 179360.0 96860.0 180705.0 ;
      RECT  96155.0 182050.0 96860.0 180705.0 ;
      RECT  96155.0 182050.0 96860.0 183395.0 ;
      RECT  96155.0 184740.0 96860.0 183395.0 ;
      RECT  96155.0 184740.0 96860.0 186085.0 ;
      RECT  96155.0 187430.0 96860.0 186085.0 ;
      RECT  96155.0 187430.0 96860.0 188775.0 ;
      RECT  96155.0 190120.0 96860.0 188775.0 ;
      RECT  96155.0 190120.0 96860.0 191465.0 ;
      RECT  96155.0 192810.0 96860.0 191465.0 ;
      RECT  96155.0 192810.0 96860.0 194155.0 ;
      RECT  96155.0 195500.0 96860.0 194155.0 ;
      RECT  96155.0 195500.0 96860.0 196845.0 ;
      RECT  96155.0 198190.0 96860.0 196845.0 ;
      RECT  96155.0 198190.0 96860.0 199535.0 ;
      RECT  96155.0 200880.0 96860.0 199535.0 ;
      RECT  96155.0 200880.0 96860.0 202225.0 ;
      RECT  96155.0 203570.0 96860.0 202225.0 ;
      RECT  96155.0 203570.0 96860.0 204915.0 ;
      RECT  96155.0 206260.0 96860.0 204915.0 ;
      RECT  96860.0 34100.0 97565.0 35445.0 ;
      RECT  96860.0 36790.0 97565.0 35445.0 ;
      RECT  96860.0 36790.0 97565.0 38135.0 ;
      RECT  96860.0 39480.0 97565.0 38135.0 ;
      RECT  96860.0 39480.0 97565.0 40825.0 ;
      RECT  96860.0 42170.0 97565.0 40825.0 ;
      RECT  96860.0 42170.0 97565.0 43515.0 ;
      RECT  96860.0 44860.0 97565.0 43515.0 ;
      RECT  96860.0 44860.0 97565.0 46205.0 ;
      RECT  96860.0 47550.0 97565.0 46205.0 ;
      RECT  96860.0 47550.0 97565.0 48895.0 ;
      RECT  96860.0 50240.0 97565.0 48895.0 ;
      RECT  96860.0 50240.0 97565.0 51585.0 ;
      RECT  96860.0 52930.0 97565.0 51585.0 ;
      RECT  96860.0 52930.0 97565.0 54275.0 ;
      RECT  96860.0 55620.0 97565.0 54275.0 ;
      RECT  96860.0 55620.0 97565.0 56965.0 ;
      RECT  96860.0 58310.0 97565.0 56965.0 ;
      RECT  96860.0 58310.0 97565.0 59655.0 ;
      RECT  96860.0 61000.0 97565.0 59655.0 ;
      RECT  96860.0 61000.0 97565.0 62345.0 ;
      RECT  96860.0 63690.0 97565.0 62345.0 ;
      RECT  96860.0 63690.0 97565.0 65035.0 ;
      RECT  96860.0 66380.0 97565.0 65035.0 ;
      RECT  96860.0 66380.0 97565.0 67725.0 ;
      RECT  96860.0 69070.0 97565.0 67725.0 ;
      RECT  96860.0 69070.0 97565.0 70415.0 ;
      RECT  96860.0 71760.0 97565.0 70415.0 ;
      RECT  96860.0 71760.0 97565.0 73105.0 ;
      RECT  96860.0 74450.0 97565.0 73105.0 ;
      RECT  96860.0 74450.0 97565.0 75795.0 ;
      RECT  96860.0 77140.0 97565.0 75795.0 ;
      RECT  96860.0 77140.0 97565.0 78485.0 ;
      RECT  96860.0 79830.0 97565.0 78485.0 ;
      RECT  96860.0 79830.0 97565.0 81175.0 ;
      RECT  96860.0 82520.0 97565.0 81175.0 ;
      RECT  96860.0 82520.0 97565.0 83865.0 ;
      RECT  96860.0 85210.0 97565.0 83865.0 ;
      RECT  96860.0 85210.0 97565.0 86555.0 ;
      RECT  96860.0 87900.0 97565.0 86555.0 ;
      RECT  96860.0 87900.0 97565.0 89245.0 ;
      RECT  96860.0 90590.0 97565.0 89245.0 ;
      RECT  96860.0 90590.0 97565.0 91935.0 ;
      RECT  96860.0 93280.0 97565.0 91935.0 ;
      RECT  96860.0 93280.0 97565.0 94625.0 ;
      RECT  96860.0 95970.0 97565.0 94625.0 ;
      RECT  96860.0 95970.0 97565.0 97315.0 ;
      RECT  96860.0 98660.0 97565.0 97315.0 ;
      RECT  96860.0 98660.0 97565.0 100005.0 ;
      RECT  96860.0 101350.0 97565.0 100005.0 ;
      RECT  96860.0 101350.0 97565.0 102695.0 ;
      RECT  96860.0 104040.0 97565.0 102695.0 ;
      RECT  96860.0 104040.0 97565.0 105385.0 ;
      RECT  96860.0 106730.0 97565.0 105385.0 ;
      RECT  96860.0 106730.0 97565.0 108075.0 ;
      RECT  96860.0 109420.0 97565.0 108075.0 ;
      RECT  96860.0 109420.0 97565.0 110765.0 ;
      RECT  96860.0 112110.0 97565.0 110765.0 ;
      RECT  96860.0 112110.0 97565.0 113455.0 ;
      RECT  96860.0 114800.0 97565.0 113455.0 ;
      RECT  96860.0 114800.0 97565.0 116145.0 ;
      RECT  96860.0 117490.0 97565.0 116145.0 ;
      RECT  96860.0 117490.0 97565.0 118835.0 ;
      RECT  96860.0 120180.0 97565.0 118835.0 ;
      RECT  96860.0 120180.0 97565.0 121525.0 ;
      RECT  96860.0 122870.0 97565.0 121525.0 ;
      RECT  96860.0 122870.0 97565.0 124215.0 ;
      RECT  96860.0 125560.0 97565.0 124215.0 ;
      RECT  96860.0 125560.0 97565.0 126905.0 ;
      RECT  96860.0 128250.0 97565.0 126905.0 ;
      RECT  96860.0 128250.0 97565.0 129595.0 ;
      RECT  96860.0 130940.0 97565.0 129595.0 ;
      RECT  96860.0 130940.0 97565.0 132285.0 ;
      RECT  96860.0 133630.0 97565.0 132285.0 ;
      RECT  96860.0 133630.0 97565.0 134975.0 ;
      RECT  96860.0 136320.0 97565.0 134975.0 ;
      RECT  96860.0 136320.0 97565.0 137665.0 ;
      RECT  96860.0 139010.0 97565.0 137665.0 ;
      RECT  96860.0 139010.0 97565.0 140355.0 ;
      RECT  96860.0 141700.0 97565.0 140355.0 ;
      RECT  96860.0 141700.0 97565.0 143045.0 ;
      RECT  96860.0 144390.0 97565.0 143045.0 ;
      RECT  96860.0 144390.0 97565.0 145735.0 ;
      RECT  96860.0 147080.0 97565.0 145735.0 ;
      RECT  96860.0 147080.0 97565.0 148425.0 ;
      RECT  96860.0 149770.0 97565.0 148425.0 ;
      RECT  96860.0 149770.0 97565.0 151115.0 ;
      RECT  96860.0 152460.0 97565.0 151115.0 ;
      RECT  96860.0 152460.0 97565.0 153805.0 ;
      RECT  96860.0 155150.0 97565.0 153805.0 ;
      RECT  96860.0 155150.0 97565.0 156495.0 ;
      RECT  96860.0 157840.0 97565.0 156495.0 ;
      RECT  96860.0 157840.0 97565.0 159185.0 ;
      RECT  96860.0 160530.0 97565.0 159185.0 ;
      RECT  96860.0 160530.0 97565.0 161875.0 ;
      RECT  96860.0 163220.0 97565.0 161875.0 ;
      RECT  96860.0 163220.0 97565.0 164565.0 ;
      RECT  96860.0 165910.0 97565.0 164565.0 ;
      RECT  96860.0 165910.0 97565.0 167255.0 ;
      RECT  96860.0 168600.0 97565.0 167255.0 ;
      RECT  96860.0 168600.0 97565.0 169945.0 ;
      RECT  96860.0 171290.0 97565.0 169945.0 ;
      RECT  96860.0 171290.0 97565.0 172635.0 ;
      RECT  96860.0 173980.0 97565.0 172635.0 ;
      RECT  96860.0 173980.0 97565.0 175325.0 ;
      RECT  96860.0 176670.0 97565.0 175325.0 ;
      RECT  96860.0 176670.0 97565.0 178015.0 ;
      RECT  96860.0 179360.0 97565.0 178015.0 ;
      RECT  96860.0 179360.0 97565.0 180705.0 ;
      RECT  96860.0 182050.0 97565.0 180705.0 ;
      RECT  96860.0 182050.0 97565.0 183395.0 ;
      RECT  96860.0 184740.0 97565.0 183395.0 ;
      RECT  96860.0 184740.0 97565.0 186085.0 ;
      RECT  96860.0 187430.0 97565.0 186085.0 ;
      RECT  96860.0 187430.0 97565.0 188775.0 ;
      RECT  96860.0 190120.0 97565.0 188775.0 ;
      RECT  96860.0 190120.0 97565.0 191465.0 ;
      RECT  96860.0 192810.0 97565.0 191465.0 ;
      RECT  96860.0 192810.0 97565.0 194155.0 ;
      RECT  96860.0 195500.0 97565.0 194155.0 ;
      RECT  96860.0 195500.0 97565.0 196845.0 ;
      RECT  96860.0 198190.0 97565.0 196845.0 ;
      RECT  96860.0 198190.0 97565.0 199535.0 ;
      RECT  96860.0 200880.0 97565.0 199535.0 ;
      RECT  96860.0 200880.0 97565.0 202225.0 ;
      RECT  96860.0 203570.0 97565.0 202225.0 ;
      RECT  96860.0 203570.0 97565.0 204915.0 ;
      RECT  96860.0 206260.0 97565.0 204915.0 ;
      RECT  97565.0 34100.0 98270.0 35445.0 ;
      RECT  97565.0 36790.0 98270.0 35445.0 ;
      RECT  97565.0 36790.0 98270.0 38135.0 ;
      RECT  97565.0 39480.0 98270.0 38135.0 ;
      RECT  97565.0 39480.0 98270.0 40825.0 ;
      RECT  97565.0 42170.0 98270.0 40825.0 ;
      RECT  97565.0 42170.0 98270.0 43515.0 ;
      RECT  97565.0 44860.0 98270.0 43515.0 ;
      RECT  97565.0 44860.0 98270.0 46205.0 ;
      RECT  97565.0 47550.0 98270.0 46205.0 ;
      RECT  97565.0 47550.0 98270.0 48895.0 ;
      RECT  97565.0 50240.0 98270.0 48895.0 ;
      RECT  97565.0 50240.0 98270.0 51585.0 ;
      RECT  97565.0 52930.0 98270.0 51585.0 ;
      RECT  97565.0 52930.0 98270.0 54275.0 ;
      RECT  97565.0 55620.0 98270.0 54275.0 ;
      RECT  97565.0 55620.0 98270.0 56965.0 ;
      RECT  97565.0 58310.0 98270.0 56965.0 ;
      RECT  97565.0 58310.0 98270.0 59655.0 ;
      RECT  97565.0 61000.0 98270.0 59655.0 ;
      RECT  97565.0 61000.0 98270.0 62345.0 ;
      RECT  97565.0 63690.0 98270.0 62345.0 ;
      RECT  97565.0 63690.0 98270.0 65035.0 ;
      RECT  97565.0 66380.0 98270.0 65035.0 ;
      RECT  97565.0 66380.0 98270.0 67725.0 ;
      RECT  97565.0 69070.0 98270.0 67725.0 ;
      RECT  97565.0 69070.0 98270.0 70415.0 ;
      RECT  97565.0 71760.0 98270.0 70415.0 ;
      RECT  97565.0 71760.0 98270.0 73105.0 ;
      RECT  97565.0 74450.0 98270.0 73105.0 ;
      RECT  97565.0 74450.0 98270.0 75795.0 ;
      RECT  97565.0 77140.0 98270.0 75795.0 ;
      RECT  97565.0 77140.0 98270.0 78485.0 ;
      RECT  97565.0 79830.0 98270.0 78485.0 ;
      RECT  97565.0 79830.0 98270.0 81175.0 ;
      RECT  97565.0 82520.0 98270.0 81175.0 ;
      RECT  97565.0 82520.0 98270.0 83865.0 ;
      RECT  97565.0 85210.0 98270.0 83865.0 ;
      RECT  97565.0 85210.0 98270.0 86555.0 ;
      RECT  97565.0 87900.0 98270.0 86555.0 ;
      RECT  97565.0 87900.0 98270.0 89245.0 ;
      RECT  97565.0 90590.0 98270.0 89245.0 ;
      RECT  97565.0 90590.0 98270.0 91935.0 ;
      RECT  97565.0 93280.0 98270.0 91935.0 ;
      RECT  97565.0 93280.0 98270.0 94625.0 ;
      RECT  97565.0 95970.0 98270.0 94625.0 ;
      RECT  97565.0 95970.0 98270.0 97315.0 ;
      RECT  97565.0 98660.0 98270.0 97315.0 ;
      RECT  97565.0 98660.0 98270.0 100005.0 ;
      RECT  97565.0 101350.0 98270.0 100005.0 ;
      RECT  97565.0 101350.0 98270.0 102695.0 ;
      RECT  97565.0 104040.0 98270.0 102695.0 ;
      RECT  97565.0 104040.0 98270.0 105385.0 ;
      RECT  97565.0 106730.0 98270.0 105385.0 ;
      RECT  97565.0 106730.0 98270.0 108075.0 ;
      RECT  97565.0 109420.0 98270.0 108075.0 ;
      RECT  97565.0 109420.0 98270.0 110765.0 ;
      RECT  97565.0 112110.0 98270.0 110765.0 ;
      RECT  97565.0 112110.0 98270.0 113455.0 ;
      RECT  97565.0 114800.0 98270.0 113455.0 ;
      RECT  97565.0 114800.0 98270.0 116145.0 ;
      RECT  97565.0 117490.0 98270.0 116145.0 ;
      RECT  97565.0 117490.0 98270.0 118835.0 ;
      RECT  97565.0 120180.0 98270.0 118835.0 ;
      RECT  97565.0 120180.0 98270.0 121525.0 ;
      RECT  97565.0 122870.0 98270.0 121525.0 ;
      RECT  97565.0 122870.0 98270.0 124215.0 ;
      RECT  97565.0 125560.0 98270.0 124215.0 ;
      RECT  97565.0 125560.0 98270.0 126905.0 ;
      RECT  97565.0 128250.0 98270.0 126905.0 ;
      RECT  97565.0 128250.0 98270.0 129595.0 ;
      RECT  97565.0 130940.0 98270.0 129595.0 ;
      RECT  97565.0 130940.0 98270.0 132285.0 ;
      RECT  97565.0 133630.0 98270.0 132285.0 ;
      RECT  97565.0 133630.0 98270.0 134975.0 ;
      RECT  97565.0 136320.0 98270.0 134975.0 ;
      RECT  97565.0 136320.0 98270.0 137665.0 ;
      RECT  97565.0 139010.0 98270.0 137665.0 ;
      RECT  97565.0 139010.0 98270.0 140355.0 ;
      RECT  97565.0 141700.0 98270.0 140355.0 ;
      RECT  97565.0 141700.0 98270.0 143045.0 ;
      RECT  97565.0 144390.0 98270.0 143045.0 ;
      RECT  97565.0 144390.0 98270.0 145735.0 ;
      RECT  97565.0 147080.0 98270.0 145735.0 ;
      RECT  97565.0 147080.0 98270.0 148425.0 ;
      RECT  97565.0 149770.0 98270.0 148425.0 ;
      RECT  97565.0 149770.0 98270.0 151115.0 ;
      RECT  97565.0 152460.0 98270.0 151115.0 ;
      RECT  97565.0 152460.0 98270.0 153805.0 ;
      RECT  97565.0 155150.0 98270.0 153805.0 ;
      RECT  97565.0 155150.0 98270.0 156495.0 ;
      RECT  97565.0 157840.0 98270.0 156495.0 ;
      RECT  97565.0 157840.0 98270.0 159185.0 ;
      RECT  97565.0 160530.0 98270.0 159185.0 ;
      RECT  97565.0 160530.0 98270.0 161875.0 ;
      RECT  97565.0 163220.0 98270.0 161875.0 ;
      RECT  97565.0 163220.0 98270.0 164565.0 ;
      RECT  97565.0 165910.0 98270.0 164565.0 ;
      RECT  97565.0 165910.0 98270.0 167255.0 ;
      RECT  97565.0 168600.0 98270.0 167255.0 ;
      RECT  97565.0 168600.0 98270.0 169945.0 ;
      RECT  97565.0 171290.0 98270.0 169945.0 ;
      RECT  97565.0 171290.0 98270.0 172635.0 ;
      RECT  97565.0 173980.0 98270.0 172635.0 ;
      RECT  97565.0 173980.0 98270.0 175325.0 ;
      RECT  97565.0 176670.0 98270.0 175325.0 ;
      RECT  97565.0 176670.0 98270.0 178015.0 ;
      RECT  97565.0 179360.0 98270.0 178015.0 ;
      RECT  97565.0 179360.0 98270.0 180705.0 ;
      RECT  97565.0 182050.0 98270.0 180705.0 ;
      RECT  97565.0 182050.0 98270.0 183395.0 ;
      RECT  97565.0 184740.0 98270.0 183395.0 ;
      RECT  97565.0 184740.0 98270.0 186085.0 ;
      RECT  97565.0 187430.0 98270.0 186085.0 ;
      RECT  97565.0 187430.0 98270.0 188775.0 ;
      RECT  97565.0 190120.0 98270.0 188775.0 ;
      RECT  97565.0 190120.0 98270.0 191465.0 ;
      RECT  97565.0 192810.0 98270.0 191465.0 ;
      RECT  97565.0 192810.0 98270.0 194155.0 ;
      RECT  97565.0 195500.0 98270.0 194155.0 ;
      RECT  97565.0 195500.0 98270.0 196845.0 ;
      RECT  97565.0 198190.0 98270.0 196845.0 ;
      RECT  97565.0 198190.0 98270.0 199535.0 ;
      RECT  97565.0 200880.0 98270.0 199535.0 ;
      RECT  97565.0 200880.0 98270.0 202225.0 ;
      RECT  97565.0 203570.0 98270.0 202225.0 ;
      RECT  97565.0 203570.0 98270.0 204915.0 ;
      RECT  97565.0 206260.0 98270.0 204915.0 ;
      RECT  98270.0 34100.0 98975.0 35445.0 ;
      RECT  98270.0 36790.0 98975.0 35445.0 ;
      RECT  98270.0 36790.0 98975.0 38135.0 ;
      RECT  98270.0 39480.0 98975.0 38135.0 ;
      RECT  98270.0 39480.0 98975.0 40825.0 ;
      RECT  98270.0 42170.0 98975.0 40825.0 ;
      RECT  98270.0 42170.0 98975.0 43515.0 ;
      RECT  98270.0 44860.0 98975.0 43515.0 ;
      RECT  98270.0 44860.0 98975.0 46205.0 ;
      RECT  98270.0 47550.0 98975.0 46205.0 ;
      RECT  98270.0 47550.0 98975.0 48895.0 ;
      RECT  98270.0 50240.0 98975.0 48895.0 ;
      RECT  98270.0 50240.0 98975.0 51585.0 ;
      RECT  98270.0 52930.0 98975.0 51585.0 ;
      RECT  98270.0 52930.0 98975.0 54275.0 ;
      RECT  98270.0 55620.0 98975.0 54275.0 ;
      RECT  98270.0 55620.0 98975.0 56965.0 ;
      RECT  98270.0 58310.0 98975.0 56965.0 ;
      RECT  98270.0 58310.0 98975.0 59655.0 ;
      RECT  98270.0 61000.0 98975.0 59655.0 ;
      RECT  98270.0 61000.0 98975.0 62345.0 ;
      RECT  98270.0 63690.0 98975.0 62345.0 ;
      RECT  98270.0 63690.0 98975.0 65035.0 ;
      RECT  98270.0 66380.0 98975.0 65035.0 ;
      RECT  98270.0 66380.0 98975.0 67725.0 ;
      RECT  98270.0 69070.0 98975.0 67725.0 ;
      RECT  98270.0 69070.0 98975.0 70415.0 ;
      RECT  98270.0 71760.0 98975.0 70415.0 ;
      RECT  98270.0 71760.0 98975.0 73105.0 ;
      RECT  98270.0 74450.0 98975.0 73105.0 ;
      RECT  98270.0 74450.0 98975.0 75795.0 ;
      RECT  98270.0 77140.0 98975.0 75795.0 ;
      RECT  98270.0 77140.0 98975.0 78485.0 ;
      RECT  98270.0 79830.0 98975.0 78485.0 ;
      RECT  98270.0 79830.0 98975.0 81175.0 ;
      RECT  98270.0 82520.0 98975.0 81175.0 ;
      RECT  98270.0 82520.0 98975.0 83865.0 ;
      RECT  98270.0 85210.0 98975.0 83865.0 ;
      RECT  98270.0 85210.0 98975.0 86555.0 ;
      RECT  98270.0 87900.0 98975.0 86555.0 ;
      RECT  98270.0 87900.0 98975.0 89245.0 ;
      RECT  98270.0 90590.0 98975.0 89245.0 ;
      RECT  98270.0 90590.0 98975.0 91935.0 ;
      RECT  98270.0 93280.0 98975.0 91935.0 ;
      RECT  98270.0 93280.0 98975.0 94625.0 ;
      RECT  98270.0 95970.0 98975.0 94625.0 ;
      RECT  98270.0 95970.0 98975.0 97315.0 ;
      RECT  98270.0 98660.0 98975.0 97315.0 ;
      RECT  98270.0 98660.0 98975.0 100005.0 ;
      RECT  98270.0 101350.0 98975.0 100005.0 ;
      RECT  98270.0 101350.0 98975.0 102695.0 ;
      RECT  98270.0 104040.0 98975.0 102695.0 ;
      RECT  98270.0 104040.0 98975.0 105385.0 ;
      RECT  98270.0 106730.0 98975.0 105385.0 ;
      RECT  98270.0 106730.0 98975.0 108075.0 ;
      RECT  98270.0 109420.0 98975.0 108075.0 ;
      RECT  98270.0 109420.0 98975.0 110765.0 ;
      RECT  98270.0 112110.0 98975.0 110765.0 ;
      RECT  98270.0 112110.0 98975.0 113455.0 ;
      RECT  98270.0 114800.0 98975.0 113455.0 ;
      RECT  98270.0 114800.0 98975.0 116145.0 ;
      RECT  98270.0 117490.0 98975.0 116145.0 ;
      RECT  98270.0 117490.0 98975.0 118835.0 ;
      RECT  98270.0 120180.0 98975.0 118835.0 ;
      RECT  98270.0 120180.0 98975.0 121525.0 ;
      RECT  98270.0 122870.0 98975.0 121525.0 ;
      RECT  98270.0 122870.0 98975.0 124215.0 ;
      RECT  98270.0 125560.0 98975.0 124215.0 ;
      RECT  98270.0 125560.0 98975.0 126905.0 ;
      RECT  98270.0 128250.0 98975.0 126905.0 ;
      RECT  98270.0 128250.0 98975.0 129595.0 ;
      RECT  98270.0 130940.0 98975.0 129595.0 ;
      RECT  98270.0 130940.0 98975.0 132285.0 ;
      RECT  98270.0 133630.0 98975.0 132285.0 ;
      RECT  98270.0 133630.0 98975.0 134975.0 ;
      RECT  98270.0 136320.0 98975.0 134975.0 ;
      RECT  98270.0 136320.0 98975.0 137665.0 ;
      RECT  98270.0 139010.0 98975.0 137665.0 ;
      RECT  98270.0 139010.0 98975.0 140355.0 ;
      RECT  98270.0 141700.0 98975.0 140355.0 ;
      RECT  98270.0 141700.0 98975.0 143045.0 ;
      RECT  98270.0 144390.0 98975.0 143045.0 ;
      RECT  98270.0 144390.0 98975.0 145735.0 ;
      RECT  98270.0 147080.0 98975.0 145735.0 ;
      RECT  98270.0 147080.0 98975.0 148425.0 ;
      RECT  98270.0 149770.0 98975.0 148425.0 ;
      RECT  98270.0 149770.0 98975.0 151115.0 ;
      RECT  98270.0 152460.0 98975.0 151115.0 ;
      RECT  98270.0 152460.0 98975.0 153805.0 ;
      RECT  98270.0 155150.0 98975.0 153805.0 ;
      RECT  98270.0 155150.0 98975.0 156495.0 ;
      RECT  98270.0 157840.0 98975.0 156495.0 ;
      RECT  98270.0 157840.0 98975.0 159185.0 ;
      RECT  98270.0 160530.0 98975.0 159185.0 ;
      RECT  98270.0 160530.0 98975.0 161875.0 ;
      RECT  98270.0 163220.0 98975.0 161875.0 ;
      RECT  98270.0 163220.0 98975.0 164565.0 ;
      RECT  98270.0 165910.0 98975.0 164565.0 ;
      RECT  98270.0 165910.0 98975.0 167255.0 ;
      RECT  98270.0 168600.0 98975.0 167255.0 ;
      RECT  98270.0 168600.0 98975.0 169945.0 ;
      RECT  98270.0 171290.0 98975.0 169945.0 ;
      RECT  98270.0 171290.0 98975.0 172635.0 ;
      RECT  98270.0 173980.0 98975.0 172635.0 ;
      RECT  98270.0 173980.0 98975.0 175325.0 ;
      RECT  98270.0 176670.0 98975.0 175325.0 ;
      RECT  98270.0 176670.0 98975.0 178015.0 ;
      RECT  98270.0 179360.0 98975.0 178015.0 ;
      RECT  98270.0 179360.0 98975.0 180705.0 ;
      RECT  98270.0 182050.0 98975.0 180705.0 ;
      RECT  98270.0 182050.0 98975.0 183395.0 ;
      RECT  98270.0 184740.0 98975.0 183395.0 ;
      RECT  98270.0 184740.0 98975.0 186085.0 ;
      RECT  98270.0 187430.0 98975.0 186085.0 ;
      RECT  98270.0 187430.0 98975.0 188775.0 ;
      RECT  98270.0 190120.0 98975.0 188775.0 ;
      RECT  98270.0 190120.0 98975.0 191465.0 ;
      RECT  98270.0 192810.0 98975.0 191465.0 ;
      RECT  98270.0 192810.0 98975.0 194155.0 ;
      RECT  98270.0 195500.0 98975.0 194155.0 ;
      RECT  98270.0 195500.0 98975.0 196845.0 ;
      RECT  98270.0 198190.0 98975.0 196845.0 ;
      RECT  98270.0 198190.0 98975.0 199535.0 ;
      RECT  98270.0 200880.0 98975.0 199535.0 ;
      RECT  98270.0 200880.0 98975.0 202225.0 ;
      RECT  98270.0 203570.0 98975.0 202225.0 ;
      RECT  98270.0 203570.0 98975.0 204915.0 ;
      RECT  98270.0 206260.0 98975.0 204915.0 ;
      RECT  98975.0 34100.0 99680.0 35445.0 ;
      RECT  98975.0 36790.0 99680.0 35445.0 ;
      RECT  98975.0 36790.0 99680.0 38135.0 ;
      RECT  98975.0 39480.0 99680.0 38135.0 ;
      RECT  98975.0 39480.0 99680.0 40825.0 ;
      RECT  98975.0 42170.0 99680.0 40825.0 ;
      RECT  98975.0 42170.0 99680.0 43515.0 ;
      RECT  98975.0 44860.0 99680.0 43515.0 ;
      RECT  98975.0 44860.0 99680.0 46205.0 ;
      RECT  98975.0 47550.0 99680.0 46205.0 ;
      RECT  98975.0 47550.0 99680.0 48895.0 ;
      RECT  98975.0 50240.0 99680.0 48895.0 ;
      RECT  98975.0 50240.0 99680.0 51585.0 ;
      RECT  98975.0 52930.0 99680.0 51585.0 ;
      RECT  98975.0 52930.0 99680.0 54275.0 ;
      RECT  98975.0 55620.0 99680.0 54275.0 ;
      RECT  98975.0 55620.0 99680.0 56965.0 ;
      RECT  98975.0 58310.0 99680.0 56965.0 ;
      RECT  98975.0 58310.0 99680.0 59655.0 ;
      RECT  98975.0 61000.0 99680.0 59655.0 ;
      RECT  98975.0 61000.0 99680.0 62345.0 ;
      RECT  98975.0 63690.0 99680.0 62345.0 ;
      RECT  98975.0 63690.0 99680.0 65035.0 ;
      RECT  98975.0 66380.0 99680.0 65035.0 ;
      RECT  98975.0 66380.0 99680.0 67725.0 ;
      RECT  98975.0 69070.0 99680.0 67725.0 ;
      RECT  98975.0 69070.0 99680.0 70415.0 ;
      RECT  98975.0 71760.0 99680.0 70415.0 ;
      RECT  98975.0 71760.0 99680.0 73105.0 ;
      RECT  98975.0 74450.0 99680.0 73105.0 ;
      RECT  98975.0 74450.0 99680.0 75795.0 ;
      RECT  98975.0 77140.0 99680.0 75795.0 ;
      RECT  98975.0 77140.0 99680.0 78485.0 ;
      RECT  98975.0 79830.0 99680.0 78485.0 ;
      RECT  98975.0 79830.0 99680.0 81175.0 ;
      RECT  98975.0 82520.0 99680.0 81175.0 ;
      RECT  98975.0 82520.0 99680.0 83865.0 ;
      RECT  98975.0 85210.0 99680.0 83865.0 ;
      RECT  98975.0 85210.0 99680.0 86555.0 ;
      RECT  98975.0 87900.0 99680.0 86555.0 ;
      RECT  98975.0 87900.0 99680.0 89245.0 ;
      RECT  98975.0 90590.0 99680.0 89245.0 ;
      RECT  98975.0 90590.0 99680.0 91935.0 ;
      RECT  98975.0 93280.0 99680.0 91935.0 ;
      RECT  98975.0 93280.0 99680.0 94625.0 ;
      RECT  98975.0 95970.0 99680.0 94625.0 ;
      RECT  98975.0 95970.0 99680.0 97315.0 ;
      RECT  98975.0 98660.0 99680.0 97315.0 ;
      RECT  98975.0 98660.0 99680.0 100005.0 ;
      RECT  98975.0 101350.0 99680.0 100005.0 ;
      RECT  98975.0 101350.0 99680.0 102695.0 ;
      RECT  98975.0 104040.0 99680.0 102695.0 ;
      RECT  98975.0 104040.0 99680.0 105385.0 ;
      RECT  98975.0 106730.0 99680.0 105385.0 ;
      RECT  98975.0 106730.0 99680.0 108075.0 ;
      RECT  98975.0 109420.0 99680.0 108075.0 ;
      RECT  98975.0 109420.0 99680.0 110765.0 ;
      RECT  98975.0 112110.0 99680.0 110765.0 ;
      RECT  98975.0 112110.0 99680.0 113455.0 ;
      RECT  98975.0 114800.0 99680.0 113455.0 ;
      RECT  98975.0 114800.0 99680.0 116145.0 ;
      RECT  98975.0 117490.0 99680.0 116145.0 ;
      RECT  98975.0 117490.0 99680.0 118835.0 ;
      RECT  98975.0 120180.0 99680.0 118835.0 ;
      RECT  98975.0 120180.0 99680.0 121525.0 ;
      RECT  98975.0 122870.0 99680.0 121525.0 ;
      RECT  98975.0 122870.0 99680.0 124215.0 ;
      RECT  98975.0 125560.0 99680.0 124215.0 ;
      RECT  98975.0 125560.0 99680.0 126905.0 ;
      RECT  98975.0 128250.0 99680.0 126905.0 ;
      RECT  98975.0 128250.0 99680.0 129595.0 ;
      RECT  98975.0 130940.0 99680.0 129595.0 ;
      RECT  98975.0 130940.0 99680.0 132285.0 ;
      RECT  98975.0 133630.0 99680.0 132285.0 ;
      RECT  98975.0 133630.0 99680.0 134975.0 ;
      RECT  98975.0 136320.0 99680.0 134975.0 ;
      RECT  98975.0 136320.0 99680.0 137665.0 ;
      RECT  98975.0 139010.0 99680.0 137665.0 ;
      RECT  98975.0 139010.0 99680.0 140355.0 ;
      RECT  98975.0 141700.0 99680.0 140355.0 ;
      RECT  98975.0 141700.0 99680.0 143045.0 ;
      RECT  98975.0 144390.0 99680.0 143045.0 ;
      RECT  98975.0 144390.0 99680.0 145735.0 ;
      RECT  98975.0 147080.0 99680.0 145735.0 ;
      RECT  98975.0 147080.0 99680.0 148425.0 ;
      RECT  98975.0 149770.0 99680.0 148425.0 ;
      RECT  98975.0 149770.0 99680.0 151115.0 ;
      RECT  98975.0 152460.0 99680.0 151115.0 ;
      RECT  98975.0 152460.0 99680.0 153805.0 ;
      RECT  98975.0 155150.0 99680.0 153805.0 ;
      RECT  98975.0 155150.0 99680.0 156495.0 ;
      RECT  98975.0 157840.0 99680.0 156495.0 ;
      RECT  98975.0 157840.0 99680.0 159185.0 ;
      RECT  98975.0 160530.0 99680.0 159185.0 ;
      RECT  98975.0 160530.0 99680.0 161875.0 ;
      RECT  98975.0 163220.0 99680.0 161875.0 ;
      RECT  98975.0 163220.0 99680.0 164565.0 ;
      RECT  98975.0 165910.0 99680.0 164565.0 ;
      RECT  98975.0 165910.0 99680.0 167255.0 ;
      RECT  98975.0 168600.0 99680.0 167255.0 ;
      RECT  98975.0 168600.0 99680.0 169945.0 ;
      RECT  98975.0 171290.0 99680.0 169945.0 ;
      RECT  98975.0 171290.0 99680.0 172635.0 ;
      RECT  98975.0 173980.0 99680.0 172635.0 ;
      RECT  98975.0 173980.0 99680.0 175325.0 ;
      RECT  98975.0 176670.0 99680.0 175325.0 ;
      RECT  98975.0 176670.0 99680.0 178015.0 ;
      RECT  98975.0 179360.0 99680.0 178015.0 ;
      RECT  98975.0 179360.0 99680.0 180705.0 ;
      RECT  98975.0 182050.0 99680.0 180705.0 ;
      RECT  98975.0 182050.0 99680.0 183395.0 ;
      RECT  98975.0 184740.0 99680.0 183395.0 ;
      RECT  98975.0 184740.0 99680.0 186085.0 ;
      RECT  98975.0 187430.0 99680.0 186085.0 ;
      RECT  98975.0 187430.0 99680.0 188775.0 ;
      RECT  98975.0 190120.0 99680.0 188775.0 ;
      RECT  98975.0 190120.0 99680.0 191465.0 ;
      RECT  98975.0 192810.0 99680.0 191465.0 ;
      RECT  98975.0 192810.0 99680.0 194155.0 ;
      RECT  98975.0 195500.0 99680.0 194155.0 ;
      RECT  98975.0 195500.0 99680.0 196845.0 ;
      RECT  98975.0 198190.0 99680.0 196845.0 ;
      RECT  98975.0 198190.0 99680.0 199535.0 ;
      RECT  98975.0 200880.0 99680.0 199535.0 ;
      RECT  98975.0 200880.0 99680.0 202225.0 ;
      RECT  98975.0 203570.0 99680.0 202225.0 ;
      RECT  98975.0 203570.0 99680.0 204915.0 ;
      RECT  98975.0 206260.0 99680.0 204915.0 ;
      RECT  99680.0 34100.0 100385.0 35445.0 ;
      RECT  99680.0 36790.0 100385.0 35445.0 ;
      RECT  99680.0 36790.0 100385.0 38135.0 ;
      RECT  99680.0 39480.0 100385.0 38135.0 ;
      RECT  99680.0 39480.0 100385.0 40825.0 ;
      RECT  99680.0 42170.0 100385.0 40825.0 ;
      RECT  99680.0 42170.0 100385.0 43515.0 ;
      RECT  99680.0 44860.0 100385.0 43515.0 ;
      RECT  99680.0 44860.0 100385.0 46205.0 ;
      RECT  99680.0 47550.0 100385.0 46205.0 ;
      RECT  99680.0 47550.0 100385.0 48895.0 ;
      RECT  99680.0 50240.0 100385.0 48895.0 ;
      RECT  99680.0 50240.0 100385.0 51585.0 ;
      RECT  99680.0 52930.0 100385.0 51585.0 ;
      RECT  99680.0 52930.0 100385.0 54275.0 ;
      RECT  99680.0 55620.0 100385.0 54275.0 ;
      RECT  99680.0 55620.0 100385.0 56965.0 ;
      RECT  99680.0 58310.0 100385.0 56965.0 ;
      RECT  99680.0 58310.0 100385.0 59655.0 ;
      RECT  99680.0 61000.0 100385.0 59655.0 ;
      RECT  99680.0 61000.0 100385.0 62345.0 ;
      RECT  99680.0 63690.0 100385.0 62345.0 ;
      RECT  99680.0 63690.0 100385.0 65035.0 ;
      RECT  99680.0 66380.0 100385.0 65035.0 ;
      RECT  99680.0 66380.0 100385.0 67725.0 ;
      RECT  99680.0 69070.0 100385.0 67725.0 ;
      RECT  99680.0 69070.0 100385.0 70415.0 ;
      RECT  99680.0 71760.0 100385.0 70415.0 ;
      RECT  99680.0 71760.0 100385.0 73105.0 ;
      RECT  99680.0 74450.0 100385.0 73105.0 ;
      RECT  99680.0 74450.0 100385.0 75795.0 ;
      RECT  99680.0 77140.0 100385.0 75795.0 ;
      RECT  99680.0 77140.0 100385.0 78485.0 ;
      RECT  99680.0 79830.0 100385.0 78485.0 ;
      RECT  99680.0 79830.0 100385.0 81175.0 ;
      RECT  99680.0 82520.0 100385.0 81175.0 ;
      RECT  99680.0 82520.0 100385.0 83865.0 ;
      RECT  99680.0 85210.0 100385.0 83865.0 ;
      RECT  99680.0 85210.0 100385.0 86555.0 ;
      RECT  99680.0 87900.0 100385.0 86555.0 ;
      RECT  99680.0 87900.0 100385.0 89245.0 ;
      RECT  99680.0 90590.0 100385.0 89245.0 ;
      RECT  99680.0 90590.0 100385.0 91935.0 ;
      RECT  99680.0 93280.0 100385.0 91935.0 ;
      RECT  99680.0 93280.0 100385.0 94625.0 ;
      RECT  99680.0 95970.0 100385.0 94625.0 ;
      RECT  99680.0 95970.0 100385.0 97315.0 ;
      RECT  99680.0 98660.0 100385.0 97315.0 ;
      RECT  99680.0 98660.0 100385.0 100005.0 ;
      RECT  99680.0 101350.0 100385.0 100005.0 ;
      RECT  99680.0 101350.0 100385.0 102695.0 ;
      RECT  99680.0 104040.0 100385.0 102695.0 ;
      RECT  99680.0 104040.0 100385.0 105385.0 ;
      RECT  99680.0 106730.0 100385.0 105385.0 ;
      RECT  99680.0 106730.0 100385.0 108075.0 ;
      RECT  99680.0 109420.0 100385.0 108075.0 ;
      RECT  99680.0 109420.0 100385.0 110765.0 ;
      RECT  99680.0 112110.0 100385.0 110765.0 ;
      RECT  99680.0 112110.0 100385.0 113455.0 ;
      RECT  99680.0 114800.0 100385.0 113455.0 ;
      RECT  99680.0 114800.0 100385.0 116145.0 ;
      RECT  99680.0 117490.0 100385.0 116145.0 ;
      RECT  99680.0 117490.0 100385.0 118835.0 ;
      RECT  99680.0 120180.0 100385.0 118835.0 ;
      RECT  99680.0 120180.0 100385.0 121525.0 ;
      RECT  99680.0 122870.0 100385.0 121525.0 ;
      RECT  99680.0 122870.0 100385.0 124215.0 ;
      RECT  99680.0 125560.0 100385.0 124215.0 ;
      RECT  99680.0 125560.0 100385.0 126905.0 ;
      RECT  99680.0 128250.0 100385.0 126905.0 ;
      RECT  99680.0 128250.0 100385.0 129595.0 ;
      RECT  99680.0 130940.0 100385.0 129595.0 ;
      RECT  99680.0 130940.0 100385.0 132285.0 ;
      RECT  99680.0 133630.0 100385.0 132285.0 ;
      RECT  99680.0 133630.0 100385.0 134975.0 ;
      RECT  99680.0 136320.0 100385.0 134975.0 ;
      RECT  99680.0 136320.0 100385.0 137665.0 ;
      RECT  99680.0 139010.0 100385.0 137665.0 ;
      RECT  99680.0 139010.0 100385.0 140355.0 ;
      RECT  99680.0 141700.0 100385.0 140355.0 ;
      RECT  99680.0 141700.0 100385.0 143045.0 ;
      RECT  99680.0 144390.0 100385.0 143045.0 ;
      RECT  99680.0 144390.0 100385.0 145735.0 ;
      RECT  99680.0 147080.0 100385.0 145735.0 ;
      RECT  99680.0 147080.0 100385.0 148425.0 ;
      RECT  99680.0 149770.0 100385.0 148425.0 ;
      RECT  99680.0 149770.0 100385.0 151115.0 ;
      RECT  99680.0 152460.0 100385.0 151115.0 ;
      RECT  99680.0 152460.0 100385.0 153805.0 ;
      RECT  99680.0 155150.0 100385.0 153805.0 ;
      RECT  99680.0 155150.0 100385.0 156495.0 ;
      RECT  99680.0 157840.0 100385.0 156495.0 ;
      RECT  99680.0 157840.0 100385.0 159185.0 ;
      RECT  99680.0 160530.0 100385.0 159185.0 ;
      RECT  99680.0 160530.0 100385.0 161875.0 ;
      RECT  99680.0 163220.0 100385.0 161875.0 ;
      RECT  99680.0 163220.0 100385.0 164565.0 ;
      RECT  99680.0 165910.0 100385.0 164565.0 ;
      RECT  99680.0 165910.0 100385.0 167255.0 ;
      RECT  99680.0 168600.0 100385.0 167255.0 ;
      RECT  99680.0 168600.0 100385.0 169945.0 ;
      RECT  99680.0 171290.0 100385.0 169945.0 ;
      RECT  99680.0 171290.0 100385.0 172635.0 ;
      RECT  99680.0 173980.0 100385.0 172635.0 ;
      RECT  99680.0 173980.0 100385.0 175325.0 ;
      RECT  99680.0 176670.0 100385.0 175325.0 ;
      RECT  99680.0 176670.0 100385.0 178015.0 ;
      RECT  99680.0 179360.0 100385.0 178015.0 ;
      RECT  99680.0 179360.0 100385.0 180705.0 ;
      RECT  99680.0 182050.0 100385.0 180705.0 ;
      RECT  99680.0 182050.0 100385.0 183395.0 ;
      RECT  99680.0 184740.0 100385.0 183395.0 ;
      RECT  99680.0 184740.0 100385.0 186085.0 ;
      RECT  99680.0 187430.0 100385.0 186085.0 ;
      RECT  99680.0 187430.0 100385.0 188775.0 ;
      RECT  99680.0 190120.0 100385.0 188775.0 ;
      RECT  99680.0 190120.0 100385.0 191465.0 ;
      RECT  99680.0 192810.0 100385.0 191465.0 ;
      RECT  99680.0 192810.0 100385.0 194155.0 ;
      RECT  99680.0 195500.0 100385.0 194155.0 ;
      RECT  99680.0 195500.0 100385.0 196845.0 ;
      RECT  99680.0 198190.0 100385.0 196845.0 ;
      RECT  99680.0 198190.0 100385.0 199535.0 ;
      RECT  99680.0 200880.0 100385.0 199535.0 ;
      RECT  99680.0 200880.0 100385.0 202225.0 ;
      RECT  99680.0 203570.0 100385.0 202225.0 ;
      RECT  99680.0 203570.0 100385.0 204915.0 ;
      RECT  99680.0 206260.0 100385.0 204915.0 ;
      RECT  100385.0 34100.0 101090.0 35445.0 ;
      RECT  100385.0 36790.0 101090.0 35445.0 ;
      RECT  100385.0 36790.0 101090.0 38135.0 ;
      RECT  100385.0 39480.0 101090.0 38135.0 ;
      RECT  100385.0 39480.0 101090.0 40825.0 ;
      RECT  100385.0 42170.0 101090.0 40825.0 ;
      RECT  100385.0 42170.0 101090.0 43515.0 ;
      RECT  100385.0 44860.0 101090.0 43515.0 ;
      RECT  100385.0 44860.0 101090.0 46205.0 ;
      RECT  100385.0 47550.0 101090.0 46205.0 ;
      RECT  100385.0 47550.0 101090.0 48895.0 ;
      RECT  100385.0 50240.0 101090.0 48895.0 ;
      RECT  100385.0 50240.0 101090.0 51585.0 ;
      RECT  100385.0 52930.0 101090.0 51585.0 ;
      RECT  100385.0 52930.0 101090.0 54275.0 ;
      RECT  100385.0 55620.0 101090.0 54275.0 ;
      RECT  100385.0 55620.0 101090.0 56965.0 ;
      RECT  100385.0 58310.0 101090.0 56965.0 ;
      RECT  100385.0 58310.0 101090.0 59655.0 ;
      RECT  100385.0 61000.0 101090.0 59655.0 ;
      RECT  100385.0 61000.0 101090.0 62345.0 ;
      RECT  100385.0 63690.0 101090.0 62345.0 ;
      RECT  100385.0 63690.0 101090.0 65035.0 ;
      RECT  100385.0 66380.0 101090.0 65035.0 ;
      RECT  100385.0 66380.0 101090.0 67725.0 ;
      RECT  100385.0 69070.0 101090.0 67725.0 ;
      RECT  100385.0 69070.0 101090.0 70415.0 ;
      RECT  100385.0 71760.0 101090.0 70415.0 ;
      RECT  100385.0 71760.0 101090.0 73105.0 ;
      RECT  100385.0 74450.0 101090.0 73105.0 ;
      RECT  100385.0 74450.0 101090.0 75795.0 ;
      RECT  100385.0 77140.0 101090.0 75795.0 ;
      RECT  100385.0 77140.0 101090.0 78485.0 ;
      RECT  100385.0 79830.0 101090.0 78485.0 ;
      RECT  100385.0 79830.0 101090.0 81175.0 ;
      RECT  100385.0 82520.0 101090.0 81175.0 ;
      RECT  100385.0 82520.0 101090.0 83865.0 ;
      RECT  100385.0 85210.0 101090.0 83865.0 ;
      RECT  100385.0 85210.0 101090.0 86555.0 ;
      RECT  100385.0 87900.0 101090.0 86555.0 ;
      RECT  100385.0 87900.0 101090.0 89245.0 ;
      RECT  100385.0 90590.0 101090.0 89245.0 ;
      RECT  100385.0 90590.0 101090.0 91935.0 ;
      RECT  100385.0 93280.0 101090.0 91935.0 ;
      RECT  100385.0 93280.0 101090.0 94625.0 ;
      RECT  100385.0 95970.0 101090.0 94625.0 ;
      RECT  100385.0 95970.0 101090.0 97315.0 ;
      RECT  100385.0 98660.0 101090.0 97315.0 ;
      RECT  100385.0 98660.0 101090.0 100005.0 ;
      RECT  100385.0 101350.0 101090.0 100005.0 ;
      RECT  100385.0 101350.0 101090.0 102695.0 ;
      RECT  100385.0 104040.0 101090.0 102695.0 ;
      RECT  100385.0 104040.0 101090.0 105385.0 ;
      RECT  100385.0 106730.0 101090.0 105385.0 ;
      RECT  100385.0 106730.0 101090.0 108075.0 ;
      RECT  100385.0 109420.0 101090.0 108075.0 ;
      RECT  100385.0 109420.0 101090.0 110765.0 ;
      RECT  100385.0 112110.0 101090.0 110765.0 ;
      RECT  100385.0 112110.0 101090.0 113455.0 ;
      RECT  100385.0 114800.0 101090.0 113455.0 ;
      RECT  100385.0 114800.0 101090.0 116145.0 ;
      RECT  100385.0 117490.0 101090.0 116145.0 ;
      RECT  100385.0 117490.0 101090.0 118835.0 ;
      RECT  100385.0 120180.0 101090.0 118835.0 ;
      RECT  100385.0 120180.0 101090.0 121525.0 ;
      RECT  100385.0 122870.0 101090.0 121525.0 ;
      RECT  100385.0 122870.0 101090.0 124215.0 ;
      RECT  100385.0 125560.0 101090.0 124215.0 ;
      RECT  100385.0 125560.0 101090.0 126905.0 ;
      RECT  100385.0 128250.0 101090.0 126905.0 ;
      RECT  100385.0 128250.0 101090.0 129595.0 ;
      RECT  100385.0 130940.0 101090.0 129595.0 ;
      RECT  100385.0 130940.0 101090.0 132285.0 ;
      RECT  100385.0 133630.0 101090.0 132285.0 ;
      RECT  100385.0 133630.0 101090.0 134975.0 ;
      RECT  100385.0 136320.0 101090.0 134975.0 ;
      RECT  100385.0 136320.0 101090.0 137665.0 ;
      RECT  100385.0 139010.0 101090.0 137665.0 ;
      RECT  100385.0 139010.0 101090.0 140355.0 ;
      RECT  100385.0 141700.0 101090.0 140355.0 ;
      RECT  100385.0 141700.0 101090.0 143045.0 ;
      RECT  100385.0 144390.0 101090.0 143045.0 ;
      RECT  100385.0 144390.0 101090.0 145735.0 ;
      RECT  100385.0 147080.0 101090.0 145735.0 ;
      RECT  100385.0 147080.0 101090.0 148425.0 ;
      RECT  100385.0 149770.0 101090.0 148425.0 ;
      RECT  100385.0 149770.0 101090.0 151115.0 ;
      RECT  100385.0 152460.0 101090.0 151115.0 ;
      RECT  100385.0 152460.0 101090.0 153805.0 ;
      RECT  100385.0 155150.0 101090.0 153805.0 ;
      RECT  100385.0 155150.0 101090.0 156495.0 ;
      RECT  100385.0 157840.0 101090.0 156495.0 ;
      RECT  100385.0 157840.0 101090.0 159185.0 ;
      RECT  100385.0 160530.0 101090.0 159185.0 ;
      RECT  100385.0 160530.0 101090.0 161875.0 ;
      RECT  100385.0 163220.0 101090.0 161875.0 ;
      RECT  100385.0 163220.0 101090.0 164565.0 ;
      RECT  100385.0 165910.0 101090.0 164565.0 ;
      RECT  100385.0 165910.0 101090.0 167255.0 ;
      RECT  100385.0 168600.0 101090.0 167255.0 ;
      RECT  100385.0 168600.0 101090.0 169945.0 ;
      RECT  100385.0 171290.0 101090.0 169945.0 ;
      RECT  100385.0 171290.0 101090.0 172635.0 ;
      RECT  100385.0 173980.0 101090.0 172635.0 ;
      RECT  100385.0 173980.0 101090.0 175325.0 ;
      RECT  100385.0 176670.0 101090.0 175325.0 ;
      RECT  100385.0 176670.0 101090.0 178015.0 ;
      RECT  100385.0 179360.0 101090.0 178015.0 ;
      RECT  100385.0 179360.0 101090.0 180705.0 ;
      RECT  100385.0 182050.0 101090.0 180705.0 ;
      RECT  100385.0 182050.0 101090.0 183395.0 ;
      RECT  100385.0 184740.0 101090.0 183395.0 ;
      RECT  100385.0 184740.0 101090.0 186085.0 ;
      RECT  100385.0 187430.0 101090.0 186085.0 ;
      RECT  100385.0 187430.0 101090.0 188775.0 ;
      RECT  100385.0 190120.0 101090.0 188775.0 ;
      RECT  100385.0 190120.0 101090.0 191465.0 ;
      RECT  100385.0 192810.0 101090.0 191465.0 ;
      RECT  100385.0 192810.0 101090.0 194155.0 ;
      RECT  100385.0 195500.0 101090.0 194155.0 ;
      RECT  100385.0 195500.0 101090.0 196845.0 ;
      RECT  100385.0 198190.0 101090.0 196845.0 ;
      RECT  100385.0 198190.0 101090.0 199535.0 ;
      RECT  100385.0 200880.0 101090.0 199535.0 ;
      RECT  100385.0 200880.0 101090.0 202225.0 ;
      RECT  100385.0 203570.0 101090.0 202225.0 ;
      RECT  100385.0 203570.0 101090.0 204915.0 ;
      RECT  100385.0 206260.0 101090.0 204915.0 ;
      RECT  101090.0 34100.0 101795.0 35445.0 ;
      RECT  101090.0 36790.0 101795.0 35445.0 ;
      RECT  101090.0 36790.0 101795.0 38135.0 ;
      RECT  101090.0 39480.0 101795.0 38135.0 ;
      RECT  101090.0 39480.0 101795.0 40825.0 ;
      RECT  101090.0 42170.0 101795.0 40825.0 ;
      RECT  101090.0 42170.0 101795.0 43515.0 ;
      RECT  101090.0 44860.0 101795.0 43515.0 ;
      RECT  101090.0 44860.0 101795.0 46205.0 ;
      RECT  101090.0 47550.0 101795.0 46205.0 ;
      RECT  101090.0 47550.0 101795.0 48895.0 ;
      RECT  101090.0 50240.0 101795.0 48895.0 ;
      RECT  101090.0 50240.0 101795.0 51585.0 ;
      RECT  101090.0 52930.0 101795.0 51585.0 ;
      RECT  101090.0 52930.0 101795.0 54275.0 ;
      RECT  101090.0 55620.0 101795.0 54275.0 ;
      RECT  101090.0 55620.0 101795.0 56965.0 ;
      RECT  101090.0 58310.0 101795.0 56965.0 ;
      RECT  101090.0 58310.0 101795.0 59655.0 ;
      RECT  101090.0 61000.0 101795.0 59655.0 ;
      RECT  101090.0 61000.0 101795.0 62345.0 ;
      RECT  101090.0 63690.0 101795.0 62345.0 ;
      RECT  101090.0 63690.0 101795.0 65035.0 ;
      RECT  101090.0 66380.0 101795.0 65035.0 ;
      RECT  101090.0 66380.0 101795.0 67725.0 ;
      RECT  101090.0 69070.0 101795.0 67725.0 ;
      RECT  101090.0 69070.0 101795.0 70415.0 ;
      RECT  101090.0 71760.0 101795.0 70415.0 ;
      RECT  101090.0 71760.0 101795.0 73105.0 ;
      RECT  101090.0 74450.0 101795.0 73105.0 ;
      RECT  101090.0 74450.0 101795.0 75795.0 ;
      RECT  101090.0 77140.0 101795.0 75795.0 ;
      RECT  101090.0 77140.0 101795.0 78485.0 ;
      RECT  101090.0 79830.0 101795.0 78485.0 ;
      RECT  101090.0 79830.0 101795.0 81175.0 ;
      RECT  101090.0 82520.0 101795.0 81175.0 ;
      RECT  101090.0 82520.0 101795.0 83865.0 ;
      RECT  101090.0 85210.0 101795.0 83865.0 ;
      RECT  101090.0 85210.0 101795.0 86555.0 ;
      RECT  101090.0 87900.0 101795.0 86555.0 ;
      RECT  101090.0 87900.0 101795.0 89245.0 ;
      RECT  101090.0 90590.0 101795.0 89245.0 ;
      RECT  101090.0 90590.0 101795.0 91935.0 ;
      RECT  101090.0 93280.0 101795.0 91935.0 ;
      RECT  101090.0 93280.0 101795.0 94625.0 ;
      RECT  101090.0 95970.0 101795.0 94625.0 ;
      RECT  101090.0 95970.0 101795.0 97315.0 ;
      RECT  101090.0 98660.0 101795.0 97315.0 ;
      RECT  101090.0 98660.0 101795.0 100005.0 ;
      RECT  101090.0 101350.0 101795.0 100005.0 ;
      RECT  101090.0 101350.0 101795.0 102695.0 ;
      RECT  101090.0 104040.0 101795.0 102695.0 ;
      RECT  101090.0 104040.0 101795.0 105385.0 ;
      RECT  101090.0 106730.0 101795.0 105385.0 ;
      RECT  101090.0 106730.0 101795.0 108075.0 ;
      RECT  101090.0 109420.0 101795.0 108075.0 ;
      RECT  101090.0 109420.0 101795.0 110765.0 ;
      RECT  101090.0 112110.0 101795.0 110765.0 ;
      RECT  101090.0 112110.0 101795.0 113455.0 ;
      RECT  101090.0 114800.0 101795.0 113455.0 ;
      RECT  101090.0 114800.0 101795.0 116145.0 ;
      RECT  101090.0 117490.0 101795.0 116145.0 ;
      RECT  101090.0 117490.0 101795.0 118835.0 ;
      RECT  101090.0 120180.0 101795.0 118835.0 ;
      RECT  101090.0 120180.0 101795.0 121525.0 ;
      RECT  101090.0 122870.0 101795.0 121525.0 ;
      RECT  101090.0 122870.0 101795.0 124215.0 ;
      RECT  101090.0 125560.0 101795.0 124215.0 ;
      RECT  101090.0 125560.0 101795.0 126905.0 ;
      RECT  101090.0 128250.0 101795.0 126905.0 ;
      RECT  101090.0 128250.0 101795.0 129595.0 ;
      RECT  101090.0 130940.0 101795.0 129595.0 ;
      RECT  101090.0 130940.0 101795.0 132285.0 ;
      RECT  101090.0 133630.0 101795.0 132285.0 ;
      RECT  101090.0 133630.0 101795.0 134975.0 ;
      RECT  101090.0 136320.0 101795.0 134975.0 ;
      RECT  101090.0 136320.0 101795.0 137665.0 ;
      RECT  101090.0 139010.0 101795.0 137665.0 ;
      RECT  101090.0 139010.0 101795.0 140355.0 ;
      RECT  101090.0 141700.0 101795.0 140355.0 ;
      RECT  101090.0 141700.0 101795.0 143045.0 ;
      RECT  101090.0 144390.0 101795.0 143045.0 ;
      RECT  101090.0 144390.0 101795.0 145735.0 ;
      RECT  101090.0 147080.0 101795.0 145735.0 ;
      RECT  101090.0 147080.0 101795.0 148425.0 ;
      RECT  101090.0 149770.0 101795.0 148425.0 ;
      RECT  101090.0 149770.0 101795.0 151115.0 ;
      RECT  101090.0 152460.0 101795.0 151115.0 ;
      RECT  101090.0 152460.0 101795.0 153805.0 ;
      RECT  101090.0 155150.0 101795.0 153805.0 ;
      RECT  101090.0 155150.0 101795.0 156495.0 ;
      RECT  101090.0 157840.0 101795.0 156495.0 ;
      RECT  101090.0 157840.0 101795.0 159185.0 ;
      RECT  101090.0 160530.0 101795.0 159185.0 ;
      RECT  101090.0 160530.0 101795.0 161875.0 ;
      RECT  101090.0 163220.0 101795.0 161875.0 ;
      RECT  101090.0 163220.0 101795.0 164565.0 ;
      RECT  101090.0 165910.0 101795.0 164565.0 ;
      RECT  101090.0 165910.0 101795.0 167255.0 ;
      RECT  101090.0 168600.0 101795.0 167255.0 ;
      RECT  101090.0 168600.0 101795.0 169945.0 ;
      RECT  101090.0 171290.0 101795.0 169945.0 ;
      RECT  101090.0 171290.0 101795.0 172635.0 ;
      RECT  101090.0 173980.0 101795.0 172635.0 ;
      RECT  101090.0 173980.0 101795.0 175325.0 ;
      RECT  101090.0 176670.0 101795.0 175325.0 ;
      RECT  101090.0 176670.0 101795.0 178015.0 ;
      RECT  101090.0 179360.0 101795.0 178015.0 ;
      RECT  101090.0 179360.0 101795.0 180705.0 ;
      RECT  101090.0 182050.0 101795.0 180705.0 ;
      RECT  101090.0 182050.0 101795.0 183395.0 ;
      RECT  101090.0 184740.0 101795.0 183395.0 ;
      RECT  101090.0 184740.0 101795.0 186085.0 ;
      RECT  101090.0 187430.0 101795.0 186085.0 ;
      RECT  101090.0 187430.0 101795.0 188775.0 ;
      RECT  101090.0 190120.0 101795.0 188775.0 ;
      RECT  101090.0 190120.0 101795.0 191465.0 ;
      RECT  101090.0 192810.0 101795.0 191465.0 ;
      RECT  101090.0 192810.0 101795.0 194155.0 ;
      RECT  101090.0 195500.0 101795.0 194155.0 ;
      RECT  101090.0 195500.0 101795.0 196845.0 ;
      RECT  101090.0 198190.0 101795.0 196845.0 ;
      RECT  101090.0 198190.0 101795.0 199535.0 ;
      RECT  101090.0 200880.0 101795.0 199535.0 ;
      RECT  101090.0 200880.0 101795.0 202225.0 ;
      RECT  101090.0 203570.0 101795.0 202225.0 ;
      RECT  101090.0 203570.0 101795.0 204915.0 ;
      RECT  101090.0 206260.0 101795.0 204915.0 ;
      RECT  101795.0 34100.0 102500.0 35445.0 ;
      RECT  101795.0 36790.0 102500.0 35445.0 ;
      RECT  101795.0 36790.0 102500.0 38135.0 ;
      RECT  101795.0 39480.0 102500.0 38135.0 ;
      RECT  101795.0 39480.0 102500.0 40825.0 ;
      RECT  101795.0 42170.0 102500.0 40825.0 ;
      RECT  101795.0 42170.0 102500.0 43515.0 ;
      RECT  101795.0 44860.0 102500.0 43515.0 ;
      RECT  101795.0 44860.0 102500.0 46205.0 ;
      RECT  101795.0 47550.0 102500.0 46205.0 ;
      RECT  101795.0 47550.0 102500.0 48895.0 ;
      RECT  101795.0 50240.0 102500.0 48895.0 ;
      RECT  101795.0 50240.0 102500.0 51585.0 ;
      RECT  101795.0 52930.0 102500.0 51585.0 ;
      RECT  101795.0 52930.0 102500.0 54275.0 ;
      RECT  101795.0 55620.0 102500.0 54275.0 ;
      RECT  101795.0 55620.0 102500.0 56965.0 ;
      RECT  101795.0 58310.0 102500.0 56965.0 ;
      RECT  101795.0 58310.0 102500.0 59655.0 ;
      RECT  101795.0 61000.0 102500.0 59655.0 ;
      RECT  101795.0 61000.0 102500.0 62345.0 ;
      RECT  101795.0 63690.0 102500.0 62345.0 ;
      RECT  101795.0 63690.0 102500.0 65035.0 ;
      RECT  101795.0 66380.0 102500.0 65035.0 ;
      RECT  101795.0 66380.0 102500.0 67725.0 ;
      RECT  101795.0 69070.0 102500.0 67725.0 ;
      RECT  101795.0 69070.0 102500.0 70415.0 ;
      RECT  101795.0 71760.0 102500.0 70415.0 ;
      RECT  101795.0 71760.0 102500.0 73105.0 ;
      RECT  101795.0 74450.0 102500.0 73105.0 ;
      RECT  101795.0 74450.0 102500.0 75795.0 ;
      RECT  101795.0 77140.0 102500.0 75795.0 ;
      RECT  101795.0 77140.0 102500.0 78485.0 ;
      RECT  101795.0 79830.0 102500.0 78485.0 ;
      RECT  101795.0 79830.0 102500.0 81175.0 ;
      RECT  101795.0 82520.0 102500.0 81175.0 ;
      RECT  101795.0 82520.0 102500.0 83865.0 ;
      RECT  101795.0 85210.0 102500.0 83865.0 ;
      RECT  101795.0 85210.0 102500.0 86555.0 ;
      RECT  101795.0 87900.0 102500.0 86555.0 ;
      RECT  101795.0 87900.0 102500.0 89245.0 ;
      RECT  101795.0 90590.0 102500.0 89245.0 ;
      RECT  101795.0 90590.0 102500.0 91935.0 ;
      RECT  101795.0 93280.0 102500.0 91935.0 ;
      RECT  101795.0 93280.0 102500.0 94625.0 ;
      RECT  101795.0 95970.0 102500.0 94625.0 ;
      RECT  101795.0 95970.0 102500.0 97315.0 ;
      RECT  101795.0 98660.0 102500.0 97315.0 ;
      RECT  101795.0 98660.0 102500.0 100005.0 ;
      RECT  101795.0 101350.0 102500.0 100005.0 ;
      RECT  101795.0 101350.0 102500.0 102695.0 ;
      RECT  101795.0 104040.0 102500.0 102695.0 ;
      RECT  101795.0 104040.0 102500.0 105385.0 ;
      RECT  101795.0 106730.0 102500.0 105385.0 ;
      RECT  101795.0 106730.0 102500.0 108075.0 ;
      RECT  101795.0 109420.0 102500.0 108075.0 ;
      RECT  101795.0 109420.0 102500.0 110765.0 ;
      RECT  101795.0 112110.0 102500.0 110765.0 ;
      RECT  101795.0 112110.0 102500.0 113455.0 ;
      RECT  101795.0 114800.0 102500.0 113455.0 ;
      RECT  101795.0 114800.0 102500.0 116145.0 ;
      RECT  101795.0 117490.0 102500.0 116145.0 ;
      RECT  101795.0 117490.0 102500.0 118835.0 ;
      RECT  101795.0 120180.0 102500.0 118835.0 ;
      RECT  101795.0 120180.0 102500.0 121525.0 ;
      RECT  101795.0 122870.0 102500.0 121525.0 ;
      RECT  101795.0 122870.0 102500.0 124215.0 ;
      RECT  101795.0 125560.0 102500.0 124215.0 ;
      RECT  101795.0 125560.0 102500.0 126905.0 ;
      RECT  101795.0 128250.0 102500.0 126905.0 ;
      RECT  101795.0 128250.0 102500.0 129595.0 ;
      RECT  101795.0 130940.0 102500.0 129595.0 ;
      RECT  101795.0 130940.0 102500.0 132285.0 ;
      RECT  101795.0 133630.0 102500.0 132285.0 ;
      RECT  101795.0 133630.0 102500.0 134975.0 ;
      RECT  101795.0 136320.0 102500.0 134975.0 ;
      RECT  101795.0 136320.0 102500.0 137665.0 ;
      RECT  101795.0 139010.0 102500.0 137665.0 ;
      RECT  101795.0 139010.0 102500.0 140355.0 ;
      RECT  101795.0 141700.0 102500.0 140355.0 ;
      RECT  101795.0 141700.0 102500.0 143045.0 ;
      RECT  101795.0 144390.0 102500.0 143045.0 ;
      RECT  101795.0 144390.0 102500.0 145735.0 ;
      RECT  101795.0 147080.0 102500.0 145735.0 ;
      RECT  101795.0 147080.0 102500.0 148425.0 ;
      RECT  101795.0 149770.0 102500.0 148425.0 ;
      RECT  101795.0 149770.0 102500.0 151115.0 ;
      RECT  101795.0 152460.0 102500.0 151115.0 ;
      RECT  101795.0 152460.0 102500.0 153805.0 ;
      RECT  101795.0 155150.0 102500.0 153805.0 ;
      RECT  101795.0 155150.0 102500.0 156495.0 ;
      RECT  101795.0 157840.0 102500.0 156495.0 ;
      RECT  101795.0 157840.0 102500.0 159185.0 ;
      RECT  101795.0 160530.0 102500.0 159185.0 ;
      RECT  101795.0 160530.0 102500.0 161875.0 ;
      RECT  101795.0 163220.0 102500.0 161875.0 ;
      RECT  101795.0 163220.0 102500.0 164565.0 ;
      RECT  101795.0 165910.0 102500.0 164565.0 ;
      RECT  101795.0 165910.0 102500.0 167255.0 ;
      RECT  101795.0 168600.0 102500.0 167255.0 ;
      RECT  101795.0 168600.0 102500.0 169945.0 ;
      RECT  101795.0 171290.0 102500.0 169945.0 ;
      RECT  101795.0 171290.0 102500.0 172635.0 ;
      RECT  101795.0 173980.0 102500.0 172635.0 ;
      RECT  101795.0 173980.0 102500.0 175325.0 ;
      RECT  101795.0 176670.0 102500.0 175325.0 ;
      RECT  101795.0 176670.0 102500.0 178015.0 ;
      RECT  101795.0 179360.0 102500.0 178015.0 ;
      RECT  101795.0 179360.0 102500.0 180705.0 ;
      RECT  101795.0 182050.0 102500.0 180705.0 ;
      RECT  101795.0 182050.0 102500.0 183395.0 ;
      RECT  101795.0 184740.0 102500.0 183395.0 ;
      RECT  101795.0 184740.0 102500.0 186085.0 ;
      RECT  101795.0 187430.0 102500.0 186085.0 ;
      RECT  101795.0 187430.0 102500.0 188775.0 ;
      RECT  101795.0 190120.0 102500.0 188775.0 ;
      RECT  101795.0 190120.0 102500.0 191465.0 ;
      RECT  101795.0 192810.0 102500.0 191465.0 ;
      RECT  101795.0 192810.0 102500.0 194155.0 ;
      RECT  101795.0 195500.0 102500.0 194155.0 ;
      RECT  101795.0 195500.0 102500.0 196845.0 ;
      RECT  101795.0 198190.0 102500.0 196845.0 ;
      RECT  101795.0 198190.0 102500.0 199535.0 ;
      RECT  101795.0 200880.0 102500.0 199535.0 ;
      RECT  101795.0 200880.0 102500.0 202225.0 ;
      RECT  101795.0 203570.0 102500.0 202225.0 ;
      RECT  101795.0 203570.0 102500.0 204915.0 ;
      RECT  101795.0 206260.0 102500.0 204915.0 ;
      RECT  102500.0 34100.0 103205.0 35445.0 ;
      RECT  102500.0 36790.0 103205.0 35445.0 ;
      RECT  102500.0 36790.0 103205.0 38135.0 ;
      RECT  102500.0 39480.0 103205.0 38135.0 ;
      RECT  102500.0 39480.0 103205.0 40825.0 ;
      RECT  102500.0 42170.0 103205.0 40825.0 ;
      RECT  102500.0 42170.0 103205.0 43515.0 ;
      RECT  102500.0 44860.0 103205.0 43515.0 ;
      RECT  102500.0 44860.0 103205.0 46205.0 ;
      RECT  102500.0 47550.0 103205.0 46205.0 ;
      RECT  102500.0 47550.0 103205.0 48895.0 ;
      RECT  102500.0 50240.0 103205.0 48895.0 ;
      RECT  102500.0 50240.0 103205.0 51585.0 ;
      RECT  102500.0 52930.0 103205.0 51585.0 ;
      RECT  102500.0 52930.0 103205.0 54275.0 ;
      RECT  102500.0 55620.0 103205.0 54275.0 ;
      RECT  102500.0 55620.0 103205.0 56965.0 ;
      RECT  102500.0 58310.0 103205.0 56965.0 ;
      RECT  102500.0 58310.0 103205.0 59655.0 ;
      RECT  102500.0 61000.0 103205.0 59655.0 ;
      RECT  102500.0 61000.0 103205.0 62345.0 ;
      RECT  102500.0 63690.0 103205.0 62345.0 ;
      RECT  102500.0 63690.0 103205.0 65035.0 ;
      RECT  102500.0 66380.0 103205.0 65035.0 ;
      RECT  102500.0 66380.0 103205.0 67725.0 ;
      RECT  102500.0 69070.0 103205.0 67725.0 ;
      RECT  102500.0 69070.0 103205.0 70415.0 ;
      RECT  102500.0 71760.0 103205.0 70415.0 ;
      RECT  102500.0 71760.0 103205.0 73105.0 ;
      RECT  102500.0 74450.0 103205.0 73105.0 ;
      RECT  102500.0 74450.0 103205.0 75795.0 ;
      RECT  102500.0 77140.0 103205.0 75795.0 ;
      RECT  102500.0 77140.0 103205.0 78485.0 ;
      RECT  102500.0 79830.0 103205.0 78485.0 ;
      RECT  102500.0 79830.0 103205.0 81175.0 ;
      RECT  102500.0 82520.0 103205.0 81175.0 ;
      RECT  102500.0 82520.0 103205.0 83865.0 ;
      RECT  102500.0 85210.0 103205.0 83865.0 ;
      RECT  102500.0 85210.0 103205.0 86555.0 ;
      RECT  102500.0 87900.0 103205.0 86555.0 ;
      RECT  102500.0 87900.0 103205.0 89245.0 ;
      RECT  102500.0 90590.0 103205.0 89245.0 ;
      RECT  102500.0 90590.0 103205.0 91935.0 ;
      RECT  102500.0 93280.0 103205.0 91935.0 ;
      RECT  102500.0 93280.0 103205.0 94625.0 ;
      RECT  102500.0 95970.0 103205.0 94625.0 ;
      RECT  102500.0 95970.0 103205.0 97315.0 ;
      RECT  102500.0 98660.0 103205.0 97315.0 ;
      RECT  102500.0 98660.0 103205.0 100005.0 ;
      RECT  102500.0 101350.0 103205.0 100005.0 ;
      RECT  102500.0 101350.0 103205.0 102695.0 ;
      RECT  102500.0 104040.0 103205.0 102695.0 ;
      RECT  102500.0 104040.0 103205.0 105385.0 ;
      RECT  102500.0 106730.0 103205.0 105385.0 ;
      RECT  102500.0 106730.0 103205.0 108075.0 ;
      RECT  102500.0 109420.0 103205.0 108075.0 ;
      RECT  102500.0 109420.0 103205.0 110765.0 ;
      RECT  102500.0 112110.0 103205.0 110765.0 ;
      RECT  102500.0 112110.0 103205.0 113455.0 ;
      RECT  102500.0 114800.0 103205.0 113455.0 ;
      RECT  102500.0 114800.0 103205.0 116145.0 ;
      RECT  102500.0 117490.0 103205.0 116145.0 ;
      RECT  102500.0 117490.0 103205.0 118835.0 ;
      RECT  102500.0 120180.0 103205.0 118835.0 ;
      RECT  102500.0 120180.0 103205.0 121525.0 ;
      RECT  102500.0 122870.0 103205.0 121525.0 ;
      RECT  102500.0 122870.0 103205.0 124215.0 ;
      RECT  102500.0 125560.0 103205.0 124215.0 ;
      RECT  102500.0 125560.0 103205.0 126905.0 ;
      RECT  102500.0 128250.0 103205.0 126905.0 ;
      RECT  102500.0 128250.0 103205.0 129595.0 ;
      RECT  102500.0 130940.0 103205.0 129595.0 ;
      RECT  102500.0 130940.0 103205.0 132285.0 ;
      RECT  102500.0 133630.0 103205.0 132285.0 ;
      RECT  102500.0 133630.0 103205.0 134975.0 ;
      RECT  102500.0 136320.0 103205.0 134975.0 ;
      RECT  102500.0 136320.0 103205.0 137665.0 ;
      RECT  102500.0 139010.0 103205.0 137665.0 ;
      RECT  102500.0 139010.0 103205.0 140355.0 ;
      RECT  102500.0 141700.0 103205.0 140355.0 ;
      RECT  102500.0 141700.0 103205.0 143045.0 ;
      RECT  102500.0 144390.0 103205.0 143045.0 ;
      RECT  102500.0 144390.0 103205.0 145735.0 ;
      RECT  102500.0 147080.0 103205.0 145735.0 ;
      RECT  102500.0 147080.0 103205.0 148425.0 ;
      RECT  102500.0 149770.0 103205.0 148425.0 ;
      RECT  102500.0 149770.0 103205.0 151115.0 ;
      RECT  102500.0 152460.0 103205.0 151115.0 ;
      RECT  102500.0 152460.0 103205.0 153805.0 ;
      RECT  102500.0 155150.0 103205.0 153805.0 ;
      RECT  102500.0 155150.0 103205.0 156495.0 ;
      RECT  102500.0 157840.0 103205.0 156495.0 ;
      RECT  102500.0 157840.0 103205.0 159185.0 ;
      RECT  102500.0 160530.0 103205.0 159185.0 ;
      RECT  102500.0 160530.0 103205.0 161875.0 ;
      RECT  102500.0 163220.0 103205.0 161875.0 ;
      RECT  102500.0 163220.0 103205.0 164565.0 ;
      RECT  102500.0 165910.0 103205.0 164565.0 ;
      RECT  102500.0 165910.0 103205.0 167255.0 ;
      RECT  102500.0 168600.0 103205.0 167255.0 ;
      RECT  102500.0 168600.0 103205.0 169945.0 ;
      RECT  102500.0 171290.0 103205.0 169945.0 ;
      RECT  102500.0 171290.0 103205.0 172635.0 ;
      RECT  102500.0 173980.0 103205.0 172635.0 ;
      RECT  102500.0 173980.0 103205.0 175325.0 ;
      RECT  102500.0 176670.0 103205.0 175325.0 ;
      RECT  102500.0 176670.0 103205.0 178015.0 ;
      RECT  102500.0 179360.0 103205.0 178015.0 ;
      RECT  102500.0 179360.0 103205.0 180705.0 ;
      RECT  102500.0 182050.0 103205.0 180705.0 ;
      RECT  102500.0 182050.0 103205.0 183395.0 ;
      RECT  102500.0 184740.0 103205.0 183395.0 ;
      RECT  102500.0 184740.0 103205.0 186085.0 ;
      RECT  102500.0 187430.0 103205.0 186085.0 ;
      RECT  102500.0 187430.0 103205.0 188775.0 ;
      RECT  102500.0 190120.0 103205.0 188775.0 ;
      RECT  102500.0 190120.0 103205.0 191465.0 ;
      RECT  102500.0 192810.0 103205.0 191465.0 ;
      RECT  102500.0 192810.0 103205.0 194155.0 ;
      RECT  102500.0 195500.0 103205.0 194155.0 ;
      RECT  102500.0 195500.0 103205.0 196845.0 ;
      RECT  102500.0 198190.0 103205.0 196845.0 ;
      RECT  102500.0 198190.0 103205.0 199535.0 ;
      RECT  102500.0 200880.0 103205.0 199535.0 ;
      RECT  102500.0 200880.0 103205.0 202225.0 ;
      RECT  102500.0 203570.0 103205.0 202225.0 ;
      RECT  102500.0 203570.0 103205.0 204915.0 ;
      RECT  102500.0 206260.0 103205.0 204915.0 ;
      RECT  103205.0 34100.0 103910.0 35445.0 ;
      RECT  103205.0 36790.0 103910.0 35445.0 ;
      RECT  103205.0 36790.0 103910.0 38135.0 ;
      RECT  103205.0 39480.0 103910.0 38135.0 ;
      RECT  103205.0 39480.0 103910.0 40825.0 ;
      RECT  103205.0 42170.0 103910.0 40825.0 ;
      RECT  103205.0 42170.0 103910.0 43515.0 ;
      RECT  103205.0 44860.0 103910.0 43515.0 ;
      RECT  103205.0 44860.0 103910.0 46205.0 ;
      RECT  103205.0 47550.0 103910.0 46205.0 ;
      RECT  103205.0 47550.0 103910.0 48895.0 ;
      RECT  103205.0 50240.0 103910.0 48895.0 ;
      RECT  103205.0 50240.0 103910.0 51585.0 ;
      RECT  103205.0 52930.0 103910.0 51585.0 ;
      RECT  103205.0 52930.0 103910.0 54275.0 ;
      RECT  103205.0 55620.0 103910.0 54275.0 ;
      RECT  103205.0 55620.0 103910.0 56965.0 ;
      RECT  103205.0 58310.0 103910.0 56965.0 ;
      RECT  103205.0 58310.0 103910.0 59655.0 ;
      RECT  103205.0 61000.0 103910.0 59655.0 ;
      RECT  103205.0 61000.0 103910.0 62345.0 ;
      RECT  103205.0 63690.0 103910.0 62345.0 ;
      RECT  103205.0 63690.0 103910.0 65035.0 ;
      RECT  103205.0 66380.0 103910.0 65035.0 ;
      RECT  103205.0 66380.0 103910.0 67725.0 ;
      RECT  103205.0 69070.0 103910.0 67725.0 ;
      RECT  103205.0 69070.0 103910.0 70415.0 ;
      RECT  103205.0 71760.0 103910.0 70415.0 ;
      RECT  103205.0 71760.0 103910.0 73105.0 ;
      RECT  103205.0 74450.0 103910.0 73105.0 ;
      RECT  103205.0 74450.0 103910.0 75795.0 ;
      RECT  103205.0 77140.0 103910.0 75795.0 ;
      RECT  103205.0 77140.0 103910.0 78485.0 ;
      RECT  103205.0 79830.0 103910.0 78485.0 ;
      RECT  103205.0 79830.0 103910.0 81175.0 ;
      RECT  103205.0 82520.0 103910.0 81175.0 ;
      RECT  103205.0 82520.0 103910.0 83865.0 ;
      RECT  103205.0 85210.0 103910.0 83865.0 ;
      RECT  103205.0 85210.0 103910.0 86555.0 ;
      RECT  103205.0 87900.0 103910.0 86555.0 ;
      RECT  103205.0 87900.0 103910.0 89245.0 ;
      RECT  103205.0 90590.0 103910.0 89245.0 ;
      RECT  103205.0 90590.0 103910.0 91935.0 ;
      RECT  103205.0 93280.0 103910.0 91935.0 ;
      RECT  103205.0 93280.0 103910.0 94625.0 ;
      RECT  103205.0 95970.0 103910.0 94625.0 ;
      RECT  103205.0 95970.0 103910.0 97315.0 ;
      RECT  103205.0 98660.0 103910.0 97315.0 ;
      RECT  103205.0 98660.0 103910.0 100005.0 ;
      RECT  103205.0 101350.0 103910.0 100005.0 ;
      RECT  103205.0 101350.0 103910.0 102695.0 ;
      RECT  103205.0 104040.0 103910.0 102695.0 ;
      RECT  103205.0 104040.0 103910.0 105385.0 ;
      RECT  103205.0 106730.0 103910.0 105385.0 ;
      RECT  103205.0 106730.0 103910.0 108075.0 ;
      RECT  103205.0 109420.0 103910.0 108075.0 ;
      RECT  103205.0 109420.0 103910.0 110765.0 ;
      RECT  103205.0 112110.0 103910.0 110765.0 ;
      RECT  103205.0 112110.0 103910.0 113455.0 ;
      RECT  103205.0 114800.0 103910.0 113455.0 ;
      RECT  103205.0 114800.0 103910.0 116145.0 ;
      RECT  103205.0 117490.0 103910.0 116145.0 ;
      RECT  103205.0 117490.0 103910.0 118835.0 ;
      RECT  103205.0 120180.0 103910.0 118835.0 ;
      RECT  103205.0 120180.0 103910.0 121525.0 ;
      RECT  103205.0 122870.0 103910.0 121525.0 ;
      RECT  103205.0 122870.0 103910.0 124215.0 ;
      RECT  103205.0 125560.0 103910.0 124215.0 ;
      RECT  103205.0 125560.0 103910.0 126905.0 ;
      RECT  103205.0 128250.0 103910.0 126905.0 ;
      RECT  103205.0 128250.0 103910.0 129595.0 ;
      RECT  103205.0 130940.0 103910.0 129595.0 ;
      RECT  103205.0 130940.0 103910.0 132285.0 ;
      RECT  103205.0 133630.0 103910.0 132285.0 ;
      RECT  103205.0 133630.0 103910.0 134975.0 ;
      RECT  103205.0 136320.0 103910.0 134975.0 ;
      RECT  103205.0 136320.0 103910.0 137665.0 ;
      RECT  103205.0 139010.0 103910.0 137665.0 ;
      RECT  103205.0 139010.0 103910.0 140355.0 ;
      RECT  103205.0 141700.0 103910.0 140355.0 ;
      RECT  103205.0 141700.0 103910.0 143045.0 ;
      RECT  103205.0 144390.0 103910.0 143045.0 ;
      RECT  103205.0 144390.0 103910.0 145735.0 ;
      RECT  103205.0 147080.0 103910.0 145735.0 ;
      RECT  103205.0 147080.0 103910.0 148425.0 ;
      RECT  103205.0 149770.0 103910.0 148425.0 ;
      RECT  103205.0 149770.0 103910.0 151115.0 ;
      RECT  103205.0 152460.0 103910.0 151115.0 ;
      RECT  103205.0 152460.0 103910.0 153805.0 ;
      RECT  103205.0 155150.0 103910.0 153805.0 ;
      RECT  103205.0 155150.0 103910.0 156495.0 ;
      RECT  103205.0 157840.0 103910.0 156495.0 ;
      RECT  103205.0 157840.0 103910.0 159185.0 ;
      RECT  103205.0 160530.0 103910.0 159185.0 ;
      RECT  103205.0 160530.0 103910.0 161875.0 ;
      RECT  103205.0 163220.0 103910.0 161875.0 ;
      RECT  103205.0 163220.0 103910.0 164565.0 ;
      RECT  103205.0 165910.0 103910.0 164565.0 ;
      RECT  103205.0 165910.0 103910.0 167255.0 ;
      RECT  103205.0 168600.0 103910.0 167255.0 ;
      RECT  103205.0 168600.0 103910.0 169945.0 ;
      RECT  103205.0 171290.0 103910.0 169945.0 ;
      RECT  103205.0 171290.0 103910.0 172635.0 ;
      RECT  103205.0 173980.0 103910.0 172635.0 ;
      RECT  103205.0 173980.0 103910.0 175325.0 ;
      RECT  103205.0 176670.0 103910.0 175325.0 ;
      RECT  103205.0 176670.0 103910.0 178015.0 ;
      RECT  103205.0 179360.0 103910.0 178015.0 ;
      RECT  103205.0 179360.0 103910.0 180705.0 ;
      RECT  103205.0 182050.0 103910.0 180705.0 ;
      RECT  103205.0 182050.0 103910.0 183395.0 ;
      RECT  103205.0 184740.0 103910.0 183395.0 ;
      RECT  103205.0 184740.0 103910.0 186085.0 ;
      RECT  103205.0 187430.0 103910.0 186085.0 ;
      RECT  103205.0 187430.0 103910.0 188775.0 ;
      RECT  103205.0 190120.0 103910.0 188775.0 ;
      RECT  103205.0 190120.0 103910.0 191465.0 ;
      RECT  103205.0 192810.0 103910.0 191465.0 ;
      RECT  103205.0 192810.0 103910.0 194155.0 ;
      RECT  103205.0 195500.0 103910.0 194155.0 ;
      RECT  103205.0 195500.0 103910.0 196845.0 ;
      RECT  103205.0 198190.0 103910.0 196845.0 ;
      RECT  103205.0 198190.0 103910.0 199535.0 ;
      RECT  103205.0 200880.0 103910.0 199535.0 ;
      RECT  103205.0 200880.0 103910.0 202225.0 ;
      RECT  103205.0 203570.0 103910.0 202225.0 ;
      RECT  103205.0 203570.0 103910.0 204915.0 ;
      RECT  103205.0 206260.0 103910.0 204915.0 ;
      RECT  103910.0 34100.0 104615.0 35445.0 ;
      RECT  103910.0 36790.0 104615.0 35445.0 ;
      RECT  103910.0 36790.0 104615.0 38135.0 ;
      RECT  103910.0 39480.0 104615.0 38135.0 ;
      RECT  103910.0 39480.0 104615.0 40825.0 ;
      RECT  103910.0 42170.0 104615.0 40825.0 ;
      RECT  103910.0 42170.0 104615.0 43515.0 ;
      RECT  103910.0 44860.0 104615.0 43515.0 ;
      RECT  103910.0 44860.0 104615.0 46205.0 ;
      RECT  103910.0 47550.0 104615.0 46205.0 ;
      RECT  103910.0 47550.0 104615.0 48895.0 ;
      RECT  103910.0 50240.0 104615.0 48895.0 ;
      RECT  103910.0 50240.0 104615.0 51585.0 ;
      RECT  103910.0 52930.0 104615.0 51585.0 ;
      RECT  103910.0 52930.0 104615.0 54275.0 ;
      RECT  103910.0 55620.0 104615.0 54275.0 ;
      RECT  103910.0 55620.0 104615.0 56965.0 ;
      RECT  103910.0 58310.0 104615.0 56965.0 ;
      RECT  103910.0 58310.0 104615.0 59655.0 ;
      RECT  103910.0 61000.0 104615.0 59655.0 ;
      RECT  103910.0 61000.0 104615.0 62345.0 ;
      RECT  103910.0 63690.0 104615.0 62345.0 ;
      RECT  103910.0 63690.0 104615.0 65035.0 ;
      RECT  103910.0 66380.0 104615.0 65035.0 ;
      RECT  103910.0 66380.0 104615.0 67725.0 ;
      RECT  103910.0 69070.0 104615.0 67725.0 ;
      RECT  103910.0 69070.0 104615.0 70415.0 ;
      RECT  103910.0 71760.0 104615.0 70415.0 ;
      RECT  103910.0 71760.0 104615.0 73105.0 ;
      RECT  103910.0 74450.0 104615.0 73105.0 ;
      RECT  103910.0 74450.0 104615.0 75795.0 ;
      RECT  103910.0 77140.0 104615.0 75795.0 ;
      RECT  103910.0 77140.0 104615.0 78485.0 ;
      RECT  103910.0 79830.0 104615.0 78485.0 ;
      RECT  103910.0 79830.0 104615.0 81175.0 ;
      RECT  103910.0 82520.0 104615.0 81175.0 ;
      RECT  103910.0 82520.0 104615.0 83865.0 ;
      RECT  103910.0 85210.0 104615.0 83865.0 ;
      RECT  103910.0 85210.0 104615.0 86555.0 ;
      RECT  103910.0 87900.0 104615.0 86555.0 ;
      RECT  103910.0 87900.0 104615.0 89245.0 ;
      RECT  103910.0 90590.0 104615.0 89245.0 ;
      RECT  103910.0 90590.0 104615.0 91935.0 ;
      RECT  103910.0 93280.0 104615.0 91935.0 ;
      RECT  103910.0 93280.0 104615.0 94625.0 ;
      RECT  103910.0 95970.0 104615.0 94625.0 ;
      RECT  103910.0 95970.0 104615.0 97315.0 ;
      RECT  103910.0 98660.0 104615.0 97315.0 ;
      RECT  103910.0 98660.0 104615.0 100005.0 ;
      RECT  103910.0 101350.0 104615.0 100005.0 ;
      RECT  103910.0 101350.0 104615.0 102695.0 ;
      RECT  103910.0 104040.0 104615.0 102695.0 ;
      RECT  103910.0 104040.0 104615.0 105385.0 ;
      RECT  103910.0 106730.0 104615.0 105385.0 ;
      RECT  103910.0 106730.0 104615.0 108075.0 ;
      RECT  103910.0 109420.0 104615.0 108075.0 ;
      RECT  103910.0 109420.0 104615.0 110765.0 ;
      RECT  103910.0 112110.0 104615.0 110765.0 ;
      RECT  103910.0 112110.0 104615.0 113455.0 ;
      RECT  103910.0 114800.0 104615.0 113455.0 ;
      RECT  103910.0 114800.0 104615.0 116145.0 ;
      RECT  103910.0 117490.0 104615.0 116145.0 ;
      RECT  103910.0 117490.0 104615.0 118835.0 ;
      RECT  103910.0 120180.0 104615.0 118835.0 ;
      RECT  103910.0 120180.0 104615.0 121525.0 ;
      RECT  103910.0 122870.0 104615.0 121525.0 ;
      RECT  103910.0 122870.0 104615.0 124215.0 ;
      RECT  103910.0 125560.0 104615.0 124215.0 ;
      RECT  103910.0 125560.0 104615.0 126905.0 ;
      RECT  103910.0 128250.0 104615.0 126905.0 ;
      RECT  103910.0 128250.0 104615.0 129595.0 ;
      RECT  103910.0 130940.0 104615.0 129595.0 ;
      RECT  103910.0 130940.0 104615.0 132285.0 ;
      RECT  103910.0 133630.0 104615.0 132285.0 ;
      RECT  103910.0 133630.0 104615.0 134975.0 ;
      RECT  103910.0 136320.0 104615.0 134975.0 ;
      RECT  103910.0 136320.0 104615.0 137665.0 ;
      RECT  103910.0 139010.0 104615.0 137665.0 ;
      RECT  103910.0 139010.0 104615.0 140355.0 ;
      RECT  103910.0 141700.0 104615.0 140355.0 ;
      RECT  103910.0 141700.0 104615.0 143045.0 ;
      RECT  103910.0 144390.0 104615.0 143045.0 ;
      RECT  103910.0 144390.0 104615.0 145735.0 ;
      RECT  103910.0 147080.0 104615.0 145735.0 ;
      RECT  103910.0 147080.0 104615.0 148425.0 ;
      RECT  103910.0 149770.0 104615.0 148425.0 ;
      RECT  103910.0 149770.0 104615.0 151115.0 ;
      RECT  103910.0 152460.0 104615.0 151115.0 ;
      RECT  103910.0 152460.0 104615.0 153805.0 ;
      RECT  103910.0 155150.0 104615.0 153805.0 ;
      RECT  103910.0 155150.0 104615.0 156495.0 ;
      RECT  103910.0 157840.0 104615.0 156495.0 ;
      RECT  103910.0 157840.0 104615.0 159185.0 ;
      RECT  103910.0 160530.0 104615.0 159185.0 ;
      RECT  103910.0 160530.0 104615.0 161875.0 ;
      RECT  103910.0 163220.0 104615.0 161875.0 ;
      RECT  103910.0 163220.0 104615.0 164565.0 ;
      RECT  103910.0 165910.0 104615.0 164565.0 ;
      RECT  103910.0 165910.0 104615.0 167255.0 ;
      RECT  103910.0 168600.0 104615.0 167255.0 ;
      RECT  103910.0 168600.0 104615.0 169945.0 ;
      RECT  103910.0 171290.0 104615.0 169945.0 ;
      RECT  103910.0 171290.0 104615.0 172635.0 ;
      RECT  103910.0 173980.0 104615.0 172635.0 ;
      RECT  103910.0 173980.0 104615.0 175325.0 ;
      RECT  103910.0 176670.0 104615.0 175325.0 ;
      RECT  103910.0 176670.0 104615.0 178015.0 ;
      RECT  103910.0 179360.0 104615.0 178015.0 ;
      RECT  103910.0 179360.0 104615.0 180705.0 ;
      RECT  103910.0 182050.0 104615.0 180705.0 ;
      RECT  103910.0 182050.0 104615.0 183395.0 ;
      RECT  103910.0 184740.0 104615.0 183395.0 ;
      RECT  103910.0 184740.0 104615.0 186085.0 ;
      RECT  103910.0 187430.0 104615.0 186085.0 ;
      RECT  103910.0 187430.0 104615.0 188775.0 ;
      RECT  103910.0 190120.0 104615.0 188775.0 ;
      RECT  103910.0 190120.0 104615.0 191465.0 ;
      RECT  103910.0 192810.0 104615.0 191465.0 ;
      RECT  103910.0 192810.0 104615.0 194155.0 ;
      RECT  103910.0 195500.0 104615.0 194155.0 ;
      RECT  103910.0 195500.0 104615.0 196845.0 ;
      RECT  103910.0 198190.0 104615.0 196845.0 ;
      RECT  103910.0 198190.0 104615.0 199535.0 ;
      RECT  103910.0 200880.0 104615.0 199535.0 ;
      RECT  103910.0 200880.0 104615.0 202225.0 ;
      RECT  103910.0 203570.0 104615.0 202225.0 ;
      RECT  103910.0 203570.0 104615.0 204915.0 ;
      RECT  103910.0 206260.0 104615.0 204915.0 ;
      RECT  104615.0 34100.0 105320.0 35445.0 ;
      RECT  104615.0 36790.0 105320.0 35445.0 ;
      RECT  104615.0 36790.0 105320.0 38135.0 ;
      RECT  104615.0 39480.0 105320.0 38135.0 ;
      RECT  104615.0 39480.0 105320.0 40825.0 ;
      RECT  104615.0 42170.0 105320.0 40825.0 ;
      RECT  104615.0 42170.0 105320.0 43515.0 ;
      RECT  104615.0 44860.0 105320.0 43515.0 ;
      RECT  104615.0 44860.0 105320.0 46205.0 ;
      RECT  104615.0 47550.0 105320.0 46205.0 ;
      RECT  104615.0 47550.0 105320.0 48895.0 ;
      RECT  104615.0 50240.0 105320.0 48895.0 ;
      RECT  104615.0 50240.0 105320.0 51585.0 ;
      RECT  104615.0 52930.0 105320.0 51585.0 ;
      RECT  104615.0 52930.0 105320.0 54275.0 ;
      RECT  104615.0 55620.0 105320.0 54275.0 ;
      RECT  104615.0 55620.0 105320.0 56965.0 ;
      RECT  104615.0 58310.0 105320.0 56965.0 ;
      RECT  104615.0 58310.0 105320.0 59655.0 ;
      RECT  104615.0 61000.0 105320.0 59655.0 ;
      RECT  104615.0 61000.0 105320.0 62345.0 ;
      RECT  104615.0 63690.0 105320.0 62345.0 ;
      RECT  104615.0 63690.0 105320.0 65035.0 ;
      RECT  104615.0 66380.0 105320.0 65035.0 ;
      RECT  104615.0 66380.0 105320.0 67725.0 ;
      RECT  104615.0 69070.0 105320.0 67725.0 ;
      RECT  104615.0 69070.0 105320.0 70415.0 ;
      RECT  104615.0 71760.0 105320.0 70415.0 ;
      RECT  104615.0 71760.0 105320.0 73105.0 ;
      RECT  104615.0 74450.0 105320.0 73105.0 ;
      RECT  104615.0 74450.0 105320.0 75795.0 ;
      RECT  104615.0 77140.0 105320.0 75795.0 ;
      RECT  104615.0 77140.0 105320.0 78485.0 ;
      RECT  104615.0 79830.0 105320.0 78485.0 ;
      RECT  104615.0 79830.0 105320.0 81175.0 ;
      RECT  104615.0 82520.0 105320.0 81175.0 ;
      RECT  104615.0 82520.0 105320.0 83865.0 ;
      RECT  104615.0 85210.0 105320.0 83865.0 ;
      RECT  104615.0 85210.0 105320.0 86555.0 ;
      RECT  104615.0 87900.0 105320.0 86555.0 ;
      RECT  104615.0 87900.0 105320.0 89245.0 ;
      RECT  104615.0 90590.0 105320.0 89245.0 ;
      RECT  104615.0 90590.0 105320.0 91935.0 ;
      RECT  104615.0 93280.0 105320.0 91935.0 ;
      RECT  104615.0 93280.0 105320.0 94625.0 ;
      RECT  104615.0 95970.0 105320.0 94625.0 ;
      RECT  104615.0 95970.0 105320.0 97315.0 ;
      RECT  104615.0 98660.0 105320.0 97315.0 ;
      RECT  104615.0 98660.0 105320.0 100005.0 ;
      RECT  104615.0 101350.0 105320.0 100005.0 ;
      RECT  104615.0 101350.0 105320.0 102695.0 ;
      RECT  104615.0 104040.0 105320.0 102695.0 ;
      RECT  104615.0 104040.0 105320.0 105385.0 ;
      RECT  104615.0 106730.0 105320.0 105385.0 ;
      RECT  104615.0 106730.0 105320.0 108075.0 ;
      RECT  104615.0 109420.0 105320.0 108075.0 ;
      RECT  104615.0 109420.0 105320.0 110765.0 ;
      RECT  104615.0 112110.0 105320.0 110765.0 ;
      RECT  104615.0 112110.0 105320.0 113455.0 ;
      RECT  104615.0 114800.0 105320.0 113455.0 ;
      RECT  104615.0 114800.0 105320.0 116145.0 ;
      RECT  104615.0 117490.0 105320.0 116145.0 ;
      RECT  104615.0 117490.0 105320.0 118835.0 ;
      RECT  104615.0 120180.0 105320.0 118835.0 ;
      RECT  104615.0 120180.0 105320.0 121525.0 ;
      RECT  104615.0 122870.0 105320.0 121525.0 ;
      RECT  104615.0 122870.0 105320.0 124215.0 ;
      RECT  104615.0 125560.0 105320.0 124215.0 ;
      RECT  104615.0 125560.0 105320.0 126905.0 ;
      RECT  104615.0 128250.0 105320.0 126905.0 ;
      RECT  104615.0 128250.0 105320.0 129595.0 ;
      RECT  104615.0 130940.0 105320.0 129595.0 ;
      RECT  104615.0 130940.0 105320.0 132285.0 ;
      RECT  104615.0 133630.0 105320.0 132285.0 ;
      RECT  104615.0 133630.0 105320.0 134975.0 ;
      RECT  104615.0 136320.0 105320.0 134975.0 ;
      RECT  104615.0 136320.0 105320.0 137665.0 ;
      RECT  104615.0 139010.0 105320.0 137665.0 ;
      RECT  104615.0 139010.0 105320.0 140355.0 ;
      RECT  104615.0 141700.0 105320.0 140355.0 ;
      RECT  104615.0 141700.0 105320.0 143045.0 ;
      RECT  104615.0 144390.0 105320.0 143045.0 ;
      RECT  104615.0 144390.0 105320.0 145735.0 ;
      RECT  104615.0 147080.0 105320.0 145735.0 ;
      RECT  104615.0 147080.0 105320.0 148425.0 ;
      RECT  104615.0 149770.0 105320.0 148425.0 ;
      RECT  104615.0 149770.0 105320.0 151115.0 ;
      RECT  104615.0 152460.0 105320.0 151115.0 ;
      RECT  104615.0 152460.0 105320.0 153805.0 ;
      RECT  104615.0 155150.0 105320.0 153805.0 ;
      RECT  104615.0 155150.0 105320.0 156495.0 ;
      RECT  104615.0 157840.0 105320.0 156495.0 ;
      RECT  104615.0 157840.0 105320.0 159185.0 ;
      RECT  104615.0 160530.0 105320.0 159185.0 ;
      RECT  104615.0 160530.0 105320.0 161875.0 ;
      RECT  104615.0 163220.0 105320.0 161875.0 ;
      RECT  104615.0 163220.0 105320.0 164565.0 ;
      RECT  104615.0 165910.0 105320.0 164565.0 ;
      RECT  104615.0 165910.0 105320.0 167255.0 ;
      RECT  104615.0 168600.0 105320.0 167255.0 ;
      RECT  104615.0 168600.0 105320.0 169945.0 ;
      RECT  104615.0 171290.0 105320.0 169945.0 ;
      RECT  104615.0 171290.0 105320.0 172635.0 ;
      RECT  104615.0 173980.0 105320.0 172635.0 ;
      RECT  104615.0 173980.0 105320.0 175325.0 ;
      RECT  104615.0 176670.0 105320.0 175325.0 ;
      RECT  104615.0 176670.0 105320.0 178015.0 ;
      RECT  104615.0 179360.0 105320.0 178015.0 ;
      RECT  104615.0 179360.0 105320.0 180705.0 ;
      RECT  104615.0 182050.0 105320.0 180705.0 ;
      RECT  104615.0 182050.0 105320.0 183395.0 ;
      RECT  104615.0 184740.0 105320.0 183395.0 ;
      RECT  104615.0 184740.0 105320.0 186085.0 ;
      RECT  104615.0 187430.0 105320.0 186085.0 ;
      RECT  104615.0 187430.0 105320.0 188775.0 ;
      RECT  104615.0 190120.0 105320.0 188775.0 ;
      RECT  104615.0 190120.0 105320.0 191465.0 ;
      RECT  104615.0 192810.0 105320.0 191465.0 ;
      RECT  104615.0 192810.0 105320.0 194155.0 ;
      RECT  104615.0 195500.0 105320.0 194155.0 ;
      RECT  104615.0 195500.0 105320.0 196845.0 ;
      RECT  104615.0 198190.0 105320.0 196845.0 ;
      RECT  104615.0 198190.0 105320.0 199535.0 ;
      RECT  104615.0 200880.0 105320.0 199535.0 ;
      RECT  104615.0 200880.0 105320.0 202225.0 ;
      RECT  104615.0 203570.0 105320.0 202225.0 ;
      RECT  104615.0 203570.0 105320.0 204915.0 ;
      RECT  104615.0 206260.0 105320.0 204915.0 ;
      RECT  105320.0 34100.0 106025.0 35445.0 ;
      RECT  105320.0 36790.0 106025.0 35445.0 ;
      RECT  105320.0 36790.0 106025.0 38135.0 ;
      RECT  105320.0 39480.0 106025.0 38135.0 ;
      RECT  105320.0 39480.0 106025.0 40825.0 ;
      RECT  105320.0 42170.0 106025.0 40825.0 ;
      RECT  105320.0 42170.0 106025.0 43515.0 ;
      RECT  105320.0 44860.0 106025.0 43515.0 ;
      RECT  105320.0 44860.0 106025.0 46205.0 ;
      RECT  105320.0 47550.0 106025.0 46205.0 ;
      RECT  105320.0 47550.0 106025.0 48895.0 ;
      RECT  105320.0 50240.0 106025.0 48895.0 ;
      RECT  105320.0 50240.0 106025.0 51585.0 ;
      RECT  105320.0 52930.0 106025.0 51585.0 ;
      RECT  105320.0 52930.0 106025.0 54275.0 ;
      RECT  105320.0 55620.0 106025.0 54275.0 ;
      RECT  105320.0 55620.0 106025.0 56965.0 ;
      RECT  105320.0 58310.0 106025.0 56965.0 ;
      RECT  105320.0 58310.0 106025.0 59655.0 ;
      RECT  105320.0 61000.0 106025.0 59655.0 ;
      RECT  105320.0 61000.0 106025.0 62345.0 ;
      RECT  105320.0 63690.0 106025.0 62345.0 ;
      RECT  105320.0 63690.0 106025.0 65035.0 ;
      RECT  105320.0 66380.0 106025.0 65035.0 ;
      RECT  105320.0 66380.0 106025.0 67725.0 ;
      RECT  105320.0 69070.0 106025.0 67725.0 ;
      RECT  105320.0 69070.0 106025.0 70415.0 ;
      RECT  105320.0 71760.0 106025.0 70415.0 ;
      RECT  105320.0 71760.0 106025.0 73105.0 ;
      RECT  105320.0 74450.0 106025.0 73105.0 ;
      RECT  105320.0 74450.0 106025.0 75795.0 ;
      RECT  105320.0 77140.0 106025.0 75795.0 ;
      RECT  105320.0 77140.0 106025.0 78485.0 ;
      RECT  105320.0 79830.0 106025.0 78485.0 ;
      RECT  105320.0 79830.0 106025.0 81175.0 ;
      RECT  105320.0 82520.0 106025.0 81175.0 ;
      RECT  105320.0 82520.0 106025.0 83865.0 ;
      RECT  105320.0 85210.0 106025.0 83865.0 ;
      RECT  105320.0 85210.0 106025.0 86555.0 ;
      RECT  105320.0 87900.0 106025.0 86555.0 ;
      RECT  105320.0 87900.0 106025.0 89245.0 ;
      RECT  105320.0 90590.0 106025.0 89245.0 ;
      RECT  105320.0 90590.0 106025.0 91935.0 ;
      RECT  105320.0 93280.0 106025.0 91935.0 ;
      RECT  105320.0 93280.0 106025.0 94625.0 ;
      RECT  105320.0 95970.0 106025.0 94625.0 ;
      RECT  105320.0 95970.0 106025.0 97315.0 ;
      RECT  105320.0 98660.0 106025.0 97315.0 ;
      RECT  105320.0 98660.0 106025.0 100005.0 ;
      RECT  105320.0 101350.0 106025.0 100005.0 ;
      RECT  105320.0 101350.0 106025.0 102695.0 ;
      RECT  105320.0 104040.0 106025.0 102695.0 ;
      RECT  105320.0 104040.0 106025.0 105385.0 ;
      RECT  105320.0 106730.0 106025.0 105385.0 ;
      RECT  105320.0 106730.0 106025.0 108075.0 ;
      RECT  105320.0 109420.0 106025.0 108075.0 ;
      RECT  105320.0 109420.0 106025.0 110765.0 ;
      RECT  105320.0 112110.0 106025.0 110765.0 ;
      RECT  105320.0 112110.0 106025.0 113455.0 ;
      RECT  105320.0 114800.0 106025.0 113455.0 ;
      RECT  105320.0 114800.0 106025.0 116145.0 ;
      RECT  105320.0 117490.0 106025.0 116145.0 ;
      RECT  105320.0 117490.0 106025.0 118835.0 ;
      RECT  105320.0 120180.0 106025.0 118835.0 ;
      RECT  105320.0 120180.0 106025.0 121525.0 ;
      RECT  105320.0 122870.0 106025.0 121525.0 ;
      RECT  105320.0 122870.0 106025.0 124215.0 ;
      RECT  105320.0 125560.0 106025.0 124215.0 ;
      RECT  105320.0 125560.0 106025.0 126905.0 ;
      RECT  105320.0 128250.0 106025.0 126905.0 ;
      RECT  105320.0 128250.0 106025.0 129595.0 ;
      RECT  105320.0 130940.0 106025.0 129595.0 ;
      RECT  105320.0 130940.0 106025.0 132285.0 ;
      RECT  105320.0 133630.0 106025.0 132285.0 ;
      RECT  105320.0 133630.0 106025.0 134975.0 ;
      RECT  105320.0 136320.0 106025.0 134975.0 ;
      RECT  105320.0 136320.0 106025.0 137665.0 ;
      RECT  105320.0 139010.0 106025.0 137665.0 ;
      RECT  105320.0 139010.0 106025.0 140355.0 ;
      RECT  105320.0 141700.0 106025.0 140355.0 ;
      RECT  105320.0 141700.0 106025.0 143045.0 ;
      RECT  105320.0 144390.0 106025.0 143045.0 ;
      RECT  105320.0 144390.0 106025.0 145735.0 ;
      RECT  105320.0 147080.0 106025.0 145735.0 ;
      RECT  105320.0 147080.0 106025.0 148425.0 ;
      RECT  105320.0 149770.0 106025.0 148425.0 ;
      RECT  105320.0 149770.0 106025.0 151115.0 ;
      RECT  105320.0 152460.0 106025.0 151115.0 ;
      RECT  105320.0 152460.0 106025.0 153805.0 ;
      RECT  105320.0 155150.0 106025.0 153805.0 ;
      RECT  105320.0 155150.0 106025.0 156495.0 ;
      RECT  105320.0 157840.0 106025.0 156495.0 ;
      RECT  105320.0 157840.0 106025.0 159185.0 ;
      RECT  105320.0 160530.0 106025.0 159185.0 ;
      RECT  105320.0 160530.0 106025.0 161875.0 ;
      RECT  105320.0 163220.0 106025.0 161875.0 ;
      RECT  105320.0 163220.0 106025.0 164565.0 ;
      RECT  105320.0 165910.0 106025.0 164565.0 ;
      RECT  105320.0 165910.0 106025.0 167255.0 ;
      RECT  105320.0 168600.0 106025.0 167255.0 ;
      RECT  105320.0 168600.0 106025.0 169945.0 ;
      RECT  105320.0 171290.0 106025.0 169945.0 ;
      RECT  105320.0 171290.0 106025.0 172635.0 ;
      RECT  105320.0 173980.0 106025.0 172635.0 ;
      RECT  105320.0 173980.0 106025.0 175325.0 ;
      RECT  105320.0 176670.0 106025.0 175325.0 ;
      RECT  105320.0 176670.0 106025.0 178015.0 ;
      RECT  105320.0 179360.0 106025.0 178015.0 ;
      RECT  105320.0 179360.0 106025.0 180705.0 ;
      RECT  105320.0 182050.0 106025.0 180705.0 ;
      RECT  105320.0 182050.0 106025.0 183395.0 ;
      RECT  105320.0 184740.0 106025.0 183395.0 ;
      RECT  105320.0 184740.0 106025.0 186085.0 ;
      RECT  105320.0 187430.0 106025.0 186085.0 ;
      RECT  105320.0 187430.0 106025.0 188775.0 ;
      RECT  105320.0 190120.0 106025.0 188775.0 ;
      RECT  105320.0 190120.0 106025.0 191465.0 ;
      RECT  105320.0 192810.0 106025.0 191465.0 ;
      RECT  105320.0 192810.0 106025.0 194155.0 ;
      RECT  105320.0 195500.0 106025.0 194155.0 ;
      RECT  105320.0 195500.0 106025.0 196845.0 ;
      RECT  105320.0 198190.0 106025.0 196845.0 ;
      RECT  105320.0 198190.0 106025.0 199535.0 ;
      RECT  105320.0 200880.0 106025.0 199535.0 ;
      RECT  105320.0 200880.0 106025.0 202225.0 ;
      RECT  105320.0 203570.0 106025.0 202225.0 ;
      RECT  105320.0 203570.0 106025.0 204915.0 ;
      RECT  105320.0 206260.0 106025.0 204915.0 ;
      RECT  106025.0 34100.0 106730.0 35445.0 ;
      RECT  106025.0 36790.0 106730.0 35445.0 ;
      RECT  106025.0 36790.0 106730.0 38135.0 ;
      RECT  106025.0 39480.0 106730.0 38135.0 ;
      RECT  106025.0 39480.0 106730.0 40825.0 ;
      RECT  106025.0 42170.0 106730.0 40825.0 ;
      RECT  106025.0 42170.0 106730.0 43515.0 ;
      RECT  106025.0 44860.0 106730.0 43515.0 ;
      RECT  106025.0 44860.0 106730.0 46205.0 ;
      RECT  106025.0 47550.0 106730.0 46205.0 ;
      RECT  106025.0 47550.0 106730.0 48895.0 ;
      RECT  106025.0 50240.0 106730.0 48895.0 ;
      RECT  106025.0 50240.0 106730.0 51585.0 ;
      RECT  106025.0 52930.0 106730.0 51585.0 ;
      RECT  106025.0 52930.0 106730.0 54275.0 ;
      RECT  106025.0 55620.0 106730.0 54275.0 ;
      RECT  106025.0 55620.0 106730.0 56965.0 ;
      RECT  106025.0 58310.0 106730.0 56965.0 ;
      RECT  106025.0 58310.0 106730.0 59655.0 ;
      RECT  106025.0 61000.0 106730.0 59655.0 ;
      RECT  106025.0 61000.0 106730.0 62345.0 ;
      RECT  106025.0 63690.0 106730.0 62345.0 ;
      RECT  106025.0 63690.0 106730.0 65035.0 ;
      RECT  106025.0 66380.0 106730.0 65035.0 ;
      RECT  106025.0 66380.0 106730.0 67725.0 ;
      RECT  106025.0 69070.0 106730.0 67725.0 ;
      RECT  106025.0 69070.0 106730.0 70415.0 ;
      RECT  106025.0 71760.0 106730.0 70415.0 ;
      RECT  106025.0 71760.0 106730.0 73105.0 ;
      RECT  106025.0 74450.0 106730.0 73105.0 ;
      RECT  106025.0 74450.0 106730.0 75795.0 ;
      RECT  106025.0 77140.0 106730.0 75795.0 ;
      RECT  106025.0 77140.0 106730.0 78485.0 ;
      RECT  106025.0 79830.0 106730.0 78485.0 ;
      RECT  106025.0 79830.0 106730.0 81175.0 ;
      RECT  106025.0 82520.0 106730.0 81175.0 ;
      RECT  106025.0 82520.0 106730.0 83865.0 ;
      RECT  106025.0 85210.0 106730.0 83865.0 ;
      RECT  106025.0 85210.0 106730.0 86555.0 ;
      RECT  106025.0 87900.0 106730.0 86555.0 ;
      RECT  106025.0 87900.0 106730.0 89245.0 ;
      RECT  106025.0 90590.0 106730.0 89245.0 ;
      RECT  106025.0 90590.0 106730.0 91935.0 ;
      RECT  106025.0 93280.0 106730.0 91935.0 ;
      RECT  106025.0 93280.0 106730.0 94625.0 ;
      RECT  106025.0 95970.0 106730.0 94625.0 ;
      RECT  106025.0 95970.0 106730.0 97315.0 ;
      RECT  106025.0 98660.0 106730.0 97315.0 ;
      RECT  106025.0 98660.0 106730.0 100005.0 ;
      RECT  106025.0 101350.0 106730.0 100005.0 ;
      RECT  106025.0 101350.0 106730.0 102695.0 ;
      RECT  106025.0 104040.0 106730.0 102695.0 ;
      RECT  106025.0 104040.0 106730.0 105385.0 ;
      RECT  106025.0 106730.0 106730.0 105385.0 ;
      RECT  106025.0 106730.0 106730.0 108075.0 ;
      RECT  106025.0 109420.0 106730.0 108075.0 ;
      RECT  106025.0 109420.0 106730.0 110765.0 ;
      RECT  106025.0 112110.0 106730.0 110765.0 ;
      RECT  106025.0 112110.0 106730.0 113455.0 ;
      RECT  106025.0 114800.0 106730.0 113455.0 ;
      RECT  106025.0 114800.0 106730.0 116145.0 ;
      RECT  106025.0 117490.0 106730.0 116145.0 ;
      RECT  106025.0 117490.0 106730.0 118835.0 ;
      RECT  106025.0 120180.0 106730.0 118835.0 ;
      RECT  106025.0 120180.0 106730.0 121525.0 ;
      RECT  106025.0 122870.0 106730.0 121525.0 ;
      RECT  106025.0 122870.0 106730.0 124215.0 ;
      RECT  106025.0 125560.0 106730.0 124215.0 ;
      RECT  106025.0 125560.0 106730.0 126905.0 ;
      RECT  106025.0 128250.0 106730.0 126905.0 ;
      RECT  106025.0 128250.0 106730.0 129595.0 ;
      RECT  106025.0 130940.0 106730.0 129595.0 ;
      RECT  106025.0 130940.0 106730.0 132285.0 ;
      RECT  106025.0 133630.0 106730.0 132285.0 ;
      RECT  106025.0 133630.0 106730.0 134975.0 ;
      RECT  106025.0 136320.0 106730.0 134975.0 ;
      RECT  106025.0 136320.0 106730.0 137665.0 ;
      RECT  106025.0 139010.0 106730.0 137665.0 ;
      RECT  106025.0 139010.0 106730.0 140355.0 ;
      RECT  106025.0 141700.0 106730.0 140355.0 ;
      RECT  106025.0 141700.0 106730.0 143045.0 ;
      RECT  106025.0 144390.0 106730.0 143045.0 ;
      RECT  106025.0 144390.0 106730.0 145735.0 ;
      RECT  106025.0 147080.0 106730.0 145735.0 ;
      RECT  106025.0 147080.0 106730.0 148425.0 ;
      RECT  106025.0 149770.0 106730.0 148425.0 ;
      RECT  106025.0 149770.0 106730.0 151115.0 ;
      RECT  106025.0 152460.0 106730.0 151115.0 ;
      RECT  106025.0 152460.0 106730.0 153805.0 ;
      RECT  106025.0 155150.0 106730.0 153805.0 ;
      RECT  106025.0 155150.0 106730.0 156495.0 ;
      RECT  106025.0 157840.0 106730.0 156495.0 ;
      RECT  106025.0 157840.0 106730.0 159185.0 ;
      RECT  106025.0 160530.0 106730.0 159185.0 ;
      RECT  106025.0 160530.0 106730.0 161875.0 ;
      RECT  106025.0 163220.0 106730.0 161875.0 ;
      RECT  106025.0 163220.0 106730.0 164565.0 ;
      RECT  106025.0 165910.0 106730.0 164565.0 ;
      RECT  106025.0 165910.0 106730.0 167255.0 ;
      RECT  106025.0 168600.0 106730.0 167255.0 ;
      RECT  106025.0 168600.0 106730.0 169945.0 ;
      RECT  106025.0 171290.0 106730.0 169945.0 ;
      RECT  106025.0 171290.0 106730.0 172635.0 ;
      RECT  106025.0 173980.0 106730.0 172635.0 ;
      RECT  106025.0 173980.0 106730.0 175325.0 ;
      RECT  106025.0 176670.0 106730.0 175325.0 ;
      RECT  106025.0 176670.0 106730.0 178015.0 ;
      RECT  106025.0 179360.0 106730.0 178015.0 ;
      RECT  106025.0 179360.0 106730.0 180705.0 ;
      RECT  106025.0 182050.0 106730.0 180705.0 ;
      RECT  106025.0 182050.0 106730.0 183395.0 ;
      RECT  106025.0 184740.0 106730.0 183395.0 ;
      RECT  106025.0 184740.0 106730.0 186085.0 ;
      RECT  106025.0 187430.0 106730.0 186085.0 ;
      RECT  106025.0 187430.0 106730.0 188775.0 ;
      RECT  106025.0 190120.0 106730.0 188775.0 ;
      RECT  106025.0 190120.0 106730.0 191465.0 ;
      RECT  106025.0 192810.0 106730.0 191465.0 ;
      RECT  106025.0 192810.0 106730.0 194155.0 ;
      RECT  106025.0 195500.0 106730.0 194155.0 ;
      RECT  106025.0 195500.0 106730.0 196845.0 ;
      RECT  106025.0 198190.0 106730.0 196845.0 ;
      RECT  106025.0 198190.0 106730.0 199535.0 ;
      RECT  106025.0 200880.0 106730.0 199535.0 ;
      RECT  106025.0 200880.0 106730.0 202225.0 ;
      RECT  106025.0 203570.0 106730.0 202225.0 ;
      RECT  106025.0 203570.0 106730.0 204915.0 ;
      RECT  106025.0 206260.0 106730.0 204915.0 ;
      RECT  106730.0 34100.0 107435.0 35445.0 ;
      RECT  106730.0 36790.0 107435.0 35445.0 ;
      RECT  106730.0 36790.0 107435.0 38135.0 ;
      RECT  106730.0 39480.0 107435.0 38135.0 ;
      RECT  106730.0 39480.0 107435.0 40825.0 ;
      RECT  106730.0 42170.0 107435.0 40825.0 ;
      RECT  106730.0 42170.0 107435.0 43515.0 ;
      RECT  106730.0 44860.0 107435.0 43515.0 ;
      RECT  106730.0 44860.0 107435.0 46205.0 ;
      RECT  106730.0 47550.0 107435.0 46205.0 ;
      RECT  106730.0 47550.0 107435.0 48895.0 ;
      RECT  106730.0 50240.0 107435.0 48895.0 ;
      RECT  106730.0 50240.0 107435.0 51585.0 ;
      RECT  106730.0 52930.0 107435.0 51585.0 ;
      RECT  106730.0 52930.0 107435.0 54275.0 ;
      RECT  106730.0 55620.0 107435.0 54275.0 ;
      RECT  106730.0 55620.0 107435.0 56965.0 ;
      RECT  106730.0 58310.0 107435.0 56965.0 ;
      RECT  106730.0 58310.0 107435.0 59655.0 ;
      RECT  106730.0 61000.0 107435.0 59655.0 ;
      RECT  106730.0 61000.0 107435.0 62345.0 ;
      RECT  106730.0 63690.0 107435.0 62345.0 ;
      RECT  106730.0 63690.0 107435.0 65035.0 ;
      RECT  106730.0 66380.0 107435.0 65035.0 ;
      RECT  106730.0 66380.0 107435.0 67725.0 ;
      RECT  106730.0 69070.0 107435.0 67725.0 ;
      RECT  106730.0 69070.0 107435.0 70415.0 ;
      RECT  106730.0 71760.0 107435.0 70415.0 ;
      RECT  106730.0 71760.0 107435.0 73105.0 ;
      RECT  106730.0 74450.0 107435.0 73105.0 ;
      RECT  106730.0 74450.0 107435.0 75795.0 ;
      RECT  106730.0 77140.0 107435.0 75795.0 ;
      RECT  106730.0 77140.0 107435.0 78485.0 ;
      RECT  106730.0 79830.0 107435.0 78485.0 ;
      RECT  106730.0 79830.0 107435.0 81175.0 ;
      RECT  106730.0 82520.0 107435.0 81175.0 ;
      RECT  106730.0 82520.0 107435.0 83865.0 ;
      RECT  106730.0 85210.0 107435.0 83865.0 ;
      RECT  106730.0 85210.0 107435.0 86555.0 ;
      RECT  106730.0 87900.0 107435.0 86555.0 ;
      RECT  106730.0 87900.0 107435.0 89245.0 ;
      RECT  106730.0 90590.0 107435.0 89245.0 ;
      RECT  106730.0 90590.0 107435.0 91935.0 ;
      RECT  106730.0 93280.0 107435.0 91935.0 ;
      RECT  106730.0 93280.0 107435.0 94625.0 ;
      RECT  106730.0 95970.0 107435.0 94625.0 ;
      RECT  106730.0 95970.0 107435.0 97315.0 ;
      RECT  106730.0 98660.0 107435.0 97315.0 ;
      RECT  106730.0 98660.0 107435.0 100005.0 ;
      RECT  106730.0 101350.0 107435.0 100005.0 ;
      RECT  106730.0 101350.0 107435.0 102695.0 ;
      RECT  106730.0 104040.0 107435.0 102695.0 ;
      RECT  106730.0 104040.0 107435.0 105385.0 ;
      RECT  106730.0 106730.0 107435.0 105385.0 ;
      RECT  106730.0 106730.0 107435.0 108075.0 ;
      RECT  106730.0 109420.0 107435.0 108075.0 ;
      RECT  106730.0 109420.0 107435.0 110765.0 ;
      RECT  106730.0 112110.0 107435.0 110765.0 ;
      RECT  106730.0 112110.0 107435.0 113455.0 ;
      RECT  106730.0 114800.0 107435.0 113455.0 ;
      RECT  106730.0 114800.0 107435.0 116145.0 ;
      RECT  106730.0 117490.0 107435.0 116145.0 ;
      RECT  106730.0 117490.0 107435.0 118835.0 ;
      RECT  106730.0 120180.0 107435.0 118835.0 ;
      RECT  106730.0 120180.0 107435.0 121525.0 ;
      RECT  106730.0 122870.0 107435.0 121525.0 ;
      RECT  106730.0 122870.0 107435.0 124215.0 ;
      RECT  106730.0 125560.0 107435.0 124215.0 ;
      RECT  106730.0 125560.0 107435.0 126905.0 ;
      RECT  106730.0 128250.0 107435.0 126905.0 ;
      RECT  106730.0 128250.0 107435.0 129595.0 ;
      RECT  106730.0 130940.0 107435.0 129595.0 ;
      RECT  106730.0 130940.0 107435.0 132285.0 ;
      RECT  106730.0 133630.0 107435.0 132285.0 ;
      RECT  106730.0 133630.0 107435.0 134975.0 ;
      RECT  106730.0 136320.0 107435.0 134975.0 ;
      RECT  106730.0 136320.0 107435.0 137665.0 ;
      RECT  106730.0 139010.0 107435.0 137665.0 ;
      RECT  106730.0 139010.0 107435.0 140355.0 ;
      RECT  106730.0 141700.0 107435.0 140355.0 ;
      RECT  106730.0 141700.0 107435.0 143045.0 ;
      RECT  106730.0 144390.0 107435.0 143045.0 ;
      RECT  106730.0 144390.0 107435.0 145735.0 ;
      RECT  106730.0 147080.0 107435.0 145735.0 ;
      RECT  106730.0 147080.0 107435.0 148425.0 ;
      RECT  106730.0 149770.0 107435.0 148425.0 ;
      RECT  106730.0 149770.0 107435.0 151115.0 ;
      RECT  106730.0 152460.0 107435.0 151115.0 ;
      RECT  106730.0 152460.0 107435.0 153805.0 ;
      RECT  106730.0 155150.0 107435.0 153805.0 ;
      RECT  106730.0 155150.0 107435.0 156495.0 ;
      RECT  106730.0 157840.0 107435.0 156495.0 ;
      RECT  106730.0 157840.0 107435.0 159185.0 ;
      RECT  106730.0 160530.0 107435.0 159185.0 ;
      RECT  106730.0 160530.0 107435.0 161875.0 ;
      RECT  106730.0 163220.0 107435.0 161875.0 ;
      RECT  106730.0 163220.0 107435.0 164565.0 ;
      RECT  106730.0 165910.0 107435.0 164565.0 ;
      RECT  106730.0 165910.0 107435.0 167255.0 ;
      RECT  106730.0 168600.0 107435.0 167255.0 ;
      RECT  106730.0 168600.0 107435.0 169945.0 ;
      RECT  106730.0 171290.0 107435.0 169945.0 ;
      RECT  106730.0 171290.0 107435.0 172635.0 ;
      RECT  106730.0 173980.0 107435.0 172635.0 ;
      RECT  106730.0 173980.0 107435.0 175325.0 ;
      RECT  106730.0 176670.0 107435.0 175325.0 ;
      RECT  106730.0 176670.0 107435.0 178015.0 ;
      RECT  106730.0 179360.0 107435.0 178015.0 ;
      RECT  106730.0 179360.0 107435.0 180705.0 ;
      RECT  106730.0 182050.0 107435.0 180705.0 ;
      RECT  106730.0 182050.0 107435.0 183395.0 ;
      RECT  106730.0 184740.0 107435.0 183395.0 ;
      RECT  106730.0 184740.0 107435.0 186085.0 ;
      RECT  106730.0 187430.0 107435.0 186085.0 ;
      RECT  106730.0 187430.0 107435.0 188775.0 ;
      RECT  106730.0 190120.0 107435.0 188775.0 ;
      RECT  106730.0 190120.0 107435.0 191465.0 ;
      RECT  106730.0 192810.0 107435.0 191465.0 ;
      RECT  106730.0 192810.0 107435.0 194155.0 ;
      RECT  106730.0 195500.0 107435.0 194155.0 ;
      RECT  106730.0 195500.0 107435.0 196845.0 ;
      RECT  106730.0 198190.0 107435.0 196845.0 ;
      RECT  106730.0 198190.0 107435.0 199535.0 ;
      RECT  106730.0 200880.0 107435.0 199535.0 ;
      RECT  106730.0 200880.0 107435.0 202225.0 ;
      RECT  106730.0 203570.0 107435.0 202225.0 ;
      RECT  106730.0 203570.0 107435.0 204915.0 ;
      RECT  106730.0 206260.0 107435.0 204915.0 ;
      RECT  17105.0 34207.5 107525.0 34272.5 ;
      RECT  17105.0 36617.5 107525.0 36682.5 ;
      RECT  17105.0 36897.5 107525.0 36962.5 ;
      RECT  17105.0 39307.5 107525.0 39372.5 ;
      RECT  17105.0 39587.5 107525.0 39652.5 ;
      RECT  17105.0 41997.5 107525.0 42062.5 ;
      RECT  17105.0 42277.5 107525.0 42342.5 ;
      RECT  17105.0 44687.5 107525.0 44752.5 ;
      RECT  17105.0 44967.5 107525.0 45032.5 ;
      RECT  17105.0 47377.5 107525.0 47442.5 ;
      RECT  17105.0 47657.5 107525.0 47722.5 ;
      RECT  17105.0 50067.5 107525.0 50132.5 ;
      RECT  17105.0 50347.5 107525.0 50412.5 ;
      RECT  17105.0 52757.5 107525.0 52822.5 ;
      RECT  17105.0 53037.5 107525.0 53102.5 ;
      RECT  17105.0 55447.5 107525.0 55512.5 ;
      RECT  17105.0 55727.5 107525.0 55792.5 ;
      RECT  17105.0 58137.5 107525.0 58202.5 ;
      RECT  17105.0 58417.5 107525.0 58482.5 ;
      RECT  17105.0 60827.5 107525.0 60892.5 ;
      RECT  17105.0 61107.5 107525.0 61172.5 ;
      RECT  17105.0 63517.5 107525.0 63582.5 ;
      RECT  17105.0 63797.5 107525.0 63862.5 ;
      RECT  17105.0 66207.5 107525.0 66272.5 ;
      RECT  17105.0 66487.5 107525.0 66552.5 ;
      RECT  17105.0 68897.5 107525.0 68962.5 ;
      RECT  17105.0 69177.5 107525.0 69242.5 ;
      RECT  17105.0 71587.5 107525.0 71652.5 ;
      RECT  17105.0 71867.5 107525.0 71932.5 ;
      RECT  17105.0 74277.5 107525.0 74342.5 ;
      RECT  17105.0 74557.5 107525.0 74622.5 ;
      RECT  17105.0 76967.5 107525.0 77032.5 ;
      RECT  17105.0 77247.5 107525.0 77312.5 ;
      RECT  17105.0 79657.5 107525.0 79722.5 ;
      RECT  17105.0 79937.5 107525.0 80002.5 ;
      RECT  17105.0 82347.5 107525.0 82412.5 ;
      RECT  17105.0 82627.5 107525.0 82692.5 ;
      RECT  17105.0 85037.5 107525.0 85102.5 ;
      RECT  17105.0 85317.5 107525.0 85382.5 ;
      RECT  17105.0 87727.5 107525.0 87792.5 ;
      RECT  17105.0 88007.5 107525.0 88072.5 ;
      RECT  17105.0 90417.5 107525.0 90482.5 ;
      RECT  17105.0 90697.5 107525.0 90762.5 ;
      RECT  17105.0 93107.5 107525.0 93172.5 ;
      RECT  17105.0 93387.5 107525.0 93452.5 ;
      RECT  17105.0 95797.5 107525.0 95862.5 ;
      RECT  17105.0 96077.5 107525.0 96142.5 ;
      RECT  17105.0 98487.5 107525.0 98552.5 ;
      RECT  17105.0 98767.5 107525.0 98832.5 ;
      RECT  17105.0 101177.5 107525.0 101242.5 ;
      RECT  17105.0 101457.5 107525.0 101522.5 ;
      RECT  17105.0 103867.5 107525.0 103932.5 ;
      RECT  17105.0 104147.5 107525.0 104212.5 ;
      RECT  17105.0 106557.5 107525.0 106622.5 ;
      RECT  17105.0 106837.5 107525.0 106902.5 ;
      RECT  17105.0 109247.5 107525.0 109312.5 ;
      RECT  17105.0 109527.5 107525.0 109592.5 ;
      RECT  17105.0 111937.5 107525.0 112002.5 ;
      RECT  17105.0 112217.5 107525.0 112282.5 ;
      RECT  17105.0 114627.5 107525.0 114692.5 ;
      RECT  17105.0 114907.5 107525.0 114972.5 ;
      RECT  17105.0 117317.5 107525.0 117382.5 ;
      RECT  17105.0 117597.5 107525.0 117662.5 ;
      RECT  17105.0 120007.5 107525.0 120072.5 ;
      RECT  17105.0 120287.5 107525.0 120352.5 ;
      RECT  17105.0 122697.5 107525.0 122762.5 ;
      RECT  17105.0 122977.5 107525.0 123042.5 ;
      RECT  17105.0 125387.5 107525.0 125452.5 ;
      RECT  17105.0 125667.5 107525.0 125732.5 ;
      RECT  17105.0 128077.5 107525.0 128142.5 ;
      RECT  17105.0 128357.5 107525.0 128422.5 ;
      RECT  17105.0 130767.5 107525.0 130832.5 ;
      RECT  17105.0 131047.5 107525.0 131112.5 ;
      RECT  17105.0 133457.5 107525.0 133522.5 ;
      RECT  17105.0 133737.5 107525.0 133802.5 ;
      RECT  17105.0 136147.5 107525.0 136212.5 ;
      RECT  17105.0 136427.5 107525.0 136492.5 ;
      RECT  17105.0 138837.5 107525.0 138902.5 ;
      RECT  17105.0 139117.5 107525.0 139182.5 ;
      RECT  17105.0 141527.5 107525.0 141592.5 ;
      RECT  17105.0 141807.5 107525.0 141872.5 ;
      RECT  17105.0 144217.5 107525.0 144282.5 ;
      RECT  17105.0 144497.5 107525.0 144562.5 ;
      RECT  17105.0 146907.5 107525.0 146972.5 ;
      RECT  17105.0 147187.5 107525.0 147252.5 ;
      RECT  17105.0 149597.5 107525.0 149662.5 ;
      RECT  17105.0 149877.5 107525.0 149942.5 ;
      RECT  17105.0 152287.5 107525.0 152352.5 ;
      RECT  17105.0 152567.5 107525.0 152632.5 ;
      RECT  17105.0 154977.5 107525.0 155042.5 ;
      RECT  17105.0 155257.5 107525.0 155322.5 ;
      RECT  17105.0 157667.5 107525.0 157732.5 ;
      RECT  17105.0 157947.5 107525.0 158012.5 ;
      RECT  17105.0 160357.5 107525.0 160422.5 ;
      RECT  17105.0 160637.5 107525.0 160702.5 ;
      RECT  17105.0 163047.5 107525.0 163112.5 ;
      RECT  17105.0 163327.5 107525.0 163392.5 ;
      RECT  17105.0 165737.5 107525.0 165802.5 ;
      RECT  17105.0 166017.5 107525.0 166082.5 ;
      RECT  17105.0 168427.5 107525.0 168492.5 ;
      RECT  17105.0 168707.5 107525.0 168772.5 ;
      RECT  17105.0 171117.5 107525.0 171182.5 ;
      RECT  17105.0 171397.5 107525.0 171462.5 ;
      RECT  17105.0 173807.5 107525.0 173872.5 ;
      RECT  17105.0 174087.5 107525.0 174152.5 ;
      RECT  17105.0 176497.5 107525.0 176562.5 ;
      RECT  17105.0 176777.5 107525.0 176842.5 ;
      RECT  17105.0 179187.5 107525.0 179252.5 ;
      RECT  17105.0 179467.5 107525.0 179532.5 ;
      RECT  17105.0 181877.5 107525.0 181942.5 ;
      RECT  17105.0 182157.5 107525.0 182222.5 ;
      RECT  17105.0 184567.5 107525.0 184632.5 ;
      RECT  17105.0 184847.5 107525.0 184912.5 ;
      RECT  17105.0 187257.5 107525.0 187322.5 ;
      RECT  17105.0 187537.5 107525.0 187602.5 ;
      RECT  17105.0 189947.5 107525.0 190012.5 ;
      RECT  17105.0 190227.5 107525.0 190292.5 ;
      RECT  17105.0 192637.5 107525.0 192702.5 ;
      RECT  17105.0 192917.5 107525.0 192982.5 ;
      RECT  17105.0 195327.5 107525.0 195392.5 ;
      RECT  17105.0 195607.5 107525.0 195672.5 ;
      RECT  17105.0 198017.5 107525.0 198082.5 ;
      RECT  17105.0 198297.5 107525.0 198362.5 ;
      RECT  17105.0 200707.5 107525.0 200772.5 ;
      RECT  17105.0 200987.5 107525.0 201052.5 ;
      RECT  17105.0 203397.5 107525.0 203462.5 ;
      RECT  17105.0 203677.5 107525.0 203742.5 ;
      RECT  17105.0 206087.5 107525.0 206152.5 ;
      RECT  17105.0 35412.5 107525.0 35477.5 ;
      RECT  17105.0 38102.5 107525.0 38167.5 ;
      RECT  17105.0 40792.5 107525.0 40857.5 ;
      RECT  17105.0 43482.5 107525.0 43547.5 ;
      RECT  17105.0 46172.5 107525.0 46237.5 ;
      RECT  17105.0 48862.5 107525.0 48927.5 ;
      RECT  17105.0 51552.5 107525.0 51617.5 ;
      RECT  17105.0 54242.5 107525.0 54307.5 ;
      RECT  17105.0 56932.5 107525.0 56997.5 ;
      RECT  17105.0 59622.5 107525.0 59687.5 ;
      RECT  17105.0 62312.5 107525.0 62377.5 ;
      RECT  17105.0 65002.5 107525.0 65067.5 ;
      RECT  17105.0 67692.5 107525.0 67757.5 ;
      RECT  17105.0 70382.5 107525.0 70447.5 ;
      RECT  17105.0 73072.5 107525.0 73137.5 ;
      RECT  17105.0 75762.5 107525.0 75827.5 ;
      RECT  17105.0 78452.5 107525.0 78517.5 ;
      RECT  17105.0 81142.5 107525.0 81207.5 ;
      RECT  17105.0 83832.5 107525.0 83897.5 ;
      RECT  17105.0 86522.5 107525.0 86587.5 ;
      RECT  17105.0 89212.5 107525.0 89277.5 ;
      RECT  17105.0 91902.5 107525.0 91967.5 ;
      RECT  17105.0 94592.5 107525.0 94657.5 ;
      RECT  17105.0 97282.5 107525.0 97347.5 ;
      RECT  17105.0 99972.5 107525.0 100037.5 ;
      RECT  17105.0 102662.5 107525.0 102727.5 ;
      RECT  17105.0 105352.5 107525.0 105417.5 ;
      RECT  17105.0 108042.5 107525.0 108107.5 ;
      RECT  17105.0 110732.5 107525.0 110797.5 ;
      RECT  17105.0 113422.5 107525.0 113487.5 ;
      RECT  17105.0 116112.5 107525.0 116177.5 ;
      RECT  17105.0 118802.5 107525.0 118867.5 ;
      RECT  17105.0 121492.5 107525.0 121557.5 ;
      RECT  17105.0 124182.5 107525.0 124247.5 ;
      RECT  17105.0 126872.5 107525.0 126937.5 ;
      RECT  17105.0 129562.5 107525.0 129627.5 ;
      RECT  17105.0 132252.5 107525.0 132317.5 ;
      RECT  17105.0 134942.5 107525.0 135007.5 ;
      RECT  17105.0 137632.5 107525.0 137697.5 ;
      RECT  17105.0 140322.5 107525.0 140387.5 ;
      RECT  17105.0 143012.5 107525.0 143077.5 ;
      RECT  17105.0 145702.5 107525.0 145767.5 ;
      RECT  17105.0 148392.5 107525.0 148457.5 ;
      RECT  17105.0 151082.5 107525.0 151147.5 ;
      RECT  17105.0 153772.5 107525.0 153837.5 ;
      RECT  17105.0 156462.5 107525.0 156527.5 ;
      RECT  17105.0 159152.5 107525.0 159217.5 ;
      RECT  17105.0 161842.5 107525.0 161907.5 ;
      RECT  17105.0 164532.5 107525.0 164597.5 ;
      RECT  17105.0 167222.5 107525.0 167287.5 ;
      RECT  17105.0 169912.5 107525.0 169977.5 ;
      RECT  17105.0 172602.5 107525.0 172667.5 ;
      RECT  17105.0 175292.5 107525.0 175357.5 ;
      RECT  17105.0 177982.5 107525.0 178047.5 ;
      RECT  17105.0 180672.5 107525.0 180737.5 ;
      RECT  17105.0 183362.5 107525.0 183427.5 ;
      RECT  17105.0 186052.5 107525.0 186117.5 ;
      RECT  17105.0 188742.5 107525.0 188807.5 ;
      RECT  17105.0 191432.5 107525.0 191497.5 ;
      RECT  17105.0 194122.5 107525.0 194187.5 ;
      RECT  17105.0 196812.5 107525.0 196877.5 ;
      RECT  17105.0 199502.5 107525.0 199567.5 ;
      RECT  17105.0 202192.5 107525.0 202257.5 ;
      RECT  17105.0 204882.5 107525.0 204947.5 ;
      RECT  17105.0 34067.5 107525.0 34132.5 ;
      RECT  17105.0 36757.5 107525.0 36822.5 ;
      RECT  17105.0 39447.5 107525.0 39512.5 ;
      RECT  17105.0 42137.5 107525.0 42202.5 ;
      RECT  17105.0 44827.5 107525.0 44892.5 ;
      RECT  17105.0 47517.5 107525.0 47582.5 ;
      RECT  17105.0 50207.5 107525.0 50272.5 ;
      RECT  17105.0 52897.5 107525.0 52962.5 ;
      RECT  17105.0 55587.5 107525.0 55652.5 ;
      RECT  17105.0 58277.5 107525.0 58342.5 ;
      RECT  17105.0 60967.5 107525.0 61032.5 ;
      RECT  17105.0 63657.5 107525.0 63722.5 ;
      RECT  17105.0 66347.5 107525.0 66412.5 ;
      RECT  17105.0 69037.5 107525.0 69102.5 ;
      RECT  17105.0 71727.5 107525.0 71792.5 ;
      RECT  17105.0 74417.5 107525.0 74482.5 ;
      RECT  17105.0 77107.5 107525.0 77172.5 ;
      RECT  17105.0 79797.5 107525.0 79862.5 ;
      RECT  17105.0 82487.5 107525.0 82552.5 ;
      RECT  17105.0 85177.5 107525.0 85242.5 ;
      RECT  17105.0 87867.5 107525.0 87932.5 ;
      RECT  17105.0 90557.5 107525.0 90622.5 ;
      RECT  17105.0 93247.5 107525.0 93312.5 ;
      RECT  17105.0 95937.5 107525.0 96002.5 ;
      RECT  17105.0 98627.5 107525.0 98692.5 ;
      RECT  17105.0 101317.5 107525.0 101382.5 ;
      RECT  17105.0 104007.5 107525.0 104072.5 ;
      RECT  17105.0 106697.5 107525.0 106762.5 ;
      RECT  17105.0 109387.5 107525.0 109452.5 ;
      RECT  17105.0 112077.5 107525.0 112142.5 ;
      RECT  17105.0 114767.5 107525.0 114832.5 ;
      RECT  17105.0 117457.5 107525.0 117522.5 ;
      RECT  17105.0 120147.5 107525.0 120212.5 ;
      RECT  17105.0 122837.5 107525.0 122902.5 ;
      RECT  17105.0 125527.5 107525.0 125592.5 ;
      RECT  17105.0 128217.5 107525.0 128282.5 ;
      RECT  17105.0 130907.5 107525.0 130972.5 ;
      RECT  17105.0 133597.5 107525.0 133662.5 ;
      RECT  17105.0 136287.5 107525.0 136352.5 ;
      RECT  17105.0 138977.5 107525.0 139042.5 ;
      RECT  17105.0 141667.5 107525.0 141732.5 ;
      RECT  17105.0 144357.5 107525.0 144422.5 ;
      RECT  17105.0 147047.5 107525.0 147112.5 ;
      RECT  17105.0 149737.5 107525.0 149802.5 ;
      RECT  17105.0 152427.5 107525.0 152492.5 ;
      RECT  17105.0 155117.5 107525.0 155182.5 ;
      RECT  17105.0 157807.5 107525.0 157872.5 ;
      RECT  17105.0 160497.5 107525.0 160562.5 ;
      RECT  17105.0 163187.5 107525.0 163252.5 ;
      RECT  17105.0 165877.5 107525.0 165942.5 ;
      RECT  17105.0 168567.5 107525.0 168632.5 ;
      RECT  17105.0 171257.5 107525.0 171322.5 ;
      RECT  17105.0 173947.5 107525.0 174012.5 ;
      RECT  17105.0 176637.5 107525.0 176702.5 ;
      RECT  17105.0 179327.5 107525.0 179392.5 ;
      RECT  17105.0 182017.5 107525.0 182082.5 ;
      RECT  17105.0 184707.5 107525.0 184772.5 ;
      RECT  17105.0 187397.5 107525.0 187462.5 ;
      RECT  17105.0 190087.5 107525.0 190152.5 ;
      RECT  17105.0 192777.5 107525.0 192842.5 ;
      RECT  17105.0 195467.5 107525.0 195532.5 ;
      RECT  17105.0 198157.5 107525.0 198222.5 ;
      RECT  17105.0 200847.5 107525.0 200912.5 ;
      RECT  17105.0 203537.5 107525.0 203602.5 ;
      RECT  17105.0 206227.5 107525.0 206292.5 ;
      RECT  17547.5 207472.5 17612.5 207987.5 ;
      RECT  17357.5 206942.5 17422.5 207077.5 ;
      RECT  17547.5 206942.5 17612.5 207077.5 ;
      RECT  17547.5 206942.5 17612.5 207077.5 ;
      RECT  17357.5 206942.5 17422.5 207077.5 ;
      RECT  17357.5 207472.5 17422.5 207607.5 ;
      RECT  17547.5 207472.5 17612.5 207607.5 ;
      RECT  17547.5 207472.5 17612.5 207607.5 ;
      RECT  17357.5 207472.5 17422.5 207607.5 ;
      RECT  17547.5 207472.5 17612.5 207607.5 ;
      RECT  17737.5 207472.5 17802.5 207607.5 ;
      RECT  17737.5 207472.5 17802.5 207607.5 ;
      RECT  17547.5 207472.5 17612.5 207607.5 ;
      RECT  17527.5 207237.5 17392.5 207302.5 ;
      RECT  17547.5 207785.0 17612.5 207920.0 ;
      RECT  17357.5 206942.5 17422.5 207077.5 ;
      RECT  17547.5 206942.5 17612.5 207077.5 ;
      RECT  17357.5 207472.5 17422.5 207607.5 ;
      RECT  17737.5 207472.5 17802.5 207607.5 ;
      RECT  17195.0 207237.5 17900.0 207302.5 ;
      RECT  17195.0 207922.5 17900.0 207987.5 ;
      RECT  18252.5 207472.5 18317.5 207987.5 ;
      RECT  18062.5 206942.5 18127.5 207077.5 ;
      RECT  18252.5 206942.5 18317.5 207077.5 ;
      RECT  18252.5 206942.5 18317.5 207077.5 ;
      RECT  18062.5 206942.5 18127.5 207077.5 ;
      RECT  18062.5 207472.5 18127.5 207607.5 ;
      RECT  18252.5 207472.5 18317.5 207607.5 ;
      RECT  18252.5 207472.5 18317.5 207607.5 ;
      RECT  18062.5 207472.5 18127.5 207607.5 ;
      RECT  18252.5 207472.5 18317.5 207607.5 ;
      RECT  18442.5 207472.5 18507.5 207607.5 ;
      RECT  18442.5 207472.5 18507.5 207607.5 ;
      RECT  18252.5 207472.5 18317.5 207607.5 ;
      RECT  18232.5 207237.5 18097.5 207302.5 ;
      RECT  18252.5 207785.0 18317.5 207920.0 ;
      RECT  18062.5 206942.5 18127.5 207077.5 ;
      RECT  18252.5 206942.5 18317.5 207077.5 ;
      RECT  18062.5 207472.5 18127.5 207607.5 ;
      RECT  18442.5 207472.5 18507.5 207607.5 ;
      RECT  17900.0 207237.5 18605.0 207302.5 ;
      RECT  17900.0 207922.5 18605.0 207987.5 ;
      RECT  18957.5 207472.5 19022.5 207987.5 ;
      RECT  18767.5 206942.5 18832.5 207077.5 ;
      RECT  18957.5 206942.5 19022.5 207077.5 ;
      RECT  18957.5 206942.5 19022.5 207077.5 ;
      RECT  18767.5 206942.5 18832.5 207077.5 ;
      RECT  18767.5 207472.5 18832.5 207607.5 ;
      RECT  18957.5 207472.5 19022.5 207607.5 ;
      RECT  18957.5 207472.5 19022.5 207607.5 ;
      RECT  18767.5 207472.5 18832.5 207607.5 ;
      RECT  18957.5 207472.5 19022.5 207607.5 ;
      RECT  19147.5 207472.5 19212.5 207607.5 ;
      RECT  19147.5 207472.5 19212.5 207607.5 ;
      RECT  18957.5 207472.5 19022.5 207607.5 ;
      RECT  18937.5 207237.5 18802.5 207302.5 ;
      RECT  18957.5 207785.0 19022.5 207920.0 ;
      RECT  18767.5 206942.5 18832.5 207077.5 ;
      RECT  18957.5 206942.5 19022.5 207077.5 ;
      RECT  18767.5 207472.5 18832.5 207607.5 ;
      RECT  19147.5 207472.5 19212.5 207607.5 ;
      RECT  18605.0 207237.5 19310.0 207302.5 ;
      RECT  18605.0 207922.5 19310.0 207987.5 ;
      RECT  19662.5 207472.5 19727.5 207987.5 ;
      RECT  19472.5 206942.5 19537.5 207077.5 ;
      RECT  19662.5 206942.5 19727.5 207077.5 ;
      RECT  19662.5 206942.5 19727.5 207077.5 ;
      RECT  19472.5 206942.5 19537.5 207077.5 ;
      RECT  19472.5 207472.5 19537.5 207607.5 ;
      RECT  19662.5 207472.5 19727.5 207607.5 ;
      RECT  19662.5 207472.5 19727.5 207607.5 ;
      RECT  19472.5 207472.5 19537.5 207607.5 ;
      RECT  19662.5 207472.5 19727.5 207607.5 ;
      RECT  19852.5 207472.5 19917.5 207607.5 ;
      RECT  19852.5 207472.5 19917.5 207607.5 ;
      RECT  19662.5 207472.5 19727.5 207607.5 ;
      RECT  19642.5 207237.5 19507.5 207302.5 ;
      RECT  19662.5 207785.0 19727.5 207920.0 ;
      RECT  19472.5 206942.5 19537.5 207077.5 ;
      RECT  19662.5 206942.5 19727.5 207077.5 ;
      RECT  19472.5 207472.5 19537.5 207607.5 ;
      RECT  19852.5 207472.5 19917.5 207607.5 ;
      RECT  19310.0 207237.5 20015.0 207302.5 ;
      RECT  19310.0 207922.5 20015.0 207987.5 ;
      RECT  20367.5 207472.5 20432.5 207987.5 ;
      RECT  20177.5 206942.5 20242.5 207077.5 ;
      RECT  20367.5 206942.5 20432.5 207077.5 ;
      RECT  20367.5 206942.5 20432.5 207077.5 ;
      RECT  20177.5 206942.5 20242.5 207077.5 ;
      RECT  20177.5 207472.5 20242.5 207607.5 ;
      RECT  20367.5 207472.5 20432.5 207607.5 ;
      RECT  20367.5 207472.5 20432.5 207607.5 ;
      RECT  20177.5 207472.5 20242.5 207607.5 ;
      RECT  20367.5 207472.5 20432.5 207607.5 ;
      RECT  20557.5 207472.5 20622.5 207607.5 ;
      RECT  20557.5 207472.5 20622.5 207607.5 ;
      RECT  20367.5 207472.5 20432.5 207607.5 ;
      RECT  20347.5 207237.5 20212.5 207302.5 ;
      RECT  20367.5 207785.0 20432.5 207920.0 ;
      RECT  20177.5 206942.5 20242.5 207077.5 ;
      RECT  20367.5 206942.5 20432.5 207077.5 ;
      RECT  20177.5 207472.5 20242.5 207607.5 ;
      RECT  20557.5 207472.5 20622.5 207607.5 ;
      RECT  20015.0 207237.5 20720.0 207302.5 ;
      RECT  20015.0 207922.5 20720.0 207987.5 ;
      RECT  21072.5 207472.5 21137.5 207987.5 ;
      RECT  20882.5 206942.5 20947.5 207077.5 ;
      RECT  21072.5 206942.5 21137.5 207077.5 ;
      RECT  21072.5 206942.5 21137.5 207077.5 ;
      RECT  20882.5 206942.5 20947.5 207077.5 ;
      RECT  20882.5 207472.5 20947.5 207607.5 ;
      RECT  21072.5 207472.5 21137.5 207607.5 ;
      RECT  21072.5 207472.5 21137.5 207607.5 ;
      RECT  20882.5 207472.5 20947.5 207607.5 ;
      RECT  21072.5 207472.5 21137.5 207607.5 ;
      RECT  21262.5 207472.5 21327.5 207607.5 ;
      RECT  21262.5 207472.5 21327.5 207607.5 ;
      RECT  21072.5 207472.5 21137.5 207607.5 ;
      RECT  21052.5 207237.5 20917.5 207302.5 ;
      RECT  21072.5 207785.0 21137.5 207920.0 ;
      RECT  20882.5 206942.5 20947.5 207077.5 ;
      RECT  21072.5 206942.5 21137.5 207077.5 ;
      RECT  20882.5 207472.5 20947.5 207607.5 ;
      RECT  21262.5 207472.5 21327.5 207607.5 ;
      RECT  20720.0 207237.5 21425.0 207302.5 ;
      RECT  20720.0 207922.5 21425.0 207987.5 ;
      RECT  21777.5 207472.5 21842.5 207987.5 ;
      RECT  21587.5 206942.5 21652.5 207077.5 ;
      RECT  21777.5 206942.5 21842.5 207077.5 ;
      RECT  21777.5 206942.5 21842.5 207077.5 ;
      RECT  21587.5 206942.5 21652.5 207077.5 ;
      RECT  21587.5 207472.5 21652.5 207607.5 ;
      RECT  21777.5 207472.5 21842.5 207607.5 ;
      RECT  21777.5 207472.5 21842.5 207607.5 ;
      RECT  21587.5 207472.5 21652.5 207607.5 ;
      RECT  21777.5 207472.5 21842.5 207607.5 ;
      RECT  21967.5 207472.5 22032.5 207607.5 ;
      RECT  21967.5 207472.5 22032.5 207607.5 ;
      RECT  21777.5 207472.5 21842.5 207607.5 ;
      RECT  21757.5 207237.5 21622.5 207302.5 ;
      RECT  21777.5 207785.0 21842.5 207920.0 ;
      RECT  21587.5 206942.5 21652.5 207077.5 ;
      RECT  21777.5 206942.5 21842.5 207077.5 ;
      RECT  21587.5 207472.5 21652.5 207607.5 ;
      RECT  21967.5 207472.5 22032.5 207607.5 ;
      RECT  21425.0 207237.5 22130.0 207302.5 ;
      RECT  21425.0 207922.5 22130.0 207987.5 ;
      RECT  22482.5 207472.5 22547.5 207987.5 ;
      RECT  22292.5 206942.5 22357.5 207077.5 ;
      RECT  22482.5 206942.5 22547.5 207077.5 ;
      RECT  22482.5 206942.5 22547.5 207077.5 ;
      RECT  22292.5 206942.5 22357.5 207077.5 ;
      RECT  22292.5 207472.5 22357.5 207607.5 ;
      RECT  22482.5 207472.5 22547.5 207607.5 ;
      RECT  22482.5 207472.5 22547.5 207607.5 ;
      RECT  22292.5 207472.5 22357.5 207607.5 ;
      RECT  22482.5 207472.5 22547.5 207607.5 ;
      RECT  22672.5 207472.5 22737.5 207607.5 ;
      RECT  22672.5 207472.5 22737.5 207607.5 ;
      RECT  22482.5 207472.5 22547.5 207607.5 ;
      RECT  22462.5 207237.5 22327.5 207302.5 ;
      RECT  22482.5 207785.0 22547.5 207920.0 ;
      RECT  22292.5 206942.5 22357.5 207077.5 ;
      RECT  22482.5 206942.5 22547.5 207077.5 ;
      RECT  22292.5 207472.5 22357.5 207607.5 ;
      RECT  22672.5 207472.5 22737.5 207607.5 ;
      RECT  22130.0 207237.5 22835.0 207302.5 ;
      RECT  22130.0 207922.5 22835.0 207987.5 ;
      RECT  23187.5 207472.5 23252.5 207987.5 ;
      RECT  22997.5 206942.5 23062.5 207077.5 ;
      RECT  23187.5 206942.5 23252.5 207077.5 ;
      RECT  23187.5 206942.5 23252.5 207077.5 ;
      RECT  22997.5 206942.5 23062.5 207077.5 ;
      RECT  22997.5 207472.5 23062.5 207607.5 ;
      RECT  23187.5 207472.5 23252.5 207607.5 ;
      RECT  23187.5 207472.5 23252.5 207607.5 ;
      RECT  22997.5 207472.5 23062.5 207607.5 ;
      RECT  23187.5 207472.5 23252.5 207607.5 ;
      RECT  23377.5 207472.5 23442.5 207607.5 ;
      RECT  23377.5 207472.5 23442.5 207607.5 ;
      RECT  23187.5 207472.5 23252.5 207607.5 ;
      RECT  23167.5 207237.5 23032.5 207302.5 ;
      RECT  23187.5 207785.0 23252.5 207920.0 ;
      RECT  22997.5 206942.5 23062.5 207077.5 ;
      RECT  23187.5 206942.5 23252.5 207077.5 ;
      RECT  22997.5 207472.5 23062.5 207607.5 ;
      RECT  23377.5 207472.5 23442.5 207607.5 ;
      RECT  22835.0 207237.5 23540.0 207302.5 ;
      RECT  22835.0 207922.5 23540.0 207987.5 ;
      RECT  23892.5 207472.5 23957.5 207987.5 ;
      RECT  23702.5 206942.5 23767.5 207077.5 ;
      RECT  23892.5 206942.5 23957.5 207077.5 ;
      RECT  23892.5 206942.5 23957.5 207077.5 ;
      RECT  23702.5 206942.5 23767.5 207077.5 ;
      RECT  23702.5 207472.5 23767.5 207607.5 ;
      RECT  23892.5 207472.5 23957.5 207607.5 ;
      RECT  23892.5 207472.5 23957.5 207607.5 ;
      RECT  23702.5 207472.5 23767.5 207607.5 ;
      RECT  23892.5 207472.5 23957.5 207607.5 ;
      RECT  24082.5 207472.5 24147.5 207607.5 ;
      RECT  24082.5 207472.5 24147.5 207607.5 ;
      RECT  23892.5 207472.5 23957.5 207607.5 ;
      RECT  23872.5 207237.5 23737.5 207302.5 ;
      RECT  23892.5 207785.0 23957.5 207920.0 ;
      RECT  23702.5 206942.5 23767.5 207077.5 ;
      RECT  23892.5 206942.5 23957.5 207077.5 ;
      RECT  23702.5 207472.5 23767.5 207607.5 ;
      RECT  24082.5 207472.5 24147.5 207607.5 ;
      RECT  23540.0 207237.5 24245.0 207302.5 ;
      RECT  23540.0 207922.5 24245.0 207987.5 ;
      RECT  24597.5 207472.5 24662.5 207987.5 ;
      RECT  24407.5 206942.5 24472.5 207077.5 ;
      RECT  24597.5 206942.5 24662.5 207077.5 ;
      RECT  24597.5 206942.5 24662.5 207077.5 ;
      RECT  24407.5 206942.5 24472.5 207077.5 ;
      RECT  24407.5 207472.5 24472.5 207607.5 ;
      RECT  24597.5 207472.5 24662.5 207607.5 ;
      RECT  24597.5 207472.5 24662.5 207607.5 ;
      RECT  24407.5 207472.5 24472.5 207607.5 ;
      RECT  24597.5 207472.5 24662.5 207607.5 ;
      RECT  24787.5 207472.5 24852.5 207607.5 ;
      RECT  24787.5 207472.5 24852.5 207607.5 ;
      RECT  24597.5 207472.5 24662.5 207607.5 ;
      RECT  24577.5 207237.5 24442.5 207302.5 ;
      RECT  24597.5 207785.0 24662.5 207920.0 ;
      RECT  24407.5 206942.5 24472.5 207077.5 ;
      RECT  24597.5 206942.5 24662.5 207077.5 ;
      RECT  24407.5 207472.5 24472.5 207607.5 ;
      RECT  24787.5 207472.5 24852.5 207607.5 ;
      RECT  24245.0 207237.5 24950.0 207302.5 ;
      RECT  24245.0 207922.5 24950.0 207987.5 ;
      RECT  25302.5 207472.5 25367.5 207987.5 ;
      RECT  25112.5 206942.5 25177.5 207077.5 ;
      RECT  25302.5 206942.5 25367.5 207077.5 ;
      RECT  25302.5 206942.5 25367.5 207077.5 ;
      RECT  25112.5 206942.5 25177.5 207077.5 ;
      RECT  25112.5 207472.5 25177.5 207607.5 ;
      RECT  25302.5 207472.5 25367.5 207607.5 ;
      RECT  25302.5 207472.5 25367.5 207607.5 ;
      RECT  25112.5 207472.5 25177.5 207607.5 ;
      RECT  25302.5 207472.5 25367.5 207607.5 ;
      RECT  25492.5 207472.5 25557.5 207607.5 ;
      RECT  25492.5 207472.5 25557.5 207607.5 ;
      RECT  25302.5 207472.5 25367.5 207607.5 ;
      RECT  25282.5 207237.5 25147.5 207302.5 ;
      RECT  25302.5 207785.0 25367.5 207920.0 ;
      RECT  25112.5 206942.5 25177.5 207077.5 ;
      RECT  25302.5 206942.5 25367.5 207077.5 ;
      RECT  25112.5 207472.5 25177.5 207607.5 ;
      RECT  25492.5 207472.5 25557.5 207607.5 ;
      RECT  24950.0 207237.5 25655.0 207302.5 ;
      RECT  24950.0 207922.5 25655.0 207987.5 ;
      RECT  26007.5 207472.5 26072.5 207987.5 ;
      RECT  25817.5 206942.5 25882.5 207077.5 ;
      RECT  26007.5 206942.5 26072.5 207077.5 ;
      RECT  26007.5 206942.5 26072.5 207077.5 ;
      RECT  25817.5 206942.5 25882.5 207077.5 ;
      RECT  25817.5 207472.5 25882.5 207607.5 ;
      RECT  26007.5 207472.5 26072.5 207607.5 ;
      RECT  26007.5 207472.5 26072.5 207607.5 ;
      RECT  25817.5 207472.5 25882.5 207607.5 ;
      RECT  26007.5 207472.5 26072.5 207607.5 ;
      RECT  26197.5 207472.5 26262.5 207607.5 ;
      RECT  26197.5 207472.5 26262.5 207607.5 ;
      RECT  26007.5 207472.5 26072.5 207607.5 ;
      RECT  25987.5 207237.5 25852.5 207302.5 ;
      RECT  26007.5 207785.0 26072.5 207920.0 ;
      RECT  25817.5 206942.5 25882.5 207077.5 ;
      RECT  26007.5 206942.5 26072.5 207077.5 ;
      RECT  25817.5 207472.5 25882.5 207607.5 ;
      RECT  26197.5 207472.5 26262.5 207607.5 ;
      RECT  25655.0 207237.5 26360.0 207302.5 ;
      RECT  25655.0 207922.5 26360.0 207987.5 ;
      RECT  26712.5 207472.5 26777.5 207987.5 ;
      RECT  26522.5 206942.5 26587.5 207077.5 ;
      RECT  26712.5 206942.5 26777.5 207077.5 ;
      RECT  26712.5 206942.5 26777.5 207077.5 ;
      RECT  26522.5 206942.5 26587.5 207077.5 ;
      RECT  26522.5 207472.5 26587.5 207607.5 ;
      RECT  26712.5 207472.5 26777.5 207607.5 ;
      RECT  26712.5 207472.5 26777.5 207607.5 ;
      RECT  26522.5 207472.5 26587.5 207607.5 ;
      RECT  26712.5 207472.5 26777.5 207607.5 ;
      RECT  26902.5 207472.5 26967.5 207607.5 ;
      RECT  26902.5 207472.5 26967.5 207607.5 ;
      RECT  26712.5 207472.5 26777.5 207607.5 ;
      RECT  26692.5 207237.5 26557.5 207302.5 ;
      RECT  26712.5 207785.0 26777.5 207920.0 ;
      RECT  26522.5 206942.5 26587.5 207077.5 ;
      RECT  26712.5 206942.5 26777.5 207077.5 ;
      RECT  26522.5 207472.5 26587.5 207607.5 ;
      RECT  26902.5 207472.5 26967.5 207607.5 ;
      RECT  26360.0 207237.5 27065.0 207302.5 ;
      RECT  26360.0 207922.5 27065.0 207987.5 ;
      RECT  27417.5 207472.5 27482.5 207987.5 ;
      RECT  27227.5 206942.5 27292.5 207077.5 ;
      RECT  27417.5 206942.5 27482.5 207077.5 ;
      RECT  27417.5 206942.5 27482.5 207077.5 ;
      RECT  27227.5 206942.5 27292.5 207077.5 ;
      RECT  27227.5 207472.5 27292.5 207607.5 ;
      RECT  27417.5 207472.5 27482.5 207607.5 ;
      RECT  27417.5 207472.5 27482.5 207607.5 ;
      RECT  27227.5 207472.5 27292.5 207607.5 ;
      RECT  27417.5 207472.5 27482.5 207607.5 ;
      RECT  27607.5 207472.5 27672.5 207607.5 ;
      RECT  27607.5 207472.5 27672.5 207607.5 ;
      RECT  27417.5 207472.5 27482.5 207607.5 ;
      RECT  27397.5 207237.5 27262.5 207302.5 ;
      RECT  27417.5 207785.0 27482.5 207920.0 ;
      RECT  27227.5 206942.5 27292.5 207077.5 ;
      RECT  27417.5 206942.5 27482.5 207077.5 ;
      RECT  27227.5 207472.5 27292.5 207607.5 ;
      RECT  27607.5 207472.5 27672.5 207607.5 ;
      RECT  27065.0 207237.5 27770.0 207302.5 ;
      RECT  27065.0 207922.5 27770.0 207987.5 ;
      RECT  28122.5 207472.5 28187.5 207987.5 ;
      RECT  27932.5 206942.5 27997.5 207077.5 ;
      RECT  28122.5 206942.5 28187.5 207077.5 ;
      RECT  28122.5 206942.5 28187.5 207077.5 ;
      RECT  27932.5 206942.5 27997.5 207077.5 ;
      RECT  27932.5 207472.5 27997.5 207607.5 ;
      RECT  28122.5 207472.5 28187.5 207607.5 ;
      RECT  28122.5 207472.5 28187.5 207607.5 ;
      RECT  27932.5 207472.5 27997.5 207607.5 ;
      RECT  28122.5 207472.5 28187.5 207607.5 ;
      RECT  28312.5 207472.5 28377.5 207607.5 ;
      RECT  28312.5 207472.5 28377.5 207607.5 ;
      RECT  28122.5 207472.5 28187.5 207607.5 ;
      RECT  28102.5 207237.5 27967.5 207302.5 ;
      RECT  28122.5 207785.0 28187.5 207920.0 ;
      RECT  27932.5 206942.5 27997.5 207077.5 ;
      RECT  28122.5 206942.5 28187.5 207077.5 ;
      RECT  27932.5 207472.5 27997.5 207607.5 ;
      RECT  28312.5 207472.5 28377.5 207607.5 ;
      RECT  27770.0 207237.5 28475.0 207302.5 ;
      RECT  27770.0 207922.5 28475.0 207987.5 ;
      RECT  28827.5 207472.5 28892.5 207987.5 ;
      RECT  28637.5 206942.5 28702.5 207077.5 ;
      RECT  28827.5 206942.5 28892.5 207077.5 ;
      RECT  28827.5 206942.5 28892.5 207077.5 ;
      RECT  28637.5 206942.5 28702.5 207077.5 ;
      RECT  28637.5 207472.5 28702.5 207607.5 ;
      RECT  28827.5 207472.5 28892.5 207607.5 ;
      RECT  28827.5 207472.5 28892.5 207607.5 ;
      RECT  28637.5 207472.5 28702.5 207607.5 ;
      RECT  28827.5 207472.5 28892.5 207607.5 ;
      RECT  29017.5 207472.5 29082.5 207607.5 ;
      RECT  29017.5 207472.5 29082.5 207607.5 ;
      RECT  28827.5 207472.5 28892.5 207607.5 ;
      RECT  28807.5 207237.5 28672.5 207302.5 ;
      RECT  28827.5 207785.0 28892.5 207920.0 ;
      RECT  28637.5 206942.5 28702.5 207077.5 ;
      RECT  28827.5 206942.5 28892.5 207077.5 ;
      RECT  28637.5 207472.5 28702.5 207607.5 ;
      RECT  29017.5 207472.5 29082.5 207607.5 ;
      RECT  28475.0 207237.5 29180.0 207302.5 ;
      RECT  28475.0 207922.5 29180.0 207987.5 ;
      RECT  29532.5 207472.5 29597.5 207987.5 ;
      RECT  29342.5 206942.5 29407.5 207077.5 ;
      RECT  29532.5 206942.5 29597.5 207077.5 ;
      RECT  29532.5 206942.5 29597.5 207077.5 ;
      RECT  29342.5 206942.5 29407.5 207077.5 ;
      RECT  29342.5 207472.5 29407.5 207607.5 ;
      RECT  29532.5 207472.5 29597.5 207607.5 ;
      RECT  29532.5 207472.5 29597.5 207607.5 ;
      RECT  29342.5 207472.5 29407.5 207607.5 ;
      RECT  29532.5 207472.5 29597.5 207607.5 ;
      RECT  29722.5 207472.5 29787.5 207607.5 ;
      RECT  29722.5 207472.5 29787.5 207607.5 ;
      RECT  29532.5 207472.5 29597.5 207607.5 ;
      RECT  29512.5 207237.5 29377.5 207302.5 ;
      RECT  29532.5 207785.0 29597.5 207920.0 ;
      RECT  29342.5 206942.5 29407.5 207077.5 ;
      RECT  29532.5 206942.5 29597.5 207077.5 ;
      RECT  29342.5 207472.5 29407.5 207607.5 ;
      RECT  29722.5 207472.5 29787.5 207607.5 ;
      RECT  29180.0 207237.5 29885.0 207302.5 ;
      RECT  29180.0 207922.5 29885.0 207987.5 ;
      RECT  30237.5 207472.5 30302.5 207987.5 ;
      RECT  30047.5 206942.5 30112.5 207077.5 ;
      RECT  30237.5 206942.5 30302.5 207077.5 ;
      RECT  30237.5 206942.5 30302.5 207077.5 ;
      RECT  30047.5 206942.5 30112.5 207077.5 ;
      RECT  30047.5 207472.5 30112.5 207607.5 ;
      RECT  30237.5 207472.5 30302.5 207607.5 ;
      RECT  30237.5 207472.5 30302.5 207607.5 ;
      RECT  30047.5 207472.5 30112.5 207607.5 ;
      RECT  30237.5 207472.5 30302.5 207607.5 ;
      RECT  30427.5 207472.5 30492.5 207607.5 ;
      RECT  30427.5 207472.5 30492.5 207607.5 ;
      RECT  30237.5 207472.5 30302.5 207607.5 ;
      RECT  30217.5 207237.5 30082.5 207302.5 ;
      RECT  30237.5 207785.0 30302.5 207920.0 ;
      RECT  30047.5 206942.5 30112.5 207077.5 ;
      RECT  30237.5 206942.5 30302.5 207077.5 ;
      RECT  30047.5 207472.5 30112.5 207607.5 ;
      RECT  30427.5 207472.5 30492.5 207607.5 ;
      RECT  29885.0 207237.5 30590.0 207302.5 ;
      RECT  29885.0 207922.5 30590.0 207987.5 ;
      RECT  30942.5 207472.5 31007.5 207987.5 ;
      RECT  30752.5 206942.5 30817.5 207077.5 ;
      RECT  30942.5 206942.5 31007.5 207077.5 ;
      RECT  30942.5 206942.5 31007.5 207077.5 ;
      RECT  30752.5 206942.5 30817.5 207077.5 ;
      RECT  30752.5 207472.5 30817.5 207607.5 ;
      RECT  30942.5 207472.5 31007.5 207607.5 ;
      RECT  30942.5 207472.5 31007.5 207607.5 ;
      RECT  30752.5 207472.5 30817.5 207607.5 ;
      RECT  30942.5 207472.5 31007.5 207607.5 ;
      RECT  31132.5 207472.5 31197.5 207607.5 ;
      RECT  31132.5 207472.5 31197.5 207607.5 ;
      RECT  30942.5 207472.5 31007.5 207607.5 ;
      RECT  30922.5 207237.5 30787.5 207302.5 ;
      RECT  30942.5 207785.0 31007.5 207920.0 ;
      RECT  30752.5 206942.5 30817.5 207077.5 ;
      RECT  30942.5 206942.5 31007.5 207077.5 ;
      RECT  30752.5 207472.5 30817.5 207607.5 ;
      RECT  31132.5 207472.5 31197.5 207607.5 ;
      RECT  30590.0 207237.5 31295.0 207302.5 ;
      RECT  30590.0 207922.5 31295.0 207987.5 ;
      RECT  31647.5 207472.5 31712.5 207987.5 ;
      RECT  31457.5 206942.5 31522.5 207077.5 ;
      RECT  31647.5 206942.5 31712.5 207077.5 ;
      RECT  31647.5 206942.5 31712.5 207077.5 ;
      RECT  31457.5 206942.5 31522.5 207077.5 ;
      RECT  31457.5 207472.5 31522.5 207607.5 ;
      RECT  31647.5 207472.5 31712.5 207607.5 ;
      RECT  31647.5 207472.5 31712.5 207607.5 ;
      RECT  31457.5 207472.5 31522.5 207607.5 ;
      RECT  31647.5 207472.5 31712.5 207607.5 ;
      RECT  31837.5 207472.5 31902.5 207607.5 ;
      RECT  31837.5 207472.5 31902.5 207607.5 ;
      RECT  31647.5 207472.5 31712.5 207607.5 ;
      RECT  31627.5 207237.5 31492.5 207302.5 ;
      RECT  31647.5 207785.0 31712.5 207920.0 ;
      RECT  31457.5 206942.5 31522.5 207077.5 ;
      RECT  31647.5 206942.5 31712.5 207077.5 ;
      RECT  31457.5 207472.5 31522.5 207607.5 ;
      RECT  31837.5 207472.5 31902.5 207607.5 ;
      RECT  31295.0 207237.5 32000.0 207302.5 ;
      RECT  31295.0 207922.5 32000.0 207987.5 ;
      RECT  32352.5 207472.5 32417.5 207987.5 ;
      RECT  32162.5 206942.5 32227.5 207077.5 ;
      RECT  32352.5 206942.5 32417.5 207077.5 ;
      RECT  32352.5 206942.5 32417.5 207077.5 ;
      RECT  32162.5 206942.5 32227.5 207077.5 ;
      RECT  32162.5 207472.5 32227.5 207607.5 ;
      RECT  32352.5 207472.5 32417.5 207607.5 ;
      RECT  32352.5 207472.5 32417.5 207607.5 ;
      RECT  32162.5 207472.5 32227.5 207607.5 ;
      RECT  32352.5 207472.5 32417.5 207607.5 ;
      RECT  32542.5 207472.5 32607.5 207607.5 ;
      RECT  32542.5 207472.5 32607.5 207607.5 ;
      RECT  32352.5 207472.5 32417.5 207607.5 ;
      RECT  32332.5 207237.5 32197.5 207302.5 ;
      RECT  32352.5 207785.0 32417.5 207920.0 ;
      RECT  32162.5 206942.5 32227.5 207077.5 ;
      RECT  32352.5 206942.5 32417.5 207077.5 ;
      RECT  32162.5 207472.5 32227.5 207607.5 ;
      RECT  32542.5 207472.5 32607.5 207607.5 ;
      RECT  32000.0 207237.5 32705.0 207302.5 ;
      RECT  32000.0 207922.5 32705.0 207987.5 ;
      RECT  33057.5 207472.5 33122.5 207987.5 ;
      RECT  32867.5 206942.5 32932.5 207077.5 ;
      RECT  33057.5 206942.5 33122.5 207077.5 ;
      RECT  33057.5 206942.5 33122.5 207077.5 ;
      RECT  32867.5 206942.5 32932.5 207077.5 ;
      RECT  32867.5 207472.5 32932.5 207607.5 ;
      RECT  33057.5 207472.5 33122.5 207607.5 ;
      RECT  33057.5 207472.5 33122.5 207607.5 ;
      RECT  32867.5 207472.5 32932.5 207607.5 ;
      RECT  33057.5 207472.5 33122.5 207607.5 ;
      RECT  33247.5 207472.5 33312.5 207607.5 ;
      RECT  33247.5 207472.5 33312.5 207607.5 ;
      RECT  33057.5 207472.5 33122.5 207607.5 ;
      RECT  33037.5 207237.5 32902.5 207302.5 ;
      RECT  33057.5 207785.0 33122.5 207920.0 ;
      RECT  32867.5 206942.5 32932.5 207077.5 ;
      RECT  33057.5 206942.5 33122.5 207077.5 ;
      RECT  32867.5 207472.5 32932.5 207607.5 ;
      RECT  33247.5 207472.5 33312.5 207607.5 ;
      RECT  32705.0 207237.5 33410.0 207302.5 ;
      RECT  32705.0 207922.5 33410.0 207987.5 ;
      RECT  33762.5 207472.5 33827.5 207987.5 ;
      RECT  33572.5 206942.5 33637.5 207077.5 ;
      RECT  33762.5 206942.5 33827.5 207077.5 ;
      RECT  33762.5 206942.5 33827.5 207077.5 ;
      RECT  33572.5 206942.5 33637.5 207077.5 ;
      RECT  33572.5 207472.5 33637.5 207607.5 ;
      RECT  33762.5 207472.5 33827.5 207607.5 ;
      RECT  33762.5 207472.5 33827.5 207607.5 ;
      RECT  33572.5 207472.5 33637.5 207607.5 ;
      RECT  33762.5 207472.5 33827.5 207607.5 ;
      RECT  33952.5 207472.5 34017.5 207607.5 ;
      RECT  33952.5 207472.5 34017.5 207607.5 ;
      RECT  33762.5 207472.5 33827.5 207607.5 ;
      RECT  33742.5 207237.5 33607.5 207302.5 ;
      RECT  33762.5 207785.0 33827.5 207920.0 ;
      RECT  33572.5 206942.5 33637.5 207077.5 ;
      RECT  33762.5 206942.5 33827.5 207077.5 ;
      RECT  33572.5 207472.5 33637.5 207607.5 ;
      RECT  33952.5 207472.5 34017.5 207607.5 ;
      RECT  33410.0 207237.5 34115.0 207302.5 ;
      RECT  33410.0 207922.5 34115.0 207987.5 ;
      RECT  34467.5 207472.5 34532.5 207987.5 ;
      RECT  34277.5 206942.5 34342.5 207077.5 ;
      RECT  34467.5 206942.5 34532.5 207077.5 ;
      RECT  34467.5 206942.5 34532.5 207077.5 ;
      RECT  34277.5 206942.5 34342.5 207077.5 ;
      RECT  34277.5 207472.5 34342.5 207607.5 ;
      RECT  34467.5 207472.5 34532.5 207607.5 ;
      RECT  34467.5 207472.5 34532.5 207607.5 ;
      RECT  34277.5 207472.5 34342.5 207607.5 ;
      RECT  34467.5 207472.5 34532.5 207607.5 ;
      RECT  34657.5 207472.5 34722.5 207607.5 ;
      RECT  34657.5 207472.5 34722.5 207607.5 ;
      RECT  34467.5 207472.5 34532.5 207607.5 ;
      RECT  34447.5 207237.5 34312.5 207302.5 ;
      RECT  34467.5 207785.0 34532.5 207920.0 ;
      RECT  34277.5 206942.5 34342.5 207077.5 ;
      RECT  34467.5 206942.5 34532.5 207077.5 ;
      RECT  34277.5 207472.5 34342.5 207607.5 ;
      RECT  34657.5 207472.5 34722.5 207607.5 ;
      RECT  34115.0 207237.5 34820.0 207302.5 ;
      RECT  34115.0 207922.5 34820.0 207987.5 ;
      RECT  35172.5 207472.5 35237.5 207987.5 ;
      RECT  34982.5 206942.5 35047.5 207077.5 ;
      RECT  35172.5 206942.5 35237.5 207077.5 ;
      RECT  35172.5 206942.5 35237.5 207077.5 ;
      RECT  34982.5 206942.5 35047.5 207077.5 ;
      RECT  34982.5 207472.5 35047.5 207607.5 ;
      RECT  35172.5 207472.5 35237.5 207607.5 ;
      RECT  35172.5 207472.5 35237.5 207607.5 ;
      RECT  34982.5 207472.5 35047.5 207607.5 ;
      RECT  35172.5 207472.5 35237.5 207607.5 ;
      RECT  35362.5 207472.5 35427.5 207607.5 ;
      RECT  35362.5 207472.5 35427.5 207607.5 ;
      RECT  35172.5 207472.5 35237.5 207607.5 ;
      RECT  35152.5 207237.5 35017.5 207302.5 ;
      RECT  35172.5 207785.0 35237.5 207920.0 ;
      RECT  34982.5 206942.5 35047.5 207077.5 ;
      RECT  35172.5 206942.5 35237.5 207077.5 ;
      RECT  34982.5 207472.5 35047.5 207607.5 ;
      RECT  35362.5 207472.5 35427.5 207607.5 ;
      RECT  34820.0 207237.5 35525.0 207302.5 ;
      RECT  34820.0 207922.5 35525.0 207987.5 ;
      RECT  35877.5 207472.5 35942.5 207987.5 ;
      RECT  35687.5 206942.5 35752.5 207077.5 ;
      RECT  35877.5 206942.5 35942.5 207077.5 ;
      RECT  35877.5 206942.5 35942.5 207077.5 ;
      RECT  35687.5 206942.5 35752.5 207077.5 ;
      RECT  35687.5 207472.5 35752.5 207607.5 ;
      RECT  35877.5 207472.5 35942.5 207607.5 ;
      RECT  35877.5 207472.5 35942.5 207607.5 ;
      RECT  35687.5 207472.5 35752.5 207607.5 ;
      RECT  35877.5 207472.5 35942.5 207607.5 ;
      RECT  36067.5 207472.5 36132.5 207607.5 ;
      RECT  36067.5 207472.5 36132.5 207607.5 ;
      RECT  35877.5 207472.5 35942.5 207607.5 ;
      RECT  35857.5 207237.5 35722.5 207302.5 ;
      RECT  35877.5 207785.0 35942.5 207920.0 ;
      RECT  35687.5 206942.5 35752.5 207077.5 ;
      RECT  35877.5 206942.5 35942.5 207077.5 ;
      RECT  35687.5 207472.5 35752.5 207607.5 ;
      RECT  36067.5 207472.5 36132.5 207607.5 ;
      RECT  35525.0 207237.5 36230.0 207302.5 ;
      RECT  35525.0 207922.5 36230.0 207987.5 ;
      RECT  36582.5 207472.5 36647.5 207987.5 ;
      RECT  36392.5 206942.5 36457.5 207077.5 ;
      RECT  36582.5 206942.5 36647.5 207077.5 ;
      RECT  36582.5 206942.5 36647.5 207077.5 ;
      RECT  36392.5 206942.5 36457.5 207077.5 ;
      RECT  36392.5 207472.5 36457.5 207607.5 ;
      RECT  36582.5 207472.5 36647.5 207607.5 ;
      RECT  36582.5 207472.5 36647.5 207607.5 ;
      RECT  36392.5 207472.5 36457.5 207607.5 ;
      RECT  36582.5 207472.5 36647.5 207607.5 ;
      RECT  36772.5 207472.5 36837.5 207607.5 ;
      RECT  36772.5 207472.5 36837.5 207607.5 ;
      RECT  36582.5 207472.5 36647.5 207607.5 ;
      RECT  36562.5 207237.5 36427.5 207302.5 ;
      RECT  36582.5 207785.0 36647.5 207920.0 ;
      RECT  36392.5 206942.5 36457.5 207077.5 ;
      RECT  36582.5 206942.5 36647.5 207077.5 ;
      RECT  36392.5 207472.5 36457.5 207607.5 ;
      RECT  36772.5 207472.5 36837.5 207607.5 ;
      RECT  36230.0 207237.5 36935.0 207302.5 ;
      RECT  36230.0 207922.5 36935.0 207987.5 ;
      RECT  37287.5 207472.5 37352.5 207987.5 ;
      RECT  37097.5 206942.5 37162.5 207077.5 ;
      RECT  37287.5 206942.5 37352.5 207077.5 ;
      RECT  37287.5 206942.5 37352.5 207077.5 ;
      RECT  37097.5 206942.5 37162.5 207077.5 ;
      RECT  37097.5 207472.5 37162.5 207607.5 ;
      RECT  37287.5 207472.5 37352.5 207607.5 ;
      RECT  37287.5 207472.5 37352.5 207607.5 ;
      RECT  37097.5 207472.5 37162.5 207607.5 ;
      RECT  37287.5 207472.5 37352.5 207607.5 ;
      RECT  37477.5 207472.5 37542.5 207607.5 ;
      RECT  37477.5 207472.5 37542.5 207607.5 ;
      RECT  37287.5 207472.5 37352.5 207607.5 ;
      RECT  37267.5 207237.5 37132.5 207302.5 ;
      RECT  37287.5 207785.0 37352.5 207920.0 ;
      RECT  37097.5 206942.5 37162.5 207077.5 ;
      RECT  37287.5 206942.5 37352.5 207077.5 ;
      RECT  37097.5 207472.5 37162.5 207607.5 ;
      RECT  37477.5 207472.5 37542.5 207607.5 ;
      RECT  36935.0 207237.5 37640.0 207302.5 ;
      RECT  36935.0 207922.5 37640.0 207987.5 ;
      RECT  37992.5 207472.5 38057.5 207987.5 ;
      RECT  37802.5 206942.5 37867.5 207077.5 ;
      RECT  37992.5 206942.5 38057.5 207077.5 ;
      RECT  37992.5 206942.5 38057.5 207077.5 ;
      RECT  37802.5 206942.5 37867.5 207077.5 ;
      RECT  37802.5 207472.5 37867.5 207607.5 ;
      RECT  37992.5 207472.5 38057.5 207607.5 ;
      RECT  37992.5 207472.5 38057.5 207607.5 ;
      RECT  37802.5 207472.5 37867.5 207607.5 ;
      RECT  37992.5 207472.5 38057.5 207607.5 ;
      RECT  38182.5 207472.5 38247.5 207607.5 ;
      RECT  38182.5 207472.5 38247.5 207607.5 ;
      RECT  37992.5 207472.5 38057.5 207607.5 ;
      RECT  37972.5 207237.5 37837.5 207302.5 ;
      RECT  37992.5 207785.0 38057.5 207920.0 ;
      RECT  37802.5 206942.5 37867.5 207077.5 ;
      RECT  37992.5 206942.5 38057.5 207077.5 ;
      RECT  37802.5 207472.5 37867.5 207607.5 ;
      RECT  38182.5 207472.5 38247.5 207607.5 ;
      RECT  37640.0 207237.5 38345.0 207302.5 ;
      RECT  37640.0 207922.5 38345.0 207987.5 ;
      RECT  38697.5 207472.5 38762.5 207987.5 ;
      RECT  38507.5 206942.5 38572.5 207077.5 ;
      RECT  38697.5 206942.5 38762.5 207077.5 ;
      RECT  38697.5 206942.5 38762.5 207077.5 ;
      RECT  38507.5 206942.5 38572.5 207077.5 ;
      RECT  38507.5 207472.5 38572.5 207607.5 ;
      RECT  38697.5 207472.5 38762.5 207607.5 ;
      RECT  38697.5 207472.5 38762.5 207607.5 ;
      RECT  38507.5 207472.5 38572.5 207607.5 ;
      RECT  38697.5 207472.5 38762.5 207607.5 ;
      RECT  38887.5 207472.5 38952.5 207607.5 ;
      RECT  38887.5 207472.5 38952.5 207607.5 ;
      RECT  38697.5 207472.5 38762.5 207607.5 ;
      RECT  38677.5 207237.5 38542.5 207302.5 ;
      RECT  38697.5 207785.0 38762.5 207920.0 ;
      RECT  38507.5 206942.5 38572.5 207077.5 ;
      RECT  38697.5 206942.5 38762.5 207077.5 ;
      RECT  38507.5 207472.5 38572.5 207607.5 ;
      RECT  38887.5 207472.5 38952.5 207607.5 ;
      RECT  38345.0 207237.5 39050.0 207302.5 ;
      RECT  38345.0 207922.5 39050.0 207987.5 ;
      RECT  39402.5 207472.5 39467.5 207987.5 ;
      RECT  39212.5 206942.5 39277.5 207077.5 ;
      RECT  39402.5 206942.5 39467.5 207077.5 ;
      RECT  39402.5 206942.5 39467.5 207077.5 ;
      RECT  39212.5 206942.5 39277.5 207077.5 ;
      RECT  39212.5 207472.5 39277.5 207607.5 ;
      RECT  39402.5 207472.5 39467.5 207607.5 ;
      RECT  39402.5 207472.5 39467.5 207607.5 ;
      RECT  39212.5 207472.5 39277.5 207607.5 ;
      RECT  39402.5 207472.5 39467.5 207607.5 ;
      RECT  39592.5 207472.5 39657.5 207607.5 ;
      RECT  39592.5 207472.5 39657.5 207607.5 ;
      RECT  39402.5 207472.5 39467.5 207607.5 ;
      RECT  39382.5 207237.5 39247.5 207302.5 ;
      RECT  39402.5 207785.0 39467.5 207920.0 ;
      RECT  39212.5 206942.5 39277.5 207077.5 ;
      RECT  39402.5 206942.5 39467.5 207077.5 ;
      RECT  39212.5 207472.5 39277.5 207607.5 ;
      RECT  39592.5 207472.5 39657.5 207607.5 ;
      RECT  39050.0 207237.5 39755.0 207302.5 ;
      RECT  39050.0 207922.5 39755.0 207987.5 ;
      RECT  40107.5 207472.5 40172.5 207987.5 ;
      RECT  39917.5 206942.5 39982.5 207077.5 ;
      RECT  40107.5 206942.5 40172.5 207077.5 ;
      RECT  40107.5 206942.5 40172.5 207077.5 ;
      RECT  39917.5 206942.5 39982.5 207077.5 ;
      RECT  39917.5 207472.5 39982.5 207607.5 ;
      RECT  40107.5 207472.5 40172.5 207607.5 ;
      RECT  40107.5 207472.5 40172.5 207607.5 ;
      RECT  39917.5 207472.5 39982.5 207607.5 ;
      RECT  40107.5 207472.5 40172.5 207607.5 ;
      RECT  40297.5 207472.5 40362.5 207607.5 ;
      RECT  40297.5 207472.5 40362.5 207607.5 ;
      RECT  40107.5 207472.5 40172.5 207607.5 ;
      RECT  40087.5 207237.5 39952.5 207302.5 ;
      RECT  40107.5 207785.0 40172.5 207920.0 ;
      RECT  39917.5 206942.5 39982.5 207077.5 ;
      RECT  40107.5 206942.5 40172.5 207077.5 ;
      RECT  39917.5 207472.5 39982.5 207607.5 ;
      RECT  40297.5 207472.5 40362.5 207607.5 ;
      RECT  39755.0 207237.5 40460.0 207302.5 ;
      RECT  39755.0 207922.5 40460.0 207987.5 ;
      RECT  40812.5 207472.5 40877.5 207987.5 ;
      RECT  40622.5 206942.5 40687.5 207077.5 ;
      RECT  40812.5 206942.5 40877.5 207077.5 ;
      RECT  40812.5 206942.5 40877.5 207077.5 ;
      RECT  40622.5 206942.5 40687.5 207077.5 ;
      RECT  40622.5 207472.5 40687.5 207607.5 ;
      RECT  40812.5 207472.5 40877.5 207607.5 ;
      RECT  40812.5 207472.5 40877.5 207607.5 ;
      RECT  40622.5 207472.5 40687.5 207607.5 ;
      RECT  40812.5 207472.5 40877.5 207607.5 ;
      RECT  41002.5 207472.5 41067.5 207607.5 ;
      RECT  41002.5 207472.5 41067.5 207607.5 ;
      RECT  40812.5 207472.5 40877.5 207607.5 ;
      RECT  40792.5 207237.5 40657.5 207302.5 ;
      RECT  40812.5 207785.0 40877.5 207920.0 ;
      RECT  40622.5 206942.5 40687.5 207077.5 ;
      RECT  40812.5 206942.5 40877.5 207077.5 ;
      RECT  40622.5 207472.5 40687.5 207607.5 ;
      RECT  41002.5 207472.5 41067.5 207607.5 ;
      RECT  40460.0 207237.5 41165.0 207302.5 ;
      RECT  40460.0 207922.5 41165.0 207987.5 ;
      RECT  41517.5 207472.5 41582.5 207987.5 ;
      RECT  41327.5 206942.5 41392.5 207077.5 ;
      RECT  41517.5 206942.5 41582.5 207077.5 ;
      RECT  41517.5 206942.5 41582.5 207077.5 ;
      RECT  41327.5 206942.5 41392.5 207077.5 ;
      RECT  41327.5 207472.5 41392.5 207607.5 ;
      RECT  41517.5 207472.5 41582.5 207607.5 ;
      RECT  41517.5 207472.5 41582.5 207607.5 ;
      RECT  41327.5 207472.5 41392.5 207607.5 ;
      RECT  41517.5 207472.5 41582.5 207607.5 ;
      RECT  41707.5 207472.5 41772.5 207607.5 ;
      RECT  41707.5 207472.5 41772.5 207607.5 ;
      RECT  41517.5 207472.5 41582.5 207607.5 ;
      RECT  41497.5 207237.5 41362.5 207302.5 ;
      RECT  41517.5 207785.0 41582.5 207920.0 ;
      RECT  41327.5 206942.5 41392.5 207077.5 ;
      RECT  41517.5 206942.5 41582.5 207077.5 ;
      RECT  41327.5 207472.5 41392.5 207607.5 ;
      RECT  41707.5 207472.5 41772.5 207607.5 ;
      RECT  41165.0 207237.5 41870.0 207302.5 ;
      RECT  41165.0 207922.5 41870.0 207987.5 ;
      RECT  42222.5 207472.5 42287.5 207987.5 ;
      RECT  42032.5 206942.5 42097.5 207077.5 ;
      RECT  42222.5 206942.5 42287.5 207077.5 ;
      RECT  42222.5 206942.5 42287.5 207077.5 ;
      RECT  42032.5 206942.5 42097.5 207077.5 ;
      RECT  42032.5 207472.5 42097.5 207607.5 ;
      RECT  42222.5 207472.5 42287.5 207607.5 ;
      RECT  42222.5 207472.5 42287.5 207607.5 ;
      RECT  42032.5 207472.5 42097.5 207607.5 ;
      RECT  42222.5 207472.5 42287.5 207607.5 ;
      RECT  42412.5 207472.5 42477.5 207607.5 ;
      RECT  42412.5 207472.5 42477.5 207607.5 ;
      RECT  42222.5 207472.5 42287.5 207607.5 ;
      RECT  42202.5 207237.5 42067.5 207302.5 ;
      RECT  42222.5 207785.0 42287.5 207920.0 ;
      RECT  42032.5 206942.5 42097.5 207077.5 ;
      RECT  42222.5 206942.5 42287.5 207077.5 ;
      RECT  42032.5 207472.5 42097.5 207607.5 ;
      RECT  42412.5 207472.5 42477.5 207607.5 ;
      RECT  41870.0 207237.5 42575.0 207302.5 ;
      RECT  41870.0 207922.5 42575.0 207987.5 ;
      RECT  42927.5 207472.5 42992.5 207987.5 ;
      RECT  42737.5 206942.5 42802.5 207077.5 ;
      RECT  42927.5 206942.5 42992.5 207077.5 ;
      RECT  42927.5 206942.5 42992.5 207077.5 ;
      RECT  42737.5 206942.5 42802.5 207077.5 ;
      RECT  42737.5 207472.5 42802.5 207607.5 ;
      RECT  42927.5 207472.5 42992.5 207607.5 ;
      RECT  42927.5 207472.5 42992.5 207607.5 ;
      RECT  42737.5 207472.5 42802.5 207607.5 ;
      RECT  42927.5 207472.5 42992.5 207607.5 ;
      RECT  43117.5 207472.5 43182.5 207607.5 ;
      RECT  43117.5 207472.5 43182.5 207607.5 ;
      RECT  42927.5 207472.5 42992.5 207607.5 ;
      RECT  42907.5 207237.5 42772.5 207302.5 ;
      RECT  42927.5 207785.0 42992.5 207920.0 ;
      RECT  42737.5 206942.5 42802.5 207077.5 ;
      RECT  42927.5 206942.5 42992.5 207077.5 ;
      RECT  42737.5 207472.5 42802.5 207607.5 ;
      RECT  43117.5 207472.5 43182.5 207607.5 ;
      RECT  42575.0 207237.5 43280.0 207302.5 ;
      RECT  42575.0 207922.5 43280.0 207987.5 ;
      RECT  43632.5 207472.5 43697.5 207987.5 ;
      RECT  43442.5 206942.5 43507.5 207077.5 ;
      RECT  43632.5 206942.5 43697.5 207077.5 ;
      RECT  43632.5 206942.5 43697.5 207077.5 ;
      RECT  43442.5 206942.5 43507.5 207077.5 ;
      RECT  43442.5 207472.5 43507.5 207607.5 ;
      RECT  43632.5 207472.5 43697.5 207607.5 ;
      RECT  43632.5 207472.5 43697.5 207607.5 ;
      RECT  43442.5 207472.5 43507.5 207607.5 ;
      RECT  43632.5 207472.5 43697.5 207607.5 ;
      RECT  43822.5 207472.5 43887.5 207607.5 ;
      RECT  43822.5 207472.5 43887.5 207607.5 ;
      RECT  43632.5 207472.5 43697.5 207607.5 ;
      RECT  43612.5 207237.5 43477.5 207302.5 ;
      RECT  43632.5 207785.0 43697.5 207920.0 ;
      RECT  43442.5 206942.5 43507.5 207077.5 ;
      RECT  43632.5 206942.5 43697.5 207077.5 ;
      RECT  43442.5 207472.5 43507.5 207607.5 ;
      RECT  43822.5 207472.5 43887.5 207607.5 ;
      RECT  43280.0 207237.5 43985.0 207302.5 ;
      RECT  43280.0 207922.5 43985.0 207987.5 ;
      RECT  44337.5 207472.5 44402.5 207987.5 ;
      RECT  44147.5 206942.5 44212.5 207077.5 ;
      RECT  44337.5 206942.5 44402.5 207077.5 ;
      RECT  44337.5 206942.5 44402.5 207077.5 ;
      RECT  44147.5 206942.5 44212.5 207077.5 ;
      RECT  44147.5 207472.5 44212.5 207607.5 ;
      RECT  44337.5 207472.5 44402.5 207607.5 ;
      RECT  44337.5 207472.5 44402.5 207607.5 ;
      RECT  44147.5 207472.5 44212.5 207607.5 ;
      RECT  44337.5 207472.5 44402.5 207607.5 ;
      RECT  44527.5 207472.5 44592.5 207607.5 ;
      RECT  44527.5 207472.5 44592.5 207607.5 ;
      RECT  44337.5 207472.5 44402.5 207607.5 ;
      RECT  44317.5 207237.5 44182.5 207302.5 ;
      RECT  44337.5 207785.0 44402.5 207920.0 ;
      RECT  44147.5 206942.5 44212.5 207077.5 ;
      RECT  44337.5 206942.5 44402.5 207077.5 ;
      RECT  44147.5 207472.5 44212.5 207607.5 ;
      RECT  44527.5 207472.5 44592.5 207607.5 ;
      RECT  43985.0 207237.5 44690.0 207302.5 ;
      RECT  43985.0 207922.5 44690.0 207987.5 ;
      RECT  45042.5 207472.5 45107.5 207987.5 ;
      RECT  44852.5 206942.5 44917.5 207077.5 ;
      RECT  45042.5 206942.5 45107.5 207077.5 ;
      RECT  45042.5 206942.5 45107.5 207077.5 ;
      RECT  44852.5 206942.5 44917.5 207077.5 ;
      RECT  44852.5 207472.5 44917.5 207607.5 ;
      RECT  45042.5 207472.5 45107.5 207607.5 ;
      RECT  45042.5 207472.5 45107.5 207607.5 ;
      RECT  44852.5 207472.5 44917.5 207607.5 ;
      RECT  45042.5 207472.5 45107.5 207607.5 ;
      RECT  45232.5 207472.5 45297.5 207607.5 ;
      RECT  45232.5 207472.5 45297.5 207607.5 ;
      RECT  45042.5 207472.5 45107.5 207607.5 ;
      RECT  45022.5 207237.5 44887.5 207302.5 ;
      RECT  45042.5 207785.0 45107.5 207920.0 ;
      RECT  44852.5 206942.5 44917.5 207077.5 ;
      RECT  45042.5 206942.5 45107.5 207077.5 ;
      RECT  44852.5 207472.5 44917.5 207607.5 ;
      RECT  45232.5 207472.5 45297.5 207607.5 ;
      RECT  44690.0 207237.5 45395.0 207302.5 ;
      RECT  44690.0 207922.5 45395.0 207987.5 ;
      RECT  45747.5 207472.5 45812.5 207987.5 ;
      RECT  45557.5 206942.5 45622.5 207077.5 ;
      RECT  45747.5 206942.5 45812.5 207077.5 ;
      RECT  45747.5 206942.5 45812.5 207077.5 ;
      RECT  45557.5 206942.5 45622.5 207077.5 ;
      RECT  45557.5 207472.5 45622.5 207607.5 ;
      RECT  45747.5 207472.5 45812.5 207607.5 ;
      RECT  45747.5 207472.5 45812.5 207607.5 ;
      RECT  45557.5 207472.5 45622.5 207607.5 ;
      RECT  45747.5 207472.5 45812.5 207607.5 ;
      RECT  45937.5 207472.5 46002.5 207607.5 ;
      RECT  45937.5 207472.5 46002.5 207607.5 ;
      RECT  45747.5 207472.5 45812.5 207607.5 ;
      RECT  45727.5 207237.5 45592.5 207302.5 ;
      RECT  45747.5 207785.0 45812.5 207920.0 ;
      RECT  45557.5 206942.5 45622.5 207077.5 ;
      RECT  45747.5 206942.5 45812.5 207077.5 ;
      RECT  45557.5 207472.5 45622.5 207607.5 ;
      RECT  45937.5 207472.5 46002.5 207607.5 ;
      RECT  45395.0 207237.5 46100.0 207302.5 ;
      RECT  45395.0 207922.5 46100.0 207987.5 ;
      RECT  46452.5 207472.5 46517.5 207987.5 ;
      RECT  46262.5 206942.5 46327.5 207077.5 ;
      RECT  46452.5 206942.5 46517.5 207077.5 ;
      RECT  46452.5 206942.5 46517.5 207077.5 ;
      RECT  46262.5 206942.5 46327.5 207077.5 ;
      RECT  46262.5 207472.5 46327.5 207607.5 ;
      RECT  46452.5 207472.5 46517.5 207607.5 ;
      RECT  46452.5 207472.5 46517.5 207607.5 ;
      RECT  46262.5 207472.5 46327.5 207607.5 ;
      RECT  46452.5 207472.5 46517.5 207607.5 ;
      RECT  46642.5 207472.5 46707.5 207607.5 ;
      RECT  46642.5 207472.5 46707.5 207607.5 ;
      RECT  46452.5 207472.5 46517.5 207607.5 ;
      RECT  46432.5 207237.5 46297.5 207302.5 ;
      RECT  46452.5 207785.0 46517.5 207920.0 ;
      RECT  46262.5 206942.5 46327.5 207077.5 ;
      RECT  46452.5 206942.5 46517.5 207077.5 ;
      RECT  46262.5 207472.5 46327.5 207607.5 ;
      RECT  46642.5 207472.5 46707.5 207607.5 ;
      RECT  46100.0 207237.5 46805.0 207302.5 ;
      RECT  46100.0 207922.5 46805.0 207987.5 ;
      RECT  47157.5 207472.5 47222.5 207987.5 ;
      RECT  46967.5 206942.5 47032.5 207077.5 ;
      RECT  47157.5 206942.5 47222.5 207077.5 ;
      RECT  47157.5 206942.5 47222.5 207077.5 ;
      RECT  46967.5 206942.5 47032.5 207077.5 ;
      RECT  46967.5 207472.5 47032.5 207607.5 ;
      RECT  47157.5 207472.5 47222.5 207607.5 ;
      RECT  47157.5 207472.5 47222.5 207607.5 ;
      RECT  46967.5 207472.5 47032.5 207607.5 ;
      RECT  47157.5 207472.5 47222.5 207607.5 ;
      RECT  47347.5 207472.5 47412.5 207607.5 ;
      RECT  47347.5 207472.5 47412.5 207607.5 ;
      RECT  47157.5 207472.5 47222.5 207607.5 ;
      RECT  47137.5 207237.5 47002.5 207302.5 ;
      RECT  47157.5 207785.0 47222.5 207920.0 ;
      RECT  46967.5 206942.5 47032.5 207077.5 ;
      RECT  47157.5 206942.5 47222.5 207077.5 ;
      RECT  46967.5 207472.5 47032.5 207607.5 ;
      RECT  47347.5 207472.5 47412.5 207607.5 ;
      RECT  46805.0 207237.5 47510.0 207302.5 ;
      RECT  46805.0 207922.5 47510.0 207987.5 ;
      RECT  47862.5 207472.5 47927.5 207987.5 ;
      RECT  47672.5 206942.5 47737.5 207077.5 ;
      RECT  47862.5 206942.5 47927.5 207077.5 ;
      RECT  47862.5 206942.5 47927.5 207077.5 ;
      RECT  47672.5 206942.5 47737.5 207077.5 ;
      RECT  47672.5 207472.5 47737.5 207607.5 ;
      RECT  47862.5 207472.5 47927.5 207607.5 ;
      RECT  47862.5 207472.5 47927.5 207607.5 ;
      RECT  47672.5 207472.5 47737.5 207607.5 ;
      RECT  47862.5 207472.5 47927.5 207607.5 ;
      RECT  48052.5 207472.5 48117.5 207607.5 ;
      RECT  48052.5 207472.5 48117.5 207607.5 ;
      RECT  47862.5 207472.5 47927.5 207607.5 ;
      RECT  47842.5 207237.5 47707.5 207302.5 ;
      RECT  47862.5 207785.0 47927.5 207920.0 ;
      RECT  47672.5 206942.5 47737.5 207077.5 ;
      RECT  47862.5 206942.5 47927.5 207077.5 ;
      RECT  47672.5 207472.5 47737.5 207607.5 ;
      RECT  48052.5 207472.5 48117.5 207607.5 ;
      RECT  47510.0 207237.5 48215.0 207302.5 ;
      RECT  47510.0 207922.5 48215.0 207987.5 ;
      RECT  48567.5 207472.5 48632.5 207987.5 ;
      RECT  48377.5 206942.5 48442.5 207077.5 ;
      RECT  48567.5 206942.5 48632.5 207077.5 ;
      RECT  48567.5 206942.5 48632.5 207077.5 ;
      RECT  48377.5 206942.5 48442.5 207077.5 ;
      RECT  48377.5 207472.5 48442.5 207607.5 ;
      RECT  48567.5 207472.5 48632.5 207607.5 ;
      RECT  48567.5 207472.5 48632.5 207607.5 ;
      RECT  48377.5 207472.5 48442.5 207607.5 ;
      RECT  48567.5 207472.5 48632.5 207607.5 ;
      RECT  48757.5 207472.5 48822.5 207607.5 ;
      RECT  48757.5 207472.5 48822.5 207607.5 ;
      RECT  48567.5 207472.5 48632.5 207607.5 ;
      RECT  48547.5 207237.5 48412.5 207302.5 ;
      RECT  48567.5 207785.0 48632.5 207920.0 ;
      RECT  48377.5 206942.5 48442.5 207077.5 ;
      RECT  48567.5 206942.5 48632.5 207077.5 ;
      RECT  48377.5 207472.5 48442.5 207607.5 ;
      RECT  48757.5 207472.5 48822.5 207607.5 ;
      RECT  48215.0 207237.5 48920.0 207302.5 ;
      RECT  48215.0 207922.5 48920.0 207987.5 ;
      RECT  49272.5 207472.5 49337.5 207987.5 ;
      RECT  49082.5 206942.5 49147.5 207077.5 ;
      RECT  49272.5 206942.5 49337.5 207077.5 ;
      RECT  49272.5 206942.5 49337.5 207077.5 ;
      RECT  49082.5 206942.5 49147.5 207077.5 ;
      RECT  49082.5 207472.5 49147.5 207607.5 ;
      RECT  49272.5 207472.5 49337.5 207607.5 ;
      RECT  49272.5 207472.5 49337.5 207607.5 ;
      RECT  49082.5 207472.5 49147.5 207607.5 ;
      RECT  49272.5 207472.5 49337.5 207607.5 ;
      RECT  49462.5 207472.5 49527.5 207607.5 ;
      RECT  49462.5 207472.5 49527.5 207607.5 ;
      RECT  49272.5 207472.5 49337.5 207607.5 ;
      RECT  49252.5 207237.5 49117.5 207302.5 ;
      RECT  49272.5 207785.0 49337.5 207920.0 ;
      RECT  49082.5 206942.5 49147.5 207077.5 ;
      RECT  49272.5 206942.5 49337.5 207077.5 ;
      RECT  49082.5 207472.5 49147.5 207607.5 ;
      RECT  49462.5 207472.5 49527.5 207607.5 ;
      RECT  48920.0 207237.5 49625.0 207302.5 ;
      RECT  48920.0 207922.5 49625.0 207987.5 ;
      RECT  49977.5 207472.5 50042.5 207987.5 ;
      RECT  49787.5 206942.5 49852.5 207077.5 ;
      RECT  49977.5 206942.5 50042.5 207077.5 ;
      RECT  49977.5 206942.5 50042.5 207077.5 ;
      RECT  49787.5 206942.5 49852.5 207077.5 ;
      RECT  49787.5 207472.5 49852.5 207607.5 ;
      RECT  49977.5 207472.5 50042.5 207607.5 ;
      RECT  49977.5 207472.5 50042.5 207607.5 ;
      RECT  49787.5 207472.5 49852.5 207607.5 ;
      RECT  49977.5 207472.5 50042.5 207607.5 ;
      RECT  50167.5 207472.5 50232.5 207607.5 ;
      RECT  50167.5 207472.5 50232.5 207607.5 ;
      RECT  49977.5 207472.5 50042.5 207607.5 ;
      RECT  49957.5 207237.5 49822.5 207302.5 ;
      RECT  49977.5 207785.0 50042.5 207920.0 ;
      RECT  49787.5 206942.5 49852.5 207077.5 ;
      RECT  49977.5 206942.5 50042.5 207077.5 ;
      RECT  49787.5 207472.5 49852.5 207607.5 ;
      RECT  50167.5 207472.5 50232.5 207607.5 ;
      RECT  49625.0 207237.5 50330.0 207302.5 ;
      RECT  49625.0 207922.5 50330.0 207987.5 ;
      RECT  50682.5 207472.5 50747.5 207987.5 ;
      RECT  50492.5 206942.5 50557.5 207077.5 ;
      RECT  50682.5 206942.5 50747.5 207077.5 ;
      RECT  50682.5 206942.5 50747.5 207077.5 ;
      RECT  50492.5 206942.5 50557.5 207077.5 ;
      RECT  50492.5 207472.5 50557.5 207607.5 ;
      RECT  50682.5 207472.5 50747.5 207607.5 ;
      RECT  50682.5 207472.5 50747.5 207607.5 ;
      RECT  50492.5 207472.5 50557.5 207607.5 ;
      RECT  50682.5 207472.5 50747.5 207607.5 ;
      RECT  50872.5 207472.5 50937.5 207607.5 ;
      RECT  50872.5 207472.5 50937.5 207607.5 ;
      RECT  50682.5 207472.5 50747.5 207607.5 ;
      RECT  50662.5 207237.5 50527.5 207302.5 ;
      RECT  50682.5 207785.0 50747.5 207920.0 ;
      RECT  50492.5 206942.5 50557.5 207077.5 ;
      RECT  50682.5 206942.5 50747.5 207077.5 ;
      RECT  50492.5 207472.5 50557.5 207607.5 ;
      RECT  50872.5 207472.5 50937.5 207607.5 ;
      RECT  50330.0 207237.5 51035.0 207302.5 ;
      RECT  50330.0 207922.5 51035.0 207987.5 ;
      RECT  51387.5 207472.5 51452.5 207987.5 ;
      RECT  51197.5 206942.5 51262.5 207077.5 ;
      RECT  51387.5 206942.5 51452.5 207077.5 ;
      RECT  51387.5 206942.5 51452.5 207077.5 ;
      RECT  51197.5 206942.5 51262.5 207077.5 ;
      RECT  51197.5 207472.5 51262.5 207607.5 ;
      RECT  51387.5 207472.5 51452.5 207607.5 ;
      RECT  51387.5 207472.5 51452.5 207607.5 ;
      RECT  51197.5 207472.5 51262.5 207607.5 ;
      RECT  51387.5 207472.5 51452.5 207607.5 ;
      RECT  51577.5 207472.5 51642.5 207607.5 ;
      RECT  51577.5 207472.5 51642.5 207607.5 ;
      RECT  51387.5 207472.5 51452.5 207607.5 ;
      RECT  51367.5 207237.5 51232.5 207302.5 ;
      RECT  51387.5 207785.0 51452.5 207920.0 ;
      RECT  51197.5 206942.5 51262.5 207077.5 ;
      RECT  51387.5 206942.5 51452.5 207077.5 ;
      RECT  51197.5 207472.5 51262.5 207607.5 ;
      RECT  51577.5 207472.5 51642.5 207607.5 ;
      RECT  51035.0 207237.5 51740.0 207302.5 ;
      RECT  51035.0 207922.5 51740.0 207987.5 ;
      RECT  52092.5 207472.5 52157.5 207987.5 ;
      RECT  51902.5 206942.5 51967.5 207077.5 ;
      RECT  52092.5 206942.5 52157.5 207077.5 ;
      RECT  52092.5 206942.5 52157.5 207077.5 ;
      RECT  51902.5 206942.5 51967.5 207077.5 ;
      RECT  51902.5 207472.5 51967.5 207607.5 ;
      RECT  52092.5 207472.5 52157.5 207607.5 ;
      RECT  52092.5 207472.5 52157.5 207607.5 ;
      RECT  51902.5 207472.5 51967.5 207607.5 ;
      RECT  52092.5 207472.5 52157.5 207607.5 ;
      RECT  52282.5 207472.5 52347.5 207607.5 ;
      RECT  52282.5 207472.5 52347.5 207607.5 ;
      RECT  52092.5 207472.5 52157.5 207607.5 ;
      RECT  52072.5 207237.5 51937.5 207302.5 ;
      RECT  52092.5 207785.0 52157.5 207920.0 ;
      RECT  51902.5 206942.5 51967.5 207077.5 ;
      RECT  52092.5 206942.5 52157.5 207077.5 ;
      RECT  51902.5 207472.5 51967.5 207607.5 ;
      RECT  52282.5 207472.5 52347.5 207607.5 ;
      RECT  51740.0 207237.5 52445.0 207302.5 ;
      RECT  51740.0 207922.5 52445.0 207987.5 ;
      RECT  52797.5 207472.5 52862.5 207987.5 ;
      RECT  52607.5 206942.5 52672.5 207077.5 ;
      RECT  52797.5 206942.5 52862.5 207077.5 ;
      RECT  52797.5 206942.5 52862.5 207077.5 ;
      RECT  52607.5 206942.5 52672.5 207077.5 ;
      RECT  52607.5 207472.5 52672.5 207607.5 ;
      RECT  52797.5 207472.5 52862.5 207607.5 ;
      RECT  52797.5 207472.5 52862.5 207607.5 ;
      RECT  52607.5 207472.5 52672.5 207607.5 ;
      RECT  52797.5 207472.5 52862.5 207607.5 ;
      RECT  52987.5 207472.5 53052.5 207607.5 ;
      RECT  52987.5 207472.5 53052.5 207607.5 ;
      RECT  52797.5 207472.5 52862.5 207607.5 ;
      RECT  52777.5 207237.5 52642.5 207302.5 ;
      RECT  52797.5 207785.0 52862.5 207920.0 ;
      RECT  52607.5 206942.5 52672.5 207077.5 ;
      RECT  52797.5 206942.5 52862.5 207077.5 ;
      RECT  52607.5 207472.5 52672.5 207607.5 ;
      RECT  52987.5 207472.5 53052.5 207607.5 ;
      RECT  52445.0 207237.5 53150.0 207302.5 ;
      RECT  52445.0 207922.5 53150.0 207987.5 ;
      RECT  53502.5 207472.5 53567.5 207987.5 ;
      RECT  53312.5 206942.5 53377.5 207077.5 ;
      RECT  53502.5 206942.5 53567.5 207077.5 ;
      RECT  53502.5 206942.5 53567.5 207077.5 ;
      RECT  53312.5 206942.5 53377.5 207077.5 ;
      RECT  53312.5 207472.5 53377.5 207607.5 ;
      RECT  53502.5 207472.5 53567.5 207607.5 ;
      RECT  53502.5 207472.5 53567.5 207607.5 ;
      RECT  53312.5 207472.5 53377.5 207607.5 ;
      RECT  53502.5 207472.5 53567.5 207607.5 ;
      RECT  53692.5 207472.5 53757.5 207607.5 ;
      RECT  53692.5 207472.5 53757.5 207607.5 ;
      RECT  53502.5 207472.5 53567.5 207607.5 ;
      RECT  53482.5 207237.5 53347.5 207302.5 ;
      RECT  53502.5 207785.0 53567.5 207920.0 ;
      RECT  53312.5 206942.5 53377.5 207077.5 ;
      RECT  53502.5 206942.5 53567.5 207077.5 ;
      RECT  53312.5 207472.5 53377.5 207607.5 ;
      RECT  53692.5 207472.5 53757.5 207607.5 ;
      RECT  53150.0 207237.5 53855.0 207302.5 ;
      RECT  53150.0 207922.5 53855.0 207987.5 ;
      RECT  54207.5 207472.5 54272.5 207987.5 ;
      RECT  54017.5 206942.5 54082.5 207077.5 ;
      RECT  54207.5 206942.5 54272.5 207077.5 ;
      RECT  54207.5 206942.5 54272.5 207077.5 ;
      RECT  54017.5 206942.5 54082.5 207077.5 ;
      RECT  54017.5 207472.5 54082.5 207607.5 ;
      RECT  54207.5 207472.5 54272.5 207607.5 ;
      RECT  54207.5 207472.5 54272.5 207607.5 ;
      RECT  54017.5 207472.5 54082.5 207607.5 ;
      RECT  54207.5 207472.5 54272.5 207607.5 ;
      RECT  54397.5 207472.5 54462.5 207607.5 ;
      RECT  54397.5 207472.5 54462.5 207607.5 ;
      RECT  54207.5 207472.5 54272.5 207607.5 ;
      RECT  54187.5 207237.5 54052.5 207302.5 ;
      RECT  54207.5 207785.0 54272.5 207920.0 ;
      RECT  54017.5 206942.5 54082.5 207077.5 ;
      RECT  54207.5 206942.5 54272.5 207077.5 ;
      RECT  54017.5 207472.5 54082.5 207607.5 ;
      RECT  54397.5 207472.5 54462.5 207607.5 ;
      RECT  53855.0 207237.5 54560.0 207302.5 ;
      RECT  53855.0 207922.5 54560.0 207987.5 ;
      RECT  54912.5 207472.5 54977.5 207987.5 ;
      RECT  54722.5 206942.5 54787.5 207077.5 ;
      RECT  54912.5 206942.5 54977.5 207077.5 ;
      RECT  54912.5 206942.5 54977.5 207077.5 ;
      RECT  54722.5 206942.5 54787.5 207077.5 ;
      RECT  54722.5 207472.5 54787.5 207607.5 ;
      RECT  54912.5 207472.5 54977.5 207607.5 ;
      RECT  54912.5 207472.5 54977.5 207607.5 ;
      RECT  54722.5 207472.5 54787.5 207607.5 ;
      RECT  54912.5 207472.5 54977.5 207607.5 ;
      RECT  55102.5 207472.5 55167.5 207607.5 ;
      RECT  55102.5 207472.5 55167.5 207607.5 ;
      RECT  54912.5 207472.5 54977.5 207607.5 ;
      RECT  54892.5 207237.5 54757.5 207302.5 ;
      RECT  54912.5 207785.0 54977.5 207920.0 ;
      RECT  54722.5 206942.5 54787.5 207077.5 ;
      RECT  54912.5 206942.5 54977.5 207077.5 ;
      RECT  54722.5 207472.5 54787.5 207607.5 ;
      RECT  55102.5 207472.5 55167.5 207607.5 ;
      RECT  54560.0 207237.5 55265.0 207302.5 ;
      RECT  54560.0 207922.5 55265.0 207987.5 ;
      RECT  55617.5 207472.5 55682.5 207987.5 ;
      RECT  55427.5 206942.5 55492.5 207077.5 ;
      RECT  55617.5 206942.5 55682.5 207077.5 ;
      RECT  55617.5 206942.5 55682.5 207077.5 ;
      RECT  55427.5 206942.5 55492.5 207077.5 ;
      RECT  55427.5 207472.5 55492.5 207607.5 ;
      RECT  55617.5 207472.5 55682.5 207607.5 ;
      RECT  55617.5 207472.5 55682.5 207607.5 ;
      RECT  55427.5 207472.5 55492.5 207607.5 ;
      RECT  55617.5 207472.5 55682.5 207607.5 ;
      RECT  55807.5 207472.5 55872.5 207607.5 ;
      RECT  55807.5 207472.5 55872.5 207607.5 ;
      RECT  55617.5 207472.5 55682.5 207607.5 ;
      RECT  55597.5 207237.5 55462.5 207302.5 ;
      RECT  55617.5 207785.0 55682.5 207920.0 ;
      RECT  55427.5 206942.5 55492.5 207077.5 ;
      RECT  55617.5 206942.5 55682.5 207077.5 ;
      RECT  55427.5 207472.5 55492.5 207607.5 ;
      RECT  55807.5 207472.5 55872.5 207607.5 ;
      RECT  55265.0 207237.5 55970.0 207302.5 ;
      RECT  55265.0 207922.5 55970.0 207987.5 ;
      RECT  56322.5 207472.5 56387.5 207987.5 ;
      RECT  56132.5 206942.5 56197.5 207077.5 ;
      RECT  56322.5 206942.5 56387.5 207077.5 ;
      RECT  56322.5 206942.5 56387.5 207077.5 ;
      RECT  56132.5 206942.5 56197.5 207077.5 ;
      RECT  56132.5 207472.5 56197.5 207607.5 ;
      RECT  56322.5 207472.5 56387.5 207607.5 ;
      RECT  56322.5 207472.5 56387.5 207607.5 ;
      RECT  56132.5 207472.5 56197.5 207607.5 ;
      RECT  56322.5 207472.5 56387.5 207607.5 ;
      RECT  56512.5 207472.5 56577.5 207607.5 ;
      RECT  56512.5 207472.5 56577.5 207607.5 ;
      RECT  56322.5 207472.5 56387.5 207607.5 ;
      RECT  56302.5 207237.5 56167.5 207302.5 ;
      RECT  56322.5 207785.0 56387.5 207920.0 ;
      RECT  56132.5 206942.5 56197.5 207077.5 ;
      RECT  56322.5 206942.5 56387.5 207077.5 ;
      RECT  56132.5 207472.5 56197.5 207607.5 ;
      RECT  56512.5 207472.5 56577.5 207607.5 ;
      RECT  55970.0 207237.5 56675.0 207302.5 ;
      RECT  55970.0 207922.5 56675.0 207987.5 ;
      RECT  57027.5 207472.5 57092.5 207987.5 ;
      RECT  56837.5 206942.5 56902.5 207077.5 ;
      RECT  57027.5 206942.5 57092.5 207077.5 ;
      RECT  57027.5 206942.5 57092.5 207077.5 ;
      RECT  56837.5 206942.5 56902.5 207077.5 ;
      RECT  56837.5 207472.5 56902.5 207607.5 ;
      RECT  57027.5 207472.5 57092.5 207607.5 ;
      RECT  57027.5 207472.5 57092.5 207607.5 ;
      RECT  56837.5 207472.5 56902.5 207607.5 ;
      RECT  57027.5 207472.5 57092.5 207607.5 ;
      RECT  57217.5 207472.5 57282.5 207607.5 ;
      RECT  57217.5 207472.5 57282.5 207607.5 ;
      RECT  57027.5 207472.5 57092.5 207607.5 ;
      RECT  57007.5 207237.5 56872.5 207302.5 ;
      RECT  57027.5 207785.0 57092.5 207920.0 ;
      RECT  56837.5 206942.5 56902.5 207077.5 ;
      RECT  57027.5 206942.5 57092.5 207077.5 ;
      RECT  56837.5 207472.5 56902.5 207607.5 ;
      RECT  57217.5 207472.5 57282.5 207607.5 ;
      RECT  56675.0 207237.5 57380.0 207302.5 ;
      RECT  56675.0 207922.5 57380.0 207987.5 ;
      RECT  57732.5 207472.5 57797.5 207987.5 ;
      RECT  57542.5 206942.5 57607.5 207077.5 ;
      RECT  57732.5 206942.5 57797.5 207077.5 ;
      RECT  57732.5 206942.5 57797.5 207077.5 ;
      RECT  57542.5 206942.5 57607.5 207077.5 ;
      RECT  57542.5 207472.5 57607.5 207607.5 ;
      RECT  57732.5 207472.5 57797.5 207607.5 ;
      RECT  57732.5 207472.5 57797.5 207607.5 ;
      RECT  57542.5 207472.5 57607.5 207607.5 ;
      RECT  57732.5 207472.5 57797.5 207607.5 ;
      RECT  57922.5 207472.5 57987.5 207607.5 ;
      RECT  57922.5 207472.5 57987.5 207607.5 ;
      RECT  57732.5 207472.5 57797.5 207607.5 ;
      RECT  57712.5 207237.5 57577.5 207302.5 ;
      RECT  57732.5 207785.0 57797.5 207920.0 ;
      RECT  57542.5 206942.5 57607.5 207077.5 ;
      RECT  57732.5 206942.5 57797.5 207077.5 ;
      RECT  57542.5 207472.5 57607.5 207607.5 ;
      RECT  57922.5 207472.5 57987.5 207607.5 ;
      RECT  57380.0 207237.5 58085.0 207302.5 ;
      RECT  57380.0 207922.5 58085.0 207987.5 ;
      RECT  58437.5 207472.5 58502.5 207987.5 ;
      RECT  58247.5 206942.5 58312.5 207077.5 ;
      RECT  58437.5 206942.5 58502.5 207077.5 ;
      RECT  58437.5 206942.5 58502.5 207077.5 ;
      RECT  58247.5 206942.5 58312.5 207077.5 ;
      RECT  58247.5 207472.5 58312.5 207607.5 ;
      RECT  58437.5 207472.5 58502.5 207607.5 ;
      RECT  58437.5 207472.5 58502.5 207607.5 ;
      RECT  58247.5 207472.5 58312.5 207607.5 ;
      RECT  58437.5 207472.5 58502.5 207607.5 ;
      RECT  58627.5 207472.5 58692.5 207607.5 ;
      RECT  58627.5 207472.5 58692.5 207607.5 ;
      RECT  58437.5 207472.5 58502.5 207607.5 ;
      RECT  58417.5 207237.5 58282.5 207302.5 ;
      RECT  58437.5 207785.0 58502.5 207920.0 ;
      RECT  58247.5 206942.5 58312.5 207077.5 ;
      RECT  58437.5 206942.5 58502.5 207077.5 ;
      RECT  58247.5 207472.5 58312.5 207607.5 ;
      RECT  58627.5 207472.5 58692.5 207607.5 ;
      RECT  58085.0 207237.5 58790.0 207302.5 ;
      RECT  58085.0 207922.5 58790.0 207987.5 ;
      RECT  59142.5 207472.5 59207.5 207987.5 ;
      RECT  58952.5 206942.5 59017.5 207077.5 ;
      RECT  59142.5 206942.5 59207.5 207077.5 ;
      RECT  59142.5 206942.5 59207.5 207077.5 ;
      RECT  58952.5 206942.5 59017.5 207077.5 ;
      RECT  58952.5 207472.5 59017.5 207607.5 ;
      RECT  59142.5 207472.5 59207.5 207607.5 ;
      RECT  59142.5 207472.5 59207.5 207607.5 ;
      RECT  58952.5 207472.5 59017.5 207607.5 ;
      RECT  59142.5 207472.5 59207.5 207607.5 ;
      RECT  59332.5 207472.5 59397.5 207607.5 ;
      RECT  59332.5 207472.5 59397.5 207607.5 ;
      RECT  59142.5 207472.5 59207.5 207607.5 ;
      RECT  59122.5 207237.5 58987.5 207302.5 ;
      RECT  59142.5 207785.0 59207.5 207920.0 ;
      RECT  58952.5 206942.5 59017.5 207077.5 ;
      RECT  59142.5 206942.5 59207.5 207077.5 ;
      RECT  58952.5 207472.5 59017.5 207607.5 ;
      RECT  59332.5 207472.5 59397.5 207607.5 ;
      RECT  58790.0 207237.5 59495.0 207302.5 ;
      RECT  58790.0 207922.5 59495.0 207987.5 ;
      RECT  59847.5 207472.5 59912.5 207987.5 ;
      RECT  59657.5 206942.5 59722.5 207077.5 ;
      RECT  59847.5 206942.5 59912.5 207077.5 ;
      RECT  59847.5 206942.5 59912.5 207077.5 ;
      RECT  59657.5 206942.5 59722.5 207077.5 ;
      RECT  59657.5 207472.5 59722.5 207607.5 ;
      RECT  59847.5 207472.5 59912.5 207607.5 ;
      RECT  59847.5 207472.5 59912.5 207607.5 ;
      RECT  59657.5 207472.5 59722.5 207607.5 ;
      RECT  59847.5 207472.5 59912.5 207607.5 ;
      RECT  60037.5 207472.5 60102.5 207607.5 ;
      RECT  60037.5 207472.5 60102.5 207607.5 ;
      RECT  59847.5 207472.5 59912.5 207607.5 ;
      RECT  59827.5 207237.5 59692.5 207302.5 ;
      RECT  59847.5 207785.0 59912.5 207920.0 ;
      RECT  59657.5 206942.5 59722.5 207077.5 ;
      RECT  59847.5 206942.5 59912.5 207077.5 ;
      RECT  59657.5 207472.5 59722.5 207607.5 ;
      RECT  60037.5 207472.5 60102.5 207607.5 ;
      RECT  59495.0 207237.5 60200.0 207302.5 ;
      RECT  59495.0 207922.5 60200.0 207987.5 ;
      RECT  60552.5 207472.5 60617.5 207987.5 ;
      RECT  60362.5 206942.5 60427.5 207077.5 ;
      RECT  60552.5 206942.5 60617.5 207077.5 ;
      RECT  60552.5 206942.5 60617.5 207077.5 ;
      RECT  60362.5 206942.5 60427.5 207077.5 ;
      RECT  60362.5 207472.5 60427.5 207607.5 ;
      RECT  60552.5 207472.5 60617.5 207607.5 ;
      RECT  60552.5 207472.5 60617.5 207607.5 ;
      RECT  60362.5 207472.5 60427.5 207607.5 ;
      RECT  60552.5 207472.5 60617.5 207607.5 ;
      RECT  60742.5 207472.5 60807.5 207607.5 ;
      RECT  60742.5 207472.5 60807.5 207607.5 ;
      RECT  60552.5 207472.5 60617.5 207607.5 ;
      RECT  60532.5 207237.5 60397.5 207302.5 ;
      RECT  60552.5 207785.0 60617.5 207920.0 ;
      RECT  60362.5 206942.5 60427.5 207077.5 ;
      RECT  60552.5 206942.5 60617.5 207077.5 ;
      RECT  60362.5 207472.5 60427.5 207607.5 ;
      RECT  60742.5 207472.5 60807.5 207607.5 ;
      RECT  60200.0 207237.5 60905.0 207302.5 ;
      RECT  60200.0 207922.5 60905.0 207987.5 ;
      RECT  61257.5 207472.5 61322.5 207987.5 ;
      RECT  61067.5 206942.5 61132.5 207077.5 ;
      RECT  61257.5 206942.5 61322.5 207077.5 ;
      RECT  61257.5 206942.5 61322.5 207077.5 ;
      RECT  61067.5 206942.5 61132.5 207077.5 ;
      RECT  61067.5 207472.5 61132.5 207607.5 ;
      RECT  61257.5 207472.5 61322.5 207607.5 ;
      RECT  61257.5 207472.5 61322.5 207607.5 ;
      RECT  61067.5 207472.5 61132.5 207607.5 ;
      RECT  61257.5 207472.5 61322.5 207607.5 ;
      RECT  61447.5 207472.5 61512.5 207607.5 ;
      RECT  61447.5 207472.5 61512.5 207607.5 ;
      RECT  61257.5 207472.5 61322.5 207607.5 ;
      RECT  61237.5 207237.5 61102.5 207302.5 ;
      RECT  61257.5 207785.0 61322.5 207920.0 ;
      RECT  61067.5 206942.5 61132.5 207077.5 ;
      RECT  61257.5 206942.5 61322.5 207077.5 ;
      RECT  61067.5 207472.5 61132.5 207607.5 ;
      RECT  61447.5 207472.5 61512.5 207607.5 ;
      RECT  60905.0 207237.5 61610.0 207302.5 ;
      RECT  60905.0 207922.5 61610.0 207987.5 ;
      RECT  61962.5 207472.5 62027.5 207987.5 ;
      RECT  61772.5 206942.5 61837.5 207077.5 ;
      RECT  61962.5 206942.5 62027.5 207077.5 ;
      RECT  61962.5 206942.5 62027.5 207077.5 ;
      RECT  61772.5 206942.5 61837.5 207077.5 ;
      RECT  61772.5 207472.5 61837.5 207607.5 ;
      RECT  61962.5 207472.5 62027.5 207607.5 ;
      RECT  61962.5 207472.5 62027.5 207607.5 ;
      RECT  61772.5 207472.5 61837.5 207607.5 ;
      RECT  61962.5 207472.5 62027.5 207607.5 ;
      RECT  62152.5 207472.5 62217.5 207607.5 ;
      RECT  62152.5 207472.5 62217.5 207607.5 ;
      RECT  61962.5 207472.5 62027.5 207607.5 ;
      RECT  61942.5 207237.5 61807.5 207302.5 ;
      RECT  61962.5 207785.0 62027.5 207920.0 ;
      RECT  61772.5 206942.5 61837.5 207077.5 ;
      RECT  61962.5 206942.5 62027.5 207077.5 ;
      RECT  61772.5 207472.5 61837.5 207607.5 ;
      RECT  62152.5 207472.5 62217.5 207607.5 ;
      RECT  61610.0 207237.5 62315.0 207302.5 ;
      RECT  61610.0 207922.5 62315.0 207987.5 ;
      RECT  62667.5 207472.5 62732.5 207987.5 ;
      RECT  62477.5 206942.5 62542.5 207077.5 ;
      RECT  62667.5 206942.5 62732.5 207077.5 ;
      RECT  62667.5 206942.5 62732.5 207077.5 ;
      RECT  62477.5 206942.5 62542.5 207077.5 ;
      RECT  62477.5 207472.5 62542.5 207607.5 ;
      RECT  62667.5 207472.5 62732.5 207607.5 ;
      RECT  62667.5 207472.5 62732.5 207607.5 ;
      RECT  62477.5 207472.5 62542.5 207607.5 ;
      RECT  62667.5 207472.5 62732.5 207607.5 ;
      RECT  62857.5 207472.5 62922.5 207607.5 ;
      RECT  62857.5 207472.5 62922.5 207607.5 ;
      RECT  62667.5 207472.5 62732.5 207607.5 ;
      RECT  62647.5 207237.5 62512.5 207302.5 ;
      RECT  62667.5 207785.0 62732.5 207920.0 ;
      RECT  62477.5 206942.5 62542.5 207077.5 ;
      RECT  62667.5 206942.5 62732.5 207077.5 ;
      RECT  62477.5 207472.5 62542.5 207607.5 ;
      RECT  62857.5 207472.5 62922.5 207607.5 ;
      RECT  62315.0 207237.5 63020.0 207302.5 ;
      RECT  62315.0 207922.5 63020.0 207987.5 ;
      RECT  63372.5 207472.5 63437.5 207987.5 ;
      RECT  63182.5 206942.5 63247.5 207077.5 ;
      RECT  63372.5 206942.5 63437.5 207077.5 ;
      RECT  63372.5 206942.5 63437.5 207077.5 ;
      RECT  63182.5 206942.5 63247.5 207077.5 ;
      RECT  63182.5 207472.5 63247.5 207607.5 ;
      RECT  63372.5 207472.5 63437.5 207607.5 ;
      RECT  63372.5 207472.5 63437.5 207607.5 ;
      RECT  63182.5 207472.5 63247.5 207607.5 ;
      RECT  63372.5 207472.5 63437.5 207607.5 ;
      RECT  63562.5 207472.5 63627.5 207607.5 ;
      RECT  63562.5 207472.5 63627.5 207607.5 ;
      RECT  63372.5 207472.5 63437.5 207607.5 ;
      RECT  63352.5 207237.5 63217.5 207302.5 ;
      RECT  63372.5 207785.0 63437.5 207920.0 ;
      RECT  63182.5 206942.5 63247.5 207077.5 ;
      RECT  63372.5 206942.5 63437.5 207077.5 ;
      RECT  63182.5 207472.5 63247.5 207607.5 ;
      RECT  63562.5 207472.5 63627.5 207607.5 ;
      RECT  63020.0 207237.5 63725.0 207302.5 ;
      RECT  63020.0 207922.5 63725.0 207987.5 ;
      RECT  64077.5 207472.5 64142.5 207987.5 ;
      RECT  63887.5 206942.5 63952.5 207077.5 ;
      RECT  64077.5 206942.5 64142.5 207077.5 ;
      RECT  64077.5 206942.5 64142.5 207077.5 ;
      RECT  63887.5 206942.5 63952.5 207077.5 ;
      RECT  63887.5 207472.5 63952.5 207607.5 ;
      RECT  64077.5 207472.5 64142.5 207607.5 ;
      RECT  64077.5 207472.5 64142.5 207607.5 ;
      RECT  63887.5 207472.5 63952.5 207607.5 ;
      RECT  64077.5 207472.5 64142.5 207607.5 ;
      RECT  64267.5 207472.5 64332.5 207607.5 ;
      RECT  64267.5 207472.5 64332.5 207607.5 ;
      RECT  64077.5 207472.5 64142.5 207607.5 ;
      RECT  64057.5 207237.5 63922.5 207302.5 ;
      RECT  64077.5 207785.0 64142.5 207920.0 ;
      RECT  63887.5 206942.5 63952.5 207077.5 ;
      RECT  64077.5 206942.5 64142.5 207077.5 ;
      RECT  63887.5 207472.5 63952.5 207607.5 ;
      RECT  64267.5 207472.5 64332.5 207607.5 ;
      RECT  63725.0 207237.5 64430.0 207302.5 ;
      RECT  63725.0 207922.5 64430.0 207987.5 ;
      RECT  64782.5 207472.5 64847.5 207987.5 ;
      RECT  64592.5 206942.5 64657.5 207077.5 ;
      RECT  64782.5 206942.5 64847.5 207077.5 ;
      RECT  64782.5 206942.5 64847.5 207077.5 ;
      RECT  64592.5 206942.5 64657.5 207077.5 ;
      RECT  64592.5 207472.5 64657.5 207607.5 ;
      RECT  64782.5 207472.5 64847.5 207607.5 ;
      RECT  64782.5 207472.5 64847.5 207607.5 ;
      RECT  64592.5 207472.5 64657.5 207607.5 ;
      RECT  64782.5 207472.5 64847.5 207607.5 ;
      RECT  64972.5 207472.5 65037.5 207607.5 ;
      RECT  64972.5 207472.5 65037.5 207607.5 ;
      RECT  64782.5 207472.5 64847.5 207607.5 ;
      RECT  64762.5 207237.5 64627.5 207302.5 ;
      RECT  64782.5 207785.0 64847.5 207920.0 ;
      RECT  64592.5 206942.5 64657.5 207077.5 ;
      RECT  64782.5 206942.5 64847.5 207077.5 ;
      RECT  64592.5 207472.5 64657.5 207607.5 ;
      RECT  64972.5 207472.5 65037.5 207607.5 ;
      RECT  64430.0 207237.5 65135.0 207302.5 ;
      RECT  64430.0 207922.5 65135.0 207987.5 ;
      RECT  65487.5 207472.5 65552.5 207987.5 ;
      RECT  65297.5 206942.5 65362.5 207077.5 ;
      RECT  65487.5 206942.5 65552.5 207077.5 ;
      RECT  65487.5 206942.5 65552.5 207077.5 ;
      RECT  65297.5 206942.5 65362.5 207077.5 ;
      RECT  65297.5 207472.5 65362.5 207607.5 ;
      RECT  65487.5 207472.5 65552.5 207607.5 ;
      RECT  65487.5 207472.5 65552.5 207607.5 ;
      RECT  65297.5 207472.5 65362.5 207607.5 ;
      RECT  65487.5 207472.5 65552.5 207607.5 ;
      RECT  65677.5 207472.5 65742.5 207607.5 ;
      RECT  65677.5 207472.5 65742.5 207607.5 ;
      RECT  65487.5 207472.5 65552.5 207607.5 ;
      RECT  65467.5 207237.5 65332.5 207302.5 ;
      RECT  65487.5 207785.0 65552.5 207920.0 ;
      RECT  65297.5 206942.5 65362.5 207077.5 ;
      RECT  65487.5 206942.5 65552.5 207077.5 ;
      RECT  65297.5 207472.5 65362.5 207607.5 ;
      RECT  65677.5 207472.5 65742.5 207607.5 ;
      RECT  65135.0 207237.5 65840.0 207302.5 ;
      RECT  65135.0 207922.5 65840.0 207987.5 ;
      RECT  66192.5 207472.5 66257.5 207987.5 ;
      RECT  66002.5 206942.5 66067.5 207077.5 ;
      RECT  66192.5 206942.5 66257.5 207077.5 ;
      RECT  66192.5 206942.5 66257.5 207077.5 ;
      RECT  66002.5 206942.5 66067.5 207077.5 ;
      RECT  66002.5 207472.5 66067.5 207607.5 ;
      RECT  66192.5 207472.5 66257.5 207607.5 ;
      RECT  66192.5 207472.5 66257.5 207607.5 ;
      RECT  66002.5 207472.5 66067.5 207607.5 ;
      RECT  66192.5 207472.5 66257.5 207607.5 ;
      RECT  66382.5 207472.5 66447.5 207607.5 ;
      RECT  66382.5 207472.5 66447.5 207607.5 ;
      RECT  66192.5 207472.5 66257.5 207607.5 ;
      RECT  66172.5 207237.5 66037.5 207302.5 ;
      RECT  66192.5 207785.0 66257.5 207920.0 ;
      RECT  66002.5 206942.5 66067.5 207077.5 ;
      RECT  66192.5 206942.5 66257.5 207077.5 ;
      RECT  66002.5 207472.5 66067.5 207607.5 ;
      RECT  66382.5 207472.5 66447.5 207607.5 ;
      RECT  65840.0 207237.5 66545.0 207302.5 ;
      RECT  65840.0 207922.5 66545.0 207987.5 ;
      RECT  66897.5 207472.5 66962.5 207987.5 ;
      RECT  66707.5 206942.5 66772.5 207077.5 ;
      RECT  66897.5 206942.5 66962.5 207077.5 ;
      RECT  66897.5 206942.5 66962.5 207077.5 ;
      RECT  66707.5 206942.5 66772.5 207077.5 ;
      RECT  66707.5 207472.5 66772.5 207607.5 ;
      RECT  66897.5 207472.5 66962.5 207607.5 ;
      RECT  66897.5 207472.5 66962.5 207607.5 ;
      RECT  66707.5 207472.5 66772.5 207607.5 ;
      RECT  66897.5 207472.5 66962.5 207607.5 ;
      RECT  67087.5 207472.5 67152.5 207607.5 ;
      RECT  67087.5 207472.5 67152.5 207607.5 ;
      RECT  66897.5 207472.5 66962.5 207607.5 ;
      RECT  66877.5 207237.5 66742.5 207302.5 ;
      RECT  66897.5 207785.0 66962.5 207920.0 ;
      RECT  66707.5 206942.5 66772.5 207077.5 ;
      RECT  66897.5 206942.5 66962.5 207077.5 ;
      RECT  66707.5 207472.5 66772.5 207607.5 ;
      RECT  67087.5 207472.5 67152.5 207607.5 ;
      RECT  66545.0 207237.5 67250.0 207302.5 ;
      RECT  66545.0 207922.5 67250.0 207987.5 ;
      RECT  67602.5 207472.5 67667.5 207987.5 ;
      RECT  67412.5 206942.5 67477.5 207077.5 ;
      RECT  67602.5 206942.5 67667.5 207077.5 ;
      RECT  67602.5 206942.5 67667.5 207077.5 ;
      RECT  67412.5 206942.5 67477.5 207077.5 ;
      RECT  67412.5 207472.5 67477.5 207607.5 ;
      RECT  67602.5 207472.5 67667.5 207607.5 ;
      RECT  67602.5 207472.5 67667.5 207607.5 ;
      RECT  67412.5 207472.5 67477.5 207607.5 ;
      RECT  67602.5 207472.5 67667.5 207607.5 ;
      RECT  67792.5 207472.5 67857.5 207607.5 ;
      RECT  67792.5 207472.5 67857.5 207607.5 ;
      RECT  67602.5 207472.5 67667.5 207607.5 ;
      RECT  67582.5 207237.5 67447.5 207302.5 ;
      RECT  67602.5 207785.0 67667.5 207920.0 ;
      RECT  67412.5 206942.5 67477.5 207077.5 ;
      RECT  67602.5 206942.5 67667.5 207077.5 ;
      RECT  67412.5 207472.5 67477.5 207607.5 ;
      RECT  67792.5 207472.5 67857.5 207607.5 ;
      RECT  67250.0 207237.5 67955.0 207302.5 ;
      RECT  67250.0 207922.5 67955.0 207987.5 ;
      RECT  68307.5 207472.5 68372.5 207987.5 ;
      RECT  68117.5 206942.5 68182.5 207077.5 ;
      RECT  68307.5 206942.5 68372.5 207077.5 ;
      RECT  68307.5 206942.5 68372.5 207077.5 ;
      RECT  68117.5 206942.5 68182.5 207077.5 ;
      RECT  68117.5 207472.5 68182.5 207607.5 ;
      RECT  68307.5 207472.5 68372.5 207607.5 ;
      RECT  68307.5 207472.5 68372.5 207607.5 ;
      RECT  68117.5 207472.5 68182.5 207607.5 ;
      RECT  68307.5 207472.5 68372.5 207607.5 ;
      RECT  68497.5 207472.5 68562.5 207607.5 ;
      RECT  68497.5 207472.5 68562.5 207607.5 ;
      RECT  68307.5 207472.5 68372.5 207607.5 ;
      RECT  68287.5 207237.5 68152.5 207302.5 ;
      RECT  68307.5 207785.0 68372.5 207920.0 ;
      RECT  68117.5 206942.5 68182.5 207077.5 ;
      RECT  68307.5 206942.5 68372.5 207077.5 ;
      RECT  68117.5 207472.5 68182.5 207607.5 ;
      RECT  68497.5 207472.5 68562.5 207607.5 ;
      RECT  67955.0 207237.5 68660.0 207302.5 ;
      RECT  67955.0 207922.5 68660.0 207987.5 ;
      RECT  69012.5 207472.5 69077.5 207987.5 ;
      RECT  68822.5 206942.5 68887.5 207077.5 ;
      RECT  69012.5 206942.5 69077.5 207077.5 ;
      RECT  69012.5 206942.5 69077.5 207077.5 ;
      RECT  68822.5 206942.5 68887.5 207077.5 ;
      RECT  68822.5 207472.5 68887.5 207607.5 ;
      RECT  69012.5 207472.5 69077.5 207607.5 ;
      RECT  69012.5 207472.5 69077.5 207607.5 ;
      RECT  68822.5 207472.5 68887.5 207607.5 ;
      RECT  69012.5 207472.5 69077.5 207607.5 ;
      RECT  69202.5 207472.5 69267.5 207607.5 ;
      RECT  69202.5 207472.5 69267.5 207607.5 ;
      RECT  69012.5 207472.5 69077.5 207607.5 ;
      RECT  68992.5 207237.5 68857.5 207302.5 ;
      RECT  69012.5 207785.0 69077.5 207920.0 ;
      RECT  68822.5 206942.5 68887.5 207077.5 ;
      RECT  69012.5 206942.5 69077.5 207077.5 ;
      RECT  68822.5 207472.5 68887.5 207607.5 ;
      RECT  69202.5 207472.5 69267.5 207607.5 ;
      RECT  68660.0 207237.5 69365.0 207302.5 ;
      RECT  68660.0 207922.5 69365.0 207987.5 ;
      RECT  69717.5 207472.5 69782.5 207987.5 ;
      RECT  69527.5 206942.5 69592.5 207077.5 ;
      RECT  69717.5 206942.5 69782.5 207077.5 ;
      RECT  69717.5 206942.5 69782.5 207077.5 ;
      RECT  69527.5 206942.5 69592.5 207077.5 ;
      RECT  69527.5 207472.5 69592.5 207607.5 ;
      RECT  69717.5 207472.5 69782.5 207607.5 ;
      RECT  69717.5 207472.5 69782.5 207607.5 ;
      RECT  69527.5 207472.5 69592.5 207607.5 ;
      RECT  69717.5 207472.5 69782.5 207607.5 ;
      RECT  69907.5 207472.5 69972.5 207607.5 ;
      RECT  69907.5 207472.5 69972.5 207607.5 ;
      RECT  69717.5 207472.5 69782.5 207607.5 ;
      RECT  69697.5 207237.5 69562.5 207302.5 ;
      RECT  69717.5 207785.0 69782.5 207920.0 ;
      RECT  69527.5 206942.5 69592.5 207077.5 ;
      RECT  69717.5 206942.5 69782.5 207077.5 ;
      RECT  69527.5 207472.5 69592.5 207607.5 ;
      RECT  69907.5 207472.5 69972.5 207607.5 ;
      RECT  69365.0 207237.5 70070.0 207302.5 ;
      RECT  69365.0 207922.5 70070.0 207987.5 ;
      RECT  70422.5 207472.5 70487.5 207987.5 ;
      RECT  70232.5 206942.5 70297.5 207077.5 ;
      RECT  70422.5 206942.5 70487.5 207077.5 ;
      RECT  70422.5 206942.5 70487.5 207077.5 ;
      RECT  70232.5 206942.5 70297.5 207077.5 ;
      RECT  70232.5 207472.5 70297.5 207607.5 ;
      RECT  70422.5 207472.5 70487.5 207607.5 ;
      RECT  70422.5 207472.5 70487.5 207607.5 ;
      RECT  70232.5 207472.5 70297.5 207607.5 ;
      RECT  70422.5 207472.5 70487.5 207607.5 ;
      RECT  70612.5 207472.5 70677.5 207607.5 ;
      RECT  70612.5 207472.5 70677.5 207607.5 ;
      RECT  70422.5 207472.5 70487.5 207607.5 ;
      RECT  70402.5 207237.5 70267.5 207302.5 ;
      RECT  70422.5 207785.0 70487.5 207920.0 ;
      RECT  70232.5 206942.5 70297.5 207077.5 ;
      RECT  70422.5 206942.5 70487.5 207077.5 ;
      RECT  70232.5 207472.5 70297.5 207607.5 ;
      RECT  70612.5 207472.5 70677.5 207607.5 ;
      RECT  70070.0 207237.5 70775.0 207302.5 ;
      RECT  70070.0 207922.5 70775.0 207987.5 ;
      RECT  71127.5 207472.5 71192.5 207987.5 ;
      RECT  70937.5 206942.5 71002.5 207077.5 ;
      RECT  71127.5 206942.5 71192.5 207077.5 ;
      RECT  71127.5 206942.5 71192.5 207077.5 ;
      RECT  70937.5 206942.5 71002.5 207077.5 ;
      RECT  70937.5 207472.5 71002.5 207607.5 ;
      RECT  71127.5 207472.5 71192.5 207607.5 ;
      RECT  71127.5 207472.5 71192.5 207607.5 ;
      RECT  70937.5 207472.5 71002.5 207607.5 ;
      RECT  71127.5 207472.5 71192.5 207607.5 ;
      RECT  71317.5 207472.5 71382.5 207607.5 ;
      RECT  71317.5 207472.5 71382.5 207607.5 ;
      RECT  71127.5 207472.5 71192.5 207607.5 ;
      RECT  71107.5 207237.5 70972.5 207302.5 ;
      RECT  71127.5 207785.0 71192.5 207920.0 ;
      RECT  70937.5 206942.5 71002.5 207077.5 ;
      RECT  71127.5 206942.5 71192.5 207077.5 ;
      RECT  70937.5 207472.5 71002.5 207607.5 ;
      RECT  71317.5 207472.5 71382.5 207607.5 ;
      RECT  70775.0 207237.5 71480.0 207302.5 ;
      RECT  70775.0 207922.5 71480.0 207987.5 ;
      RECT  71832.5 207472.5 71897.5 207987.5 ;
      RECT  71642.5 206942.5 71707.5 207077.5 ;
      RECT  71832.5 206942.5 71897.5 207077.5 ;
      RECT  71832.5 206942.5 71897.5 207077.5 ;
      RECT  71642.5 206942.5 71707.5 207077.5 ;
      RECT  71642.5 207472.5 71707.5 207607.5 ;
      RECT  71832.5 207472.5 71897.5 207607.5 ;
      RECT  71832.5 207472.5 71897.5 207607.5 ;
      RECT  71642.5 207472.5 71707.5 207607.5 ;
      RECT  71832.5 207472.5 71897.5 207607.5 ;
      RECT  72022.5 207472.5 72087.5 207607.5 ;
      RECT  72022.5 207472.5 72087.5 207607.5 ;
      RECT  71832.5 207472.5 71897.5 207607.5 ;
      RECT  71812.5 207237.5 71677.5 207302.5 ;
      RECT  71832.5 207785.0 71897.5 207920.0 ;
      RECT  71642.5 206942.5 71707.5 207077.5 ;
      RECT  71832.5 206942.5 71897.5 207077.5 ;
      RECT  71642.5 207472.5 71707.5 207607.5 ;
      RECT  72022.5 207472.5 72087.5 207607.5 ;
      RECT  71480.0 207237.5 72185.0 207302.5 ;
      RECT  71480.0 207922.5 72185.0 207987.5 ;
      RECT  72537.5 207472.5 72602.5 207987.5 ;
      RECT  72347.5 206942.5 72412.5 207077.5 ;
      RECT  72537.5 206942.5 72602.5 207077.5 ;
      RECT  72537.5 206942.5 72602.5 207077.5 ;
      RECT  72347.5 206942.5 72412.5 207077.5 ;
      RECT  72347.5 207472.5 72412.5 207607.5 ;
      RECT  72537.5 207472.5 72602.5 207607.5 ;
      RECT  72537.5 207472.5 72602.5 207607.5 ;
      RECT  72347.5 207472.5 72412.5 207607.5 ;
      RECT  72537.5 207472.5 72602.5 207607.5 ;
      RECT  72727.5 207472.5 72792.5 207607.5 ;
      RECT  72727.5 207472.5 72792.5 207607.5 ;
      RECT  72537.5 207472.5 72602.5 207607.5 ;
      RECT  72517.5 207237.5 72382.5 207302.5 ;
      RECT  72537.5 207785.0 72602.5 207920.0 ;
      RECT  72347.5 206942.5 72412.5 207077.5 ;
      RECT  72537.5 206942.5 72602.5 207077.5 ;
      RECT  72347.5 207472.5 72412.5 207607.5 ;
      RECT  72727.5 207472.5 72792.5 207607.5 ;
      RECT  72185.0 207237.5 72890.0 207302.5 ;
      RECT  72185.0 207922.5 72890.0 207987.5 ;
      RECT  73242.5 207472.5 73307.5 207987.5 ;
      RECT  73052.5 206942.5 73117.5 207077.5 ;
      RECT  73242.5 206942.5 73307.5 207077.5 ;
      RECT  73242.5 206942.5 73307.5 207077.5 ;
      RECT  73052.5 206942.5 73117.5 207077.5 ;
      RECT  73052.5 207472.5 73117.5 207607.5 ;
      RECT  73242.5 207472.5 73307.5 207607.5 ;
      RECT  73242.5 207472.5 73307.5 207607.5 ;
      RECT  73052.5 207472.5 73117.5 207607.5 ;
      RECT  73242.5 207472.5 73307.5 207607.5 ;
      RECT  73432.5 207472.5 73497.5 207607.5 ;
      RECT  73432.5 207472.5 73497.5 207607.5 ;
      RECT  73242.5 207472.5 73307.5 207607.5 ;
      RECT  73222.5 207237.5 73087.5 207302.5 ;
      RECT  73242.5 207785.0 73307.5 207920.0 ;
      RECT  73052.5 206942.5 73117.5 207077.5 ;
      RECT  73242.5 206942.5 73307.5 207077.5 ;
      RECT  73052.5 207472.5 73117.5 207607.5 ;
      RECT  73432.5 207472.5 73497.5 207607.5 ;
      RECT  72890.0 207237.5 73595.0 207302.5 ;
      RECT  72890.0 207922.5 73595.0 207987.5 ;
      RECT  73947.5 207472.5 74012.5 207987.5 ;
      RECT  73757.5 206942.5 73822.5 207077.5 ;
      RECT  73947.5 206942.5 74012.5 207077.5 ;
      RECT  73947.5 206942.5 74012.5 207077.5 ;
      RECT  73757.5 206942.5 73822.5 207077.5 ;
      RECT  73757.5 207472.5 73822.5 207607.5 ;
      RECT  73947.5 207472.5 74012.5 207607.5 ;
      RECT  73947.5 207472.5 74012.5 207607.5 ;
      RECT  73757.5 207472.5 73822.5 207607.5 ;
      RECT  73947.5 207472.5 74012.5 207607.5 ;
      RECT  74137.5 207472.5 74202.5 207607.5 ;
      RECT  74137.5 207472.5 74202.5 207607.5 ;
      RECT  73947.5 207472.5 74012.5 207607.5 ;
      RECT  73927.5 207237.5 73792.5 207302.5 ;
      RECT  73947.5 207785.0 74012.5 207920.0 ;
      RECT  73757.5 206942.5 73822.5 207077.5 ;
      RECT  73947.5 206942.5 74012.5 207077.5 ;
      RECT  73757.5 207472.5 73822.5 207607.5 ;
      RECT  74137.5 207472.5 74202.5 207607.5 ;
      RECT  73595.0 207237.5 74300.0 207302.5 ;
      RECT  73595.0 207922.5 74300.0 207987.5 ;
      RECT  74652.5 207472.5 74717.5 207987.5 ;
      RECT  74462.5 206942.5 74527.5 207077.5 ;
      RECT  74652.5 206942.5 74717.5 207077.5 ;
      RECT  74652.5 206942.5 74717.5 207077.5 ;
      RECT  74462.5 206942.5 74527.5 207077.5 ;
      RECT  74462.5 207472.5 74527.5 207607.5 ;
      RECT  74652.5 207472.5 74717.5 207607.5 ;
      RECT  74652.5 207472.5 74717.5 207607.5 ;
      RECT  74462.5 207472.5 74527.5 207607.5 ;
      RECT  74652.5 207472.5 74717.5 207607.5 ;
      RECT  74842.5 207472.5 74907.5 207607.5 ;
      RECT  74842.5 207472.5 74907.5 207607.5 ;
      RECT  74652.5 207472.5 74717.5 207607.5 ;
      RECT  74632.5 207237.5 74497.5 207302.5 ;
      RECT  74652.5 207785.0 74717.5 207920.0 ;
      RECT  74462.5 206942.5 74527.5 207077.5 ;
      RECT  74652.5 206942.5 74717.5 207077.5 ;
      RECT  74462.5 207472.5 74527.5 207607.5 ;
      RECT  74842.5 207472.5 74907.5 207607.5 ;
      RECT  74300.0 207237.5 75005.0 207302.5 ;
      RECT  74300.0 207922.5 75005.0 207987.5 ;
      RECT  75357.5 207472.5 75422.5 207987.5 ;
      RECT  75167.5 206942.5 75232.5 207077.5 ;
      RECT  75357.5 206942.5 75422.5 207077.5 ;
      RECT  75357.5 206942.5 75422.5 207077.5 ;
      RECT  75167.5 206942.5 75232.5 207077.5 ;
      RECT  75167.5 207472.5 75232.5 207607.5 ;
      RECT  75357.5 207472.5 75422.5 207607.5 ;
      RECT  75357.5 207472.5 75422.5 207607.5 ;
      RECT  75167.5 207472.5 75232.5 207607.5 ;
      RECT  75357.5 207472.5 75422.5 207607.5 ;
      RECT  75547.5 207472.5 75612.5 207607.5 ;
      RECT  75547.5 207472.5 75612.5 207607.5 ;
      RECT  75357.5 207472.5 75422.5 207607.5 ;
      RECT  75337.5 207237.5 75202.5 207302.5 ;
      RECT  75357.5 207785.0 75422.5 207920.0 ;
      RECT  75167.5 206942.5 75232.5 207077.5 ;
      RECT  75357.5 206942.5 75422.5 207077.5 ;
      RECT  75167.5 207472.5 75232.5 207607.5 ;
      RECT  75547.5 207472.5 75612.5 207607.5 ;
      RECT  75005.0 207237.5 75710.0 207302.5 ;
      RECT  75005.0 207922.5 75710.0 207987.5 ;
      RECT  76062.5 207472.5 76127.5 207987.5 ;
      RECT  75872.5 206942.5 75937.5 207077.5 ;
      RECT  76062.5 206942.5 76127.5 207077.5 ;
      RECT  76062.5 206942.5 76127.5 207077.5 ;
      RECT  75872.5 206942.5 75937.5 207077.5 ;
      RECT  75872.5 207472.5 75937.5 207607.5 ;
      RECT  76062.5 207472.5 76127.5 207607.5 ;
      RECT  76062.5 207472.5 76127.5 207607.5 ;
      RECT  75872.5 207472.5 75937.5 207607.5 ;
      RECT  76062.5 207472.5 76127.5 207607.5 ;
      RECT  76252.5 207472.5 76317.5 207607.5 ;
      RECT  76252.5 207472.5 76317.5 207607.5 ;
      RECT  76062.5 207472.5 76127.5 207607.5 ;
      RECT  76042.5 207237.5 75907.5 207302.5 ;
      RECT  76062.5 207785.0 76127.5 207920.0 ;
      RECT  75872.5 206942.5 75937.5 207077.5 ;
      RECT  76062.5 206942.5 76127.5 207077.5 ;
      RECT  75872.5 207472.5 75937.5 207607.5 ;
      RECT  76252.5 207472.5 76317.5 207607.5 ;
      RECT  75710.0 207237.5 76415.0 207302.5 ;
      RECT  75710.0 207922.5 76415.0 207987.5 ;
      RECT  76767.5 207472.5 76832.5 207987.5 ;
      RECT  76577.5 206942.5 76642.5 207077.5 ;
      RECT  76767.5 206942.5 76832.5 207077.5 ;
      RECT  76767.5 206942.5 76832.5 207077.5 ;
      RECT  76577.5 206942.5 76642.5 207077.5 ;
      RECT  76577.5 207472.5 76642.5 207607.5 ;
      RECT  76767.5 207472.5 76832.5 207607.5 ;
      RECT  76767.5 207472.5 76832.5 207607.5 ;
      RECT  76577.5 207472.5 76642.5 207607.5 ;
      RECT  76767.5 207472.5 76832.5 207607.5 ;
      RECT  76957.5 207472.5 77022.5 207607.5 ;
      RECT  76957.5 207472.5 77022.5 207607.5 ;
      RECT  76767.5 207472.5 76832.5 207607.5 ;
      RECT  76747.5 207237.5 76612.5 207302.5 ;
      RECT  76767.5 207785.0 76832.5 207920.0 ;
      RECT  76577.5 206942.5 76642.5 207077.5 ;
      RECT  76767.5 206942.5 76832.5 207077.5 ;
      RECT  76577.5 207472.5 76642.5 207607.5 ;
      RECT  76957.5 207472.5 77022.5 207607.5 ;
      RECT  76415.0 207237.5 77120.0 207302.5 ;
      RECT  76415.0 207922.5 77120.0 207987.5 ;
      RECT  77472.5 207472.5 77537.5 207987.5 ;
      RECT  77282.5 206942.5 77347.5 207077.5 ;
      RECT  77472.5 206942.5 77537.5 207077.5 ;
      RECT  77472.5 206942.5 77537.5 207077.5 ;
      RECT  77282.5 206942.5 77347.5 207077.5 ;
      RECT  77282.5 207472.5 77347.5 207607.5 ;
      RECT  77472.5 207472.5 77537.5 207607.5 ;
      RECT  77472.5 207472.5 77537.5 207607.5 ;
      RECT  77282.5 207472.5 77347.5 207607.5 ;
      RECT  77472.5 207472.5 77537.5 207607.5 ;
      RECT  77662.5 207472.5 77727.5 207607.5 ;
      RECT  77662.5 207472.5 77727.5 207607.5 ;
      RECT  77472.5 207472.5 77537.5 207607.5 ;
      RECT  77452.5 207237.5 77317.5 207302.5 ;
      RECT  77472.5 207785.0 77537.5 207920.0 ;
      RECT  77282.5 206942.5 77347.5 207077.5 ;
      RECT  77472.5 206942.5 77537.5 207077.5 ;
      RECT  77282.5 207472.5 77347.5 207607.5 ;
      RECT  77662.5 207472.5 77727.5 207607.5 ;
      RECT  77120.0 207237.5 77825.0 207302.5 ;
      RECT  77120.0 207922.5 77825.0 207987.5 ;
      RECT  78177.5 207472.5 78242.5 207987.5 ;
      RECT  77987.5 206942.5 78052.5 207077.5 ;
      RECT  78177.5 206942.5 78242.5 207077.5 ;
      RECT  78177.5 206942.5 78242.5 207077.5 ;
      RECT  77987.5 206942.5 78052.5 207077.5 ;
      RECT  77987.5 207472.5 78052.5 207607.5 ;
      RECT  78177.5 207472.5 78242.5 207607.5 ;
      RECT  78177.5 207472.5 78242.5 207607.5 ;
      RECT  77987.5 207472.5 78052.5 207607.5 ;
      RECT  78177.5 207472.5 78242.5 207607.5 ;
      RECT  78367.5 207472.5 78432.5 207607.5 ;
      RECT  78367.5 207472.5 78432.5 207607.5 ;
      RECT  78177.5 207472.5 78242.5 207607.5 ;
      RECT  78157.5 207237.5 78022.5 207302.5 ;
      RECT  78177.5 207785.0 78242.5 207920.0 ;
      RECT  77987.5 206942.5 78052.5 207077.5 ;
      RECT  78177.5 206942.5 78242.5 207077.5 ;
      RECT  77987.5 207472.5 78052.5 207607.5 ;
      RECT  78367.5 207472.5 78432.5 207607.5 ;
      RECT  77825.0 207237.5 78530.0 207302.5 ;
      RECT  77825.0 207922.5 78530.0 207987.5 ;
      RECT  78882.5 207472.5 78947.5 207987.5 ;
      RECT  78692.5 206942.5 78757.5 207077.5 ;
      RECT  78882.5 206942.5 78947.5 207077.5 ;
      RECT  78882.5 206942.5 78947.5 207077.5 ;
      RECT  78692.5 206942.5 78757.5 207077.5 ;
      RECT  78692.5 207472.5 78757.5 207607.5 ;
      RECT  78882.5 207472.5 78947.5 207607.5 ;
      RECT  78882.5 207472.5 78947.5 207607.5 ;
      RECT  78692.5 207472.5 78757.5 207607.5 ;
      RECT  78882.5 207472.5 78947.5 207607.5 ;
      RECT  79072.5 207472.5 79137.5 207607.5 ;
      RECT  79072.5 207472.5 79137.5 207607.5 ;
      RECT  78882.5 207472.5 78947.5 207607.5 ;
      RECT  78862.5 207237.5 78727.5 207302.5 ;
      RECT  78882.5 207785.0 78947.5 207920.0 ;
      RECT  78692.5 206942.5 78757.5 207077.5 ;
      RECT  78882.5 206942.5 78947.5 207077.5 ;
      RECT  78692.5 207472.5 78757.5 207607.5 ;
      RECT  79072.5 207472.5 79137.5 207607.5 ;
      RECT  78530.0 207237.5 79235.0 207302.5 ;
      RECT  78530.0 207922.5 79235.0 207987.5 ;
      RECT  79587.5 207472.5 79652.5 207987.5 ;
      RECT  79397.5 206942.5 79462.5 207077.5 ;
      RECT  79587.5 206942.5 79652.5 207077.5 ;
      RECT  79587.5 206942.5 79652.5 207077.5 ;
      RECT  79397.5 206942.5 79462.5 207077.5 ;
      RECT  79397.5 207472.5 79462.5 207607.5 ;
      RECT  79587.5 207472.5 79652.5 207607.5 ;
      RECT  79587.5 207472.5 79652.5 207607.5 ;
      RECT  79397.5 207472.5 79462.5 207607.5 ;
      RECT  79587.5 207472.5 79652.5 207607.5 ;
      RECT  79777.5 207472.5 79842.5 207607.5 ;
      RECT  79777.5 207472.5 79842.5 207607.5 ;
      RECT  79587.5 207472.5 79652.5 207607.5 ;
      RECT  79567.5 207237.5 79432.5 207302.5 ;
      RECT  79587.5 207785.0 79652.5 207920.0 ;
      RECT  79397.5 206942.5 79462.5 207077.5 ;
      RECT  79587.5 206942.5 79652.5 207077.5 ;
      RECT  79397.5 207472.5 79462.5 207607.5 ;
      RECT  79777.5 207472.5 79842.5 207607.5 ;
      RECT  79235.0 207237.5 79940.0 207302.5 ;
      RECT  79235.0 207922.5 79940.0 207987.5 ;
      RECT  80292.5 207472.5 80357.5 207987.5 ;
      RECT  80102.5 206942.5 80167.5 207077.5 ;
      RECT  80292.5 206942.5 80357.5 207077.5 ;
      RECT  80292.5 206942.5 80357.5 207077.5 ;
      RECT  80102.5 206942.5 80167.5 207077.5 ;
      RECT  80102.5 207472.5 80167.5 207607.5 ;
      RECT  80292.5 207472.5 80357.5 207607.5 ;
      RECT  80292.5 207472.5 80357.5 207607.5 ;
      RECT  80102.5 207472.5 80167.5 207607.5 ;
      RECT  80292.5 207472.5 80357.5 207607.5 ;
      RECT  80482.5 207472.5 80547.5 207607.5 ;
      RECT  80482.5 207472.5 80547.5 207607.5 ;
      RECT  80292.5 207472.5 80357.5 207607.5 ;
      RECT  80272.5 207237.5 80137.5 207302.5 ;
      RECT  80292.5 207785.0 80357.5 207920.0 ;
      RECT  80102.5 206942.5 80167.5 207077.5 ;
      RECT  80292.5 206942.5 80357.5 207077.5 ;
      RECT  80102.5 207472.5 80167.5 207607.5 ;
      RECT  80482.5 207472.5 80547.5 207607.5 ;
      RECT  79940.0 207237.5 80645.0 207302.5 ;
      RECT  79940.0 207922.5 80645.0 207987.5 ;
      RECT  80997.5 207472.5 81062.5 207987.5 ;
      RECT  80807.5 206942.5 80872.5 207077.5 ;
      RECT  80997.5 206942.5 81062.5 207077.5 ;
      RECT  80997.5 206942.5 81062.5 207077.5 ;
      RECT  80807.5 206942.5 80872.5 207077.5 ;
      RECT  80807.5 207472.5 80872.5 207607.5 ;
      RECT  80997.5 207472.5 81062.5 207607.5 ;
      RECT  80997.5 207472.5 81062.5 207607.5 ;
      RECT  80807.5 207472.5 80872.5 207607.5 ;
      RECT  80997.5 207472.5 81062.5 207607.5 ;
      RECT  81187.5 207472.5 81252.5 207607.5 ;
      RECT  81187.5 207472.5 81252.5 207607.5 ;
      RECT  80997.5 207472.5 81062.5 207607.5 ;
      RECT  80977.5 207237.5 80842.5 207302.5 ;
      RECT  80997.5 207785.0 81062.5 207920.0 ;
      RECT  80807.5 206942.5 80872.5 207077.5 ;
      RECT  80997.5 206942.5 81062.5 207077.5 ;
      RECT  80807.5 207472.5 80872.5 207607.5 ;
      RECT  81187.5 207472.5 81252.5 207607.5 ;
      RECT  80645.0 207237.5 81350.0 207302.5 ;
      RECT  80645.0 207922.5 81350.0 207987.5 ;
      RECT  81702.5 207472.5 81767.5 207987.5 ;
      RECT  81512.5 206942.5 81577.5 207077.5 ;
      RECT  81702.5 206942.5 81767.5 207077.5 ;
      RECT  81702.5 206942.5 81767.5 207077.5 ;
      RECT  81512.5 206942.5 81577.5 207077.5 ;
      RECT  81512.5 207472.5 81577.5 207607.5 ;
      RECT  81702.5 207472.5 81767.5 207607.5 ;
      RECT  81702.5 207472.5 81767.5 207607.5 ;
      RECT  81512.5 207472.5 81577.5 207607.5 ;
      RECT  81702.5 207472.5 81767.5 207607.5 ;
      RECT  81892.5 207472.5 81957.5 207607.5 ;
      RECT  81892.5 207472.5 81957.5 207607.5 ;
      RECT  81702.5 207472.5 81767.5 207607.5 ;
      RECT  81682.5 207237.5 81547.5 207302.5 ;
      RECT  81702.5 207785.0 81767.5 207920.0 ;
      RECT  81512.5 206942.5 81577.5 207077.5 ;
      RECT  81702.5 206942.5 81767.5 207077.5 ;
      RECT  81512.5 207472.5 81577.5 207607.5 ;
      RECT  81892.5 207472.5 81957.5 207607.5 ;
      RECT  81350.0 207237.5 82055.0 207302.5 ;
      RECT  81350.0 207922.5 82055.0 207987.5 ;
      RECT  82407.5 207472.5 82472.5 207987.5 ;
      RECT  82217.5 206942.5 82282.5 207077.5 ;
      RECT  82407.5 206942.5 82472.5 207077.5 ;
      RECT  82407.5 206942.5 82472.5 207077.5 ;
      RECT  82217.5 206942.5 82282.5 207077.5 ;
      RECT  82217.5 207472.5 82282.5 207607.5 ;
      RECT  82407.5 207472.5 82472.5 207607.5 ;
      RECT  82407.5 207472.5 82472.5 207607.5 ;
      RECT  82217.5 207472.5 82282.5 207607.5 ;
      RECT  82407.5 207472.5 82472.5 207607.5 ;
      RECT  82597.5 207472.5 82662.5 207607.5 ;
      RECT  82597.5 207472.5 82662.5 207607.5 ;
      RECT  82407.5 207472.5 82472.5 207607.5 ;
      RECT  82387.5 207237.5 82252.5 207302.5 ;
      RECT  82407.5 207785.0 82472.5 207920.0 ;
      RECT  82217.5 206942.5 82282.5 207077.5 ;
      RECT  82407.5 206942.5 82472.5 207077.5 ;
      RECT  82217.5 207472.5 82282.5 207607.5 ;
      RECT  82597.5 207472.5 82662.5 207607.5 ;
      RECT  82055.0 207237.5 82760.0 207302.5 ;
      RECT  82055.0 207922.5 82760.0 207987.5 ;
      RECT  83112.5 207472.5 83177.5 207987.5 ;
      RECT  82922.5 206942.5 82987.5 207077.5 ;
      RECT  83112.5 206942.5 83177.5 207077.5 ;
      RECT  83112.5 206942.5 83177.5 207077.5 ;
      RECT  82922.5 206942.5 82987.5 207077.5 ;
      RECT  82922.5 207472.5 82987.5 207607.5 ;
      RECT  83112.5 207472.5 83177.5 207607.5 ;
      RECT  83112.5 207472.5 83177.5 207607.5 ;
      RECT  82922.5 207472.5 82987.5 207607.5 ;
      RECT  83112.5 207472.5 83177.5 207607.5 ;
      RECT  83302.5 207472.5 83367.5 207607.5 ;
      RECT  83302.5 207472.5 83367.5 207607.5 ;
      RECT  83112.5 207472.5 83177.5 207607.5 ;
      RECT  83092.5 207237.5 82957.5 207302.5 ;
      RECT  83112.5 207785.0 83177.5 207920.0 ;
      RECT  82922.5 206942.5 82987.5 207077.5 ;
      RECT  83112.5 206942.5 83177.5 207077.5 ;
      RECT  82922.5 207472.5 82987.5 207607.5 ;
      RECT  83302.5 207472.5 83367.5 207607.5 ;
      RECT  82760.0 207237.5 83465.0 207302.5 ;
      RECT  82760.0 207922.5 83465.0 207987.5 ;
      RECT  83817.5 207472.5 83882.5 207987.5 ;
      RECT  83627.5 206942.5 83692.5 207077.5 ;
      RECT  83817.5 206942.5 83882.5 207077.5 ;
      RECT  83817.5 206942.5 83882.5 207077.5 ;
      RECT  83627.5 206942.5 83692.5 207077.5 ;
      RECT  83627.5 207472.5 83692.5 207607.5 ;
      RECT  83817.5 207472.5 83882.5 207607.5 ;
      RECT  83817.5 207472.5 83882.5 207607.5 ;
      RECT  83627.5 207472.5 83692.5 207607.5 ;
      RECT  83817.5 207472.5 83882.5 207607.5 ;
      RECT  84007.5 207472.5 84072.5 207607.5 ;
      RECT  84007.5 207472.5 84072.5 207607.5 ;
      RECT  83817.5 207472.5 83882.5 207607.5 ;
      RECT  83797.5 207237.5 83662.5 207302.5 ;
      RECT  83817.5 207785.0 83882.5 207920.0 ;
      RECT  83627.5 206942.5 83692.5 207077.5 ;
      RECT  83817.5 206942.5 83882.5 207077.5 ;
      RECT  83627.5 207472.5 83692.5 207607.5 ;
      RECT  84007.5 207472.5 84072.5 207607.5 ;
      RECT  83465.0 207237.5 84170.0 207302.5 ;
      RECT  83465.0 207922.5 84170.0 207987.5 ;
      RECT  84522.5 207472.5 84587.5 207987.5 ;
      RECT  84332.5 206942.5 84397.5 207077.5 ;
      RECT  84522.5 206942.5 84587.5 207077.5 ;
      RECT  84522.5 206942.5 84587.5 207077.5 ;
      RECT  84332.5 206942.5 84397.5 207077.5 ;
      RECT  84332.5 207472.5 84397.5 207607.5 ;
      RECT  84522.5 207472.5 84587.5 207607.5 ;
      RECT  84522.5 207472.5 84587.5 207607.5 ;
      RECT  84332.5 207472.5 84397.5 207607.5 ;
      RECT  84522.5 207472.5 84587.5 207607.5 ;
      RECT  84712.5 207472.5 84777.5 207607.5 ;
      RECT  84712.5 207472.5 84777.5 207607.5 ;
      RECT  84522.5 207472.5 84587.5 207607.5 ;
      RECT  84502.5 207237.5 84367.5 207302.5 ;
      RECT  84522.5 207785.0 84587.5 207920.0 ;
      RECT  84332.5 206942.5 84397.5 207077.5 ;
      RECT  84522.5 206942.5 84587.5 207077.5 ;
      RECT  84332.5 207472.5 84397.5 207607.5 ;
      RECT  84712.5 207472.5 84777.5 207607.5 ;
      RECT  84170.0 207237.5 84875.0 207302.5 ;
      RECT  84170.0 207922.5 84875.0 207987.5 ;
      RECT  85227.5 207472.5 85292.5 207987.5 ;
      RECT  85037.5 206942.5 85102.5 207077.5 ;
      RECT  85227.5 206942.5 85292.5 207077.5 ;
      RECT  85227.5 206942.5 85292.5 207077.5 ;
      RECT  85037.5 206942.5 85102.5 207077.5 ;
      RECT  85037.5 207472.5 85102.5 207607.5 ;
      RECT  85227.5 207472.5 85292.5 207607.5 ;
      RECT  85227.5 207472.5 85292.5 207607.5 ;
      RECT  85037.5 207472.5 85102.5 207607.5 ;
      RECT  85227.5 207472.5 85292.5 207607.5 ;
      RECT  85417.5 207472.5 85482.5 207607.5 ;
      RECT  85417.5 207472.5 85482.5 207607.5 ;
      RECT  85227.5 207472.5 85292.5 207607.5 ;
      RECT  85207.5 207237.5 85072.5 207302.5 ;
      RECT  85227.5 207785.0 85292.5 207920.0 ;
      RECT  85037.5 206942.5 85102.5 207077.5 ;
      RECT  85227.5 206942.5 85292.5 207077.5 ;
      RECT  85037.5 207472.5 85102.5 207607.5 ;
      RECT  85417.5 207472.5 85482.5 207607.5 ;
      RECT  84875.0 207237.5 85580.0 207302.5 ;
      RECT  84875.0 207922.5 85580.0 207987.5 ;
      RECT  85932.5 207472.5 85997.5 207987.5 ;
      RECT  85742.5 206942.5 85807.5 207077.5 ;
      RECT  85932.5 206942.5 85997.5 207077.5 ;
      RECT  85932.5 206942.5 85997.5 207077.5 ;
      RECT  85742.5 206942.5 85807.5 207077.5 ;
      RECT  85742.5 207472.5 85807.5 207607.5 ;
      RECT  85932.5 207472.5 85997.5 207607.5 ;
      RECT  85932.5 207472.5 85997.5 207607.5 ;
      RECT  85742.5 207472.5 85807.5 207607.5 ;
      RECT  85932.5 207472.5 85997.5 207607.5 ;
      RECT  86122.5 207472.5 86187.5 207607.5 ;
      RECT  86122.5 207472.5 86187.5 207607.5 ;
      RECT  85932.5 207472.5 85997.5 207607.5 ;
      RECT  85912.5 207237.5 85777.5 207302.5 ;
      RECT  85932.5 207785.0 85997.5 207920.0 ;
      RECT  85742.5 206942.5 85807.5 207077.5 ;
      RECT  85932.5 206942.5 85997.5 207077.5 ;
      RECT  85742.5 207472.5 85807.5 207607.5 ;
      RECT  86122.5 207472.5 86187.5 207607.5 ;
      RECT  85580.0 207237.5 86285.0 207302.5 ;
      RECT  85580.0 207922.5 86285.0 207987.5 ;
      RECT  86637.5 207472.5 86702.5 207987.5 ;
      RECT  86447.5 206942.5 86512.5 207077.5 ;
      RECT  86637.5 206942.5 86702.5 207077.5 ;
      RECT  86637.5 206942.5 86702.5 207077.5 ;
      RECT  86447.5 206942.5 86512.5 207077.5 ;
      RECT  86447.5 207472.5 86512.5 207607.5 ;
      RECT  86637.5 207472.5 86702.5 207607.5 ;
      RECT  86637.5 207472.5 86702.5 207607.5 ;
      RECT  86447.5 207472.5 86512.5 207607.5 ;
      RECT  86637.5 207472.5 86702.5 207607.5 ;
      RECT  86827.5 207472.5 86892.5 207607.5 ;
      RECT  86827.5 207472.5 86892.5 207607.5 ;
      RECT  86637.5 207472.5 86702.5 207607.5 ;
      RECT  86617.5 207237.5 86482.5 207302.5 ;
      RECT  86637.5 207785.0 86702.5 207920.0 ;
      RECT  86447.5 206942.5 86512.5 207077.5 ;
      RECT  86637.5 206942.5 86702.5 207077.5 ;
      RECT  86447.5 207472.5 86512.5 207607.5 ;
      RECT  86827.5 207472.5 86892.5 207607.5 ;
      RECT  86285.0 207237.5 86990.0 207302.5 ;
      RECT  86285.0 207922.5 86990.0 207987.5 ;
      RECT  87342.5 207472.5 87407.5 207987.5 ;
      RECT  87152.5 206942.5 87217.5 207077.5 ;
      RECT  87342.5 206942.5 87407.5 207077.5 ;
      RECT  87342.5 206942.5 87407.5 207077.5 ;
      RECT  87152.5 206942.5 87217.5 207077.5 ;
      RECT  87152.5 207472.5 87217.5 207607.5 ;
      RECT  87342.5 207472.5 87407.5 207607.5 ;
      RECT  87342.5 207472.5 87407.5 207607.5 ;
      RECT  87152.5 207472.5 87217.5 207607.5 ;
      RECT  87342.5 207472.5 87407.5 207607.5 ;
      RECT  87532.5 207472.5 87597.5 207607.5 ;
      RECT  87532.5 207472.5 87597.5 207607.5 ;
      RECT  87342.5 207472.5 87407.5 207607.5 ;
      RECT  87322.5 207237.5 87187.5 207302.5 ;
      RECT  87342.5 207785.0 87407.5 207920.0 ;
      RECT  87152.5 206942.5 87217.5 207077.5 ;
      RECT  87342.5 206942.5 87407.5 207077.5 ;
      RECT  87152.5 207472.5 87217.5 207607.5 ;
      RECT  87532.5 207472.5 87597.5 207607.5 ;
      RECT  86990.0 207237.5 87695.0 207302.5 ;
      RECT  86990.0 207922.5 87695.0 207987.5 ;
      RECT  88047.5 207472.5 88112.5 207987.5 ;
      RECT  87857.5 206942.5 87922.5 207077.5 ;
      RECT  88047.5 206942.5 88112.5 207077.5 ;
      RECT  88047.5 206942.5 88112.5 207077.5 ;
      RECT  87857.5 206942.5 87922.5 207077.5 ;
      RECT  87857.5 207472.5 87922.5 207607.5 ;
      RECT  88047.5 207472.5 88112.5 207607.5 ;
      RECT  88047.5 207472.5 88112.5 207607.5 ;
      RECT  87857.5 207472.5 87922.5 207607.5 ;
      RECT  88047.5 207472.5 88112.5 207607.5 ;
      RECT  88237.5 207472.5 88302.5 207607.5 ;
      RECT  88237.5 207472.5 88302.5 207607.5 ;
      RECT  88047.5 207472.5 88112.5 207607.5 ;
      RECT  88027.5 207237.5 87892.5 207302.5 ;
      RECT  88047.5 207785.0 88112.5 207920.0 ;
      RECT  87857.5 206942.5 87922.5 207077.5 ;
      RECT  88047.5 206942.5 88112.5 207077.5 ;
      RECT  87857.5 207472.5 87922.5 207607.5 ;
      RECT  88237.5 207472.5 88302.5 207607.5 ;
      RECT  87695.0 207237.5 88400.0 207302.5 ;
      RECT  87695.0 207922.5 88400.0 207987.5 ;
      RECT  88752.5 207472.5 88817.5 207987.5 ;
      RECT  88562.5 206942.5 88627.5 207077.5 ;
      RECT  88752.5 206942.5 88817.5 207077.5 ;
      RECT  88752.5 206942.5 88817.5 207077.5 ;
      RECT  88562.5 206942.5 88627.5 207077.5 ;
      RECT  88562.5 207472.5 88627.5 207607.5 ;
      RECT  88752.5 207472.5 88817.5 207607.5 ;
      RECT  88752.5 207472.5 88817.5 207607.5 ;
      RECT  88562.5 207472.5 88627.5 207607.5 ;
      RECT  88752.5 207472.5 88817.5 207607.5 ;
      RECT  88942.5 207472.5 89007.5 207607.5 ;
      RECT  88942.5 207472.5 89007.5 207607.5 ;
      RECT  88752.5 207472.5 88817.5 207607.5 ;
      RECT  88732.5 207237.5 88597.5 207302.5 ;
      RECT  88752.5 207785.0 88817.5 207920.0 ;
      RECT  88562.5 206942.5 88627.5 207077.5 ;
      RECT  88752.5 206942.5 88817.5 207077.5 ;
      RECT  88562.5 207472.5 88627.5 207607.5 ;
      RECT  88942.5 207472.5 89007.5 207607.5 ;
      RECT  88400.0 207237.5 89105.0 207302.5 ;
      RECT  88400.0 207922.5 89105.0 207987.5 ;
      RECT  89457.5 207472.5 89522.5 207987.5 ;
      RECT  89267.5 206942.5 89332.5 207077.5 ;
      RECT  89457.5 206942.5 89522.5 207077.5 ;
      RECT  89457.5 206942.5 89522.5 207077.5 ;
      RECT  89267.5 206942.5 89332.5 207077.5 ;
      RECT  89267.5 207472.5 89332.5 207607.5 ;
      RECT  89457.5 207472.5 89522.5 207607.5 ;
      RECT  89457.5 207472.5 89522.5 207607.5 ;
      RECT  89267.5 207472.5 89332.5 207607.5 ;
      RECT  89457.5 207472.5 89522.5 207607.5 ;
      RECT  89647.5 207472.5 89712.5 207607.5 ;
      RECT  89647.5 207472.5 89712.5 207607.5 ;
      RECT  89457.5 207472.5 89522.5 207607.5 ;
      RECT  89437.5 207237.5 89302.5 207302.5 ;
      RECT  89457.5 207785.0 89522.5 207920.0 ;
      RECT  89267.5 206942.5 89332.5 207077.5 ;
      RECT  89457.5 206942.5 89522.5 207077.5 ;
      RECT  89267.5 207472.5 89332.5 207607.5 ;
      RECT  89647.5 207472.5 89712.5 207607.5 ;
      RECT  89105.0 207237.5 89810.0 207302.5 ;
      RECT  89105.0 207922.5 89810.0 207987.5 ;
      RECT  90162.5 207472.5 90227.5 207987.5 ;
      RECT  89972.5 206942.5 90037.5 207077.5 ;
      RECT  90162.5 206942.5 90227.5 207077.5 ;
      RECT  90162.5 206942.5 90227.5 207077.5 ;
      RECT  89972.5 206942.5 90037.5 207077.5 ;
      RECT  89972.5 207472.5 90037.5 207607.5 ;
      RECT  90162.5 207472.5 90227.5 207607.5 ;
      RECT  90162.5 207472.5 90227.5 207607.5 ;
      RECT  89972.5 207472.5 90037.5 207607.5 ;
      RECT  90162.5 207472.5 90227.5 207607.5 ;
      RECT  90352.5 207472.5 90417.5 207607.5 ;
      RECT  90352.5 207472.5 90417.5 207607.5 ;
      RECT  90162.5 207472.5 90227.5 207607.5 ;
      RECT  90142.5 207237.5 90007.5 207302.5 ;
      RECT  90162.5 207785.0 90227.5 207920.0 ;
      RECT  89972.5 206942.5 90037.5 207077.5 ;
      RECT  90162.5 206942.5 90227.5 207077.5 ;
      RECT  89972.5 207472.5 90037.5 207607.5 ;
      RECT  90352.5 207472.5 90417.5 207607.5 ;
      RECT  89810.0 207237.5 90515.0 207302.5 ;
      RECT  89810.0 207922.5 90515.0 207987.5 ;
      RECT  90867.5 207472.5 90932.5 207987.5 ;
      RECT  90677.5 206942.5 90742.5 207077.5 ;
      RECT  90867.5 206942.5 90932.5 207077.5 ;
      RECT  90867.5 206942.5 90932.5 207077.5 ;
      RECT  90677.5 206942.5 90742.5 207077.5 ;
      RECT  90677.5 207472.5 90742.5 207607.5 ;
      RECT  90867.5 207472.5 90932.5 207607.5 ;
      RECT  90867.5 207472.5 90932.5 207607.5 ;
      RECT  90677.5 207472.5 90742.5 207607.5 ;
      RECT  90867.5 207472.5 90932.5 207607.5 ;
      RECT  91057.5 207472.5 91122.5 207607.5 ;
      RECT  91057.5 207472.5 91122.5 207607.5 ;
      RECT  90867.5 207472.5 90932.5 207607.5 ;
      RECT  90847.5 207237.5 90712.5 207302.5 ;
      RECT  90867.5 207785.0 90932.5 207920.0 ;
      RECT  90677.5 206942.5 90742.5 207077.5 ;
      RECT  90867.5 206942.5 90932.5 207077.5 ;
      RECT  90677.5 207472.5 90742.5 207607.5 ;
      RECT  91057.5 207472.5 91122.5 207607.5 ;
      RECT  90515.0 207237.5 91220.0 207302.5 ;
      RECT  90515.0 207922.5 91220.0 207987.5 ;
      RECT  91572.5 207472.5 91637.5 207987.5 ;
      RECT  91382.5 206942.5 91447.5 207077.5 ;
      RECT  91572.5 206942.5 91637.5 207077.5 ;
      RECT  91572.5 206942.5 91637.5 207077.5 ;
      RECT  91382.5 206942.5 91447.5 207077.5 ;
      RECT  91382.5 207472.5 91447.5 207607.5 ;
      RECT  91572.5 207472.5 91637.5 207607.5 ;
      RECT  91572.5 207472.5 91637.5 207607.5 ;
      RECT  91382.5 207472.5 91447.5 207607.5 ;
      RECT  91572.5 207472.5 91637.5 207607.5 ;
      RECT  91762.5 207472.5 91827.5 207607.5 ;
      RECT  91762.5 207472.5 91827.5 207607.5 ;
      RECT  91572.5 207472.5 91637.5 207607.5 ;
      RECT  91552.5 207237.5 91417.5 207302.5 ;
      RECT  91572.5 207785.0 91637.5 207920.0 ;
      RECT  91382.5 206942.5 91447.5 207077.5 ;
      RECT  91572.5 206942.5 91637.5 207077.5 ;
      RECT  91382.5 207472.5 91447.5 207607.5 ;
      RECT  91762.5 207472.5 91827.5 207607.5 ;
      RECT  91220.0 207237.5 91925.0 207302.5 ;
      RECT  91220.0 207922.5 91925.0 207987.5 ;
      RECT  92277.5 207472.5 92342.5 207987.5 ;
      RECT  92087.5 206942.5 92152.5 207077.5 ;
      RECT  92277.5 206942.5 92342.5 207077.5 ;
      RECT  92277.5 206942.5 92342.5 207077.5 ;
      RECT  92087.5 206942.5 92152.5 207077.5 ;
      RECT  92087.5 207472.5 92152.5 207607.5 ;
      RECT  92277.5 207472.5 92342.5 207607.5 ;
      RECT  92277.5 207472.5 92342.5 207607.5 ;
      RECT  92087.5 207472.5 92152.5 207607.5 ;
      RECT  92277.5 207472.5 92342.5 207607.5 ;
      RECT  92467.5 207472.5 92532.5 207607.5 ;
      RECT  92467.5 207472.5 92532.5 207607.5 ;
      RECT  92277.5 207472.5 92342.5 207607.5 ;
      RECT  92257.5 207237.5 92122.5 207302.5 ;
      RECT  92277.5 207785.0 92342.5 207920.0 ;
      RECT  92087.5 206942.5 92152.5 207077.5 ;
      RECT  92277.5 206942.5 92342.5 207077.5 ;
      RECT  92087.5 207472.5 92152.5 207607.5 ;
      RECT  92467.5 207472.5 92532.5 207607.5 ;
      RECT  91925.0 207237.5 92630.0 207302.5 ;
      RECT  91925.0 207922.5 92630.0 207987.5 ;
      RECT  92982.5 207472.5 93047.5 207987.5 ;
      RECT  92792.5 206942.5 92857.5 207077.5 ;
      RECT  92982.5 206942.5 93047.5 207077.5 ;
      RECT  92982.5 206942.5 93047.5 207077.5 ;
      RECT  92792.5 206942.5 92857.5 207077.5 ;
      RECT  92792.5 207472.5 92857.5 207607.5 ;
      RECT  92982.5 207472.5 93047.5 207607.5 ;
      RECT  92982.5 207472.5 93047.5 207607.5 ;
      RECT  92792.5 207472.5 92857.5 207607.5 ;
      RECT  92982.5 207472.5 93047.5 207607.5 ;
      RECT  93172.5 207472.5 93237.5 207607.5 ;
      RECT  93172.5 207472.5 93237.5 207607.5 ;
      RECT  92982.5 207472.5 93047.5 207607.5 ;
      RECT  92962.5 207237.5 92827.5 207302.5 ;
      RECT  92982.5 207785.0 93047.5 207920.0 ;
      RECT  92792.5 206942.5 92857.5 207077.5 ;
      RECT  92982.5 206942.5 93047.5 207077.5 ;
      RECT  92792.5 207472.5 92857.5 207607.5 ;
      RECT  93172.5 207472.5 93237.5 207607.5 ;
      RECT  92630.0 207237.5 93335.0 207302.5 ;
      RECT  92630.0 207922.5 93335.0 207987.5 ;
      RECT  93687.5 207472.5 93752.5 207987.5 ;
      RECT  93497.5 206942.5 93562.5 207077.5 ;
      RECT  93687.5 206942.5 93752.5 207077.5 ;
      RECT  93687.5 206942.5 93752.5 207077.5 ;
      RECT  93497.5 206942.5 93562.5 207077.5 ;
      RECT  93497.5 207472.5 93562.5 207607.5 ;
      RECT  93687.5 207472.5 93752.5 207607.5 ;
      RECT  93687.5 207472.5 93752.5 207607.5 ;
      RECT  93497.5 207472.5 93562.5 207607.5 ;
      RECT  93687.5 207472.5 93752.5 207607.5 ;
      RECT  93877.5 207472.5 93942.5 207607.5 ;
      RECT  93877.5 207472.5 93942.5 207607.5 ;
      RECT  93687.5 207472.5 93752.5 207607.5 ;
      RECT  93667.5 207237.5 93532.5 207302.5 ;
      RECT  93687.5 207785.0 93752.5 207920.0 ;
      RECT  93497.5 206942.5 93562.5 207077.5 ;
      RECT  93687.5 206942.5 93752.5 207077.5 ;
      RECT  93497.5 207472.5 93562.5 207607.5 ;
      RECT  93877.5 207472.5 93942.5 207607.5 ;
      RECT  93335.0 207237.5 94040.0 207302.5 ;
      RECT  93335.0 207922.5 94040.0 207987.5 ;
      RECT  94392.5 207472.5 94457.5 207987.5 ;
      RECT  94202.5 206942.5 94267.5 207077.5 ;
      RECT  94392.5 206942.5 94457.5 207077.5 ;
      RECT  94392.5 206942.5 94457.5 207077.5 ;
      RECT  94202.5 206942.5 94267.5 207077.5 ;
      RECT  94202.5 207472.5 94267.5 207607.5 ;
      RECT  94392.5 207472.5 94457.5 207607.5 ;
      RECT  94392.5 207472.5 94457.5 207607.5 ;
      RECT  94202.5 207472.5 94267.5 207607.5 ;
      RECT  94392.5 207472.5 94457.5 207607.5 ;
      RECT  94582.5 207472.5 94647.5 207607.5 ;
      RECT  94582.5 207472.5 94647.5 207607.5 ;
      RECT  94392.5 207472.5 94457.5 207607.5 ;
      RECT  94372.5 207237.5 94237.5 207302.5 ;
      RECT  94392.5 207785.0 94457.5 207920.0 ;
      RECT  94202.5 206942.5 94267.5 207077.5 ;
      RECT  94392.5 206942.5 94457.5 207077.5 ;
      RECT  94202.5 207472.5 94267.5 207607.5 ;
      RECT  94582.5 207472.5 94647.5 207607.5 ;
      RECT  94040.0 207237.5 94745.0 207302.5 ;
      RECT  94040.0 207922.5 94745.0 207987.5 ;
      RECT  95097.5 207472.5 95162.5 207987.5 ;
      RECT  94907.5 206942.5 94972.5 207077.5 ;
      RECT  95097.5 206942.5 95162.5 207077.5 ;
      RECT  95097.5 206942.5 95162.5 207077.5 ;
      RECT  94907.5 206942.5 94972.5 207077.5 ;
      RECT  94907.5 207472.5 94972.5 207607.5 ;
      RECT  95097.5 207472.5 95162.5 207607.5 ;
      RECT  95097.5 207472.5 95162.5 207607.5 ;
      RECT  94907.5 207472.5 94972.5 207607.5 ;
      RECT  95097.5 207472.5 95162.5 207607.5 ;
      RECT  95287.5 207472.5 95352.5 207607.5 ;
      RECT  95287.5 207472.5 95352.5 207607.5 ;
      RECT  95097.5 207472.5 95162.5 207607.5 ;
      RECT  95077.5 207237.5 94942.5 207302.5 ;
      RECT  95097.5 207785.0 95162.5 207920.0 ;
      RECT  94907.5 206942.5 94972.5 207077.5 ;
      RECT  95097.5 206942.5 95162.5 207077.5 ;
      RECT  94907.5 207472.5 94972.5 207607.5 ;
      RECT  95287.5 207472.5 95352.5 207607.5 ;
      RECT  94745.0 207237.5 95450.0 207302.5 ;
      RECT  94745.0 207922.5 95450.0 207987.5 ;
      RECT  95802.5 207472.5 95867.5 207987.5 ;
      RECT  95612.5 206942.5 95677.5 207077.5 ;
      RECT  95802.5 206942.5 95867.5 207077.5 ;
      RECT  95802.5 206942.5 95867.5 207077.5 ;
      RECT  95612.5 206942.5 95677.5 207077.5 ;
      RECT  95612.5 207472.5 95677.5 207607.5 ;
      RECT  95802.5 207472.5 95867.5 207607.5 ;
      RECT  95802.5 207472.5 95867.5 207607.5 ;
      RECT  95612.5 207472.5 95677.5 207607.5 ;
      RECT  95802.5 207472.5 95867.5 207607.5 ;
      RECT  95992.5 207472.5 96057.5 207607.5 ;
      RECT  95992.5 207472.5 96057.5 207607.5 ;
      RECT  95802.5 207472.5 95867.5 207607.5 ;
      RECT  95782.5 207237.5 95647.5 207302.5 ;
      RECT  95802.5 207785.0 95867.5 207920.0 ;
      RECT  95612.5 206942.5 95677.5 207077.5 ;
      RECT  95802.5 206942.5 95867.5 207077.5 ;
      RECT  95612.5 207472.5 95677.5 207607.5 ;
      RECT  95992.5 207472.5 96057.5 207607.5 ;
      RECT  95450.0 207237.5 96155.0 207302.5 ;
      RECT  95450.0 207922.5 96155.0 207987.5 ;
      RECT  96507.5 207472.5 96572.5 207987.5 ;
      RECT  96317.5 206942.5 96382.5 207077.5 ;
      RECT  96507.5 206942.5 96572.5 207077.5 ;
      RECT  96507.5 206942.5 96572.5 207077.5 ;
      RECT  96317.5 206942.5 96382.5 207077.5 ;
      RECT  96317.5 207472.5 96382.5 207607.5 ;
      RECT  96507.5 207472.5 96572.5 207607.5 ;
      RECT  96507.5 207472.5 96572.5 207607.5 ;
      RECT  96317.5 207472.5 96382.5 207607.5 ;
      RECT  96507.5 207472.5 96572.5 207607.5 ;
      RECT  96697.5 207472.5 96762.5 207607.5 ;
      RECT  96697.5 207472.5 96762.5 207607.5 ;
      RECT  96507.5 207472.5 96572.5 207607.5 ;
      RECT  96487.5 207237.5 96352.5 207302.5 ;
      RECT  96507.5 207785.0 96572.5 207920.0 ;
      RECT  96317.5 206942.5 96382.5 207077.5 ;
      RECT  96507.5 206942.5 96572.5 207077.5 ;
      RECT  96317.5 207472.5 96382.5 207607.5 ;
      RECT  96697.5 207472.5 96762.5 207607.5 ;
      RECT  96155.0 207237.5 96860.0 207302.5 ;
      RECT  96155.0 207922.5 96860.0 207987.5 ;
      RECT  97212.5 207472.5 97277.5 207987.5 ;
      RECT  97022.5 206942.5 97087.5 207077.5 ;
      RECT  97212.5 206942.5 97277.5 207077.5 ;
      RECT  97212.5 206942.5 97277.5 207077.5 ;
      RECT  97022.5 206942.5 97087.5 207077.5 ;
      RECT  97022.5 207472.5 97087.5 207607.5 ;
      RECT  97212.5 207472.5 97277.5 207607.5 ;
      RECT  97212.5 207472.5 97277.5 207607.5 ;
      RECT  97022.5 207472.5 97087.5 207607.5 ;
      RECT  97212.5 207472.5 97277.5 207607.5 ;
      RECT  97402.5 207472.5 97467.5 207607.5 ;
      RECT  97402.5 207472.5 97467.5 207607.5 ;
      RECT  97212.5 207472.5 97277.5 207607.5 ;
      RECT  97192.5 207237.5 97057.5 207302.5 ;
      RECT  97212.5 207785.0 97277.5 207920.0 ;
      RECT  97022.5 206942.5 97087.5 207077.5 ;
      RECT  97212.5 206942.5 97277.5 207077.5 ;
      RECT  97022.5 207472.5 97087.5 207607.5 ;
      RECT  97402.5 207472.5 97467.5 207607.5 ;
      RECT  96860.0 207237.5 97565.0 207302.5 ;
      RECT  96860.0 207922.5 97565.0 207987.5 ;
      RECT  97917.5 207472.5 97982.5 207987.5 ;
      RECT  97727.5 206942.5 97792.5 207077.5 ;
      RECT  97917.5 206942.5 97982.5 207077.5 ;
      RECT  97917.5 206942.5 97982.5 207077.5 ;
      RECT  97727.5 206942.5 97792.5 207077.5 ;
      RECT  97727.5 207472.5 97792.5 207607.5 ;
      RECT  97917.5 207472.5 97982.5 207607.5 ;
      RECT  97917.5 207472.5 97982.5 207607.5 ;
      RECT  97727.5 207472.5 97792.5 207607.5 ;
      RECT  97917.5 207472.5 97982.5 207607.5 ;
      RECT  98107.5 207472.5 98172.5 207607.5 ;
      RECT  98107.5 207472.5 98172.5 207607.5 ;
      RECT  97917.5 207472.5 97982.5 207607.5 ;
      RECT  97897.5 207237.5 97762.5 207302.5 ;
      RECT  97917.5 207785.0 97982.5 207920.0 ;
      RECT  97727.5 206942.5 97792.5 207077.5 ;
      RECT  97917.5 206942.5 97982.5 207077.5 ;
      RECT  97727.5 207472.5 97792.5 207607.5 ;
      RECT  98107.5 207472.5 98172.5 207607.5 ;
      RECT  97565.0 207237.5 98270.0 207302.5 ;
      RECT  97565.0 207922.5 98270.0 207987.5 ;
      RECT  98622.5 207472.5 98687.5 207987.5 ;
      RECT  98432.5 206942.5 98497.5 207077.5 ;
      RECT  98622.5 206942.5 98687.5 207077.5 ;
      RECT  98622.5 206942.5 98687.5 207077.5 ;
      RECT  98432.5 206942.5 98497.5 207077.5 ;
      RECT  98432.5 207472.5 98497.5 207607.5 ;
      RECT  98622.5 207472.5 98687.5 207607.5 ;
      RECT  98622.5 207472.5 98687.5 207607.5 ;
      RECT  98432.5 207472.5 98497.5 207607.5 ;
      RECT  98622.5 207472.5 98687.5 207607.5 ;
      RECT  98812.5 207472.5 98877.5 207607.5 ;
      RECT  98812.5 207472.5 98877.5 207607.5 ;
      RECT  98622.5 207472.5 98687.5 207607.5 ;
      RECT  98602.5 207237.5 98467.5 207302.5 ;
      RECT  98622.5 207785.0 98687.5 207920.0 ;
      RECT  98432.5 206942.5 98497.5 207077.5 ;
      RECT  98622.5 206942.5 98687.5 207077.5 ;
      RECT  98432.5 207472.5 98497.5 207607.5 ;
      RECT  98812.5 207472.5 98877.5 207607.5 ;
      RECT  98270.0 207237.5 98975.0 207302.5 ;
      RECT  98270.0 207922.5 98975.0 207987.5 ;
      RECT  99327.5 207472.5 99392.5 207987.5 ;
      RECT  99137.5 206942.5 99202.5 207077.5 ;
      RECT  99327.5 206942.5 99392.5 207077.5 ;
      RECT  99327.5 206942.5 99392.5 207077.5 ;
      RECT  99137.5 206942.5 99202.5 207077.5 ;
      RECT  99137.5 207472.5 99202.5 207607.5 ;
      RECT  99327.5 207472.5 99392.5 207607.5 ;
      RECT  99327.5 207472.5 99392.5 207607.5 ;
      RECT  99137.5 207472.5 99202.5 207607.5 ;
      RECT  99327.5 207472.5 99392.5 207607.5 ;
      RECT  99517.5 207472.5 99582.5 207607.5 ;
      RECT  99517.5 207472.5 99582.5 207607.5 ;
      RECT  99327.5 207472.5 99392.5 207607.5 ;
      RECT  99307.5 207237.5 99172.5 207302.5 ;
      RECT  99327.5 207785.0 99392.5 207920.0 ;
      RECT  99137.5 206942.5 99202.5 207077.5 ;
      RECT  99327.5 206942.5 99392.5 207077.5 ;
      RECT  99137.5 207472.5 99202.5 207607.5 ;
      RECT  99517.5 207472.5 99582.5 207607.5 ;
      RECT  98975.0 207237.5 99680.0 207302.5 ;
      RECT  98975.0 207922.5 99680.0 207987.5 ;
      RECT  100032.5 207472.5 100097.5 207987.5 ;
      RECT  99842.5 206942.5 99907.5 207077.5 ;
      RECT  100032.5 206942.5 100097.5 207077.5 ;
      RECT  100032.5 206942.5 100097.5 207077.5 ;
      RECT  99842.5 206942.5 99907.5 207077.5 ;
      RECT  99842.5 207472.5 99907.5 207607.5 ;
      RECT  100032.5 207472.5 100097.5 207607.5 ;
      RECT  100032.5 207472.5 100097.5 207607.5 ;
      RECT  99842.5 207472.5 99907.5 207607.5 ;
      RECT  100032.5 207472.5 100097.5 207607.5 ;
      RECT  100222.5 207472.5 100287.5 207607.5 ;
      RECT  100222.5 207472.5 100287.5 207607.5 ;
      RECT  100032.5 207472.5 100097.5 207607.5 ;
      RECT  100012.5 207237.5 99877.5 207302.5 ;
      RECT  100032.5 207785.0 100097.5 207920.0 ;
      RECT  99842.5 206942.5 99907.5 207077.5 ;
      RECT  100032.5 206942.5 100097.5 207077.5 ;
      RECT  99842.5 207472.5 99907.5 207607.5 ;
      RECT  100222.5 207472.5 100287.5 207607.5 ;
      RECT  99680.0 207237.5 100385.0 207302.5 ;
      RECT  99680.0 207922.5 100385.0 207987.5 ;
      RECT  100737.5 207472.5 100802.5 207987.5 ;
      RECT  100547.5 206942.5 100612.5 207077.5 ;
      RECT  100737.5 206942.5 100802.5 207077.5 ;
      RECT  100737.5 206942.5 100802.5 207077.5 ;
      RECT  100547.5 206942.5 100612.5 207077.5 ;
      RECT  100547.5 207472.5 100612.5 207607.5 ;
      RECT  100737.5 207472.5 100802.5 207607.5 ;
      RECT  100737.5 207472.5 100802.5 207607.5 ;
      RECT  100547.5 207472.5 100612.5 207607.5 ;
      RECT  100737.5 207472.5 100802.5 207607.5 ;
      RECT  100927.5 207472.5 100992.5 207607.5 ;
      RECT  100927.5 207472.5 100992.5 207607.5 ;
      RECT  100737.5 207472.5 100802.5 207607.5 ;
      RECT  100717.5 207237.5 100582.5 207302.5 ;
      RECT  100737.5 207785.0 100802.5 207920.0 ;
      RECT  100547.5 206942.5 100612.5 207077.5 ;
      RECT  100737.5 206942.5 100802.5 207077.5 ;
      RECT  100547.5 207472.5 100612.5 207607.5 ;
      RECT  100927.5 207472.5 100992.5 207607.5 ;
      RECT  100385.0 207237.5 101090.0 207302.5 ;
      RECT  100385.0 207922.5 101090.0 207987.5 ;
      RECT  101442.5 207472.5 101507.5 207987.5 ;
      RECT  101252.5 206942.5 101317.5 207077.5 ;
      RECT  101442.5 206942.5 101507.5 207077.5 ;
      RECT  101442.5 206942.5 101507.5 207077.5 ;
      RECT  101252.5 206942.5 101317.5 207077.5 ;
      RECT  101252.5 207472.5 101317.5 207607.5 ;
      RECT  101442.5 207472.5 101507.5 207607.5 ;
      RECT  101442.5 207472.5 101507.5 207607.5 ;
      RECT  101252.5 207472.5 101317.5 207607.5 ;
      RECT  101442.5 207472.5 101507.5 207607.5 ;
      RECT  101632.5 207472.5 101697.5 207607.5 ;
      RECT  101632.5 207472.5 101697.5 207607.5 ;
      RECT  101442.5 207472.5 101507.5 207607.5 ;
      RECT  101422.5 207237.5 101287.5 207302.5 ;
      RECT  101442.5 207785.0 101507.5 207920.0 ;
      RECT  101252.5 206942.5 101317.5 207077.5 ;
      RECT  101442.5 206942.5 101507.5 207077.5 ;
      RECT  101252.5 207472.5 101317.5 207607.5 ;
      RECT  101632.5 207472.5 101697.5 207607.5 ;
      RECT  101090.0 207237.5 101795.0 207302.5 ;
      RECT  101090.0 207922.5 101795.0 207987.5 ;
      RECT  102147.5 207472.5 102212.5 207987.5 ;
      RECT  101957.5 206942.5 102022.5 207077.5 ;
      RECT  102147.5 206942.5 102212.5 207077.5 ;
      RECT  102147.5 206942.5 102212.5 207077.5 ;
      RECT  101957.5 206942.5 102022.5 207077.5 ;
      RECT  101957.5 207472.5 102022.5 207607.5 ;
      RECT  102147.5 207472.5 102212.5 207607.5 ;
      RECT  102147.5 207472.5 102212.5 207607.5 ;
      RECT  101957.5 207472.5 102022.5 207607.5 ;
      RECT  102147.5 207472.5 102212.5 207607.5 ;
      RECT  102337.5 207472.5 102402.5 207607.5 ;
      RECT  102337.5 207472.5 102402.5 207607.5 ;
      RECT  102147.5 207472.5 102212.5 207607.5 ;
      RECT  102127.5 207237.5 101992.5 207302.5 ;
      RECT  102147.5 207785.0 102212.5 207920.0 ;
      RECT  101957.5 206942.5 102022.5 207077.5 ;
      RECT  102147.5 206942.5 102212.5 207077.5 ;
      RECT  101957.5 207472.5 102022.5 207607.5 ;
      RECT  102337.5 207472.5 102402.5 207607.5 ;
      RECT  101795.0 207237.5 102500.0 207302.5 ;
      RECT  101795.0 207922.5 102500.0 207987.5 ;
      RECT  102852.5 207472.5 102917.5 207987.5 ;
      RECT  102662.5 206942.5 102727.5 207077.5 ;
      RECT  102852.5 206942.5 102917.5 207077.5 ;
      RECT  102852.5 206942.5 102917.5 207077.5 ;
      RECT  102662.5 206942.5 102727.5 207077.5 ;
      RECT  102662.5 207472.5 102727.5 207607.5 ;
      RECT  102852.5 207472.5 102917.5 207607.5 ;
      RECT  102852.5 207472.5 102917.5 207607.5 ;
      RECT  102662.5 207472.5 102727.5 207607.5 ;
      RECT  102852.5 207472.5 102917.5 207607.5 ;
      RECT  103042.5 207472.5 103107.5 207607.5 ;
      RECT  103042.5 207472.5 103107.5 207607.5 ;
      RECT  102852.5 207472.5 102917.5 207607.5 ;
      RECT  102832.5 207237.5 102697.5 207302.5 ;
      RECT  102852.5 207785.0 102917.5 207920.0 ;
      RECT  102662.5 206942.5 102727.5 207077.5 ;
      RECT  102852.5 206942.5 102917.5 207077.5 ;
      RECT  102662.5 207472.5 102727.5 207607.5 ;
      RECT  103042.5 207472.5 103107.5 207607.5 ;
      RECT  102500.0 207237.5 103205.0 207302.5 ;
      RECT  102500.0 207922.5 103205.0 207987.5 ;
      RECT  103557.5 207472.5 103622.5 207987.5 ;
      RECT  103367.5 206942.5 103432.5 207077.5 ;
      RECT  103557.5 206942.5 103622.5 207077.5 ;
      RECT  103557.5 206942.5 103622.5 207077.5 ;
      RECT  103367.5 206942.5 103432.5 207077.5 ;
      RECT  103367.5 207472.5 103432.5 207607.5 ;
      RECT  103557.5 207472.5 103622.5 207607.5 ;
      RECT  103557.5 207472.5 103622.5 207607.5 ;
      RECT  103367.5 207472.5 103432.5 207607.5 ;
      RECT  103557.5 207472.5 103622.5 207607.5 ;
      RECT  103747.5 207472.5 103812.5 207607.5 ;
      RECT  103747.5 207472.5 103812.5 207607.5 ;
      RECT  103557.5 207472.5 103622.5 207607.5 ;
      RECT  103537.5 207237.5 103402.5 207302.5 ;
      RECT  103557.5 207785.0 103622.5 207920.0 ;
      RECT  103367.5 206942.5 103432.5 207077.5 ;
      RECT  103557.5 206942.5 103622.5 207077.5 ;
      RECT  103367.5 207472.5 103432.5 207607.5 ;
      RECT  103747.5 207472.5 103812.5 207607.5 ;
      RECT  103205.0 207237.5 103910.0 207302.5 ;
      RECT  103205.0 207922.5 103910.0 207987.5 ;
      RECT  104262.5 207472.5 104327.5 207987.5 ;
      RECT  104072.5 206942.5 104137.5 207077.5 ;
      RECT  104262.5 206942.5 104327.5 207077.5 ;
      RECT  104262.5 206942.5 104327.5 207077.5 ;
      RECT  104072.5 206942.5 104137.5 207077.5 ;
      RECT  104072.5 207472.5 104137.5 207607.5 ;
      RECT  104262.5 207472.5 104327.5 207607.5 ;
      RECT  104262.5 207472.5 104327.5 207607.5 ;
      RECT  104072.5 207472.5 104137.5 207607.5 ;
      RECT  104262.5 207472.5 104327.5 207607.5 ;
      RECT  104452.5 207472.5 104517.5 207607.5 ;
      RECT  104452.5 207472.5 104517.5 207607.5 ;
      RECT  104262.5 207472.5 104327.5 207607.5 ;
      RECT  104242.5 207237.5 104107.5 207302.5 ;
      RECT  104262.5 207785.0 104327.5 207920.0 ;
      RECT  104072.5 206942.5 104137.5 207077.5 ;
      RECT  104262.5 206942.5 104327.5 207077.5 ;
      RECT  104072.5 207472.5 104137.5 207607.5 ;
      RECT  104452.5 207472.5 104517.5 207607.5 ;
      RECT  103910.0 207237.5 104615.0 207302.5 ;
      RECT  103910.0 207922.5 104615.0 207987.5 ;
      RECT  104967.5 207472.5 105032.5 207987.5 ;
      RECT  104777.5 206942.5 104842.5 207077.5 ;
      RECT  104967.5 206942.5 105032.5 207077.5 ;
      RECT  104967.5 206942.5 105032.5 207077.5 ;
      RECT  104777.5 206942.5 104842.5 207077.5 ;
      RECT  104777.5 207472.5 104842.5 207607.5 ;
      RECT  104967.5 207472.5 105032.5 207607.5 ;
      RECT  104967.5 207472.5 105032.5 207607.5 ;
      RECT  104777.5 207472.5 104842.5 207607.5 ;
      RECT  104967.5 207472.5 105032.5 207607.5 ;
      RECT  105157.5 207472.5 105222.5 207607.5 ;
      RECT  105157.5 207472.5 105222.5 207607.5 ;
      RECT  104967.5 207472.5 105032.5 207607.5 ;
      RECT  104947.5 207237.5 104812.5 207302.5 ;
      RECT  104967.5 207785.0 105032.5 207920.0 ;
      RECT  104777.5 206942.5 104842.5 207077.5 ;
      RECT  104967.5 206942.5 105032.5 207077.5 ;
      RECT  104777.5 207472.5 104842.5 207607.5 ;
      RECT  105157.5 207472.5 105222.5 207607.5 ;
      RECT  104615.0 207237.5 105320.0 207302.5 ;
      RECT  104615.0 207922.5 105320.0 207987.5 ;
      RECT  105672.5 207472.5 105737.5 207987.5 ;
      RECT  105482.5 206942.5 105547.5 207077.5 ;
      RECT  105672.5 206942.5 105737.5 207077.5 ;
      RECT  105672.5 206942.5 105737.5 207077.5 ;
      RECT  105482.5 206942.5 105547.5 207077.5 ;
      RECT  105482.5 207472.5 105547.5 207607.5 ;
      RECT  105672.5 207472.5 105737.5 207607.5 ;
      RECT  105672.5 207472.5 105737.5 207607.5 ;
      RECT  105482.5 207472.5 105547.5 207607.5 ;
      RECT  105672.5 207472.5 105737.5 207607.5 ;
      RECT  105862.5 207472.5 105927.5 207607.5 ;
      RECT  105862.5 207472.5 105927.5 207607.5 ;
      RECT  105672.5 207472.5 105737.5 207607.5 ;
      RECT  105652.5 207237.5 105517.5 207302.5 ;
      RECT  105672.5 207785.0 105737.5 207920.0 ;
      RECT  105482.5 206942.5 105547.5 207077.5 ;
      RECT  105672.5 206942.5 105737.5 207077.5 ;
      RECT  105482.5 207472.5 105547.5 207607.5 ;
      RECT  105862.5 207472.5 105927.5 207607.5 ;
      RECT  105320.0 207237.5 106025.0 207302.5 ;
      RECT  105320.0 207922.5 106025.0 207987.5 ;
      RECT  106377.5 207472.5 106442.5 207987.5 ;
      RECT  106187.5 206942.5 106252.5 207077.5 ;
      RECT  106377.5 206942.5 106442.5 207077.5 ;
      RECT  106377.5 206942.5 106442.5 207077.5 ;
      RECT  106187.5 206942.5 106252.5 207077.5 ;
      RECT  106187.5 207472.5 106252.5 207607.5 ;
      RECT  106377.5 207472.5 106442.5 207607.5 ;
      RECT  106377.5 207472.5 106442.5 207607.5 ;
      RECT  106187.5 207472.5 106252.5 207607.5 ;
      RECT  106377.5 207472.5 106442.5 207607.5 ;
      RECT  106567.5 207472.5 106632.5 207607.5 ;
      RECT  106567.5 207472.5 106632.5 207607.5 ;
      RECT  106377.5 207472.5 106442.5 207607.5 ;
      RECT  106357.5 207237.5 106222.5 207302.5 ;
      RECT  106377.5 207785.0 106442.5 207920.0 ;
      RECT  106187.5 206942.5 106252.5 207077.5 ;
      RECT  106377.5 206942.5 106442.5 207077.5 ;
      RECT  106187.5 207472.5 106252.5 207607.5 ;
      RECT  106567.5 207472.5 106632.5 207607.5 ;
      RECT  106025.0 207237.5 106730.0 207302.5 ;
      RECT  106025.0 207922.5 106730.0 207987.5 ;
      RECT  107082.5 207472.5 107147.5 207987.5 ;
      RECT  106892.5 206942.5 106957.5 207077.5 ;
      RECT  107082.5 206942.5 107147.5 207077.5 ;
      RECT  107082.5 206942.5 107147.5 207077.5 ;
      RECT  106892.5 206942.5 106957.5 207077.5 ;
      RECT  106892.5 207472.5 106957.5 207607.5 ;
      RECT  107082.5 207472.5 107147.5 207607.5 ;
      RECT  107082.5 207472.5 107147.5 207607.5 ;
      RECT  106892.5 207472.5 106957.5 207607.5 ;
      RECT  107082.5 207472.5 107147.5 207607.5 ;
      RECT  107272.5 207472.5 107337.5 207607.5 ;
      RECT  107272.5 207472.5 107337.5 207607.5 ;
      RECT  107082.5 207472.5 107147.5 207607.5 ;
      RECT  107062.5 207237.5 106927.5 207302.5 ;
      RECT  107082.5 207785.0 107147.5 207920.0 ;
      RECT  106892.5 206942.5 106957.5 207077.5 ;
      RECT  107082.5 206942.5 107147.5 207077.5 ;
      RECT  106892.5 207472.5 106957.5 207607.5 ;
      RECT  107272.5 207472.5 107337.5 207607.5 ;
      RECT  106730.0 207237.5 107435.0 207302.5 ;
      RECT  106730.0 207922.5 107435.0 207987.5 ;
      RECT  17195.0 207237.5 107435.0 207302.5 ;
      RECT  17195.0 207922.5 107435.0 207987.5 ;
      RECT  17345.0 31535.0 19530.0 31605.0 ;
      RECT  17680.0 31395.0 19865.0 31465.0 ;
      RECT  20165.0 31535.0 22350.0 31605.0 ;
      RECT  20500.0 31395.0 22685.0 31465.0 ;
      RECT  22985.0 31535.0 25170.0 31605.0 ;
      RECT  23320.0 31395.0 25505.0 31465.0 ;
      RECT  25805.0 31535.0 27990.0 31605.0 ;
      RECT  26140.0 31395.0 28325.0 31465.0 ;
      RECT  28625.0 31535.0 30810.0 31605.0 ;
      RECT  28960.0 31395.0 31145.0 31465.0 ;
      RECT  31445.0 31535.0 33630.0 31605.0 ;
      RECT  31780.0 31395.0 33965.0 31465.0 ;
      RECT  34265.0 31535.0 36450.0 31605.0 ;
      RECT  34600.0 31395.0 36785.0 31465.0 ;
      RECT  37085.0 31535.0 39270.0 31605.0 ;
      RECT  37420.0 31395.0 39605.0 31465.0 ;
      RECT  39905.0 31535.0 42090.0 31605.0 ;
      RECT  40240.0 31395.0 42425.0 31465.0 ;
      RECT  42725.0 31535.0 44910.0 31605.0 ;
      RECT  43060.0 31395.0 45245.0 31465.0 ;
      RECT  45545.0 31535.0 47730.0 31605.0 ;
      RECT  45880.0 31395.0 48065.0 31465.0 ;
      RECT  48365.0 31535.0 50550.0 31605.0 ;
      RECT  48700.0 31395.0 50885.0 31465.0 ;
      RECT  51185.0 31535.0 53370.0 31605.0 ;
      RECT  51520.0 31395.0 53705.0 31465.0 ;
      RECT  54005.0 31535.0 56190.0 31605.0 ;
      RECT  54340.0 31395.0 56525.0 31465.0 ;
      RECT  56825.0 31535.0 59010.0 31605.0 ;
      RECT  57160.0 31395.0 59345.0 31465.0 ;
      RECT  59645.0 31535.0 61830.0 31605.0 ;
      RECT  59980.0 31395.0 62165.0 31465.0 ;
      RECT  62465.0 31535.0 64650.0 31605.0 ;
      RECT  62800.0 31395.0 64985.0 31465.0 ;
      RECT  65285.0 31535.0 67470.0 31605.0 ;
      RECT  65620.0 31395.0 67805.0 31465.0 ;
      RECT  68105.0 31535.0 70290.0 31605.0 ;
      RECT  68440.0 31395.0 70625.0 31465.0 ;
      RECT  70925.0 31535.0 73110.0 31605.0 ;
      RECT  71260.0 31395.0 73445.0 31465.0 ;
      RECT  73745.0 31535.0 75930.0 31605.0 ;
      RECT  74080.0 31395.0 76265.0 31465.0 ;
      RECT  76565.0 31535.0 78750.0 31605.0 ;
      RECT  76900.0 31395.0 79085.0 31465.0 ;
      RECT  79385.0 31535.0 81570.0 31605.0 ;
      RECT  79720.0 31395.0 81905.0 31465.0 ;
      RECT  82205.0 31535.0 84390.0 31605.0 ;
      RECT  82540.0 31395.0 84725.0 31465.0 ;
      RECT  85025.0 31535.0 87210.0 31605.0 ;
      RECT  85360.0 31395.0 87545.0 31465.0 ;
      RECT  87845.0 31535.0 90030.0 31605.0 ;
      RECT  88180.0 31395.0 90365.0 31465.0 ;
      RECT  90665.0 31535.0 92850.0 31605.0 ;
      RECT  91000.0 31395.0 93185.0 31465.0 ;
      RECT  93485.0 31535.0 95670.0 31605.0 ;
      RECT  93820.0 31395.0 96005.0 31465.0 ;
      RECT  96305.0 31535.0 98490.0 31605.0 ;
      RECT  96640.0 31395.0 98825.0 31465.0 ;
      RECT  99125.0 31535.0 101310.0 31605.0 ;
      RECT  99460.0 31395.0 101645.0 31465.0 ;
      RECT  101945.0 31535.0 104130.0 31605.0 ;
      RECT  102280.0 31395.0 104465.0 31465.0 ;
      RECT  104765.0 31535.0 106950.0 31605.0 ;
      RECT  105100.0 31395.0 107285.0 31465.0 ;
      RECT  17610.0 33892.5 17675.0 33957.5 ;
      RECT  17345.0 33892.5 17642.5 33957.5 ;
      RECT  17610.0 33510.0 17675.0 33925.0 ;
      RECT  17420.0 32342.5 17485.0 32407.5 ;
      RECT  17452.5 32342.5 17715.0 32407.5 ;
      RECT  17420.0 32375.0 17485.0 32650.0 ;
      RECT  17420.0 32582.5 17485.0 32717.5 ;
      RECT  17610.0 32582.5 17675.0 32717.5 ;
      RECT  17610.0 32582.5 17675.0 32717.5 ;
      RECT  17420.0 32582.5 17485.0 32717.5 ;
      RECT  17420.0 33442.5 17485.0 33577.5 ;
      RECT  17610.0 33442.5 17675.0 33577.5 ;
      RECT  17610.0 33442.5 17675.0 33577.5 ;
      RECT  17420.0 33442.5 17485.0 33577.5 ;
      RECT  17347.5 33857.5 17412.5 33992.5 ;
      RECT  17682.5 32307.5 17747.5 32442.5 ;
      RECT  17420.0 33442.5 17485.0 33577.5 ;
      RECT  17610.0 32582.5 17675.0 32717.5 ;
      RECT  17867.5 32482.5 17932.5 32617.5 ;
      RECT  17867.5 32482.5 17932.5 32617.5 ;
      RECT  18315.0 33892.5 18380.0 33957.5 ;
      RECT  18050.0 33892.5 18347.5 33957.5 ;
      RECT  18315.0 33510.0 18380.0 33925.0 ;
      RECT  18125.0 32342.5 18190.0 32407.5 ;
      RECT  18157.5 32342.5 18420.0 32407.5 ;
      RECT  18125.0 32375.0 18190.0 32650.0 ;
      RECT  18125.0 32582.5 18190.0 32717.5 ;
      RECT  18315.0 32582.5 18380.0 32717.5 ;
      RECT  18315.0 32582.5 18380.0 32717.5 ;
      RECT  18125.0 32582.5 18190.0 32717.5 ;
      RECT  18125.0 33442.5 18190.0 33577.5 ;
      RECT  18315.0 33442.5 18380.0 33577.5 ;
      RECT  18315.0 33442.5 18380.0 33577.5 ;
      RECT  18125.0 33442.5 18190.0 33577.5 ;
      RECT  18052.5 33857.5 18117.5 33992.5 ;
      RECT  18387.5 32307.5 18452.5 32442.5 ;
      RECT  18125.0 33442.5 18190.0 33577.5 ;
      RECT  18315.0 32582.5 18380.0 32717.5 ;
      RECT  18572.5 32482.5 18637.5 32617.5 ;
      RECT  18572.5 32482.5 18637.5 32617.5 ;
      RECT  19020.0 33892.5 19085.0 33957.5 ;
      RECT  18755.0 33892.5 19052.5 33957.5 ;
      RECT  19020.0 33510.0 19085.0 33925.0 ;
      RECT  18830.0 32342.5 18895.0 32407.5 ;
      RECT  18862.5 32342.5 19125.0 32407.5 ;
      RECT  18830.0 32375.0 18895.0 32650.0 ;
      RECT  18830.0 32582.5 18895.0 32717.5 ;
      RECT  19020.0 32582.5 19085.0 32717.5 ;
      RECT  19020.0 32582.5 19085.0 32717.5 ;
      RECT  18830.0 32582.5 18895.0 32717.5 ;
      RECT  18830.0 33442.5 18895.0 33577.5 ;
      RECT  19020.0 33442.5 19085.0 33577.5 ;
      RECT  19020.0 33442.5 19085.0 33577.5 ;
      RECT  18830.0 33442.5 18895.0 33577.5 ;
      RECT  18757.5 33857.5 18822.5 33992.5 ;
      RECT  19092.5 32307.5 19157.5 32442.5 ;
      RECT  18830.0 33442.5 18895.0 33577.5 ;
      RECT  19020.0 32582.5 19085.0 32717.5 ;
      RECT  19277.5 32482.5 19342.5 32617.5 ;
      RECT  19277.5 32482.5 19342.5 32617.5 ;
      RECT  19725.0 33892.5 19790.0 33957.5 ;
      RECT  19460.0 33892.5 19757.5 33957.5 ;
      RECT  19725.0 33510.0 19790.0 33925.0 ;
      RECT  19535.0 32342.5 19600.0 32407.5 ;
      RECT  19567.5 32342.5 19830.0 32407.5 ;
      RECT  19535.0 32375.0 19600.0 32650.0 ;
      RECT  19535.0 32582.5 19600.0 32717.5 ;
      RECT  19725.0 32582.5 19790.0 32717.5 ;
      RECT  19725.0 32582.5 19790.0 32717.5 ;
      RECT  19535.0 32582.5 19600.0 32717.5 ;
      RECT  19535.0 33442.5 19600.0 33577.5 ;
      RECT  19725.0 33442.5 19790.0 33577.5 ;
      RECT  19725.0 33442.5 19790.0 33577.5 ;
      RECT  19535.0 33442.5 19600.0 33577.5 ;
      RECT  19462.5 33857.5 19527.5 33992.5 ;
      RECT  19797.5 32307.5 19862.5 32442.5 ;
      RECT  19535.0 33442.5 19600.0 33577.5 ;
      RECT  19725.0 32582.5 19790.0 32717.5 ;
      RECT  19982.5 32482.5 20047.5 32617.5 ;
      RECT  19982.5 32482.5 20047.5 32617.5 ;
      RECT  20430.0 33892.5 20495.0 33957.5 ;
      RECT  20165.0 33892.5 20462.5 33957.5 ;
      RECT  20430.0 33510.0 20495.0 33925.0 ;
      RECT  20240.0 32342.5 20305.0 32407.5 ;
      RECT  20272.5 32342.5 20535.0 32407.5 ;
      RECT  20240.0 32375.0 20305.0 32650.0 ;
      RECT  20240.0 32582.5 20305.0 32717.5 ;
      RECT  20430.0 32582.5 20495.0 32717.5 ;
      RECT  20430.0 32582.5 20495.0 32717.5 ;
      RECT  20240.0 32582.5 20305.0 32717.5 ;
      RECT  20240.0 33442.5 20305.0 33577.5 ;
      RECT  20430.0 33442.5 20495.0 33577.5 ;
      RECT  20430.0 33442.5 20495.0 33577.5 ;
      RECT  20240.0 33442.5 20305.0 33577.5 ;
      RECT  20167.5 33857.5 20232.5 33992.5 ;
      RECT  20502.5 32307.5 20567.5 32442.5 ;
      RECT  20240.0 33442.5 20305.0 33577.5 ;
      RECT  20430.0 32582.5 20495.0 32717.5 ;
      RECT  20687.5 32482.5 20752.5 32617.5 ;
      RECT  20687.5 32482.5 20752.5 32617.5 ;
      RECT  21135.0 33892.5 21200.0 33957.5 ;
      RECT  20870.0 33892.5 21167.5 33957.5 ;
      RECT  21135.0 33510.0 21200.0 33925.0 ;
      RECT  20945.0 32342.5 21010.0 32407.5 ;
      RECT  20977.5 32342.5 21240.0 32407.5 ;
      RECT  20945.0 32375.0 21010.0 32650.0 ;
      RECT  20945.0 32582.5 21010.0 32717.5 ;
      RECT  21135.0 32582.5 21200.0 32717.5 ;
      RECT  21135.0 32582.5 21200.0 32717.5 ;
      RECT  20945.0 32582.5 21010.0 32717.5 ;
      RECT  20945.0 33442.5 21010.0 33577.5 ;
      RECT  21135.0 33442.5 21200.0 33577.5 ;
      RECT  21135.0 33442.5 21200.0 33577.5 ;
      RECT  20945.0 33442.5 21010.0 33577.5 ;
      RECT  20872.5 33857.5 20937.5 33992.5 ;
      RECT  21207.5 32307.5 21272.5 32442.5 ;
      RECT  20945.0 33442.5 21010.0 33577.5 ;
      RECT  21135.0 32582.5 21200.0 32717.5 ;
      RECT  21392.5 32482.5 21457.5 32617.5 ;
      RECT  21392.5 32482.5 21457.5 32617.5 ;
      RECT  21840.0 33892.5 21905.0 33957.5 ;
      RECT  21575.0 33892.5 21872.5 33957.5 ;
      RECT  21840.0 33510.0 21905.0 33925.0 ;
      RECT  21650.0 32342.5 21715.0 32407.5 ;
      RECT  21682.5 32342.5 21945.0 32407.5 ;
      RECT  21650.0 32375.0 21715.0 32650.0 ;
      RECT  21650.0 32582.5 21715.0 32717.5 ;
      RECT  21840.0 32582.5 21905.0 32717.5 ;
      RECT  21840.0 32582.5 21905.0 32717.5 ;
      RECT  21650.0 32582.5 21715.0 32717.5 ;
      RECT  21650.0 33442.5 21715.0 33577.5 ;
      RECT  21840.0 33442.5 21905.0 33577.5 ;
      RECT  21840.0 33442.5 21905.0 33577.5 ;
      RECT  21650.0 33442.5 21715.0 33577.5 ;
      RECT  21577.5 33857.5 21642.5 33992.5 ;
      RECT  21912.5 32307.5 21977.5 32442.5 ;
      RECT  21650.0 33442.5 21715.0 33577.5 ;
      RECT  21840.0 32582.5 21905.0 32717.5 ;
      RECT  22097.5 32482.5 22162.5 32617.5 ;
      RECT  22097.5 32482.5 22162.5 32617.5 ;
      RECT  22545.0 33892.5 22610.0 33957.5 ;
      RECT  22280.0 33892.5 22577.5 33957.5 ;
      RECT  22545.0 33510.0 22610.0 33925.0 ;
      RECT  22355.0 32342.5 22420.0 32407.5 ;
      RECT  22387.5 32342.5 22650.0 32407.5 ;
      RECT  22355.0 32375.0 22420.0 32650.0 ;
      RECT  22355.0 32582.5 22420.0 32717.5 ;
      RECT  22545.0 32582.5 22610.0 32717.5 ;
      RECT  22545.0 32582.5 22610.0 32717.5 ;
      RECT  22355.0 32582.5 22420.0 32717.5 ;
      RECT  22355.0 33442.5 22420.0 33577.5 ;
      RECT  22545.0 33442.5 22610.0 33577.5 ;
      RECT  22545.0 33442.5 22610.0 33577.5 ;
      RECT  22355.0 33442.5 22420.0 33577.5 ;
      RECT  22282.5 33857.5 22347.5 33992.5 ;
      RECT  22617.5 32307.5 22682.5 32442.5 ;
      RECT  22355.0 33442.5 22420.0 33577.5 ;
      RECT  22545.0 32582.5 22610.0 32717.5 ;
      RECT  22802.5 32482.5 22867.5 32617.5 ;
      RECT  22802.5 32482.5 22867.5 32617.5 ;
      RECT  23250.0 33892.5 23315.0 33957.5 ;
      RECT  22985.0 33892.5 23282.5 33957.5 ;
      RECT  23250.0 33510.0 23315.0 33925.0 ;
      RECT  23060.0 32342.5 23125.0 32407.5 ;
      RECT  23092.5 32342.5 23355.0 32407.5 ;
      RECT  23060.0 32375.0 23125.0 32650.0 ;
      RECT  23060.0 32582.5 23125.0 32717.5 ;
      RECT  23250.0 32582.5 23315.0 32717.5 ;
      RECT  23250.0 32582.5 23315.0 32717.5 ;
      RECT  23060.0 32582.5 23125.0 32717.5 ;
      RECT  23060.0 33442.5 23125.0 33577.5 ;
      RECT  23250.0 33442.5 23315.0 33577.5 ;
      RECT  23250.0 33442.5 23315.0 33577.5 ;
      RECT  23060.0 33442.5 23125.0 33577.5 ;
      RECT  22987.5 33857.5 23052.5 33992.5 ;
      RECT  23322.5 32307.5 23387.5 32442.5 ;
      RECT  23060.0 33442.5 23125.0 33577.5 ;
      RECT  23250.0 32582.5 23315.0 32717.5 ;
      RECT  23507.5 32482.5 23572.5 32617.5 ;
      RECT  23507.5 32482.5 23572.5 32617.5 ;
      RECT  23955.0 33892.5 24020.0 33957.5 ;
      RECT  23690.0 33892.5 23987.5 33957.5 ;
      RECT  23955.0 33510.0 24020.0 33925.0 ;
      RECT  23765.0 32342.5 23830.0 32407.5 ;
      RECT  23797.5 32342.5 24060.0 32407.5 ;
      RECT  23765.0 32375.0 23830.0 32650.0 ;
      RECT  23765.0 32582.5 23830.0 32717.5 ;
      RECT  23955.0 32582.5 24020.0 32717.5 ;
      RECT  23955.0 32582.5 24020.0 32717.5 ;
      RECT  23765.0 32582.5 23830.0 32717.5 ;
      RECT  23765.0 33442.5 23830.0 33577.5 ;
      RECT  23955.0 33442.5 24020.0 33577.5 ;
      RECT  23955.0 33442.5 24020.0 33577.5 ;
      RECT  23765.0 33442.5 23830.0 33577.5 ;
      RECT  23692.5 33857.5 23757.5 33992.5 ;
      RECT  24027.5 32307.5 24092.5 32442.5 ;
      RECT  23765.0 33442.5 23830.0 33577.5 ;
      RECT  23955.0 32582.5 24020.0 32717.5 ;
      RECT  24212.5 32482.5 24277.5 32617.5 ;
      RECT  24212.5 32482.5 24277.5 32617.5 ;
      RECT  24660.0 33892.5 24725.0 33957.5 ;
      RECT  24395.0 33892.5 24692.5 33957.5 ;
      RECT  24660.0 33510.0 24725.0 33925.0 ;
      RECT  24470.0 32342.5 24535.0 32407.5 ;
      RECT  24502.5 32342.5 24765.0 32407.5 ;
      RECT  24470.0 32375.0 24535.0 32650.0 ;
      RECT  24470.0 32582.5 24535.0 32717.5 ;
      RECT  24660.0 32582.5 24725.0 32717.5 ;
      RECT  24660.0 32582.5 24725.0 32717.5 ;
      RECT  24470.0 32582.5 24535.0 32717.5 ;
      RECT  24470.0 33442.5 24535.0 33577.5 ;
      RECT  24660.0 33442.5 24725.0 33577.5 ;
      RECT  24660.0 33442.5 24725.0 33577.5 ;
      RECT  24470.0 33442.5 24535.0 33577.5 ;
      RECT  24397.5 33857.5 24462.5 33992.5 ;
      RECT  24732.5 32307.5 24797.5 32442.5 ;
      RECT  24470.0 33442.5 24535.0 33577.5 ;
      RECT  24660.0 32582.5 24725.0 32717.5 ;
      RECT  24917.5 32482.5 24982.5 32617.5 ;
      RECT  24917.5 32482.5 24982.5 32617.5 ;
      RECT  25365.0 33892.5 25430.0 33957.5 ;
      RECT  25100.0 33892.5 25397.5 33957.5 ;
      RECT  25365.0 33510.0 25430.0 33925.0 ;
      RECT  25175.0 32342.5 25240.0 32407.5 ;
      RECT  25207.5 32342.5 25470.0 32407.5 ;
      RECT  25175.0 32375.0 25240.0 32650.0 ;
      RECT  25175.0 32582.5 25240.0 32717.5 ;
      RECT  25365.0 32582.5 25430.0 32717.5 ;
      RECT  25365.0 32582.5 25430.0 32717.5 ;
      RECT  25175.0 32582.5 25240.0 32717.5 ;
      RECT  25175.0 33442.5 25240.0 33577.5 ;
      RECT  25365.0 33442.5 25430.0 33577.5 ;
      RECT  25365.0 33442.5 25430.0 33577.5 ;
      RECT  25175.0 33442.5 25240.0 33577.5 ;
      RECT  25102.5 33857.5 25167.5 33992.5 ;
      RECT  25437.5 32307.5 25502.5 32442.5 ;
      RECT  25175.0 33442.5 25240.0 33577.5 ;
      RECT  25365.0 32582.5 25430.0 32717.5 ;
      RECT  25622.5 32482.5 25687.5 32617.5 ;
      RECT  25622.5 32482.5 25687.5 32617.5 ;
      RECT  26070.0 33892.5 26135.0 33957.5 ;
      RECT  25805.0 33892.5 26102.5 33957.5 ;
      RECT  26070.0 33510.0 26135.0 33925.0 ;
      RECT  25880.0 32342.5 25945.0 32407.5 ;
      RECT  25912.5 32342.5 26175.0 32407.5 ;
      RECT  25880.0 32375.0 25945.0 32650.0 ;
      RECT  25880.0 32582.5 25945.0 32717.5 ;
      RECT  26070.0 32582.5 26135.0 32717.5 ;
      RECT  26070.0 32582.5 26135.0 32717.5 ;
      RECT  25880.0 32582.5 25945.0 32717.5 ;
      RECT  25880.0 33442.5 25945.0 33577.5 ;
      RECT  26070.0 33442.5 26135.0 33577.5 ;
      RECT  26070.0 33442.5 26135.0 33577.5 ;
      RECT  25880.0 33442.5 25945.0 33577.5 ;
      RECT  25807.5 33857.5 25872.5 33992.5 ;
      RECT  26142.5 32307.5 26207.5 32442.5 ;
      RECT  25880.0 33442.5 25945.0 33577.5 ;
      RECT  26070.0 32582.5 26135.0 32717.5 ;
      RECT  26327.5 32482.5 26392.5 32617.5 ;
      RECT  26327.5 32482.5 26392.5 32617.5 ;
      RECT  26775.0 33892.5 26840.0 33957.5 ;
      RECT  26510.0 33892.5 26807.5 33957.5 ;
      RECT  26775.0 33510.0 26840.0 33925.0 ;
      RECT  26585.0 32342.5 26650.0 32407.5 ;
      RECT  26617.5 32342.5 26880.0 32407.5 ;
      RECT  26585.0 32375.0 26650.0 32650.0 ;
      RECT  26585.0 32582.5 26650.0 32717.5 ;
      RECT  26775.0 32582.5 26840.0 32717.5 ;
      RECT  26775.0 32582.5 26840.0 32717.5 ;
      RECT  26585.0 32582.5 26650.0 32717.5 ;
      RECT  26585.0 33442.5 26650.0 33577.5 ;
      RECT  26775.0 33442.5 26840.0 33577.5 ;
      RECT  26775.0 33442.5 26840.0 33577.5 ;
      RECT  26585.0 33442.5 26650.0 33577.5 ;
      RECT  26512.5 33857.5 26577.5 33992.5 ;
      RECT  26847.5 32307.5 26912.5 32442.5 ;
      RECT  26585.0 33442.5 26650.0 33577.5 ;
      RECT  26775.0 32582.5 26840.0 32717.5 ;
      RECT  27032.5 32482.5 27097.5 32617.5 ;
      RECT  27032.5 32482.5 27097.5 32617.5 ;
      RECT  27480.0 33892.5 27545.0 33957.5 ;
      RECT  27215.0 33892.5 27512.5 33957.5 ;
      RECT  27480.0 33510.0 27545.0 33925.0 ;
      RECT  27290.0 32342.5 27355.0 32407.5 ;
      RECT  27322.5 32342.5 27585.0 32407.5 ;
      RECT  27290.0 32375.0 27355.0 32650.0 ;
      RECT  27290.0 32582.5 27355.0 32717.5 ;
      RECT  27480.0 32582.5 27545.0 32717.5 ;
      RECT  27480.0 32582.5 27545.0 32717.5 ;
      RECT  27290.0 32582.5 27355.0 32717.5 ;
      RECT  27290.0 33442.5 27355.0 33577.5 ;
      RECT  27480.0 33442.5 27545.0 33577.5 ;
      RECT  27480.0 33442.5 27545.0 33577.5 ;
      RECT  27290.0 33442.5 27355.0 33577.5 ;
      RECT  27217.5 33857.5 27282.5 33992.5 ;
      RECT  27552.5 32307.5 27617.5 32442.5 ;
      RECT  27290.0 33442.5 27355.0 33577.5 ;
      RECT  27480.0 32582.5 27545.0 32717.5 ;
      RECT  27737.5 32482.5 27802.5 32617.5 ;
      RECT  27737.5 32482.5 27802.5 32617.5 ;
      RECT  28185.0 33892.5 28250.0 33957.5 ;
      RECT  27920.0 33892.5 28217.5 33957.5 ;
      RECT  28185.0 33510.0 28250.0 33925.0 ;
      RECT  27995.0 32342.5 28060.0 32407.5 ;
      RECT  28027.5 32342.5 28290.0 32407.5 ;
      RECT  27995.0 32375.0 28060.0 32650.0 ;
      RECT  27995.0 32582.5 28060.0 32717.5 ;
      RECT  28185.0 32582.5 28250.0 32717.5 ;
      RECT  28185.0 32582.5 28250.0 32717.5 ;
      RECT  27995.0 32582.5 28060.0 32717.5 ;
      RECT  27995.0 33442.5 28060.0 33577.5 ;
      RECT  28185.0 33442.5 28250.0 33577.5 ;
      RECT  28185.0 33442.5 28250.0 33577.5 ;
      RECT  27995.0 33442.5 28060.0 33577.5 ;
      RECT  27922.5 33857.5 27987.5 33992.5 ;
      RECT  28257.5 32307.5 28322.5 32442.5 ;
      RECT  27995.0 33442.5 28060.0 33577.5 ;
      RECT  28185.0 32582.5 28250.0 32717.5 ;
      RECT  28442.5 32482.5 28507.5 32617.5 ;
      RECT  28442.5 32482.5 28507.5 32617.5 ;
      RECT  28890.0 33892.5 28955.0 33957.5 ;
      RECT  28625.0 33892.5 28922.5 33957.5 ;
      RECT  28890.0 33510.0 28955.0 33925.0 ;
      RECT  28700.0 32342.5 28765.0 32407.5 ;
      RECT  28732.5 32342.5 28995.0 32407.5 ;
      RECT  28700.0 32375.0 28765.0 32650.0 ;
      RECT  28700.0 32582.5 28765.0 32717.5 ;
      RECT  28890.0 32582.5 28955.0 32717.5 ;
      RECT  28890.0 32582.5 28955.0 32717.5 ;
      RECT  28700.0 32582.5 28765.0 32717.5 ;
      RECT  28700.0 33442.5 28765.0 33577.5 ;
      RECT  28890.0 33442.5 28955.0 33577.5 ;
      RECT  28890.0 33442.5 28955.0 33577.5 ;
      RECT  28700.0 33442.5 28765.0 33577.5 ;
      RECT  28627.5 33857.5 28692.5 33992.5 ;
      RECT  28962.5 32307.5 29027.5 32442.5 ;
      RECT  28700.0 33442.5 28765.0 33577.5 ;
      RECT  28890.0 32582.5 28955.0 32717.5 ;
      RECT  29147.5 32482.5 29212.5 32617.5 ;
      RECT  29147.5 32482.5 29212.5 32617.5 ;
      RECT  29595.0 33892.5 29660.0 33957.5 ;
      RECT  29330.0 33892.5 29627.5 33957.5 ;
      RECT  29595.0 33510.0 29660.0 33925.0 ;
      RECT  29405.0 32342.5 29470.0 32407.5 ;
      RECT  29437.5 32342.5 29700.0 32407.5 ;
      RECT  29405.0 32375.0 29470.0 32650.0 ;
      RECT  29405.0 32582.5 29470.0 32717.5 ;
      RECT  29595.0 32582.5 29660.0 32717.5 ;
      RECT  29595.0 32582.5 29660.0 32717.5 ;
      RECT  29405.0 32582.5 29470.0 32717.5 ;
      RECT  29405.0 33442.5 29470.0 33577.5 ;
      RECT  29595.0 33442.5 29660.0 33577.5 ;
      RECT  29595.0 33442.5 29660.0 33577.5 ;
      RECT  29405.0 33442.5 29470.0 33577.5 ;
      RECT  29332.5 33857.5 29397.5 33992.5 ;
      RECT  29667.5 32307.5 29732.5 32442.5 ;
      RECT  29405.0 33442.5 29470.0 33577.5 ;
      RECT  29595.0 32582.5 29660.0 32717.5 ;
      RECT  29852.5 32482.5 29917.5 32617.5 ;
      RECT  29852.5 32482.5 29917.5 32617.5 ;
      RECT  30300.0 33892.5 30365.0 33957.5 ;
      RECT  30035.0 33892.5 30332.5 33957.5 ;
      RECT  30300.0 33510.0 30365.0 33925.0 ;
      RECT  30110.0 32342.5 30175.0 32407.5 ;
      RECT  30142.5 32342.5 30405.0 32407.5 ;
      RECT  30110.0 32375.0 30175.0 32650.0 ;
      RECT  30110.0 32582.5 30175.0 32717.5 ;
      RECT  30300.0 32582.5 30365.0 32717.5 ;
      RECT  30300.0 32582.5 30365.0 32717.5 ;
      RECT  30110.0 32582.5 30175.0 32717.5 ;
      RECT  30110.0 33442.5 30175.0 33577.5 ;
      RECT  30300.0 33442.5 30365.0 33577.5 ;
      RECT  30300.0 33442.5 30365.0 33577.5 ;
      RECT  30110.0 33442.5 30175.0 33577.5 ;
      RECT  30037.5 33857.5 30102.5 33992.5 ;
      RECT  30372.5 32307.5 30437.5 32442.5 ;
      RECT  30110.0 33442.5 30175.0 33577.5 ;
      RECT  30300.0 32582.5 30365.0 32717.5 ;
      RECT  30557.5 32482.5 30622.5 32617.5 ;
      RECT  30557.5 32482.5 30622.5 32617.5 ;
      RECT  31005.0 33892.5 31070.0 33957.5 ;
      RECT  30740.0 33892.5 31037.5 33957.5 ;
      RECT  31005.0 33510.0 31070.0 33925.0 ;
      RECT  30815.0 32342.5 30880.0 32407.5 ;
      RECT  30847.5 32342.5 31110.0 32407.5 ;
      RECT  30815.0 32375.0 30880.0 32650.0 ;
      RECT  30815.0 32582.5 30880.0 32717.5 ;
      RECT  31005.0 32582.5 31070.0 32717.5 ;
      RECT  31005.0 32582.5 31070.0 32717.5 ;
      RECT  30815.0 32582.5 30880.0 32717.5 ;
      RECT  30815.0 33442.5 30880.0 33577.5 ;
      RECT  31005.0 33442.5 31070.0 33577.5 ;
      RECT  31005.0 33442.5 31070.0 33577.5 ;
      RECT  30815.0 33442.5 30880.0 33577.5 ;
      RECT  30742.5 33857.5 30807.5 33992.5 ;
      RECT  31077.5 32307.5 31142.5 32442.5 ;
      RECT  30815.0 33442.5 30880.0 33577.5 ;
      RECT  31005.0 32582.5 31070.0 32717.5 ;
      RECT  31262.5 32482.5 31327.5 32617.5 ;
      RECT  31262.5 32482.5 31327.5 32617.5 ;
      RECT  31710.0 33892.5 31775.0 33957.5 ;
      RECT  31445.0 33892.5 31742.5 33957.5 ;
      RECT  31710.0 33510.0 31775.0 33925.0 ;
      RECT  31520.0 32342.5 31585.0 32407.5 ;
      RECT  31552.5 32342.5 31815.0 32407.5 ;
      RECT  31520.0 32375.0 31585.0 32650.0 ;
      RECT  31520.0 32582.5 31585.0 32717.5 ;
      RECT  31710.0 32582.5 31775.0 32717.5 ;
      RECT  31710.0 32582.5 31775.0 32717.5 ;
      RECT  31520.0 32582.5 31585.0 32717.5 ;
      RECT  31520.0 33442.5 31585.0 33577.5 ;
      RECT  31710.0 33442.5 31775.0 33577.5 ;
      RECT  31710.0 33442.5 31775.0 33577.5 ;
      RECT  31520.0 33442.5 31585.0 33577.5 ;
      RECT  31447.5 33857.5 31512.5 33992.5 ;
      RECT  31782.5 32307.5 31847.5 32442.5 ;
      RECT  31520.0 33442.5 31585.0 33577.5 ;
      RECT  31710.0 32582.5 31775.0 32717.5 ;
      RECT  31967.5 32482.5 32032.5 32617.5 ;
      RECT  31967.5 32482.5 32032.5 32617.5 ;
      RECT  32415.0 33892.5 32480.0 33957.5 ;
      RECT  32150.0 33892.5 32447.5 33957.5 ;
      RECT  32415.0 33510.0 32480.0 33925.0 ;
      RECT  32225.0 32342.5 32290.0 32407.5 ;
      RECT  32257.5 32342.5 32520.0 32407.5 ;
      RECT  32225.0 32375.0 32290.0 32650.0 ;
      RECT  32225.0 32582.5 32290.0 32717.5 ;
      RECT  32415.0 32582.5 32480.0 32717.5 ;
      RECT  32415.0 32582.5 32480.0 32717.5 ;
      RECT  32225.0 32582.5 32290.0 32717.5 ;
      RECT  32225.0 33442.5 32290.0 33577.5 ;
      RECT  32415.0 33442.5 32480.0 33577.5 ;
      RECT  32415.0 33442.5 32480.0 33577.5 ;
      RECT  32225.0 33442.5 32290.0 33577.5 ;
      RECT  32152.5 33857.5 32217.5 33992.5 ;
      RECT  32487.5 32307.5 32552.5 32442.5 ;
      RECT  32225.0 33442.5 32290.0 33577.5 ;
      RECT  32415.0 32582.5 32480.0 32717.5 ;
      RECT  32672.5 32482.5 32737.5 32617.5 ;
      RECT  32672.5 32482.5 32737.5 32617.5 ;
      RECT  33120.0 33892.5 33185.0 33957.5 ;
      RECT  32855.0 33892.5 33152.5 33957.5 ;
      RECT  33120.0 33510.0 33185.0 33925.0 ;
      RECT  32930.0 32342.5 32995.0 32407.5 ;
      RECT  32962.5 32342.5 33225.0 32407.5 ;
      RECT  32930.0 32375.0 32995.0 32650.0 ;
      RECT  32930.0 32582.5 32995.0 32717.5 ;
      RECT  33120.0 32582.5 33185.0 32717.5 ;
      RECT  33120.0 32582.5 33185.0 32717.5 ;
      RECT  32930.0 32582.5 32995.0 32717.5 ;
      RECT  32930.0 33442.5 32995.0 33577.5 ;
      RECT  33120.0 33442.5 33185.0 33577.5 ;
      RECT  33120.0 33442.5 33185.0 33577.5 ;
      RECT  32930.0 33442.5 32995.0 33577.5 ;
      RECT  32857.5 33857.5 32922.5 33992.5 ;
      RECT  33192.5 32307.5 33257.5 32442.5 ;
      RECT  32930.0 33442.5 32995.0 33577.5 ;
      RECT  33120.0 32582.5 33185.0 32717.5 ;
      RECT  33377.5 32482.5 33442.5 32617.5 ;
      RECT  33377.5 32482.5 33442.5 32617.5 ;
      RECT  33825.0 33892.5 33890.0 33957.5 ;
      RECT  33560.0 33892.5 33857.5 33957.5 ;
      RECT  33825.0 33510.0 33890.0 33925.0 ;
      RECT  33635.0 32342.5 33700.0 32407.5 ;
      RECT  33667.5 32342.5 33930.0 32407.5 ;
      RECT  33635.0 32375.0 33700.0 32650.0 ;
      RECT  33635.0 32582.5 33700.0 32717.5 ;
      RECT  33825.0 32582.5 33890.0 32717.5 ;
      RECT  33825.0 32582.5 33890.0 32717.5 ;
      RECT  33635.0 32582.5 33700.0 32717.5 ;
      RECT  33635.0 33442.5 33700.0 33577.5 ;
      RECT  33825.0 33442.5 33890.0 33577.5 ;
      RECT  33825.0 33442.5 33890.0 33577.5 ;
      RECT  33635.0 33442.5 33700.0 33577.5 ;
      RECT  33562.5 33857.5 33627.5 33992.5 ;
      RECT  33897.5 32307.5 33962.5 32442.5 ;
      RECT  33635.0 33442.5 33700.0 33577.5 ;
      RECT  33825.0 32582.5 33890.0 32717.5 ;
      RECT  34082.5 32482.5 34147.5 32617.5 ;
      RECT  34082.5 32482.5 34147.5 32617.5 ;
      RECT  34530.0 33892.5 34595.0 33957.5 ;
      RECT  34265.0 33892.5 34562.5 33957.5 ;
      RECT  34530.0 33510.0 34595.0 33925.0 ;
      RECT  34340.0 32342.5 34405.0 32407.5 ;
      RECT  34372.5 32342.5 34635.0 32407.5 ;
      RECT  34340.0 32375.0 34405.0 32650.0 ;
      RECT  34340.0 32582.5 34405.0 32717.5 ;
      RECT  34530.0 32582.5 34595.0 32717.5 ;
      RECT  34530.0 32582.5 34595.0 32717.5 ;
      RECT  34340.0 32582.5 34405.0 32717.5 ;
      RECT  34340.0 33442.5 34405.0 33577.5 ;
      RECT  34530.0 33442.5 34595.0 33577.5 ;
      RECT  34530.0 33442.5 34595.0 33577.5 ;
      RECT  34340.0 33442.5 34405.0 33577.5 ;
      RECT  34267.5 33857.5 34332.5 33992.5 ;
      RECT  34602.5 32307.5 34667.5 32442.5 ;
      RECT  34340.0 33442.5 34405.0 33577.5 ;
      RECT  34530.0 32582.5 34595.0 32717.5 ;
      RECT  34787.5 32482.5 34852.5 32617.5 ;
      RECT  34787.5 32482.5 34852.5 32617.5 ;
      RECT  35235.0 33892.5 35300.0 33957.5 ;
      RECT  34970.0 33892.5 35267.5 33957.5 ;
      RECT  35235.0 33510.0 35300.0 33925.0 ;
      RECT  35045.0 32342.5 35110.0 32407.5 ;
      RECT  35077.5 32342.5 35340.0 32407.5 ;
      RECT  35045.0 32375.0 35110.0 32650.0 ;
      RECT  35045.0 32582.5 35110.0 32717.5 ;
      RECT  35235.0 32582.5 35300.0 32717.5 ;
      RECT  35235.0 32582.5 35300.0 32717.5 ;
      RECT  35045.0 32582.5 35110.0 32717.5 ;
      RECT  35045.0 33442.5 35110.0 33577.5 ;
      RECT  35235.0 33442.5 35300.0 33577.5 ;
      RECT  35235.0 33442.5 35300.0 33577.5 ;
      RECT  35045.0 33442.5 35110.0 33577.5 ;
      RECT  34972.5 33857.5 35037.5 33992.5 ;
      RECT  35307.5 32307.5 35372.5 32442.5 ;
      RECT  35045.0 33442.5 35110.0 33577.5 ;
      RECT  35235.0 32582.5 35300.0 32717.5 ;
      RECT  35492.5 32482.5 35557.5 32617.5 ;
      RECT  35492.5 32482.5 35557.5 32617.5 ;
      RECT  35940.0 33892.5 36005.0 33957.5 ;
      RECT  35675.0 33892.5 35972.5 33957.5 ;
      RECT  35940.0 33510.0 36005.0 33925.0 ;
      RECT  35750.0 32342.5 35815.0 32407.5 ;
      RECT  35782.5 32342.5 36045.0 32407.5 ;
      RECT  35750.0 32375.0 35815.0 32650.0 ;
      RECT  35750.0 32582.5 35815.0 32717.5 ;
      RECT  35940.0 32582.5 36005.0 32717.5 ;
      RECT  35940.0 32582.5 36005.0 32717.5 ;
      RECT  35750.0 32582.5 35815.0 32717.5 ;
      RECT  35750.0 33442.5 35815.0 33577.5 ;
      RECT  35940.0 33442.5 36005.0 33577.5 ;
      RECT  35940.0 33442.5 36005.0 33577.5 ;
      RECT  35750.0 33442.5 35815.0 33577.5 ;
      RECT  35677.5 33857.5 35742.5 33992.5 ;
      RECT  36012.5 32307.5 36077.5 32442.5 ;
      RECT  35750.0 33442.5 35815.0 33577.5 ;
      RECT  35940.0 32582.5 36005.0 32717.5 ;
      RECT  36197.5 32482.5 36262.5 32617.5 ;
      RECT  36197.5 32482.5 36262.5 32617.5 ;
      RECT  36645.0 33892.5 36710.0 33957.5 ;
      RECT  36380.0 33892.5 36677.5 33957.5 ;
      RECT  36645.0 33510.0 36710.0 33925.0 ;
      RECT  36455.0 32342.5 36520.0 32407.5 ;
      RECT  36487.5 32342.5 36750.0 32407.5 ;
      RECT  36455.0 32375.0 36520.0 32650.0 ;
      RECT  36455.0 32582.5 36520.0 32717.5 ;
      RECT  36645.0 32582.5 36710.0 32717.5 ;
      RECT  36645.0 32582.5 36710.0 32717.5 ;
      RECT  36455.0 32582.5 36520.0 32717.5 ;
      RECT  36455.0 33442.5 36520.0 33577.5 ;
      RECT  36645.0 33442.5 36710.0 33577.5 ;
      RECT  36645.0 33442.5 36710.0 33577.5 ;
      RECT  36455.0 33442.5 36520.0 33577.5 ;
      RECT  36382.5 33857.5 36447.5 33992.5 ;
      RECT  36717.5 32307.5 36782.5 32442.5 ;
      RECT  36455.0 33442.5 36520.0 33577.5 ;
      RECT  36645.0 32582.5 36710.0 32717.5 ;
      RECT  36902.5 32482.5 36967.5 32617.5 ;
      RECT  36902.5 32482.5 36967.5 32617.5 ;
      RECT  37350.0 33892.5 37415.0 33957.5 ;
      RECT  37085.0 33892.5 37382.5 33957.5 ;
      RECT  37350.0 33510.0 37415.0 33925.0 ;
      RECT  37160.0 32342.5 37225.0 32407.5 ;
      RECT  37192.5 32342.5 37455.0 32407.5 ;
      RECT  37160.0 32375.0 37225.0 32650.0 ;
      RECT  37160.0 32582.5 37225.0 32717.5 ;
      RECT  37350.0 32582.5 37415.0 32717.5 ;
      RECT  37350.0 32582.5 37415.0 32717.5 ;
      RECT  37160.0 32582.5 37225.0 32717.5 ;
      RECT  37160.0 33442.5 37225.0 33577.5 ;
      RECT  37350.0 33442.5 37415.0 33577.5 ;
      RECT  37350.0 33442.5 37415.0 33577.5 ;
      RECT  37160.0 33442.5 37225.0 33577.5 ;
      RECT  37087.5 33857.5 37152.5 33992.5 ;
      RECT  37422.5 32307.5 37487.5 32442.5 ;
      RECT  37160.0 33442.5 37225.0 33577.5 ;
      RECT  37350.0 32582.5 37415.0 32717.5 ;
      RECT  37607.5 32482.5 37672.5 32617.5 ;
      RECT  37607.5 32482.5 37672.5 32617.5 ;
      RECT  38055.0 33892.5 38120.0 33957.5 ;
      RECT  37790.0 33892.5 38087.5 33957.5 ;
      RECT  38055.0 33510.0 38120.0 33925.0 ;
      RECT  37865.0 32342.5 37930.0 32407.5 ;
      RECT  37897.5 32342.5 38160.0 32407.5 ;
      RECT  37865.0 32375.0 37930.0 32650.0 ;
      RECT  37865.0 32582.5 37930.0 32717.5 ;
      RECT  38055.0 32582.5 38120.0 32717.5 ;
      RECT  38055.0 32582.5 38120.0 32717.5 ;
      RECT  37865.0 32582.5 37930.0 32717.5 ;
      RECT  37865.0 33442.5 37930.0 33577.5 ;
      RECT  38055.0 33442.5 38120.0 33577.5 ;
      RECT  38055.0 33442.5 38120.0 33577.5 ;
      RECT  37865.0 33442.5 37930.0 33577.5 ;
      RECT  37792.5 33857.5 37857.5 33992.5 ;
      RECT  38127.5 32307.5 38192.5 32442.5 ;
      RECT  37865.0 33442.5 37930.0 33577.5 ;
      RECT  38055.0 32582.5 38120.0 32717.5 ;
      RECT  38312.5 32482.5 38377.5 32617.5 ;
      RECT  38312.5 32482.5 38377.5 32617.5 ;
      RECT  38760.0 33892.5 38825.0 33957.5 ;
      RECT  38495.0 33892.5 38792.5 33957.5 ;
      RECT  38760.0 33510.0 38825.0 33925.0 ;
      RECT  38570.0 32342.5 38635.0 32407.5 ;
      RECT  38602.5 32342.5 38865.0 32407.5 ;
      RECT  38570.0 32375.0 38635.0 32650.0 ;
      RECT  38570.0 32582.5 38635.0 32717.5 ;
      RECT  38760.0 32582.5 38825.0 32717.5 ;
      RECT  38760.0 32582.5 38825.0 32717.5 ;
      RECT  38570.0 32582.5 38635.0 32717.5 ;
      RECT  38570.0 33442.5 38635.0 33577.5 ;
      RECT  38760.0 33442.5 38825.0 33577.5 ;
      RECT  38760.0 33442.5 38825.0 33577.5 ;
      RECT  38570.0 33442.5 38635.0 33577.5 ;
      RECT  38497.5 33857.5 38562.5 33992.5 ;
      RECT  38832.5 32307.5 38897.5 32442.5 ;
      RECT  38570.0 33442.5 38635.0 33577.5 ;
      RECT  38760.0 32582.5 38825.0 32717.5 ;
      RECT  39017.5 32482.5 39082.5 32617.5 ;
      RECT  39017.5 32482.5 39082.5 32617.5 ;
      RECT  39465.0 33892.5 39530.0 33957.5 ;
      RECT  39200.0 33892.5 39497.5 33957.5 ;
      RECT  39465.0 33510.0 39530.0 33925.0 ;
      RECT  39275.0 32342.5 39340.0 32407.5 ;
      RECT  39307.5 32342.5 39570.0 32407.5 ;
      RECT  39275.0 32375.0 39340.0 32650.0 ;
      RECT  39275.0 32582.5 39340.0 32717.5 ;
      RECT  39465.0 32582.5 39530.0 32717.5 ;
      RECT  39465.0 32582.5 39530.0 32717.5 ;
      RECT  39275.0 32582.5 39340.0 32717.5 ;
      RECT  39275.0 33442.5 39340.0 33577.5 ;
      RECT  39465.0 33442.5 39530.0 33577.5 ;
      RECT  39465.0 33442.5 39530.0 33577.5 ;
      RECT  39275.0 33442.5 39340.0 33577.5 ;
      RECT  39202.5 33857.5 39267.5 33992.5 ;
      RECT  39537.5 32307.5 39602.5 32442.5 ;
      RECT  39275.0 33442.5 39340.0 33577.5 ;
      RECT  39465.0 32582.5 39530.0 32717.5 ;
      RECT  39722.5 32482.5 39787.5 32617.5 ;
      RECT  39722.5 32482.5 39787.5 32617.5 ;
      RECT  40170.0 33892.5 40235.0 33957.5 ;
      RECT  39905.0 33892.5 40202.5 33957.5 ;
      RECT  40170.0 33510.0 40235.0 33925.0 ;
      RECT  39980.0 32342.5 40045.0 32407.5 ;
      RECT  40012.5 32342.5 40275.0 32407.5 ;
      RECT  39980.0 32375.0 40045.0 32650.0 ;
      RECT  39980.0 32582.5 40045.0 32717.5 ;
      RECT  40170.0 32582.5 40235.0 32717.5 ;
      RECT  40170.0 32582.5 40235.0 32717.5 ;
      RECT  39980.0 32582.5 40045.0 32717.5 ;
      RECT  39980.0 33442.5 40045.0 33577.5 ;
      RECT  40170.0 33442.5 40235.0 33577.5 ;
      RECT  40170.0 33442.5 40235.0 33577.5 ;
      RECT  39980.0 33442.5 40045.0 33577.5 ;
      RECT  39907.5 33857.5 39972.5 33992.5 ;
      RECT  40242.5 32307.5 40307.5 32442.5 ;
      RECT  39980.0 33442.5 40045.0 33577.5 ;
      RECT  40170.0 32582.5 40235.0 32717.5 ;
      RECT  40427.5 32482.5 40492.5 32617.5 ;
      RECT  40427.5 32482.5 40492.5 32617.5 ;
      RECT  40875.0 33892.5 40940.0 33957.5 ;
      RECT  40610.0 33892.5 40907.5 33957.5 ;
      RECT  40875.0 33510.0 40940.0 33925.0 ;
      RECT  40685.0 32342.5 40750.0 32407.5 ;
      RECT  40717.5 32342.5 40980.0 32407.5 ;
      RECT  40685.0 32375.0 40750.0 32650.0 ;
      RECT  40685.0 32582.5 40750.0 32717.5 ;
      RECT  40875.0 32582.5 40940.0 32717.5 ;
      RECT  40875.0 32582.5 40940.0 32717.5 ;
      RECT  40685.0 32582.5 40750.0 32717.5 ;
      RECT  40685.0 33442.5 40750.0 33577.5 ;
      RECT  40875.0 33442.5 40940.0 33577.5 ;
      RECT  40875.0 33442.5 40940.0 33577.5 ;
      RECT  40685.0 33442.5 40750.0 33577.5 ;
      RECT  40612.5 33857.5 40677.5 33992.5 ;
      RECT  40947.5 32307.5 41012.5 32442.5 ;
      RECT  40685.0 33442.5 40750.0 33577.5 ;
      RECT  40875.0 32582.5 40940.0 32717.5 ;
      RECT  41132.5 32482.5 41197.5 32617.5 ;
      RECT  41132.5 32482.5 41197.5 32617.5 ;
      RECT  41580.0 33892.5 41645.0 33957.5 ;
      RECT  41315.0 33892.5 41612.5 33957.5 ;
      RECT  41580.0 33510.0 41645.0 33925.0 ;
      RECT  41390.0 32342.5 41455.0 32407.5 ;
      RECT  41422.5 32342.5 41685.0 32407.5 ;
      RECT  41390.0 32375.0 41455.0 32650.0 ;
      RECT  41390.0 32582.5 41455.0 32717.5 ;
      RECT  41580.0 32582.5 41645.0 32717.5 ;
      RECT  41580.0 32582.5 41645.0 32717.5 ;
      RECT  41390.0 32582.5 41455.0 32717.5 ;
      RECT  41390.0 33442.5 41455.0 33577.5 ;
      RECT  41580.0 33442.5 41645.0 33577.5 ;
      RECT  41580.0 33442.5 41645.0 33577.5 ;
      RECT  41390.0 33442.5 41455.0 33577.5 ;
      RECT  41317.5 33857.5 41382.5 33992.5 ;
      RECT  41652.5 32307.5 41717.5 32442.5 ;
      RECT  41390.0 33442.5 41455.0 33577.5 ;
      RECT  41580.0 32582.5 41645.0 32717.5 ;
      RECT  41837.5 32482.5 41902.5 32617.5 ;
      RECT  41837.5 32482.5 41902.5 32617.5 ;
      RECT  42285.0 33892.5 42350.0 33957.5 ;
      RECT  42020.0 33892.5 42317.5 33957.5 ;
      RECT  42285.0 33510.0 42350.0 33925.0 ;
      RECT  42095.0 32342.5 42160.0 32407.5 ;
      RECT  42127.5 32342.5 42390.0 32407.5 ;
      RECT  42095.0 32375.0 42160.0 32650.0 ;
      RECT  42095.0 32582.5 42160.0 32717.5 ;
      RECT  42285.0 32582.5 42350.0 32717.5 ;
      RECT  42285.0 32582.5 42350.0 32717.5 ;
      RECT  42095.0 32582.5 42160.0 32717.5 ;
      RECT  42095.0 33442.5 42160.0 33577.5 ;
      RECT  42285.0 33442.5 42350.0 33577.5 ;
      RECT  42285.0 33442.5 42350.0 33577.5 ;
      RECT  42095.0 33442.5 42160.0 33577.5 ;
      RECT  42022.5 33857.5 42087.5 33992.5 ;
      RECT  42357.5 32307.5 42422.5 32442.5 ;
      RECT  42095.0 33442.5 42160.0 33577.5 ;
      RECT  42285.0 32582.5 42350.0 32717.5 ;
      RECT  42542.5 32482.5 42607.5 32617.5 ;
      RECT  42542.5 32482.5 42607.5 32617.5 ;
      RECT  42990.0 33892.5 43055.0 33957.5 ;
      RECT  42725.0 33892.5 43022.5 33957.5 ;
      RECT  42990.0 33510.0 43055.0 33925.0 ;
      RECT  42800.0 32342.5 42865.0 32407.5 ;
      RECT  42832.5 32342.5 43095.0 32407.5 ;
      RECT  42800.0 32375.0 42865.0 32650.0 ;
      RECT  42800.0 32582.5 42865.0 32717.5 ;
      RECT  42990.0 32582.5 43055.0 32717.5 ;
      RECT  42990.0 32582.5 43055.0 32717.5 ;
      RECT  42800.0 32582.5 42865.0 32717.5 ;
      RECT  42800.0 33442.5 42865.0 33577.5 ;
      RECT  42990.0 33442.5 43055.0 33577.5 ;
      RECT  42990.0 33442.5 43055.0 33577.5 ;
      RECT  42800.0 33442.5 42865.0 33577.5 ;
      RECT  42727.5 33857.5 42792.5 33992.5 ;
      RECT  43062.5 32307.5 43127.5 32442.5 ;
      RECT  42800.0 33442.5 42865.0 33577.5 ;
      RECT  42990.0 32582.5 43055.0 32717.5 ;
      RECT  43247.5 32482.5 43312.5 32617.5 ;
      RECT  43247.5 32482.5 43312.5 32617.5 ;
      RECT  43695.0 33892.5 43760.0 33957.5 ;
      RECT  43430.0 33892.5 43727.5 33957.5 ;
      RECT  43695.0 33510.0 43760.0 33925.0 ;
      RECT  43505.0 32342.5 43570.0 32407.5 ;
      RECT  43537.5 32342.5 43800.0 32407.5 ;
      RECT  43505.0 32375.0 43570.0 32650.0 ;
      RECT  43505.0 32582.5 43570.0 32717.5 ;
      RECT  43695.0 32582.5 43760.0 32717.5 ;
      RECT  43695.0 32582.5 43760.0 32717.5 ;
      RECT  43505.0 32582.5 43570.0 32717.5 ;
      RECT  43505.0 33442.5 43570.0 33577.5 ;
      RECT  43695.0 33442.5 43760.0 33577.5 ;
      RECT  43695.0 33442.5 43760.0 33577.5 ;
      RECT  43505.0 33442.5 43570.0 33577.5 ;
      RECT  43432.5 33857.5 43497.5 33992.5 ;
      RECT  43767.5 32307.5 43832.5 32442.5 ;
      RECT  43505.0 33442.5 43570.0 33577.5 ;
      RECT  43695.0 32582.5 43760.0 32717.5 ;
      RECT  43952.5 32482.5 44017.5 32617.5 ;
      RECT  43952.5 32482.5 44017.5 32617.5 ;
      RECT  44400.0 33892.5 44465.0 33957.5 ;
      RECT  44135.0 33892.5 44432.5 33957.5 ;
      RECT  44400.0 33510.0 44465.0 33925.0 ;
      RECT  44210.0 32342.5 44275.0 32407.5 ;
      RECT  44242.5 32342.5 44505.0 32407.5 ;
      RECT  44210.0 32375.0 44275.0 32650.0 ;
      RECT  44210.0 32582.5 44275.0 32717.5 ;
      RECT  44400.0 32582.5 44465.0 32717.5 ;
      RECT  44400.0 32582.5 44465.0 32717.5 ;
      RECT  44210.0 32582.5 44275.0 32717.5 ;
      RECT  44210.0 33442.5 44275.0 33577.5 ;
      RECT  44400.0 33442.5 44465.0 33577.5 ;
      RECT  44400.0 33442.5 44465.0 33577.5 ;
      RECT  44210.0 33442.5 44275.0 33577.5 ;
      RECT  44137.5 33857.5 44202.5 33992.5 ;
      RECT  44472.5 32307.5 44537.5 32442.5 ;
      RECT  44210.0 33442.5 44275.0 33577.5 ;
      RECT  44400.0 32582.5 44465.0 32717.5 ;
      RECT  44657.5 32482.5 44722.5 32617.5 ;
      RECT  44657.5 32482.5 44722.5 32617.5 ;
      RECT  45105.0 33892.5 45170.0 33957.5 ;
      RECT  44840.0 33892.5 45137.5 33957.5 ;
      RECT  45105.0 33510.0 45170.0 33925.0 ;
      RECT  44915.0 32342.5 44980.0 32407.5 ;
      RECT  44947.5 32342.5 45210.0 32407.5 ;
      RECT  44915.0 32375.0 44980.0 32650.0 ;
      RECT  44915.0 32582.5 44980.0 32717.5 ;
      RECT  45105.0 32582.5 45170.0 32717.5 ;
      RECT  45105.0 32582.5 45170.0 32717.5 ;
      RECT  44915.0 32582.5 44980.0 32717.5 ;
      RECT  44915.0 33442.5 44980.0 33577.5 ;
      RECT  45105.0 33442.5 45170.0 33577.5 ;
      RECT  45105.0 33442.5 45170.0 33577.5 ;
      RECT  44915.0 33442.5 44980.0 33577.5 ;
      RECT  44842.5 33857.5 44907.5 33992.5 ;
      RECT  45177.5 32307.5 45242.5 32442.5 ;
      RECT  44915.0 33442.5 44980.0 33577.5 ;
      RECT  45105.0 32582.5 45170.0 32717.5 ;
      RECT  45362.5 32482.5 45427.5 32617.5 ;
      RECT  45362.5 32482.5 45427.5 32617.5 ;
      RECT  45810.0 33892.5 45875.0 33957.5 ;
      RECT  45545.0 33892.5 45842.5 33957.5 ;
      RECT  45810.0 33510.0 45875.0 33925.0 ;
      RECT  45620.0 32342.5 45685.0 32407.5 ;
      RECT  45652.5 32342.5 45915.0 32407.5 ;
      RECT  45620.0 32375.0 45685.0 32650.0 ;
      RECT  45620.0 32582.5 45685.0 32717.5 ;
      RECT  45810.0 32582.5 45875.0 32717.5 ;
      RECT  45810.0 32582.5 45875.0 32717.5 ;
      RECT  45620.0 32582.5 45685.0 32717.5 ;
      RECT  45620.0 33442.5 45685.0 33577.5 ;
      RECT  45810.0 33442.5 45875.0 33577.5 ;
      RECT  45810.0 33442.5 45875.0 33577.5 ;
      RECT  45620.0 33442.5 45685.0 33577.5 ;
      RECT  45547.5 33857.5 45612.5 33992.5 ;
      RECT  45882.5 32307.5 45947.5 32442.5 ;
      RECT  45620.0 33442.5 45685.0 33577.5 ;
      RECT  45810.0 32582.5 45875.0 32717.5 ;
      RECT  46067.5 32482.5 46132.5 32617.5 ;
      RECT  46067.5 32482.5 46132.5 32617.5 ;
      RECT  46515.0 33892.5 46580.0 33957.5 ;
      RECT  46250.0 33892.5 46547.5 33957.5 ;
      RECT  46515.0 33510.0 46580.0 33925.0 ;
      RECT  46325.0 32342.5 46390.0 32407.5 ;
      RECT  46357.5 32342.5 46620.0 32407.5 ;
      RECT  46325.0 32375.0 46390.0 32650.0 ;
      RECT  46325.0 32582.5 46390.0 32717.5 ;
      RECT  46515.0 32582.5 46580.0 32717.5 ;
      RECT  46515.0 32582.5 46580.0 32717.5 ;
      RECT  46325.0 32582.5 46390.0 32717.5 ;
      RECT  46325.0 33442.5 46390.0 33577.5 ;
      RECT  46515.0 33442.5 46580.0 33577.5 ;
      RECT  46515.0 33442.5 46580.0 33577.5 ;
      RECT  46325.0 33442.5 46390.0 33577.5 ;
      RECT  46252.5 33857.5 46317.5 33992.5 ;
      RECT  46587.5 32307.5 46652.5 32442.5 ;
      RECT  46325.0 33442.5 46390.0 33577.5 ;
      RECT  46515.0 32582.5 46580.0 32717.5 ;
      RECT  46772.5 32482.5 46837.5 32617.5 ;
      RECT  46772.5 32482.5 46837.5 32617.5 ;
      RECT  47220.0 33892.5 47285.0 33957.5 ;
      RECT  46955.0 33892.5 47252.5 33957.5 ;
      RECT  47220.0 33510.0 47285.0 33925.0 ;
      RECT  47030.0 32342.5 47095.0 32407.5 ;
      RECT  47062.5 32342.5 47325.0 32407.5 ;
      RECT  47030.0 32375.0 47095.0 32650.0 ;
      RECT  47030.0 32582.5 47095.0 32717.5 ;
      RECT  47220.0 32582.5 47285.0 32717.5 ;
      RECT  47220.0 32582.5 47285.0 32717.5 ;
      RECT  47030.0 32582.5 47095.0 32717.5 ;
      RECT  47030.0 33442.5 47095.0 33577.5 ;
      RECT  47220.0 33442.5 47285.0 33577.5 ;
      RECT  47220.0 33442.5 47285.0 33577.5 ;
      RECT  47030.0 33442.5 47095.0 33577.5 ;
      RECT  46957.5 33857.5 47022.5 33992.5 ;
      RECT  47292.5 32307.5 47357.5 32442.5 ;
      RECT  47030.0 33442.5 47095.0 33577.5 ;
      RECT  47220.0 32582.5 47285.0 32717.5 ;
      RECT  47477.5 32482.5 47542.5 32617.5 ;
      RECT  47477.5 32482.5 47542.5 32617.5 ;
      RECT  47925.0 33892.5 47990.0 33957.5 ;
      RECT  47660.0 33892.5 47957.5 33957.5 ;
      RECT  47925.0 33510.0 47990.0 33925.0 ;
      RECT  47735.0 32342.5 47800.0 32407.5 ;
      RECT  47767.5 32342.5 48030.0 32407.5 ;
      RECT  47735.0 32375.0 47800.0 32650.0 ;
      RECT  47735.0 32582.5 47800.0 32717.5 ;
      RECT  47925.0 32582.5 47990.0 32717.5 ;
      RECT  47925.0 32582.5 47990.0 32717.5 ;
      RECT  47735.0 32582.5 47800.0 32717.5 ;
      RECT  47735.0 33442.5 47800.0 33577.5 ;
      RECT  47925.0 33442.5 47990.0 33577.5 ;
      RECT  47925.0 33442.5 47990.0 33577.5 ;
      RECT  47735.0 33442.5 47800.0 33577.5 ;
      RECT  47662.5 33857.5 47727.5 33992.5 ;
      RECT  47997.5 32307.5 48062.5 32442.5 ;
      RECT  47735.0 33442.5 47800.0 33577.5 ;
      RECT  47925.0 32582.5 47990.0 32717.5 ;
      RECT  48182.5 32482.5 48247.5 32617.5 ;
      RECT  48182.5 32482.5 48247.5 32617.5 ;
      RECT  48630.0 33892.5 48695.0 33957.5 ;
      RECT  48365.0 33892.5 48662.5 33957.5 ;
      RECT  48630.0 33510.0 48695.0 33925.0 ;
      RECT  48440.0 32342.5 48505.0 32407.5 ;
      RECT  48472.5 32342.5 48735.0 32407.5 ;
      RECT  48440.0 32375.0 48505.0 32650.0 ;
      RECT  48440.0 32582.5 48505.0 32717.5 ;
      RECT  48630.0 32582.5 48695.0 32717.5 ;
      RECT  48630.0 32582.5 48695.0 32717.5 ;
      RECT  48440.0 32582.5 48505.0 32717.5 ;
      RECT  48440.0 33442.5 48505.0 33577.5 ;
      RECT  48630.0 33442.5 48695.0 33577.5 ;
      RECT  48630.0 33442.5 48695.0 33577.5 ;
      RECT  48440.0 33442.5 48505.0 33577.5 ;
      RECT  48367.5 33857.5 48432.5 33992.5 ;
      RECT  48702.5 32307.5 48767.5 32442.5 ;
      RECT  48440.0 33442.5 48505.0 33577.5 ;
      RECT  48630.0 32582.5 48695.0 32717.5 ;
      RECT  48887.5 32482.5 48952.5 32617.5 ;
      RECT  48887.5 32482.5 48952.5 32617.5 ;
      RECT  49335.0 33892.5 49400.0 33957.5 ;
      RECT  49070.0 33892.5 49367.5 33957.5 ;
      RECT  49335.0 33510.0 49400.0 33925.0 ;
      RECT  49145.0 32342.5 49210.0 32407.5 ;
      RECT  49177.5 32342.5 49440.0 32407.5 ;
      RECT  49145.0 32375.0 49210.0 32650.0 ;
      RECT  49145.0 32582.5 49210.0 32717.5 ;
      RECT  49335.0 32582.5 49400.0 32717.5 ;
      RECT  49335.0 32582.5 49400.0 32717.5 ;
      RECT  49145.0 32582.5 49210.0 32717.5 ;
      RECT  49145.0 33442.5 49210.0 33577.5 ;
      RECT  49335.0 33442.5 49400.0 33577.5 ;
      RECT  49335.0 33442.5 49400.0 33577.5 ;
      RECT  49145.0 33442.5 49210.0 33577.5 ;
      RECT  49072.5 33857.5 49137.5 33992.5 ;
      RECT  49407.5 32307.5 49472.5 32442.5 ;
      RECT  49145.0 33442.5 49210.0 33577.5 ;
      RECT  49335.0 32582.5 49400.0 32717.5 ;
      RECT  49592.5 32482.5 49657.5 32617.5 ;
      RECT  49592.5 32482.5 49657.5 32617.5 ;
      RECT  50040.0 33892.5 50105.0 33957.5 ;
      RECT  49775.0 33892.5 50072.5 33957.5 ;
      RECT  50040.0 33510.0 50105.0 33925.0 ;
      RECT  49850.0 32342.5 49915.0 32407.5 ;
      RECT  49882.5 32342.5 50145.0 32407.5 ;
      RECT  49850.0 32375.0 49915.0 32650.0 ;
      RECT  49850.0 32582.5 49915.0 32717.5 ;
      RECT  50040.0 32582.5 50105.0 32717.5 ;
      RECT  50040.0 32582.5 50105.0 32717.5 ;
      RECT  49850.0 32582.5 49915.0 32717.5 ;
      RECT  49850.0 33442.5 49915.0 33577.5 ;
      RECT  50040.0 33442.5 50105.0 33577.5 ;
      RECT  50040.0 33442.5 50105.0 33577.5 ;
      RECT  49850.0 33442.5 49915.0 33577.5 ;
      RECT  49777.5 33857.5 49842.5 33992.5 ;
      RECT  50112.5 32307.5 50177.5 32442.5 ;
      RECT  49850.0 33442.5 49915.0 33577.5 ;
      RECT  50040.0 32582.5 50105.0 32717.5 ;
      RECT  50297.5 32482.5 50362.5 32617.5 ;
      RECT  50297.5 32482.5 50362.5 32617.5 ;
      RECT  50745.0 33892.5 50810.0 33957.5 ;
      RECT  50480.0 33892.5 50777.5 33957.5 ;
      RECT  50745.0 33510.0 50810.0 33925.0 ;
      RECT  50555.0 32342.5 50620.0 32407.5 ;
      RECT  50587.5 32342.5 50850.0 32407.5 ;
      RECT  50555.0 32375.0 50620.0 32650.0 ;
      RECT  50555.0 32582.5 50620.0 32717.5 ;
      RECT  50745.0 32582.5 50810.0 32717.5 ;
      RECT  50745.0 32582.5 50810.0 32717.5 ;
      RECT  50555.0 32582.5 50620.0 32717.5 ;
      RECT  50555.0 33442.5 50620.0 33577.5 ;
      RECT  50745.0 33442.5 50810.0 33577.5 ;
      RECT  50745.0 33442.5 50810.0 33577.5 ;
      RECT  50555.0 33442.5 50620.0 33577.5 ;
      RECT  50482.5 33857.5 50547.5 33992.5 ;
      RECT  50817.5 32307.5 50882.5 32442.5 ;
      RECT  50555.0 33442.5 50620.0 33577.5 ;
      RECT  50745.0 32582.5 50810.0 32717.5 ;
      RECT  51002.5 32482.5 51067.5 32617.5 ;
      RECT  51002.5 32482.5 51067.5 32617.5 ;
      RECT  51450.0 33892.5 51515.0 33957.5 ;
      RECT  51185.0 33892.5 51482.5 33957.5 ;
      RECT  51450.0 33510.0 51515.0 33925.0 ;
      RECT  51260.0 32342.5 51325.0 32407.5 ;
      RECT  51292.5 32342.5 51555.0 32407.5 ;
      RECT  51260.0 32375.0 51325.0 32650.0 ;
      RECT  51260.0 32582.5 51325.0 32717.5 ;
      RECT  51450.0 32582.5 51515.0 32717.5 ;
      RECT  51450.0 32582.5 51515.0 32717.5 ;
      RECT  51260.0 32582.5 51325.0 32717.5 ;
      RECT  51260.0 33442.5 51325.0 33577.5 ;
      RECT  51450.0 33442.5 51515.0 33577.5 ;
      RECT  51450.0 33442.5 51515.0 33577.5 ;
      RECT  51260.0 33442.5 51325.0 33577.5 ;
      RECT  51187.5 33857.5 51252.5 33992.5 ;
      RECT  51522.5 32307.5 51587.5 32442.5 ;
      RECT  51260.0 33442.5 51325.0 33577.5 ;
      RECT  51450.0 32582.5 51515.0 32717.5 ;
      RECT  51707.5 32482.5 51772.5 32617.5 ;
      RECT  51707.5 32482.5 51772.5 32617.5 ;
      RECT  52155.0 33892.5 52220.0 33957.5 ;
      RECT  51890.0 33892.5 52187.5 33957.5 ;
      RECT  52155.0 33510.0 52220.0 33925.0 ;
      RECT  51965.0 32342.5 52030.0 32407.5 ;
      RECT  51997.5 32342.5 52260.0 32407.5 ;
      RECT  51965.0 32375.0 52030.0 32650.0 ;
      RECT  51965.0 32582.5 52030.0 32717.5 ;
      RECT  52155.0 32582.5 52220.0 32717.5 ;
      RECT  52155.0 32582.5 52220.0 32717.5 ;
      RECT  51965.0 32582.5 52030.0 32717.5 ;
      RECT  51965.0 33442.5 52030.0 33577.5 ;
      RECT  52155.0 33442.5 52220.0 33577.5 ;
      RECT  52155.0 33442.5 52220.0 33577.5 ;
      RECT  51965.0 33442.5 52030.0 33577.5 ;
      RECT  51892.5 33857.5 51957.5 33992.5 ;
      RECT  52227.5 32307.5 52292.5 32442.5 ;
      RECT  51965.0 33442.5 52030.0 33577.5 ;
      RECT  52155.0 32582.5 52220.0 32717.5 ;
      RECT  52412.5 32482.5 52477.5 32617.5 ;
      RECT  52412.5 32482.5 52477.5 32617.5 ;
      RECT  52860.0 33892.5 52925.0 33957.5 ;
      RECT  52595.0 33892.5 52892.5 33957.5 ;
      RECT  52860.0 33510.0 52925.0 33925.0 ;
      RECT  52670.0 32342.5 52735.0 32407.5 ;
      RECT  52702.5 32342.5 52965.0 32407.5 ;
      RECT  52670.0 32375.0 52735.0 32650.0 ;
      RECT  52670.0 32582.5 52735.0 32717.5 ;
      RECT  52860.0 32582.5 52925.0 32717.5 ;
      RECT  52860.0 32582.5 52925.0 32717.5 ;
      RECT  52670.0 32582.5 52735.0 32717.5 ;
      RECT  52670.0 33442.5 52735.0 33577.5 ;
      RECT  52860.0 33442.5 52925.0 33577.5 ;
      RECT  52860.0 33442.5 52925.0 33577.5 ;
      RECT  52670.0 33442.5 52735.0 33577.5 ;
      RECT  52597.5 33857.5 52662.5 33992.5 ;
      RECT  52932.5 32307.5 52997.5 32442.5 ;
      RECT  52670.0 33442.5 52735.0 33577.5 ;
      RECT  52860.0 32582.5 52925.0 32717.5 ;
      RECT  53117.5 32482.5 53182.5 32617.5 ;
      RECT  53117.5 32482.5 53182.5 32617.5 ;
      RECT  53565.0 33892.5 53630.0 33957.5 ;
      RECT  53300.0 33892.5 53597.5 33957.5 ;
      RECT  53565.0 33510.0 53630.0 33925.0 ;
      RECT  53375.0 32342.5 53440.0 32407.5 ;
      RECT  53407.5 32342.5 53670.0 32407.5 ;
      RECT  53375.0 32375.0 53440.0 32650.0 ;
      RECT  53375.0 32582.5 53440.0 32717.5 ;
      RECT  53565.0 32582.5 53630.0 32717.5 ;
      RECT  53565.0 32582.5 53630.0 32717.5 ;
      RECT  53375.0 32582.5 53440.0 32717.5 ;
      RECT  53375.0 33442.5 53440.0 33577.5 ;
      RECT  53565.0 33442.5 53630.0 33577.5 ;
      RECT  53565.0 33442.5 53630.0 33577.5 ;
      RECT  53375.0 33442.5 53440.0 33577.5 ;
      RECT  53302.5 33857.5 53367.5 33992.5 ;
      RECT  53637.5 32307.5 53702.5 32442.5 ;
      RECT  53375.0 33442.5 53440.0 33577.5 ;
      RECT  53565.0 32582.5 53630.0 32717.5 ;
      RECT  53822.5 32482.5 53887.5 32617.5 ;
      RECT  53822.5 32482.5 53887.5 32617.5 ;
      RECT  54270.0 33892.5 54335.0 33957.5 ;
      RECT  54005.0 33892.5 54302.5 33957.5 ;
      RECT  54270.0 33510.0 54335.0 33925.0 ;
      RECT  54080.0 32342.5 54145.0 32407.5 ;
      RECT  54112.5 32342.5 54375.0 32407.5 ;
      RECT  54080.0 32375.0 54145.0 32650.0 ;
      RECT  54080.0 32582.5 54145.0 32717.5 ;
      RECT  54270.0 32582.5 54335.0 32717.5 ;
      RECT  54270.0 32582.5 54335.0 32717.5 ;
      RECT  54080.0 32582.5 54145.0 32717.5 ;
      RECT  54080.0 33442.5 54145.0 33577.5 ;
      RECT  54270.0 33442.5 54335.0 33577.5 ;
      RECT  54270.0 33442.5 54335.0 33577.5 ;
      RECT  54080.0 33442.5 54145.0 33577.5 ;
      RECT  54007.5 33857.5 54072.5 33992.5 ;
      RECT  54342.5 32307.5 54407.5 32442.5 ;
      RECT  54080.0 33442.5 54145.0 33577.5 ;
      RECT  54270.0 32582.5 54335.0 32717.5 ;
      RECT  54527.5 32482.5 54592.5 32617.5 ;
      RECT  54527.5 32482.5 54592.5 32617.5 ;
      RECT  54975.0 33892.5 55040.0 33957.5 ;
      RECT  54710.0 33892.5 55007.5 33957.5 ;
      RECT  54975.0 33510.0 55040.0 33925.0 ;
      RECT  54785.0 32342.5 54850.0 32407.5 ;
      RECT  54817.5 32342.5 55080.0 32407.5 ;
      RECT  54785.0 32375.0 54850.0 32650.0 ;
      RECT  54785.0 32582.5 54850.0 32717.5 ;
      RECT  54975.0 32582.5 55040.0 32717.5 ;
      RECT  54975.0 32582.5 55040.0 32717.5 ;
      RECT  54785.0 32582.5 54850.0 32717.5 ;
      RECT  54785.0 33442.5 54850.0 33577.5 ;
      RECT  54975.0 33442.5 55040.0 33577.5 ;
      RECT  54975.0 33442.5 55040.0 33577.5 ;
      RECT  54785.0 33442.5 54850.0 33577.5 ;
      RECT  54712.5 33857.5 54777.5 33992.5 ;
      RECT  55047.5 32307.5 55112.5 32442.5 ;
      RECT  54785.0 33442.5 54850.0 33577.5 ;
      RECT  54975.0 32582.5 55040.0 32717.5 ;
      RECT  55232.5 32482.5 55297.5 32617.5 ;
      RECT  55232.5 32482.5 55297.5 32617.5 ;
      RECT  55680.0 33892.5 55745.0 33957.5 ;
      RECT  55415.0 33892.5 55712.5 33957.5 ;
      RECT  55680.0 33510.0 55745.0 33925.0 ;
      RECT  55490.0 32342.5 55555.0 32407.5 ;
      RECT  55522.5 32342.5 55785.0 32407.5 ;
      RECT  55490.0 32375.0 55555.0 32650.0 ;
      RECT  55490.0 32582.5 55555.0 32717.5 ;
      RECT  55680.0 32582.5 55745.0 32717.5 ;
      RECT  55680.0 32582.5 55745.0 32717.5 ;
      RECT  55490.0 32582.5 55555.0 32717.5 ;
      RECT  55490.0 33442.5 55555.0 33577.5 ;
      RECT  55680.0 33442.5 55745.0 33577.5 ;
      RECT  55680.0 33442.5 55745.0 33577.5 ;
      RECT  55490.0 33442.5 55555.0 33577.5 ;
      RECT  55417.5 33857.5 55482.5 33992.5 ;
      RECT  55752.5 32307.5 55817.5 32442.5 ;
      RECT  55490.0 33442.5 55555.0 33577.5 ;
      RECT  55680.0 32582.5 55745.0 32717.5 ;
      RECT  55937.5 32482.5 56002.5 32617.5 ;
      RECT  55937.5 32482.5 56002.5 32617.5 ;
      RECT  56385.0 33892.5 56450.0 33957.5 ;
      RECT  56120.0 33892.5 56417.5 33957.5 ;
      RECT  56385.0 33510.0 56450.0 33925.0 ;
      RECT  56195.0 32342.5 56260.0 32407.5 ;
      RECT  56227.5 32342.5 56490.0 32407.5 ;
      RECT  56195.0 32375.0 56260.0 32650.0 ;
      RECT  56195.0 32582.5 56260.0 32717.5 ;
      RECT  56385.0 32582.5 56450.0 32717.5 ;
      RECT  56385.0 32582.5 56450.0 32717.5 ;
      RECT  56195.0 32582.5 56260.0 32717.5 ;
      RECT  56195.0 33442.5 56260.0 33577.5 ;
      RECT  56385.0 33442.5 56450.0 33577.5 ;
      RECT  56385.0 33442.5 56450.0 33577.5 ;
      RECT  56195.0 33442.5 56260.0 33577.5 ;
      RECT  56122.5 33857.5 56187.5 33992.5 ;
      RECT  56457.5 32307.5 56522.5 32442.5 ;
      RECT  56195.0 33442.5 56260.0 33577.5 ;
      RECT  56385.0 32582.5 56450.0 32717.5 ;
      RECT  56642.5 32482.5 56707.5 32617.5 ;
      RECT  56642.5 32482.5 56707.5 32617.5 ;
      RECT  57090.0 33892.5 57155.0 33957.5 ;
      RECT  56825.0 33892.5 57122.5 33957.5 ;
      RECT  57090.0 33510.0 57155.0 33925.0 ;
      RECT  56900.0 32342.5 56965.0 32407.5 ;
      RECT  56932.5 32342.5 57195.0 32407.5 ;
      RECT  56900.0 32375.0 56965.0 32650.0 ;
      RECT  56900.0 32582.5 56965.0 32717.5 ;
      RECT  57090.0 32582.5 57155.0 32717.5 ;
      RECT  57090.0 32582.5 57155.0 32717.5 ;
      RECT  56900.0 32582.5 56965.0 32717.5 ;
      RECT  56900.0 33442.5 56965.0 33577.5 ;
      RECT  57090.0 33442.5 57155.0 33577.5 ;
      RECT  57090.0 33442.5 57155.0 33577.5 ;
      RECT  56900.0 33442.5 56965.0 33577.5 ;
      RECT  56827.5 33857.5 56892.5 33992.5 ;
      RECT  57162.5 32307.5 57227.5 32442.5 ;
      RECT  56900.0 33442.5 56965.0 33577.5 ;
      RECT  57090.0 32582.5 57155.0 32717.5 ;
      RECT  57347.5 32482.5 57412.5 32617.5 ;
      RECT  57347.5 32482.5 57412.5 32617.5 ;
      RECT  57795.0 33892.5 57860.0 33957.5 ;
      RECT  57530.0 33892.5 57827.5 33957.5 ;
      RECT  57795.0 33510.0 57860.0 33925.0 ;
      RECT  57605.0 32342.5 57670.0 32407.5 ;
      RECT  57637.5 32342.5 57900.0 32407.5 ;
      RECT  57605.0 32375.0 57670.0 32650.0 ;
      RECT  57605.0 32582.5 57670.0 32717.5 ;
      RECT  57795.0 32582.5 57860.0 32717.5 ;
      RECT  57795.0 32582.5 57860.0 32717.5 ;
      RECT  57605.0 32582.5 57670.0 32717.5 ;
      RECT  57605.0 33442.5 57670.0 33577.5 ;
      RECT  57795.0 33442.5 57860.0 33577.5 ;
      RECT  57795.0 33442.5 57860.0 33577.5 ;
      RECT  57605.0 33442.5 57670.0 33577.5 ;
      RECT  57532.5 33857.5 57597.5 33992.5 ;
      RECT  57867.5 32307.5 57932.5 32442.5 ;
      RECT  57605.0 33442.5 57670.0 33577.5 ;
      RECT  57795.0 32582.5 57860.0 32717.5 ;
      RECT  58052.5 32482.5 58117.5 32617.5 ;
      RECT  58052.5 32482.5 58117.5 32617.5 ;
      RECT  58500.0 33892.5 58565.0 33957.5 ;
      RECT  58235.0 33892.5 58532.5 33957.5 ;
      RECT  58500.0 33510.0 58565.0 33925.0 ;
      RECT  58310.0 32342.5 58375.0 32407.5 ;
      RECT  58342.5 32342.5 58605.0 32407.5 ;
      RECT  58310.0 32375.0 58375.0 32650.0 ;
      RECT  58310.0 32582.5 58375.0 32717.5 ;
      RECT  58500.0 32582.5 58565.0 32717.5 ;
      RECT  58500.0 32582.5 58565.0 32717.5 ;
      RECT  58310.0 32582.5 58375.0 32717.5 ;
      RECT  58310.0 33442.5 58375.0 33577.5 ;
      RECT  58500.0 33442.5 58565.0 33577.5 ;
      RECT  58500.0 33442.5 58565.0 33577.5 ;
      RECT  58310.0 33442.5 58375.0 33577.5 ;
      RECT  58237.5 33857.5 58302.5 33992.5 ;
      RECT  58572.5 32307.5 58637.5 32442.5 ;
      RECT  58310.0 33442.5 58375.0 33577.5 ;
      RECT  58500.0 32582.5 58565.0 32717.5 ;
      RECT  58757.5 32482.5 58822.5 32617.5 ;
      RECT  58757.5 32482.5 58822.5 32617.5 ;
      RECT  59205.0 33892.5 59270.0 33957.5 ;
      RECT  58940.0 33892.5 59237.5 33957.5 ;
      RECT  59205.0 33510.0 59270.0 33925.0 ;
      RECT  59015.0 32342.5 59080.0 32407.5 ;
      RECT  59047.5 32342.5 59310.0 32407.5 ;
      RECT  59015.0 32375.0 59080.0 32650.0 ;
      RECT  59015.0 32582.5 59080.0 32717.5 ;
      RECT  59205.0 32582.5 59270.0 32717.5 ;
      RECT  59205.0 32582.5 59270.0 32717.5 ;
      RECT  59015.0 32582.5 59080.0 32717.5 ;
      RECT  59015.0 33442.5 59080.0 33577.5 ;
      RECT  59205.0 33442.5 59270.0 33577.5 ;
      RECT  59205.0 33442.5 59270.0 33577.5 ;
      RECT  59015.0 33442.5 59080.0 33577.5 ;
      RECT  58942.5 33857.5 59007.5 33992.5 ;
      RECT  59277.5 32307.5 59342.5 32442.5 ;
      RECT  59015.0 33442.5 59080.0 33577.5 ;
      RECT  59205.0 32582.5 59270.0 32717.5 ;
      RECT  59462.5 32482.5 59527.5 32617.5 ;
      RECT  59462.5 32482.5 59527.5 32617.5 ;
      RECT  59910.0 33892.5 59975.0 33957.5 ;
      RECT  59645.0 33892.5 59942.5 33957.5 ;
      RECT  59910.0 33510.0 59975.0 33925.0 ;
      RECT  59720.0 32342.5 59785.0 32407.5 ;
      RECT  59752.5 32342.5 60015.0 32407.5 ;
      RECT  59720.0 32375.0 59785.0 32650.0 ;
      RECT  59720.0 32582.5 59785.0 32717.5 ;
      RECT  59910.0 32582.5 59975.0 32717.5 ;
      RECT  59910.0 32582.5 59975.0 32717.5 ;
      RECT  59720.0 32582.5 59785.0 32717.5 ;
      RECT  59720.0 33442.5 59785.0 33577.5 ;
      RECT  59910.0 33442.5 59975.0 33577.5 ;
      RECT  59910.0 33442.5 59975.0 33577.5 ;
      RECT  59720.0 33442.5 59785.0 33577.5 ;
      RECT  59647.5 33857.5 59712.5 33992.5 ;
      RECT  59982.5 32307.5 60047.5 32442.5 ;
      RECT  59720.0 33442.5 59785.0 33577.5 ;
      RECT  59910.0 32582.5 59975.0 32717.5 ;
      RECT  60167.5 32482.5 60232.5 32617.5 ;
      RECT  60167.5 32482.5 60232.5 32617.5 ;
      RECT  60615.0 33892.5 60680.0 33957.5 ;
      RECT  60350.0 33892.5 60647.5 33957.5 ;
      RECT  60615.0 33510.0 60680.0 33925.0 ;
      RECT  60425.0 32342.5 60490.0 32407.5 ;
      RECT  60457.5 32342.5 60720.0 32407.5 ;
      RECT  60425.0 32375.0 60490.0 32650.0 ;
      RECT  60425.0 32582.5 60490.0 32717.5 ;
      RECT  60615.0 32582.5 60680.0 32717.5 ;
      RECT  60615.0 32582.5 60680.0 32717.5 ;
      RECT  60425.0 32582.5 60490.0 32717.5 ;
      RECT  60425.0 33442.5 60490.0 33577.5 ;
      RECT  60615.0 33442.5 60680.0 33577.5 ;
      RECT  60615.0 33442.5 60680.0 33577.5 ;
      RECT  60425.0 33442.5 60490.0 33577.5 ;
      RECT  60352.5 33857.5 60417.5 33992.5 ;
      RECT  60687.5 32307.5 60752.5 32442.5 ;
      RECT  60425.0 33442.5 60490.0 33577.5 ;
      RECT  60615.0 32582.5 60680.0 32717.5 ;
      RECT  60872.5 32482.5 60937.5 32617.5 ;
      RECT  60872.5 32482.5 60937.5 32617.5 ;
      RECT  61320.0 33892.5 61385.0 33957.5 ;
      RECT  61055.0 33892.5 61352.5 33957.5 ;
      RECT  61320.0 33510.0 61385.0 33925.0 ;
      RECT  61130.0 32342.5 61195.0 32407.5 ;
      RECT  61162.5 32342.5 61425.0 32407.5 ;
      RECT  61130.0 32375.0 61195.0 32650.0 ;
      RECT  61130.0 32582.5 61195.0 32717.5 ;
      RECT  61320.0 32582.5 61385.0 32717.5 ;
      RECT  61320.0 32582.5 61385.0 32717.5 ;
      RECT  61130.0 32582.5 61195.0 32717.5 ;
      RECT  61130.0 33442.5 61195.0 33577.5 ;
      RECT  61320.0 33442.5 61385.0 33577.5 ;
      RECT  61320.0 33442.5 61385.0 33577.5 ;
      RECT  61130.0 33442.5 61195.0 33577.5 ;
      RECT  61057.5 33857.5 61122.5 33992.5 ;
      RECT  61392.5 32307.5 61457.5 32442.5 ;
      RECT  61130.0 33442.5 61195.0 33577.5 ;
      RECT  61320.0 32582.5 61385.0 32717.5 ;
      RECT  61577.5 32482.5 61642.5 32617.5 ;
      RECT  61577.5 32482.5 61642.5 32617.5 ;
      RECT  62025.0 33892.5 62090.0 33957.5 ;
      RECT  61760.0 33892.5 62057.5 33957.5 ;
      RECT  62025.0 33510.0 62090.0 33925.0 ;
      RECT  61835.0 32342.5 61900.0 32407.5 ;
      RECT  61867.5 32342.5 62130.0 32407.5 ;
      RECT  61835.0 32375.0 61900.0 32650.0 ;
      RECT  61835.0 32582.5 61900.0 32717.5 ;
      RECT  62025.0 32582.5 62090.0 32717.5 ;
      RECT  62025.0 32582.5 62090.0 32717.5 ;
      RECT  61835.0 32582.5 61900.0 32717.5 ;
      RECT  61835.0 33442.5 61900.0 33577.5 ;
      RECT  62025.0 33442.5 62090.0 33577.5 ;
      RECT  62025.0 33442.5 62090.0 33577.5 ;
      RECT  61835.0 33442.5 61900.0 33577.5 ;
      RECT  61762.5 33857.5 61827.5 33992.5 ;
      RECT  62097.5 32307.5 62162.5 32442.5 ;
      RECT  61835.0 33442.5 61900.0 33577.5 ;
      RECT  62025.0 32582.5 62090.0 32717.5 ;
      RECT  62282.5 32482.5 62347.5 32617.5 ;
      RECT  62282.5 32482.5 62347.5 32617.5 ;
      RECT  62730.0 33892.5 62795.0 33957.5 ;
      RECT  62465.0 33892.5 62762.5 33957.5 ;
      RECT  62730.0 33510.0 62795.0 33925.0 ;
      RECT  62540.0 32342.5 62605.0 32407.5 ;
      RECT  62572.5 32342.5 62835.0 32407.5 ;
      RECT  62540.0 32375.0 62605.0 32650.0 ;
      RECT  62540.0 32582.5 62605.0 32717.5 ;
      RECT  62730.0 32582.5 62795.0 32717.5 ;
      RECT  62730.0 32582.5 62795.0 32717.5 ;
      RECT  62540.0 32582.5 62605.0 32717.5 ;
      RECT  62540.0 33442.5 62605.0 33577.5 ;
      RECT  62730.0 33442.5 62795.0 33577.5 ;
      RECT  62730.0 33442.5 62795.0 33577.5 ;
      RECT  62540.0 33442.5 62605.0 33577.5 ;
      RECT  62467.5 33857.5 62532.5 33992.5 ;
      RECT  62802.5 32307.5 62867.5 32442.5 ;
      RECT  62540.0 33442.5 62605.0 33577.5 ;
      RECT  62730.0 32582.5 62795.0 32717.5 ;
      RECT  62987.5 32482.5 63052.5 32617.5 ;
      RECT  62987.5 32482.5 63052.5 32617.5 ;
      RECT  63435.0 33892.5 63500.0 33957.5 ;
      RECT  63170.0 33892.5 63467.5 33957.5 ;
      RECT  63435.0 33510.0 63500.0 33925.0 ;
      RECT  63245.0 32342.5 63310.0 32407.5 ;
      RECT  63277.5 32342.5 63540.0 32407.5 ;
      RECT  63245.0 32375.0 63310.0 32650.0 ;
      RECT  63245.0 32582.5 63310.0 32717.5 ;
      RECT  63435.0 32582.5 63500.0 32717.5 ;
      RECT  63435.0 32582.5 63500.0 32717.5 ;
      RECT  63245.0 32582.5 63310.0 32717.5 ;
      RECT  63245.0 33442.5 63310.0 33577.5 ;
      RECT  63435.0 33442.5 63500.0 33577.5 ;
      RECT  63435.0 33442.5 63500.0 33577.5 ;
      RECT  63245.0 33442.5 63310.0 33577.5 ;
      RECT  63172.5 33857.5 63237.5 33992.5 ;
      RECT  63507.5 32307.5 63572.5 32442.5 ;
      RECT  63245.0 33442.5 63310.0 33577.5 ;
      RECT  63435.0 32582.5 63500.0 32717.5 ;
      RECT  63692.5 32482.5 63757.5 32617.5 ;
      RECT  63692.5 32482.5 63757.5 32617.5 ;
      RECT  64140.0 33892.5 64205.0 33957.5 ;
      RECT  63875.0 33892.5 64172.5 33957.5 ;
      RECT  64140.0 33510.0 64205.0 33925.0 ;
      RECT  63950.0 32342.5 64015.0 32407.5 ;
      RECT  63982.5 32342.5 64245.0 32407.5 ;
      RECT  63950.0 32375.0 64015.0 32650.0 ;
      RECT  63950.0 32582.5 64015.0 32717.5 ;
      RECT  64140.0 32582.5 64205.0 32717.5 ;
      RECT  64140.0 32582.5 64205.0 32717.5 ;
      RECT  63950.0 32582.5 64015.0 32717.5 ;
      RECT  63950.0 33442.5 64015.0 33577.5 ;
      RECT  64140.0 33442.5 64205.0 33577.5 ;
      RECT  64140.0 33442.5 64205.0 33577.5 ;
      RECT  63950.0 33442.5 64015.0 33577.5 ;
      RECT  63877.5 33857.5 63942.5 33992.5 ;
      RECT  64212.5 32307.5 64277.5 32442.5 ;
      RECT  63950.0 33442.5 64015.0 33577.5 ;
      RECT  64140.0 32582.5 64205.0 32717.5 ;
      RECT  64397.5 32482.5 64462.5 32617.5 ;
      RECT  64397.5 32482.5 64462.5 32617.5 ;
      RECT  64845.0 33892.5 64910.0 33957.5 ;
      RECT  64580.0 33892.5 64877.5 33957.5 ;
      RECT  64845.0 33510.0 64910.0 33925.0 ;
      RECT  64655.0 32342.5 64720.0 32407.5 ;
      RECT  64687.5 32342.5 64950.0 32407.5 ;
      RECT  64655.0 32375.0 64720.0 32650.0 ;
      RECT  64655.0 32582.5 64720.0 32717.5 ;
      RECT  64845.0 32582.5 64910.0 32717.5 ;
      RECT  64845.0 32582.5 64910.0 32717.5 ;
      RECT  64655.0 32582.5 64720.0 32717.5 ;
      RECT  64655.0 33442.5 64720.0 33577.5 ;
      RECT  64845.0 33442.5 64910.0 33577.5 ;
      RECT  64845.0 33442.5 64910.0 33577.5 ;
      RECT  64655.0 33442.5 64720.0 33577.5 ;
      RECT  64582.5 33857.5 64647.5 33992.5 ;
      RECT  64917.5 32307.5 64982.5 32442.5 ;
      RECT  64655.0 33442.5 64720.0 33577.5 ;
      RECT  64845.0 32582.5 64910.0 32717.5 ;
      RECT  65102.5 32482.5 65167.5 32617.5 ;
      RECT  65102.5 32482.5 65167.5 32617.5 ;
      RECT  65550.0 33892.5 65615.0 33957.5 ;
      RECT  65285.0 33892.5 65582.5 33957.5 ;
      RECT  65550.0 33510.0 65615.0 33925.0 ;
      RECT  65360.0 32342.5 65425.0 32407.5 ;
      RECT  65392.5 32342.5 65655.0 32407.5 ;
      RECT  65360.0 32375.0 65425.0 32650.0 ;
      RECT  65360.0 32582.5 65425.0 32717.5 ;
      RECT  65550.0 32582.5 65615.0 32717.5 ;
      RECT  65550.0 32582.5 65615.0 32717.5 ;
      RECT  65360.0 32582.5 65425.0 32717.5 ;
      RECT  65360.0 33442.5 65425.0 33577.5 ;
      RECT  65550.0 33442.5 65615.0 33577.5 ;
      RECT  65550.0 33442.5 65615.0 33577.5 ;
      RECT  65360.0 33442.5 65425.0 33577.5 ;
      RECT  65287.5 33857.5 65352.5 33992.5 ;
      RECT  65622.5 32307.5 65687.5 32442.5 ;
      RECT  65360.0 33442.5 65425.0 33577.5 ;
      RECT  65550.0 32582.5 65615.0 32717.5 ;
      RECT  65807.5 32482.5 65872.5 32617.5 ;
      RECT  65807.5 32482.5 65872.5 32617.5 ;
      RECT  66255.0 33892.5 66320.0 33957.5 ;
      RECT  65990.0 33892.5 66287.5 33957.5 ;
      RECT  66255.0 33510.0 66320.0 33925.0 ;
      RECT  66065.0 32342.5 66130.0 32407.5 ;
      RECT  66097.5 32342.5 66360.0 32407.5 ;
      RECT  66065.0 32375.0 66130.0 32650.0 ;
      RECT  66065.0 32582.5 66130.0 32717.5 ;
      RECT  66255.0 32582.5 66320.0 32717.5 ;
      RECT  66255.0 32582.5 66320.0 32717.5 ;
      RECT  66065.0 32582.5 66130.0 32717.5 ;
      RECT  66065.0 33442.5 66130.0 33577.5 ;
      RECT  66255.0 33442.5 66320.0 33577.5 ;
      RECT  66255.0 33442.5 66320.0 33577.5 ;
      RECT  66065.0 33442.5 66130.0 33577.5 ;
      RECT  65992.5 33857.5 66057.5 33992.5 ;
      RECT  66327.5 32307.5 66392.5 32442.5 ;
      RECT  66065.0 33442.5 66130.0 33577.5 ;
      RECT  66255.0 32582.5 66320.0 32717.5 ;
      RECT  66512.5 32482.5 66577.5 32617.5 ;
      RECT  66512.5 32482.5 66577.5 32617.5 ;
      RECT  66960.0 33892.5 67025.0 33957.5 ;
      RECT  66695.0 33892.5 66992.5 33957.5 ;
      RECT  66960.0 33510.0 67025.0 33925.0 ;
      RECT  66770.0 32342.5 66835.0 32407.5 ;
      RECT  66802.5 32342.5 67065.0 32407.5 ;
      RECT  66770.0 32375.0 66835.0 32650.0 ;
      RECT  66770.0 32582.5 66835.0 32717.5 ;
      RECT  66960.0 32582.5 67025.0 32717.5 ;
      RECT  66960.0 32582.5 67025.0 32717.5 ;
      RECT  66770.0 32582.5 66835.0 32717.5 ;
      RECT  66770.0 33442.5 66835.0 33577.5 ;
      RECT  66960.0 33442.5 67025.0 33577.5 ;
      RECT  66960.0 33442.5 67025.0 33577.5 ;
      RECT  66770.0 33442.5 66835.0 33577.5 ;
      RECT  66697.5 33857.5 66762.5 33992.5 ;
      RECT  67032.5 32307.5 67097.5 32442.5 ;
      RECT  66770.0 33442.5 66835.0 33577.5 ;
      RECT  66960.0 32582.5 67025.0 32717.5 ;
      RECT  67217.5 32482.5 67282.5 32617.5 ;
      RECT  67217.5 32482.5 67282.5 32617.5 ;
      RECT  67665.0 33892.5 67730.0 33957.5 ;
      RECT  67400.0 33892.5 67697.5 33957.5 ;
      RECT  67665.0 33510.0 67730.0 33925.0 ;
      RECT  67475.0 32342.5 67540.0 32407.5 ;
      RECT  67507.5 32342.5 67770.0 32407.5 ;
      RECT  67475.0 32375.0 67540.0 32650.0 ;
      RECT  67475.0 32582.5 67540.0 32717.5 ;
      RECT  67665.0 32582.5 67730.0 32717.5 ;
      RECT  67665.0 32582.5 67730.0 32717.5 ;
      RECT  67475.0 32582.5 67540.0 32717.5 ;
      RECT  67475.0 33442.5 67540.0 33577.5 ;
      RECT  67665.0 33442.5 67730.0 33577.5 ;
      RECT  67665.0 33442.5 67730.0 33577.5 ;
      RECT  67475.0 33442.5 67540.0 33577.5 ;
      RECT  67402.5 33857.5 67467.5 33992.5 ;
      RECT  67737.5 32307.5 67802.5 32442.5 ;
      RECT  67475.0 33442.5 67540.0 33577.5 ;
      RECT  67665.0 32582.5 67730.0 32717.5 ;
      RECT  67922.5 32482.5 67987.5 32617.5 ;
      RECT  67922.5 32482.5 67987.5 32617.5 ;
      RECT  68370.0 33892.5 68435.0 33957.5 ;
      RECT  68105.0 33892.5 68402.5 33957.5 ;
      RECT  68370.0 33510.0 68435.0 33925.0 ;
      RECT  68180.0 32342.5 68245.0 32407.5 ;
      RECT  68212.5 32342.5 68475.0 32407.5 ;
      RECT  68180.0 32375.0 68245.0 32650.0 ;
      RECT  68180.0 32582.5 68245.0 32717.5 ;
      RECT  68370.0 32582.5 68435.0 32717.5 ;
      RECT  68370.0 32582.5 68435.0 32717.5 ;
      RECT  68180.0 32582.5 68245.0 32717.5 ;
      RECT  68180.0 33442.5 68245.0 33577.5 ;
      RECT  68370.0 33442.5 68435.0 33577.5 ;
      RECT  68370.0 33442.5 68435.0 33577.5 ;
      RECT  68180.0 33442.5 68245.0 33577.5 ;
      RECT  68107.5 33857.5 68172.5 33992.5 ;
      RECT  68442.5 32307.5 68507.5 32442.5 ;
      RECT  68180.0 33442.5 68245.0 33577.5 ;
      RECT  68370.0 32582.5 68435.0 32717.5 ;
      RECT  68627.5 32482.5 68692.5 32617.5 ;
      RECT  68627.5 32482.5 68692.5 32617.5 ;
      RECT  69075.0 33892.5 69140.0 33957.5 ;
      RECT  68810.0 33892.5 69107.5 33957.5 ;
      RECT  69075.0 33510.0 69140.0 33925.0 ;
      RECT  68885.0 32342.5 68950.0 32407.5 ;
      RECT  68917.5 32342.5 69180.0 32407.5 ;
      RECT  68885.0 32375.0 68950.0 32650.0 ;
      RECT  68885.0 32582.5 68950.0 32717.5 ;
      RECT  69075.0 32582.5 69140.0 32717.5 ;
      RECT  69075.0 32582.5 69140.0 32717.5 ;
      RECT  68885.0 32582.5 68950.0 32717.5 ;
      RECT  68885.0 33442.5 68950.0 33577.5 ;
      RECT  69075.0 33442.5 69140.0 33577.5 ;
      RECT  69075.0 33442.5 69140.0 33577.5 ;
      RECT  68885.0 33442.5 68950.0 33577.5 ;
      RECT  68812.5 33857.5 68877.5 33992.5 ;
      RECT  69147.5 32307.5 69212.5 32442.5 ;
      RECT  68885.0 33442.5 68950.0 33577.5 ;
      RECT  69075.0 32582.5 69140.0 32717.5 ;
      RECT  69332.5 32482.5 69397.5 32617.5 ;
      RECT  69332.5 32482.5 69397.5 32617.5 ;
      RECT  69780.0 33892.5 69845.0 33957.5 ;
      RECT  69515.0 33892.5 69812.5 33957.5 ;
      RECT  69780.0 33510.0 69845.0 33925.0 ;
      RECT  69590.0 32342.5 69655.0 32407.5 ;
      RECT  69622.5 32342.5 69885.0 32407.5 ;
      RECT  69590.0 32375.0 69655.0 32650.0 ;
      RECT  69590.0 32582.5 69655.0 32717.5 ;
      RECT  69780.0 32582.5 69845.0 32717.5 ;
      RECT  69780.0 32582.5 69845.0 32717.5 ;
      RECT  69590.0 32582.5 69655.0 32717.5 ;
      RECT  69590.0 33442.5 69655.0 33577.5 ;
      RECT  69780.0 33442.5 69845.0 33577.5 ;
      RECT  69780.0 33442.5 69845.0 33577.5 ;
      RECT  69590.0 33442.5 69655.0 33577.5 ;
      RECT  69517.5 33857.5 69582.5 33992.5 ;
      RECT  69852.5 32307.5 69917.5 32442.5 ;
      RECT  69590.0 33442.5 69655.0 33577.5 ;
      RECT  69780.0 32582.5 69845.0 32717.5 ;
      RECT  70037.5 32482.5 70102.5 32617.5 ;
      RECT  70037.5 32482.5 70102.5 32617.5 ;
      RECT  70485.0 33892.5 70550.0 33957.5 ;
      RECT  70220.0 33892.5 70517.5 33957.5 ;
      RECT  70485.0 33510.0 70550.0 33925.0 ;
      RECT  70295.0 32342.5 70360.0 32407.5 ;
      RECT  70327.5 32342.5 70590.0 32407.5 ;
      RECT  70295.0 32375.0 70360.0 32650.0 ;
      RECT  70295.0 32582.5 70360.0 32717.5 ;
      RECT  70485.0 32582.5 70550.0 32717.5 ;
      RECT  70485.0 32582.5 70550.0 32717.5 ;
      RECT  70295.0 32582.5 70360.0 32717.5 ;
      RECT  70295.0 33442.5 70360.0 33577.5 ;
      RECT  70485.0 33442.5 70550.0 33577.5 ;
      RECT  70485.0 33442.5 70550.0 33577.5 ;
      RECT  70295.0 33442.5 70360.0 33577.5 ;
      RECT  70222.5 33857.5 70287.5 33992.5 ;
      RECT  70557.5 32307.5 70622.5 32442.5 ;
      RECT  70295.0 33442.5 70360.0 33577.5 ;
      RECT  70485.0 32582.5 70550.0 32717.5 ;
      RECT  70742.5 32482.5 70807.5 32617.5 ;
      RECT  70742.5 32482.5 70807.5 32617.5 ;
      RECT  71190.0 33892.5 71255.0 33957.5 ;
      RECT  70925.0 33892.5 71222.5 33957.5 ;
      RECT  71190.0 33510.0 71255.0 33925.0 ;
      RECT  71000.0 32342.5 71065.0 32407.5 ;
      RECT  71032.5 32342.5 71295.0 32407.5 ;
      RECT  71000.0 32375.0 71065.0 32650.0 ;
      RECT  71000.0 32582.5 71065.0 32717.5 ;
      RECT  71190.0 32582.5 71255.0 32717.5 ;
      RECT  71190.0 32582.5 71255.0 32717.5 ;
      RECT  71000.0 32582.5 71065.0 32717.5 ;
      RECT  71000.0 33442.5 71065.0 33577.5 ;
      RECT  71190.0 33442.5 71255.0 33577.5 ;
      RECT  71190.0 33442.5 71255.0 33577.5 ;
      RECT  71000.0 33442.5 71065.0 33577.5 ;
      RECT  70927.5 33857.5 70992.5 33992.5 ;
      RECT  71262.5 32307.5 71327.5 32442.5 ;
      RECT  71000.0 33442.5 71065.0 33577.5 ;
      RECT  71190.0 32582.5 71255.0 32717.5 ;
      RECT  71447.5 32482.5 71512.5 32617.5 ;
      RECT  71447.5 32482.5 71512.5 32617.5 ;
      RECT  71895.0 33892.5 71960.0 33957.5 ;
      RECT  71630.0 33892.5 71927.5 33957.5 ;
      RECT  71895.0 33510.0 71960.0 33925.0 ;
      RECT  71705.0 32342.5 71770.0 32407.5 ;
      RECT  71737.5 32342.5 72000.0 32407.5 ;
      RECT  71705.0 32375.0 71770.0 32650.0 ;
      RECT  71705.0 32582.5 71770.0 32717.5 ;
      RECT  71895.0 32582.5 71960.0 32717.5 ;
      RECT  71895.0 32582.5 71960.0 32717.5 ;
      RECT  71705.0 32582.5 71770.0 32717.5 ;
      RECT  71705.0 33442.5 71770.0 33577.5 ;
      RECT  71895.0 33442.5 71960.0 33577.5 ;
      RECT  71895.0 33442.5 71960.0 33577.5 ;
      RECT  71705.0 33442.5 71770.0 33577.5 ;
      RECT  71632.5 33857.5 71697.5 33992.5 ;
      RECT  71967.5 32307.5 72032.5 32442.5 ;
      RECT  71705.0 33442.5 71770.0 33577.5 ;
      RECT  71895.0 32582.5 71960.0 32717.5 ;
      RECT  72152.5 32482.5 72217.5 32617.5 ;
      RECT  72152.5 32482.5 72217.5 32617.5 ;
      RECT  72600.0 33892.5 72665.0 33957.5 ;
      RECT  72335.0 33892.5 72632.5 33957.5 ;
      RECT  72600.0 33510.0 72665.0 33925.0 ;
      RECT  72410.0 32342.5 72475.0 32407.5 ;
      RECT  72442.5 32342.5 72705.0 32407.5 ;
      RECT  72410.0 32375.0 72475.0 32650.0 ;
      RECT  72410.0 32582.5 72475.0 32717.5 ;
      RECT  72600.0 32582.5 72665.0 32717.5 ;
      RECT  72600.0 32582.5 72665.0 32717.5 ;
      RECT  72410.0 32582.5 72475.0 32717.5 ;
      RECT  72410.0 33442.5 72475.0 33577.5 ;
      RECT  72600.0 33442.5 72665.0 33577.5 ;
      RECT  72600.0 33442.5 72665.0 33577.5 ;
      RECT  72410.0 33442.5 72475.0 33577.5 ;
      RECT  72337.5 33857.5 72402.5 33992.5 ;
      RECT  72672.5 32307.5 72737.5 32442.5 ;
      RECT  72410.0 33442.5 72475.0 33577.5 ;
      RECT  72600.0 32582.5 72665.0 32717.5 ;
      RECT  72857.5 32482.5 72922.5 32617.5 ;
      RECT  72857.5 32482.5 72922.5 32617.5 ;
      RECT  73305.0 33892.5 73370.0 33957.5 ;
      RECT  73040.0 33892.5 73337.5 33957.5 ;
      RECT  73305.0 33510.0 73370.0 33925.0 ;
      RECT  73115.0 32342.5 73180.0 32407.5 ;
      RECT  73147.5 32342.5 73410.0 32407.5 ;
      RECT  73115.0 32375.0 73180.0 32650.0 ;
      RECT  73115.0 32582.5 73180.0 32717.5 ;
      RECT  73305.0 32582.5 73370.0 32717.5 ;
      RECT  73305.0 32582.5 73370.0 32717.5 ;
      RECT  73115.0 32582.5 73180.0 32717.5 ;
      RECT  73115.0 33442.5 73180.0 33577.5 ;
      RECT  73305.0 33442.5 73370.0 33577.5 ;
      RECT  73305.0 33442.5 73370.0 33577.5 ;
      RECT  73115.0 33442.5 73180.0 33577.5 ;
      RECT  73042.5 33857.5 73107.5 33992.5 ;
      RECT  73377.5 32307.5 73442.5 32442.5 ;
      RECT  73115.0 33442.5 73180.0 33577.5 ;
      RECT  73305.0 32582.5 73370.0 32717.5 ;
      RECT  73562.5 32482.5 73627.5 32617.5 ;
      RECT  73562.5 32482.5 73627.5 32617.5 ;
      RECT  74010.0 33892.5 74075.0 33957.5 ;
      RECT  73745.0 33892.5 74042.5 33957.5 ;
      RECT  74010.0 33510.0 74075.0 33925.0 ;
      RECT  73820.0 32342.5 73885.0 32407.5 ;
      RECT  73852.5 32342.5 74115.0 32407.5 ;
      RECT  73820.0 32375.0 73885.0 32650.0 ;
      RECT  73820.0 32582.5 73885.0 32717.5 ;
      RECT  74010.0 32582.5 74075.0 32717.5 ;
      RECT  74010.0 32582.5 74075.0 32717.5 ;
      RECT  73820.0 32582.5 73885.0 32717.5 ;
      RECT  73820.0 33442.5 73885.0 33577.5 ;
      RECT  74010.0 33442.5 74075.0 33577.5 ;
      RECT  74010.0 33442.5 74075.0 33577.5 ;
      RECT  73820.0 33442.5 73885.0 33577.5 ;
      RECT  73747.5 33857.5 73812.5 33992.5 ;
      RECT  74082.5 32307.5 74147.5 32442.5 ;
      RECT  73820.0 33442.5 73885.0 33577.5 ;
      RECT  74010.0 32582.5 74075.0 32717.5 ;
      RECT  74267.5 32482.5 74332.5 32617.5 ;
      RECT  74267.5 32482.5 74332.5 32617.5 ;
      RECT  74715.0 33892.5 74780.0 33957.5 ;
      RECT  74450.0 33892.5 74747.5 33957.5 ;
      RECT  74715.0 33510.0 74780.0 33925.0 ;
      RECT  74525.0 32342.5 74590.0 32407.5 ;
      RECT  74557.5 32342.5 74820.0 32407.5 ;
      RECT  74525.0 32375.0 74590.0 32650.0 ;
      RECT  74525.0 32582.5 74590.0 32717.5 ;
      RECT  74715.0 32582.5 74780.0 32717.5 ;
      RECT  74715.0 32582.5 74780.0 32717.5 ;
      RECT  74525.0 32582.5 74590.0 32717.5 ;
      RECT  74525.0 33442.5 74590.0 33577.5 ;
      RECT  74715.0 33442.5 74780.0 33577.5 ;
      RECT  74715.0 33442.5 74780.0 33577.5 ;
      RECT  74525.0 33442.5 74590.0 33577.5 ;
      RECT  74452.5 33857.5 74517.5 33992.5 ;
      RECT  74787.5 32307.5 74852.5 32442.5 ;
      RECT  74525.0 33442.5 74590.0 33577.5 ;
      RECT  74715.0 32582.5 74780.0 32717.5 ;
      RECT  74972.5 32482.5 75037.5 32617.5 ;
      RECT  74972.5 32482.5 75037.5 32617.5 ;
      RECT  75420.0 33892.5 75485.0 33957.5 ;
      RECT  75155.0 33892.5 75452.5 33957.5 ;
      RECT  75420.0 33510.0 75485.0 33925.0 ;
      RECT  75230.0 32342.5 75295.0 32407.5 ;
      RECT  75262.5 32342.5 75525.0 32407.5 ;
      RECT  75230.0 32375.0 75295.0 32650.0 ;
      RECT  75230.0 32582.5 75295.0 32717.5 ;
      RECT  75420.0 32582.5 75485.0 32717.5 ;
      RECT  75420.0 32582.5 75485.0 32717.5 ;
      RECT  75230.0 32582.5 75295.0 32717.5 ;
      RECT  75230.0 33442.5 75295.0 33577.5 ;
      RECT  75420.0 33442.5 75485.0 33577.5 ;
      RECT  75420.0 33442.5 75485.0 33577.5 ;
      RECT  75230.0 33442.5 75295.0 33577.5 ;
      RECT  75157.5 33857.5 75222.5 33992.5 ;
      RECT  75492.5 32307.5 75557.5 32442.5 ;
      RECT  75230.0 33442.5 75295.0 33577.5 ;
      RECT  75420.0 32582.5 75485.0 32717.5 ;
      RECT  75677.5 32482.5 75742.5 32617.5 ;
      RECT  75677.5 32482.5 75742.5 32617.5 ;
      RECT  76125.0 33892.5 76190.0 33957.5 ;
      RECT  75860.0 33892.5 76157.5 33957.5 ;
      RECT  76125.0 33510.0 76190.0 33925.0 ;
      RECT  75935.0 32342.5 76000.0 32407.5 ;
      RECT  75967.5 32342.5 76230.0 32407.5 ;
      RECT  75935.0 32375.0 76000.0 32650.0 ;
      RECT  75935.0 32582.5 76000.0 32717.5 ;
      RECT  76125.0 32582.5 76190.0 32717.5 ;
      RECT  76125.0 32582.5 76190.0 32717.5 ;
      RECT  75935.0 32582.5 76000.0 32717.5 ;
      RECT  75935.0 33442.5 76000.0 33577.5 ;
      RECT  76125.0 33442.5 76190.0 33577.5 ;
      RECT  76125.0 33442.5 76190.0 33577.5 ;
      RECT  75935.0 33442.5 76000.0 33577.5 ;
      RECT  75862.5 33857.5 75927.5 33992.5 ;
      RECT  76197.5 32307.5 76262.5 32442.5 ;
      RECT  75935.0 33442.5 76000.0 33577.5 ;
      RECT  76125.0 32582.5 76190.0 32717.5 ;
      RECT  76382.5 32482.5 76447.5 32617.5 ;
      RECT  76382.5 32482.5 76447.5 32617.5 ;
      RECT  76830.0 33892.5 76895.0 33957.5 ;
      RECT  76565.0 33892.5 76862.5 33957.5 ;
      RECT  76830.0 33510.0 76895.0 33925.0 ;
      RECT  76640.0 32342.5 76705.0 32407.5 ;
      RECT  76672.5 32342.5 76935.0 32407.5 ;
      RECT  76640.0 32375.0 76705.0 32650.0 ;
      RECT  76640.0 32582.5 76705.0 32717.5 ;
      RECT  76830.0 32582.5 76895.0 32717.5 ;
      RECT  76830.0 32582.5 76895.0 32717.5 ;
      RECT  76640.0 32582.5 76705.0 32717.5 ;
      RECT  76640.0 33442.5 76705.0 33577.5 ;
      RECT  76830.0 33442.5 76895.0 33577.5 ;
      RECT  76830.0 33442.5 76895.0 33577.5 ;
      RECT  76640.0 33442.5 76705.0 33577.5 ;
      RECT  76567.5 33857.5 76632.5 33992.5 ;
      RECT  76902.5 32307.5 76967.5 32442.5 ;
      RECT  76640.0 33442.5 76705.0 33577.5 ;
      RECT  76830.0 32582.5 76895.0 32717.5 ;
      RECT  77087.5 32482.5 77152.5 32617.5 ;
      RECT  77087.5 32482.5 77152.5 32617.5 ;
      RECT  77535.0 33892.5 77600.0 33957.5 ;
      RECT  77270.0 33892.5 77567.5 33957.5 ;
      RECT  77535.0 33510.0 77600.0 33925.0 ;
      RECT  77345.0 32342.5 77410.0 32407.5 ;
      RECT  77377.5 32342.5 77640.0 32407.5 ;
      RECT  77345.0 32375.0 77410.0 32650.0 ;
      RECT  77345.0 32582.5 77410.0 32717.5 ;
      RECT  77535.0 32582.5 77600.0 32717.5 ;
      RECT  77535.0 32582.5 77600.0 32717.5 ;
      RECT  77345.0 32582.5 77410.0 32717.5 ;
      RECT  77345.0 33442.5 77410.0 33577.5 ;
      RECT  77535.0 33442.5 77600.0 33577.5 ;
      RECT  77535.0 33442.5 77600.0 33577.5 ;
      RECT  77345.0 33442.5 77410.0 33577.5 ;
      RECT  77272.5 33857.5 77337.5 33992.5 ;
      RECT  77607.5 32307.5 77672.5 32442.5 ;
      RECT  77345.0 33442.5 77410.0 33577.5 ;
      RECT  77535.0 32582.5 77600.0 32717.5 ;
      RECT  77792.5 32482.5 77857.5 32617.5 ;
      RECT  77792.5 32482.5 77857.5 32617.5 ;
      RECT  78240.0 33892.5 78305.0 33957.5 ;
      RECT  77975.0 33892.5 78272.5 33957.5 ;
      RECT  78240.0 33510.0 78305.0 33925.0 ;
      RECT  78050.0 32342.5 78115.0 32407.5 ;
      RECT  78082.5 32342.5 78345.0 32407.5 ;
      RECT  78050.0 32375.0 78115.0 32650.0 ;
      RECT  78050.0 32582.5 78115.0 32717.5 ;
      RECT  78240.0 32582.5 78305.0 32717.5 ;
      RECT  78240.0 32582.5 78305.0 32717.5 ;
      RECT  78050.0 32582.5 78115.0 32717.5 ;
      RECT  78050.0 33442.5 78115.0 33577.5 ;
      RECT  78240.0 33442.5 78305.0 33577.5 ;
      RECT  78240.0 33442.5 78305.0 33577.5 ;
      RECT  78050.0 33442.5 78115.0 33577.5 ;
      RECT  77977.5 33857.5 78042.5 33992.5 ;
      RECT  78312.5 32307.5 78377.5 32442.5 ;
      RECT  78050.0 33442.5 78115.0 33577.5 ;
      RECT  78240.0 32582.5 78305.0 32717.5 ;
      RECT  78497.5 32482.5 78562.5 32617.5 ;
      RECT  78497.5 32482.5 78562.5 32617.5 ;
      RECT  78945.0 33892.5 79010.0 33957.5 ;
      RECT  78680.0 33892.5 78977.5 33957.5 ;
      RECT  78945.0 33510.0 79010.0 33925.0 ;
      RECT  78755.0 32342.5 78820.0 32407.5 ;
      RECT  78787.5 32342.5 79050.0 32407.5 ;
      RECT  78755.0 32375.0 78820.0 32650.0 ;
      RECT  78755.0 32582.5 78820.0 32717.5 ;
      RECT  78945.0 32582.5 79010.0 32717.5 ;
      RECT  78945.0 32582.5 79010.0 32717.5 ;
      RECT  78755.0 32582.5 78820.0 32717.5 ;
      RECT  78755.0 33442.5 78820.0 33577.5 ;
      RECT  78945.0 33442.5 79010.0 33577.5 ;
      RECT  78945.0 33442.5 79010.0 33577.5 ;
      RECT  78755.0 33442.5 78820.0 33577.5 ;
      RECT  78682.5 33857.5 78747.5 33992.5 ;
      RECT  79017.5 32307.5 79082.5 32442.5 ;
      RECT  78755.0 33442.5 78820.0 33577.5 ;
      RECT  78945.0 32582.5 79010.0 32717.5 ;
      RECT  79202.5 32482.5 79267.5 32617.5 ;
      RECT  79202.5 32482.5 79267.5 32617.5 ;
      RECT  79650.0 33892.5 79715.0 33957.5 ;
      RECT  79385.0 33892.5 79682.5 33957.5 ;
      RECT  79650.0 33510.0 79715.0 33925.0 ;
      RECT  79460.0 32342.5 79525.0 32407.5 ;
      RECT  79492.5 32342.5 79755.0 32407.5 ;
      RECT  79460.0 32375.0 79525.0 32650.0 ;
      RECT  79460.0 32582.5 79525.0 32717.5 ;
      RECT  79650.0 32582.5 79715.0 32717.5 ;
      RECT  79650.0 32582.5 79715.0 32717.5 ;
      RECT  79460.0 32582.5 79525.0 32717.5 ;
      RECT  79460.0 33442.5 79525.0 33577.5 ;
      RECT  79650.0 33442.5 79715.0 33577.5 ;
      RECT  79650.0 33442.5 79715.0 33577.5 ;
      RECT  79460.0 33442.5 79525.0 33577.5 ;
      RECT  79387.5 33857.5 79452.5 33992.5 ;
      RECT  79722.5 32307.5 79787.5 32442.5 ;
      RECT  79460.0 33442.5 79525.0 33577.5 ;
      RECT  79650.0 32582.5 79715.0 32717.5 ;
      RECT  79907.5 32482.5 79972.5 32617.5 ;
      RECT  79907.5 32482.5 79972.5 32617.5 ;
      RECT  80355.0 33892.5 80420.0 33957.5 ;
      RECT  80090.0 33892.5 80387.5 33957.5 ;
      RECT  80355.0 33510.0 80420.0 33925.0 ;
      RECT  80165.0 32342.5 80230.0 32407.5 ;
      RECT  80197.5 32342.5 80460.0 32407.5 ;
      RECT  80165.0 32375.0 80230.0 32650.0 ;
      RECT  80165.0 32582.5 80230.0 32717.5 ;
      RECT  80355.0 32582.5 80420.0 32717.5 ;
      RECT  80355.0 32582.5 80420.0 32717.5 ;
      RECT  80165.0 32582.5 80230.0 32717.5 ;
      RECT  80165.0 33442.5 80230.0 33577.5 ;
      RECT  80355.0 33442.5 80420.0 33577.5 ;
      RECT  80355.0 33442.5 80420.0 33577.5 ;
      RECT  80165.0 33442.5 80230.0 33577.5 ;
      RECT  80092.5 33857.5 80157.5 33992.5 ;
      RECT  80427.5 32307.5 80492.5 32442.5 ;
      RECT  80165.0 33442.5 80230.0 33577.5 ;
      RECT  80355.0 32582.5 80420.0 32717.5 ;
      RECT  80612.5 32482.5 80677.5 32617.5 ;
      RECT  80612.5 32482.5 80677.5 32617.5 ;
      RECT  81060.0 33892.5 81125.0 33957.5 ;
      RECT  80795.0 33892.5 81092.5 33957.5 ;
      RECT  81060.0 33510.0 81125.0 33925.0 ;
      RECT  80870.0 32342.5 80935.0 32407.5 ;
      RECT  80902.5 32342.5 81165.0 32407.5 ;
      RECT  80870.0 32375.0 80935.0 32650.0 ;
      RECT  80870.0 32582.5 80935.0 32717.5 ;
      RECT  81060.0 32582.5 81125.0 32717.5 ;
      RECT  81060.0 32582.5 81125.0 32717.5 ;
      RECT  80870.0 32582.5 80935.0 32717.5 ;
      RECT  80870.0 33442.5 80935.0 33577.5 ;
      RECT  81060.0 33442.5 81125.0 33577.5 ;
      RECT  81060.0 33442.5 81125.0 33577.5 ;
      RECT  80870.0 33442.5 80935.0 33577.5 ;
      RECT  80797.5 33857.5 80862.5 33992.5 ;
      RECT  81132.5 32307.5 81197.5 32442.5 ;
      RECT  80870.0 33442.5 80935.0 33577.5 ;
      RECT  81060.0 32582.5 81125.0 32717.5 ;
      RECT  81317.5 32482.5 81382.5 32617.5 ;
      RECT  81317.5 32482.5 81382.5 32617.5 ;
      RECT  81765.0 33892.5 81830.0 33957.5 ;
      RECT  81500.0 33892.5 81797.5 33957.5 ;
      RECT  81765.0 33510.0 81830.0 33925.0 ;
      RECT  81575.0 32342.5 81640.0 32407.5 ;
      RECT  81607.5 32342.5 81870.0 32407.5 ;
      RECT  81575.0 32375.0 81640.0 32650.0 ;
      RECT  81575.0 32582.5 81640.0 32717.5 ;
      RECT  81765.0 32582.5 81830.0 32717.5 ;
      RECT  81765.0 32582.5 81830.0 32717.5 ;
      RECT  81575.0 32582.5 81640.0 32717.5 ;
      RECT  81575.0 33442.5 81640.0 33577.5 ;
      RECT  81765.0 33442.5 81830.0 33577.5 ;
      RECT  81765.0 33442.5 81830.0 33577.5 ;
      RECT  81575.0 33442.5 81640.0 33577.5 ;
      RECT  81502.5 33857.5 81567.5 33992.5 ;
      RECT  81837.5 32307.5 81902.5 32442.5 ;
      RECT  81575.0 33442.5 81640.0 33577.5 ;
      RECT  81765.0 32582.5 81830.0 32717.5 ;
      RECT  82022.5 32482.5 82087.5 32617.5 ;
      RECT  82022.5 32482.5 82087.5 32617.5 ;
      RECT  82470.0 33892.5 82535.0 33957.5 ;
      RECT  82205.0 33892.5 82502.5 33957.5 ;
      RECT  82470.0 33510.0 82535.0 33925.0 ;
      RECT  82280.0 32342.5 82345.0 32407.5 ;
      RECT  82312.5 32342.5 82575.0 32407.5 ;
      RECT  82280.0 32375.0 82345.0 32650.0 ;
      RECT  82280.0 32582.5 82345.0 32717.5 ;
      RECT  82470.0 32582.5 82535.0 32717.5 ;
      RECT  82470.0 32582.5 82535.0 32717.5 ;
      RECT  82280.0 32582.5 82345.0 32717.5 ;
      RECT  82280.0 33442.5 82345.0 33577.5 ;
      RECT  82470.0 33442.5 82535.0 33577.5 ;
      RECT  82470.0 33442.5 82535.0 33577.5 ;
      RECT  82280.0 33442.5 82345.0 33577.5 ;
      RECT  82207.5 33857.5 82272.5 33992.5 ;
      RECT  82542.5 32307.5 82607.5 32442.5 ;
      RECT  82280.0 33442.5 82345.0 33577.5 ;
      RECT  82470.0 32582.5 82535.0 32717.5 ;
      RECT  82727.5 32482.5 82792.5 32617.5 ;
      RECT  82727.5 32482.5 82792.5 32617.5 ;
      RECT  83175.0 33892.5 83240.0 33957.5 ;
      RECT  82910.0 33892.5 83207.5 33957.5 ;
      RECT  83175.0 33510.0 83240.0 33925.0 ;
      RECT  82985.0 32342.5 83050.0 32407.5 ;
      RECT  83017.5 32342.5 83280.0 32407.5 ;
      RECT  82985.0 32375.0 83050.0 32650.0 ;
      RECT  82985.0 32582.5 83050.0 32717.5 ;
      RECT  83175.0 32582.5 83240.0 32717.5 ;
      RECT  83175.0 32582.5 83240.0 32717.5 ;
      RECT  82985.0 32582.5 83050.0 32717.5 ;
      RECT  82985.0 33442.5 83050.0 33577.5 ;
      RECT  83175.0 33442.5 83240.0 33577.5 ;
      RECT  83175.0 33442.5 83240.0 33577.5 ;
      RECT  82985.0 33442.5 83050.0 33577.5 ;
      RECT  82912.5 33857.5 82977.5 33992.5 ;
      RECT  83247.5 32307.5 83312.5 32442.5 ;
      RECT  82985.0 33442.5 83050.0 33577.5 ;
      RECT  83175.0 32582.5 83240.0 32717.5 ;
      RECT  83432.5 32482.5 83497.5 32617.5 ;
      RECT  83432.5 32482.5 83497.5 32617.5 ;
      RECT  83880.0 33892.5 83945.0 33957.5 ;
      RECT  83615.0 33892.5 83912.5 33957.5 ;
      RECT  83880.0 33510.0 83945.0 33925.0 ;
      RECT  83690.0 32342.5 83755.0 32407.5 ;
      RECT  83722.5 32342.5 83985.0 32407.5 ;
      RECT  83690.0 32375.0 83755.0 32650.0 ;
      RECT  83690.0 32582.5 83755.0 32717.5 ;
      RECT  83880.0 32582.5 83945.0 32717.5 ;
      RECT  83880.0 32582.5 83945.0 32717.5 ;
      RECT  83690.0 32582.5 83755.0 32717.5 ;
      RECT  83690.0 33442.5 83755.0 33577.5 ;
      RECT  83880.0 33442.5 83945.0 33577.5 ;
      RECT  83880.0 33442.5 83945.0 33577.5 ;
      RECT  83690.0 33442.5 83755.0 33577.5 ;
      RECT  83617.5 33857.5 83682.5 33992.5 ;
      RECT  83952.5 32307.5 84017.5 32442.5 ;
      RECT  83690.0 33442.5 83755.0 33577.5 ;
      RECT  83880.0 32582.5 83945.0 32717.5 ;
      RECT  84137.5 32482.5 84202.5 32617.5 ;
      RECT  84137.5 32482.5 84202.5 32617.5 ;
      RECT  84585.0 33892.5 84650.0 33957.5 ;
      RECT  84320.0 33892.5 84617.5 33957.5 ;
      RECT  84585.0 33510.0 84650.0 33925.0 ;
      RECT  84395.0 32342.5 84460.0 32407.5 ;
      RECT  84427.5 32342.5 84690.0 32407.5 ;
      RECT  84395.0 32375.0 84460.0 32650.0 ;
      RECT  84395.0 32582.5 84460.0 32717.5 ;
      RECT  84585.0 32582.5 84650.0 32717.5 ;
      RECT  84585.0 32582.5 84650.0 32717.5 ;
      RECT  84395.0 32582.5 84460.0 32717.5 ;
      RECT  84395.0 33442.5 84460.0 33577.5 ;
      RECT  84585.0 33442.5 84650.0 33577.5 ;
      RECT  84585.0 33442.5 84650.0 33577.5 ;
      RECT  84395.0 33442.5 84460.0 33577.5 ;
      RECT  84322.5 33857.5 84387.5 33992.5 ;
      RECT  84657.5 32307.5 84722.5 32442.5 ;
      RECT  84395.0 33442.5 84460.0 33577.5 ;
      RECT  84585.0 32582.5 84650.0 32717.5 ;
      RECT  84842.5 32482.5 84907.5 32617.5 ;
      RECT  84842.5 32482.5 84907.5 32617.5 ;
      RECT  85290.0 33892.5 85355.0 33957.5 ;
      RECT  85025.0 33892.5 85322.5 33957.5 ;
      RECT  85290.0 33510.0 85355.0 33925.0 ;
      RECT  85100.0 32342.5 85165.0 32407.5 ;
      RECT  85132.5 32342.5 85395.0 32407.5 ;
      RECT  85100.0 32375.0 85165.0 32650.0 ;
      RECT  85100.0 32582.5 85165.0 32717.5 ;
      RECT  85290.0 32582.5 85355.0 32717.5 ;
      RECT  85290.0 32582.5 85355.0 32717.5 ;
      RECT  85100.0 32582.5 85165.0 32717.5 ;
      RECT  85100.0 33442.5 85165.0 33577.5 ;
      RECT  85290.0 33442.5 85355.0 33577.5 ;
      RECT  85290.0 33442.5 85355.0 33577.5 ;
      RECT  85100.0 33442.5 85165.0 33577.5 ;
      RECT  85027.5 33857.5 85092.5 33992.5 ;
      RECT  85362.5 32307.5 85427.5 32442.5 ;
      RECT  85100.0 33442.5 85165.0 33577.5 ;
      RECT  85290.0 32582.5 85355.0 32717.5 ;
      RECT  85547.5 32482.5 85612.5 32617.5 ;
      RECT  85547.5 32482.5 85612.5 32617.5 ;
      RECT  85995.0 33892.5 86060.0 33957.5 ;
      RECT  85730.0 33892.5 86027.5 33957.5 ;
      RECT  85995.0 33510.0 86060.0 33925.0 ;
      RECT  85805.0 32342.5 85870.0 32407.5 ;
      RECT  85837.5 32342.5 86100.0 32407.5 ;
      RECT  85805.0 32375.0 85870.0 32650.0 ;
      RECT  85805.0 32582.5 85870.0 32717.5 ;
      RECT  85995.0 32582.5 86060.0 32717.5 ;
      RECT  85995.0 32582.5 86060.0 32717.5 ;
      RECT  85805.0 32582.5 85870.0 32717.5 ;
      RECT  85805.0 33442.5 85870.0 33577.5 ;
      RECT  85995.0 33442.5 86060.0 33577.5 ;
      RECT  85995.0 33442.5 86060.0 33577.5 ;
      RECT  85805.0 33442.5 85870.0 33577.5 ;
      RECT  85732.5 33857.5 85797.5 33992.5 ;
      RECT  86067.5 32307.5 86132.5 32442.5 ;
      RECT  85805.0 33442.5 85870.0 33577.5 ;
      RECT  85995.0 32582.5 86060.0 32717.5 ;
      RECT  86252.5 32482.5 86317.5 32617.5 ;
      RECT  86252.5 32482.5 86317.5 32617.5 ;
      RECT  86700.0 33892.5 86765.0 33957.5 ;
      RECT  86435.0 33892.5 86732.5 33957.5 ;
      RECT  86700.0 33510.0 86765.0 33925.0 ;
      RECT  86510.0 32342.5 86575.0 32407.5 ;
      RECT  86542.5 32342.5 86805.0 32407.5 ;
      RECT  86510.0 32375.0 86575.0 32650.0 ;
      RECT  86510.0 32582.5 86575.0 32717.5 ;
      RECT  86700.0 32582.5 86765.0 32717.5 ;
      RECT  86700.0 32582.5 86765.0 32717.5 ;
      RECT  86510.0 32582.5 86575.0 32717.5 ;
      RECT  86510.0 33442.5 86575.0 33577.5 ;
      RECT  86700.0 33442.5 86765.0 33577.5 ;
      RECT  86700.0 33442.5 86765.0 33577.5 ;
      RECT  86510.0 33442.5 86575.0 33577.5 ;
      RECT  86437.5 33857.5 86502.5 33992.5 ;
      RECT  86772.5 32307.5 86837.5 32442.5 ;
      RECT  86510.0 33442.5 86575.0 33577.5 ;
      RECT  86700.0 32582.5 86765.0 32717.5 ;
      RECT  86957.5 32482.5 87022.5 32617.5 ;
      RECT  86957.5 32482.5 87022.5 32617.5 ;
      RECT  87405.0 33892.5 87470.0 33957.5 ;
      RECT  87140.0 33892.5 87437.5 33957.5 ;
      RECT  87405.0 33510.0 87470.0 33925.0 ;
      RECT  87215.0 32342.5 87280.0 32407.5 ;
      RECT  87247.5 32342.5 87510.0 32407.5 ;
      RECT  87215.0 32375.0 87280.0 32650.0 ;
      RECT  87215.0 32582.5 87280.0 32717.5 ;
      RECT  87405.0 32582.5 87470.0 32717.5 ;
      RECT  87405.0 32582.5 87470.0 32717.5 ;
      RECT  87215.0 32582.5 87280.0 32717.5 ;
      RECT  87215.0 33442.5 87280.0 33577.5 ;
      RECT  87405.0 33442.5 87470.0 33577.5 ;
      RECT  87405.0 33442.5 87470.0 33577.5 ;
      RECT  87215.0 33442.5 87280.0 33577.5 ;
      RECT  87142.5 33857.5 87207.5 33992.5 ;
      RECT  87477.5 32307.5 87542.5 32442.5 ;
      RECT  87215.0 33442.5 87280.0 33577.5 ;
      RECT  87405.0 32582.5 87470.0 32717.5 ;
      RECT  87662.5 32482.5 87727.5 32617.5 ;
      RECT  87662.5 32482.5 87727.5 32617.5 ;
      RECT  88110.0 33892.5 88175.0 33957.5 ;
      RECT  87845.0 33892.5 88142.5 33957.5 ;
      RECT  88110.0 33510.0 88175.0 33925.0 ;
      RECT  87920.0 32342.5 87985.0 32407.5 ;
      RECT  87952.5 32342.5 88215.0 32407.5 ;
      RECT  87920.0 32375.0 87985.0 32650.0 ;
      RECT  87920.0 32582.5 87985.0 32717.5 ;
      RECT  88110.0 32582.5 88175.0 32717.5 ;
      RECT  88110.0 32582.5 88175.0 32717.5 ;
      RECT  87920.0 32582.5 87985.0 32717.5 ;
      RECT  87920.0 33442.5 87985.0 33577.5 ;
      RECT  88110.0 33442.5 88175.0 33577.5 ;
      RECT  88110.0 33442.5 88175.0 33577.5 ;
      RECT  87920.0 33442.5 87985.0 33577.5 ;
      RECT  87847.5 33857.5 87912.5 33992.5 ;
      RECT  88182.5 32307.5 88247.5 32442.5 ;
      RECT  87920.0 33442.5 87985.0 33577.5 ;
      RECT  88110.0 32582.5 88175.0 32717.5 ;
      RECT  88367.5 32482.5 88432.5 32617.5 ;
      RECT  88367.5 32482.5 88432.5 32617.5 ;
      RECT  88815.0 33892.5 88880.0 33957.5 ;
      RECT  88550.0 33892.5 88847.5 33957.5 ;
      RECT  88815.0 33510.0 88880.0 33925.0 ;
      RECT  88625.0 32342.5 88690.0 32407.5 ;
      RECT  88657.5 32342.5 88920.0 32407.5 ;
      RECT  88625.0 32375.0 88690.0 32650.0 ;
      RECT  88625.0 32582.5 88690.0 32717.5 ;
      RECT  88815.0 32582.5 88880.0 32717.5 ;
      RECT  88815.0 32582.5 88880.0 32717.5 ;
      RECT  88625.0 32582.5 88690.0 32717.5 ;
      RECT  88625.0 33442.5 88690.0 33577.5 ;
      RECT  88815.0 33442.5 88880.0 33577.5 ;
      RECT  88815.0 33442.5 88880.0 33577.5 ;
      RECT  88625.0 33442.5 88690.0 33577.5 ;
      RECT  88552.5 33857.5 88617.5 33992.5 ;
      RECT  88887.5 32307.5 88952.5 32442.5 ;
      RECT  88625.0 33442.5 88690.0 33577.5 ;
      RECT  88815.0 32582.5 88880.0 32717.5 ;
      RECT  89072.5 32482.5 89137.5 32617.5 ;
      RECT  89072.5 32482.5 89137.5 32617.5 ;
      RECT  89520.0 33892.5 89585.0 33957.5 ;
      RECT  89255.0 33892.5 89552.5 33957.5 ;
      RECT  89520.0 33510.0 89585.0 33925.0 ;
      RECT  89330.0 32342.5 89395.0 32407.5 ;
      RECT  89362.5 32342.5 89625.0 32407.5 ;
      RECT  89330.0 32375.0 89395.0 32650.0 ;
      RECT  89330.0 32582.5 89395.0 32717.5 ;
      RECT  89520.0 32582.5 89585.0 32717.5 ;
      RECT  89520.0 32582.5 89585.0 32717.5 ;
      RECT  89330.0 32582.5 89395.0 32717.5 ;
      RECT  89330.0 33442.5 89395.0 33577.5 ;
      RECT  89520.0 33442.5 89585.0 33577.5 ;
      RECT  89520.0 33442.5 89585.0 33577.5 ;
      RECT  89330.0 33442.5 89395.0 33577.5 ;
      RECT  89257.5 33857.5 89322.5 33992.5 ;
      RECT  89592.5 32307.5 89657.5 32442.5 ;
      RECT  89330.0 33442.5 89395.0 33577.5 ;
      RECT  89520.0 32582.5 89585.0 32717.5 ;
      RECT  89777.5 32482.5 89842.5 32617.5 ;
      RECT  89777.5 32482.5 89842.5 32617.5 ;
      RECT  90225.0 33892.5 90290.0 33957.5 ;
      RECT  89960.0 33892.5 90257.5 33957.5 ;
      RECT  90225.0 33510.0 90290.0 33925.0 ;
      RECT  90035.0 32342.5 90100.0 32407.5 ;
      RECT  90067.5 32342.5 90330.0 32407.5 ;
      RECT  90035.0 32375.0 90100.0 32650.0 ;
      RECT  90035.0 32582.5 90100.0 32717.5 ;
      RECT  90225.0 32582.5 90290.0 32717.5 ;
      RECT  90225.0 32582.5 90290.0 32717.5 ;
      RECT  90035.0 32582.5 90100.0 32717.5 ;
      RECT  90035.0 33442.5 90100.0 33577.5 ;
      RECT  90225.0 33442.5 90290.0 33577.5 ;
      RECT  90225.0 33442.5 90290.0 33577.5 ;
      RECT  90035.0 33442.5 90100.0 33577.5 ;
      RECT  89962.5 33857.5 90027.5 33992.5 ;
      RECT  90297.5 32307.5 90362.5 32442.5 ;
      RECT  90035.0 33442.5 90100.0 33577.5 ;
      RECT  90225.0 32582.5 90290.0 32717.5 ;
      RECT  90482.5 32482.5 90547.5 32617.5 ;
      RECT  90482.5 32482.5 90547.5 32617.5 ;
      RECT  90930.0 33892.5 90995.0 33957.5 ;
      RECT  90665.0 33892.5 90962.5 33957.5 ;
      RECT  90930.0 33510.0 90995.0 33925.0 ;
      RECT  90740.0 32342.5 90805.0 32407.5 ;
      RECT  90772.5 32342.5 91035.0 32407.5 ;
      RECT  90740.0 32375.0 90805.0 32650.0 ;
      RECT  90740.0 32582.5 90805.0 32717.5 ;
      RECT  90930.0 32582.5 90995.0 32717.5 ;
      RECT  90930.0 32582.5 90995.0 32717.5 ;
      RECT  90740.0 32582.5 90805.0 32717.5 ;
      RECT  90740.0 33442.5 90805.0 33577.5 ;
      RECT  90930.0 33442.5 90995.0 33577.5 ;
      RECT  90930.0 33442.5 90995.0 33577.5 ;
      RECT  90740.0 33442.5 90805.0 33577.5 ;
      RECT  90667.5 33857.5 90732.5 33992.5 ;
      RECT  91002.5 32307.5 91067.5 32442.5 ;
      RECT  90740.0 33442.5 90805.0 33577.5 ;
      RECT  90930.0 32582.5 90995.0 32717.5 ;
      RECT  91187.5 32482.5 91252.5 32617.5 ;
      RECT  91187.5 32482.5 91252.5 32617.5 ;
      RECT  91635.0 33892.5 91700.0 33957.5 ;
      RECT  91370.0 33892.5 91667.5 33957.5 ;
      RECT  91635.0 33510.0 91700.0 33925.0 ;
      RECT  91445.0 32342.5 91510.0 32407.5 ;
      RECT  91477.5 32342.5 91740.0 32407.5 ;
      RECT  91445.0 32375.0 91510.0 32650.0 ;
      RECT  91445.0 32582.5 91510.0 32717.5 ;
      RECT  91635.0 32582.5 91700.0 32717.5 ;
      RECT  91635.0 32582.5 91700.0 32717.5 ;
      RECT  91445.0 32582.5 91510.0 32717.5 ;
      RECT  91445.0 33442.5 91510.0 33577.5 ;
      RECT  91635.0 33442.5 91700.0 33577.5 ;
      RECT  91635.0 33442.5 91700.0 33577.5 ;
      RECT  91445.0 33442.5 91510.0 33577.5 ;
      RECT  91372.5 33857.5 91437.5 33992.5 ;
      RECT  91707.5 32307.5 91772.5 32442.5 ;
      RECT  91445.0 33442.5 91510.0 33577.5 ;
      RECT  91635.0 32582.5 91700.0 32717.5 ;
      RECT  91892.5 32482.5 91957.5 32617.5 ;
      RECT  91892.5 32482.5 91957.5 32617.5 ;
      RECT  92340.0 33892.5 92405.0 33957.5 ;
      RECT  92075.0 33892.5 92372.5 33957.5 ;
      RECT  92340.0 33510.0 92405.0 33925.0 ;
      RECT  92150.0 32342.5 92215.0 32407.5 ;
      RECT  92182.5 32342.5 92445.0 32407.5 ;
      RECT  92150.0 32375.0 92215.0 32650.0 ;
      RECT  92150.0 32582.5 92215.0 32717.5 ;
      RECT  92340.0 32582.5 92405.0 32717.5 ;
      RECT  92340.0 32582.5 92405.0 32717.5 ;
      RECT  92150.0 32582.5 92215.0 32717.5 ;
      RECT  92150.0 33442.5 92215.0 33577.5 ;
      RECT  92340.0 33442.5 92405.0 33577.5 ;
      RECT  92340.0 33442.5 92405.0 33577.5 ;
      RECT  92150.0 33442.5 92215.0 33577.5 ;
      RECT  92077.5 33857.5 92142.5 33992.5 ;
      RECT  92412.5 32307.5 92477.5 32442.5 ;
      RECT  92150.0 33442.5 92215.0 33577.5 ;
      RECT  92340.0 32582.5 92405.0 32717.5 ;
      RECT  92597.5 32482.5 92662.5 32617.5 ;
      RECT  92597.5 32482.5 92662.5 32617.5 ;
      RECT  93045.0 33892.5 93110.0 33957.5 ;
      RECT  92780.0 33892.5 93077.5 33957.5 ;
      RECT  93045.0 33510.0 93110.0 33925.0 ;
      RECT  92855.0 32342.5 92920.0 32407.5 ;
      RECT  92887.5 32342.5 93150.0 32407.5 ;
      RECT  92855.0 32375.0 92920.0 32650.0 ;
      RECT  92855.0 32582.5 92920.0 32717.5 ;
      RECT  93045.0 32582.5 93110.0 32717.5 ;
      RECT  93045.0 32582.5 93110.0 32717.5 ;
      RECT  92855.0 32582.5 92920.0 32717.5 ;
      RECT  92855.0 33442.5 92920.0 33577.5 ;
      RECT  93045.0 33442.5 93110.0 33577.5 ;
      RECT  93045.0 33442.5 93110.0 33577.5 ;
      RECT  92855.0 33442.5 92920.0 33577.5 ;
      RECT  92782.5 33857.5 92847.5 33992.5 ;
      RECT  93117.5 32307.5 93182.5 32442.5 ;
      RECT  92855.0 33442.5 92920.0 33577.5 ;
      RECT  93045.0 32582.5 93110.0 32717.5 ;
      RECT  93302.5 32482.5 93367.5 32617.5 ;
      RECT  93302.5 32482.5 93367.5 32617.5 ;
      RECT  93750.0 33892.5 93815.0 33957.5 ;
      RECT  93485.0 33892.5 93782.5 33957.5 ;
      RECT  93750.0 33510.0 93815.0 33925.0 ;
      RECT  93560.0 32342.5 93625.0 32407.5 ;
      RECT  93592.5 32342.5 93855.0 32407.5 ;
      RECT  93560.0 32375.0 93625.0 32650.0 ;
      RECT  93560.0 32582.5 93625.0 32717.5 ;
      RECT  93750.0 32582.5 93815.0 32717.5 ;
      RECT  93750.0 32582.5 93815.0 32717.5 ;
      RECT  93560.0 32582.5 93625.0 32717.5 ;
      RECT  93560.0 33442.5 93625.0 33577.5 ;
      RECT  93750.0 33442.5 93815.0 33577.5 ;
      RECT  93750.0 33442.5 93815.0 33577.5 ;
      RECT  93560.0 33442.5 93625.0 33577.5 ;
      RECT  93487.5 33857.5 93552.5 33992.5 ;
      RECT  93822.5 32307.5 93887.5 32442.5 ;
      RECT  93560.0 33442.5 93625.0 33577.5 ;
      RECT  93750.0 32582.5 93815.0 32717.5 ;
      RECT  94007.5 32482.5 94072.5 32617.5 ;
      RECT  94007.5 32482.5 94072.5 32617.5 ;
      RECT  94455.0 33892.5 94520.0 33957.5 ;
      RECT  94190.0 33892.5 94487.5 33957.5 ;
      RECT  94455.0 33510.0 94520.0 33925.0 ;
      RECT  94265.0 32342.5 94330.0 32407.5 ;
      RECT  94297.5 32342.5 94560.0 32407.5 ;
      RECT  94265.0 32375.0 94330.0 32650.0 ;
      RECT  94265.0 32582.5 94330.0 32717.5 ;
      RECT  94455.0 32582.5 94520.0 32717.5 ;
      RECT  94455.0 32582.5 94520.0 32717.5 ;
      RECT  94265.0 32582.5 94330.0 32717.5 ;
      RECT  94265.0 33442.5 94330.0 33577.5 ;
      RECT  94455.0 33442.5 94520.0 33577.5 ;
      RECT  94455.0 33442.5 94520.0 33577.5 ;
      RECT  94265.0 33442.5 94330.0 33577.5 ;
      RECT  94192.5 33857.5 94257.5 33992.5 ;
      RECT  94527.5 32307.5 94592.5 32442.5 ;
      RECT  94265.0 33442.5 94330.0 33577.5 ;
      RECT  94455.0 32582.5 94520.0 32717.5 ;
      RECT  94712.5 32482.5 94777.5 32617.5 ;
      RECT  94712.5 32482.5 94777.5 32617.5 ;
      RECT  95160.0 33892.5 95225.0 33957.5 ;
      RECT  94895.0 33892.5 95192.5 33957.5 ;
      RECT  95160.0 33510.0 95225.0 33925.0 ;
      RECT  94970.0 32342.5 95035.0 32407.5 ;
      RECT  95002.5 32342.5 95265.0 32407.5 ;
      RECT  94970.0 32375.0 95035.0 32650.0 ;
      RECT  94970.0 32582.5 95035.0 32717.5 ;
      RECT  95160.0 32582.5 95225.0 32717.5 ;
      RECT  95160.0 32582.5 95225.0 32717.5 ;
      RECT  94970.0 32582.5 95035.0 32717.5 ;
      RECT  94970.0 33442.5 95035.0 33577.5 ;
      RECT  95160.0 33442.5 95225.0 33577.5 ;
      RECT  95160.0 33442.5 95225.0 33577.5 ;
      RECT  94970.0 33442.5 95035.0 33577.5 ;
      RECT  94897.5 33857.5 94962.5 33992.5 ;
      RECT  95232.5 32307.5 95297.5 32442.5 ;
      RECT  94970.0 33442.5 95035.0 33577.5 ;
      RECT  95160.0 32582.5 95225.0 32717.5 ;
      RECT  95417.5 32482.5 95482.5 32617.5 ;
      RECT  95417.5 32482.5 95482.5 32617.5 ;
      RECT  95865.0 33892.5 95930.0 33957.5 ;
      RECT  95600.0 33892.5 95897.5 33957.5 ;
      RECT  95865.0 33510.0 95930.0 33925.0 ;
      RECT  95675.0 32342.5 95740.0 32407.5 ;
      RECT  95707.5 32342.5 95970.0 32407.5 ;
      RECT  95675.0 32375.0 95740.0 32650.0 ;
      RECT  95675.0 32582.5 95740.0 32717.5 ;
      RECT  95865.0 32582.5 95930.0 32717.5 ;
      RECT  95865.0 32582.5 95930.0 32717.5 ;
      RECT  95675.0 32582.5 95740.0 32717.5 ;
      RECT  95675.0 33442.5 95740.0 33577.5 ;
      RECT  95865.0 33442.5 95930.0 33577.5 ;
      RECT  95865.0 33442.5 95930.0 33577.5 ;
      RECT  95675.0 33442.5 95740.0 33577.5 ;
      RECT  95602.5 33857.5 95667.5 33992.5 ;
      RECT  95937.5 32307.5 96002.5 32442.5 ;
      RECT  95675.0 33442.5 95740.0 33577.5 ;
      RECT  95865.0 32582.5 95930.0 32717.5 ;
      RECT  96122.5 32482.5 96187.5 32617.5 ;
      RECT  96122.5 32482.5 96187.5 32617.5 ;
      RECT  96570.0 33892.5 96635.0 33957.5 ;
      RECT  96305.0 33892.5 96602.5 33957.5 ;
      RECT  96570.0 33510.0 96635.0 33925.0 ;
      RECT  96380.0 32342.5 96445.0 32407.5 ;
      RECT  96412.5 32342.5 96675.0 32407.5 ;
      RECT  96380.0 32375.0 96445.0 32650.0 ;
      RECT  96380.0 32582.5 96445.0 32717.5 ;
      RECT  96570.0 32582.5 96635.0 32717.5 ;
      RECT  96570.0 32582.5 96635.0 32717.5 ;
      RECT  96380.0 32582.5 96445.0 32717.5 ;
      RECT  96380.0 33442.5 96445.0 33577.5 ;
      RECT  96570.0 33442.5 96635.0 33577.5 ;
      RECT  96570.0 33442.5 96635.0 33577.5 ;
      RECT  96380.0 33442.5 96445.0 33577.5 ;
      RECT  96307.5 33857.5 96372.5 33992.5 ;
      RECT  96642.5 32307.5 96707.5 32442.5 ;
      RECT  96380.0 33442.5 96445.0 33577.5 ;
      RECT  96570.0 32582.5 96635.0 32717.5 ;
      RECT  96827.5 32482.5 96892.5 32617.5 ;
      RECT  96827.5 32482.5 96892.5 32617.5 ;
      RECT  97275.0 33892.5 97340.0 33957.5 ;
      RECT  97010.0 33892.5 97307.5 33957.5 ;
      RECT  97275.0 33510.0 97340.0 33925.0 ;
      RECT  97085.0 32342.5 97150.0 32407.5 ;
      RECT  97117.5 32342.5 97380.0 32407.5 ;
      RECT  97085.0 32375.0 97150.0 32650.0 ;
      RECT  97085.0 32582.5 97150.0 32717.5 ;
      RECT  97275.0 32582.5 97340.0 32717.5 ;
      RECT  97275.0 32582.5 97340.0 32717.5 ;
      RECT  97085.0 32582.5 97150.0 32717.5 ;
      RECT  97085.0 33442.5 97150.0 33577.5 ;
      RECT  97275.0 33442.5 97340.0 33577.5 ;
      RECT  97275.0 33442.5 97340.0 33577.5 ;
      RECT  97085.0 33442.5 97150.0 33577.5 ;
      RECT  97012.5 33857.5 97077.5 33992.5 ;
      RECT  97347.5 32307.5 97412.5 32442.5 ;
      RECT  97085.0 33442.5 97150.0 33577.5 ;
      RECT  97275.0 32582.5 97340.0 32717.5 ;
      RECT  97532.5 32482.5 97597.5 32617.5 ;
      RECT  97532.5 32482.5 97597.5 32617.5 ;
      RECT  97980.0 33892.5 98045.0 33957.5 ;
      RECT  97715.0 33892.5 98012.5 33957.5 ;
      RECT  97980.0 33510.0 98045.0 33925.0 ;
      RECT  97790.0 32342.5 97855.0 32407.5 ;
      RECT  97822.5 32342.5 98085.0 32407.5 ;
      RECT  97790.0 32375.0 97855.0 32650.0 ;
      RECT  97790.0 32582.5 97855.0 32717.5 ;
      RECT  97980.0 32582.5 98045.0 32717.5 ;
      RECT  97980.0 32582.5 98045.0 32717.5 ;
      RECT  97790.0 32582.5 97855.0 32717.5 ;
      RECT  97790.0 33442.5 97855.0 33577.5 ;
      RECT  97980.0 33442.5 98045.0 33577.5 ;
      RECT  97980.0 33442.5 98045.0 33577.5 ;
      RECT  97790.0 33442.5 97855.0 33577.5 ;
      RECT  97717.5 33857.5 97782.5 33992.5 ;
      RECT  98052.5 32307.5 98117.5 32442.5 ;
      RECT  97790.0 33442.5 97855.0 33577.5 ;
      RECT  97980.0 32582.5 98045.0 32717.5 ;
      RECT  98237.5 32482.5 98302.5 32617.5 ;
      RECT  98237.5 32482.5 98302.5 32617.5 ;
      RECT  98685.0 33892.5 98750.0 33957.5 ;
      RECT  98420.0 33892.5 98717.5 33957.5 ;
      RECT  98685.0 33510.0 98750.0 33925.0 ;
      RECT  98495.0 32342.5 98560.0 32407.5 ;
      RECT  98527.5 32342.5 98790.0 32407.5 ;
      RECT  98495.0 32375.0 98560.0 32650.0 ;
      RECT  98495.0 32582.5 98560.0 32717.5 ;
      RECT  98685.0 32582.5 98750.0 32717.5 ;
      RECT  98685.0 32582.5 98750.0 32717.5 ;
      RECT  98495.0 32582.5 98560.0 32717.5 ;
      RECT  98495.0 33442.5 98560.0 33577.5 ;
      RECT  98685.0 33442.5 98750.0 33577.5 ;
      RECT  98685.0 33442.5 98750.0 33577.5 ;
      RECT  98495.0 33442.5 98560.0 33577.5 ;
      RECT  98422.5 33857.5 98487.5 33992.5 ;
      RECT  98757.5 32307.5 98822.5 32442.5 ;
      RECT  98495.0 33442.5 98560.0 33577.5 ;
      RECT  98685.0 32582.5 98750.0 32717.5 ;
      RECT  98942.5 32482.5 99007.5 32617.5 ;
      RECT  98942.5 32482.5 99007.5 32617.5 ;
      RECT  99390.0 33892.5 99455.0 33957.5 ;
      RECT  99125.0 33892.5 99422.5 33957.5 ;
      RECT  99390.0 33510.0 99455.0 33925.0 ;
      RECT  99200.0 32342.5 99265.0 32407.5 ;
      RECT  99232.5 32342.5 99495.0 32407.5 ;
      RECT  99200.0 32375.0 99265.0 32650.0 ;
      RECT  99200.0 32582.5 99265.0 32717.5 ;
      RECT  99390.0 32582.5 99455.0 32717.5 ;
      RECT  99390.0 32582.5 99455.0 32717.5 ;
      RECT  99200.0 32582.5 99265.0 32717.5 ;
      RECT  99200.0 33442.5 99265.0 33577.5 ;
      RECT  99390.0 33442.5 99455.0 33577.5 ;
      RECT  99390.0 33442.5 99455.0 33577.5 ;
      RECT  99200.0 33442.5 99265.0 33577.5 ;
      RECT  99127.5 33857.5 99192.5 33992.5 ;
      RECT  99462.5 32307.5 99527.5 32442.5 ;
      RECT  99200.0 33442.5 99265.0 33577.5 ;
      RECT  99390.0 32582.5 99455.0 32717.5 ;
      RECT  99647.5 32482.5 99712.5 32617.5 ;
      RECT  99647.5 32482.5 99712.5 32617.5 ;
      RECT  100095.0 33892.5 100160.0 33957.5 ;
      RECT  99830.0 33892.5 100127.5 33957.5 ;
      RECT  100095.0 33510.0 100160.0 33925.0 ;
      RECT  99905.0 32342.5 99970.0 32407.5 ;
      RECT  99937.5 32342.5 100200.0 32407.5 ;
      RECT  99905.0 32375.0 99970.0 32650.0 ;
      RECT  99905.0 32582.5 99970.0 32717.5 ;
      RECT  100095.0 32582.5 100160.0 32717.5 ;
      RECT  100095.0 32582.5 100160.0 32717.5 ;
      RECT  99905.0 32582.5 99970.0 32717.5 ;
      RECT  99905.0 33442.5 99970.0 33577.5 ;
      RECT  100095.0 33442.5 100160.0 33577.5 ;
      RECT  100095.0 33442.5 100160.0 33577.5 ;
      RECT  99905.0 33442.5 99970.0 33577.5 ;
      RECT  99832.5 33857.5 99897.5 33992.5 ;
      RECT  100167.5 32307.5 100232.5 32442.5 ;
      RECT  99905.0 33442.5 99970.0 33577.5 ;
      RECT  100095.0 32582.5 100160.0 32717.5 ;
      RECT  100352.5 32482.5 100417.5 32617.5 ;
      RECT  100352.5 32482.5 100417.5 32617.5 ;
      RECT  100800.0 33892.5 100865.0 33957.5 ;
      RECT  100535.0 33892.5 100832.5 33957.5 ;
      RECT  100800.0 33510.0 100865.0 33925.0 ;
      RECT  100610.0 32342.5 100675.0 32407.5 ;
      RECT  100642.5 32342.5 100905.0 32407.5 ;
      RECT  100610.0 32375.0 100675.0 32650.0 ;
      RECT  100610.0 32582.5 100675.0 32717.5 ;
      RECT  100800.0 32582.5 100865.0 32717.5 ;
      RECT  100800.0 32582.5 100865.0 32717.5 ;
      RECT  100610.0 32582.5 100675.0 32717.5 ;
      RECT  100610.0 33442.5 100675.0 33577.5 ;
      RECT  100800.0 33442.5 100865.0 33577.5 ;
      RECT  100800.0 33442.5 100865.0 33577.5 ;
      RECT  100610.0 33442.5 100675.0 33577.5 ;
      RECT  100537.5 33857.5 100602.5 33992.5 ;
      RECT  100872.5 32307.5 100937.5 32442.5 ;
      RECT  100610.0 33442.5 100675.0 33577.5 ;
      RECT  100800.0 32582.5 100865.0 32717.5 ;
      RECT  101057.5 32482.5 101122.5 32617.5 ;
      RECT  101057.5 32482.5 101122.5 32617.5 ;
      RECT  101505.0 33892.5 101570.0 33957.5 ;
      RECT  101240.0 33892.5 101537.5 33957.5 ;
      RECT  101505.0 33510.0 101570.0 33925.0 ;
      RECT  101315.0 32342.5 101380.0 32407.5 ;
      RECT  101347.5 32342.5 101610.0 32407.5 ;
      RECT  101315.0 32375.0 101380.0 32650.0 ;
      RECT  101315.0 32582.5 101380.0 32717.5 ;
      RECT  101505.0 32582.5 101570.0 32717.5 ;
      RECT  101505.0 32582.5 101570.0 32717.5 ;
      RECT  101315.0 32582.5 101380.0 32717.5 ;
      RECT  101315.0 33442.5 101380.0 33577.5 ;
      RECT  101505.0 33442.5 101570.0 33577.5 ;
      RECT  101505.0 33442.5 101570.0 33577.5 ;
      RECT  101315.0 33442.5 101380.0 33577.5 ;
      RECT  101242.5 33857.5 101307.5 33992.5 ;
      RECT  101577.5 32307.5 101642.5 32442.5 ;
      RECT  101315.0 33442.5 101380.0 33577.5 ;
      RECT  101505.0 32582.5 101570.0 32717.5 ;
      RECT  101762.5 32482.5 101827.5 32617.5 ;
      RECT  101762.5 32482.5 101827.5 32617.5 ;
      RECT  102210.0 33892.5 102275.0 33957.5 ;
      RECT  101945.0 33892.5 102242.5 33957.5 ;
      RECT  102210.0 33510.0 102275.0 33925.0 ;
      RECT  102020.0 32342.5 102085.0 32407.5 ;
      RECT  102052.5 32342.5 102315.0 32407.5 ;
      RECT  102020.0 32375.0 102085.0 32650.0 ;
      RECT  102020.0 32582.5 102085.0 32717.5 ;
      RECT  102210.0 32582.5 102275.0 32717.5 ;
      RECT  102210.0 32582.5 102275.0 32717.5 ;
      RECT  102020.0 32582.5 102085.0 32717.5 ;
      RECT  102020.0 33442.5 102085.0 33577.5 ;
      RECT  102210.0 33442.5 102275.0 33577.5 ;
      RECT  102210.0 33442.5 102275.0 33577.5 ;
      RECT  102020.0 33442.5 102085.0 33577.5 ;
      RECT  101947.5 33857.5 102012.5 33992.5 ;
      RECT  102282.5 32307.5 102347.5 32442.5 ;
      RECT  102020.0 33442.5 102085.0 33577.5 ;
      RECT  102210.0 32582.5 102275.0 32717.5 ;
      RECT  102467.5 32482.5 102532.5 32617.5 ;
      RECT  102467.5 32482.5 102532.5 32617.5 ;
      RECT  102915.0 33892.5 102980.0 33957.5 ;
      RECT  102650.0 33892.5 102947.5 33957.5 ;
      RECT  102915.0 33510.0 102980.0 33925.0 ;
      RECT  102725.0 32342.5 102790.0 32407.5 ;
      RECT  102757.5 32342.5 103020.0 32407.5 ;
      RECT  102725.0 32375.0 102790.0 32650.0 ;
      RECT  102725.0 32582.5 102790.0 32717.5 ;
      RECT  102915.0 32582.5 102980.0 32717.5 ;
      RECT  102915.0 32582.5 102980.0 32717.5 ;
      RECT  102725.0 32582.5 102790.0 32717.5 ;
      RECT  102725.0 33442.5 102790.0 33577.5 ;
      RECT  102915.0 33442.5 102980.0 33577.5 ;
      RECT  102915.0 33442.5 102980.0 33577.5 ;
      RECT  102725.0 33442.5 102790.0 33577.5 ;
      RECT  102652.5 33857.5 102717.5 33992.5 ;
      RECT  102987.5 32307.5 103052.5 32442.5 ;
      RECT  102725.0 33442.5 102790.0 33577.5 ;
      RECT  102915.0 32582.5 102980.0 32717.5 ;
      RECT  103172.5 32482.5 103237.5 32617.5 ;
      RECT  103172.5 32482.5 103237.5 32617.5 ;
      RECT  103620.0 33892.5 103685.0 33957.5 ;
      RECT  103355.0 33892.5 103652.5 33957.5 ;
      RECT  103620.0 33510.0 103685.0 33925.0 ;
      RECT  103430.0 32342.5 103495.0 32407.5 ;
      RECT  103462.5 32342.5 103725.0 32407.5 ;
      RECT  103430.0 32375.0 103495.0 32650.0 ;
      RECT  103430.0 32582.5 103495.0 32717.5 ;
      RECT  103620.0 32582.5 103685.0 32717.5 ;
      RECT  103620.0 32582.5 103685.0 32717.5 ;
      RECT  103430.0 32582.5 103495.0 32717.5 ;
      RECT  103430.0 33442.5 103495.0 33577.5 ;
      RECT  103620.0 33442.5 103685.0 33577.5 ;
      RECT  103620.0 33442.5 103685.0 33577.5 ;
      RECT  103430.0 33442.5 103495.0 33577.5 ;
      RECT  103357.5 33857.5 103422.5 33992.5 ;
      RECT  103692.5 32307.5 103757.5 32442.5 ;
      RECT  103430.0 33442.5 103495.0 33577.5 ;
      RECT  103620.0 32582.5 103685.0 32717.5 ;
      RECT  103877.5 32482.5 103942.5 32617.5 ;
      RECT  103877.5 32482.5 103942.5 32617.5 ;
      RECT  104325.0 33892.5 104390.0 33957.5 ;
      RECT  104060.0 33892.5 104357.5 33957.5 ;
      RECT  104325.0 33510.0 104390.0 33925.0 ;
      RECT  104135.0 32342.5 104200.0 32407.5 ;
      RECT  104167.5 32342.5 104430.0 32407.5 ;
      RECT  104135.0 32375.0 104200.0 32650.0 ;
      RECT  104135.0 32582.5 104200.0 32717.5 ;
      RECT  104325.0 32582.5 104390.0 32717.5 ;
      RECT  104325.0 32582.5 104390.0 32717.5 ;
      RECT  104135.0 32582.5 104200.0 32717.5 ;
      RECT  104135.0 33442.5 104200.0 33577.5 ;
      RECT  104325.0 33442.5 104390.0 33577.5 ;
      RECT  104325.0 33442.5 104390.0 33577.5 ;
      RECT  104135.0 33442.5 104200.0 33577.5 ;
      RECT  104062.5 33857.5 104127.5 33992.5 ;
      RECT  104397.5 32307.5 104462.5 32442.5 ;
      RECT  104135.0 33442.5 104200.0 33577.5 ;
      RECT  104325.0 32582.5 104390.0 32717.5 ;
      RECT  104582.5 32482.5 104647.5 32617.5 ;
      RECT  104582.5 32482.5 104647.5 32617.5 ;
      RECT  105030.0 33892.5 105095.0 33957.5 ;
      RECT  104765.0 33892.5 105062.5 33957.5 ;
      RECT  105030.0 33510.0 105095.0 33925.0 ;
      RECT  104840.0 32342.5 104905.0 32407.5 ;
      RECT  104872.5 32342.5 105135.0 32407.5 ;
      RECT  104840.0 32375.0 104905.0 32650.0 ;
      RECT  104840.0 32582.5 104905.0 32717.5 ;
      RECT  105030.0 32582.5 105095.0 32717.5 ;
      RECT  105030.0 32582.5 105095.0 32717.5 ;
      RECT  104840.0 32582.5 104905.0 32717.5 ;
      RECT  104840.0 33442.5 104905.0 33577.5 ;
      RECT  105030.0 33442.5 105095.0 33577.5 ;
      RECT  105030.0 33442.5 105095.0 33577.5 ;
      RECT  104840.0 33442.5 104905.0 33577.5 ;
      RECT  104767.5 33857.5 104832.5 33992.5 ;
      RECT  105102.5 32307.5 105167.5 32442.5 ;
      RECT  104840.0 33442.5 104905.0 33577.5 ;
      RECT  105030.0 32582.5 105095.0 32717.5 ;
      RECT  105287.5 32482.5 105352.5 32617.5 ;
      RECT  105287.5 32482.5 105352.5 32617.5 ;
      RECT  105735.0 33892.5 105800.0 33957.5 ;
      RECT  105470.0 33892.5 105767.5 33957.5 ;
      RECT  105735.0 33510.0 105800.0 33925.0 ;
      RECT  105545.0 32342.5 105610.0 32407.5 ;
      RECT  105577.5 32342.5 105840.0 32407.5 ;
      RECT  105545.0 32375.0 105610.0 32650.0 ;
      RECT  105545.0 32582.5 105610.0 32717.5 ;
      RECT  105735.0 32582.5 105800.0 32717.5 ;
      RECT  105735.0 32582.5 105800.0 32717.5 ;
      RECT  105545.0 32582.5 105610.0 32717.5 ;
      RECT  105545.0 33442.5 105610.0 33577.5 ;
      RECT  105735.0 33442.5 105800.0 33577.5 ;
      RECT  105735.0 33442.5 105800.0 33577.5 ;
      RECT  105545.0 33442.5 105610.0 33577.5 ;
      RECT  105472.5 33857.5 105537.5 33992.5 ;
      RECT  105807.5 32307.5 105872.5 32442.5 ;
      RECT  105545.0 33442.5 105610.0 33577.5 ;
      RECT  105735.0 32582.5 105800.0 32717.5 ;
      RECT  105992.5 32482.5 106057.5 32617.5 ;
      RECT  105992.5 32482.5 106057.5 32617.5 ;
      RECT  106440.0 33892.5 106505.0 33957.5 ;
      RECT  106175.0 33892.5 106472.5 33957.5 ;
      RECT  106440.0 33510.0 106505.0 33925.0 ;
      RECT  106250.0 32342.5 106315.0 32407.5 ;
      RECT  106282.5 32342.5 106545.0 32407.5 ;
      RECT  106250.0 32375.0 106315.0 32650.0 ;
      RECT  106250.0 32582.5 106315.0 32717.5 ;
      RECT  106440.0 32582.5 106505.0 32717.5 ;
      RECT  106440.0 32582.5 106505.0 32717.5 ;
      RECT  106250.0 32582.5 106315.0 32717.5 ;
      RECT  106250.0 33442.5 106315.0 33577.5 ;
      RECT  106440.0 33442.5 106505.0 33577.5 ;
      RECT  106440.0 33442.5 106505.0 33577.5 ;
      RECT  106250.0 33442.5 106315.0 33577.5 ;
      RECT  106177.5 33857.5 106242.5 33992.5 ;
      RECT  106512.5 32307.5 106577.5 32442.5 ;
      RECT  106250.0 33442.5 106315.0 33577.5 ;
      RECT  106440.0 32582.5 106505.0 32717.5 ;
      RECT  106697.5 32482.5 106762.5 32617.5 ;
      RECT  106697.5 32482.5 106762.5 32617.5 ;
      RECT  107145.0 33892.5 107210.0 33957.5 ;
      RECT  106880.0 33892.5 107177.5 33957.5 ;
      RECT  107145.0 33510.0 107210.0 33925.0 ;
      RECT  106955.0 32342.5 107020.0 32407.5 ;
      RECT  106987.5 32342.5 107250.0 32407.5 ;
      RECT  106955.0 32375.0 107020.0 32650.0 ;
      RECT  106955.0 32582.5 107020.0 32717.5 ;
      RECT  107145.0 32582.5 107210.0 32717.5 ;
      RECT  107145.0 32582.5 107210.0 32717.5 ;
      RECT  106955.0 32582.5 107020.0 32717.5 ;
      RECT  106955.0 33442.5 107020.0 33577.5 ;
      RECT  107145.0 33442.5 107210.0 33577.5 ;
      RECT  107145.0 33442.5 107210.0 33577.5 ;
      RECT  106955.0 33442.5 107020.0 33577.5 ;
      RECT  106882.5 33857.5 106947.5 33992.5 ;
      RECT  107217.5 32307.5 107282.5 32442.5 ;
      RECT  106955.0 33442.5 107020.0 33577.5 ;
      RECT  107145.0 32582.5 107210.0 32717.5 ;
      RECT  107402.5 32482.5 107467.5 32617.5 ;
      RECT  107402.5 32482.5 107467.5 32617.5 ;
      RECT  17615.0 32097.5 17480.0 32162.5 ;
      RECT  18320.0 31957.5 18185.0 32022.5 ;
      RECT  19025.0 31817.5 18890.0 31882.5 ;
      RECT  19730.0 31677.5 19595.0 31742.5 ;
      RECT  20435.0 32097.5 20300.0 32162.5 ;
      RECT  21140.0 31957.5 21005.0 32022.5 ;
      RECT  21845.0 31817.5 21710.0 31882.5 ;
      RECT  22550.0 31677.5 22415.0 31742.5 ;
      RECT  23255.0 32097.5 23120.0 32162.5 ;
      RECT  23960.0 31957.5 23825.0 32022.5 ;
      RECT  24665.0 31817.5 24530.0 31882.5 ;
      RECT  25370.0 31677.5 25235.0 31742.5 ;
      RECT  26075.0 32097.5 25940.0 32162.5 ;
      RECT  26780.0 31957.5 26645.0 32022.5 ;
      RECT  27485.0 31817.5 27350.0 31882.5 ;
      RECT  28190.0 31677.5 28055.0 31742.5 ;
      RECT  28895.0 32097.5 28760.0 32162.5 ;
      RECT  29600.0 31957.5 29465.0 32022.5 ;
      RECT  30305.0 31817.5 30170.0 31882.5 ;
      RECT  31010.0 31677.5 30875.0 31742.5 ;
      RECT  31715.0 32097.5 31580.0 32162.5 ;
      RECT  32420.0 31957.5 32285.0 32022.5 ;
      RECT  33125.0 31817.5 32990.0 31882.5 ;
      RECT  33830.0 31677.5 33695.0 31742.5 ;
      RECT  34535.0 32097.5 34400.0 32162.5 ;
      RECT  35240.0 31957.5 35105.0 32022.5 ;
      RECT  35945.0 31817.5 35810.0 31882.5 ;
      RECT  36650.0 31677.5 36515.0 31742.5 ;
      RECT  37355.0 32097.5 37220.0 32162.5 ;
      RECT  38060.0 31957.5 37925.0 32022.5 ;
      RECT  38765.0 31817.5 38630.0 31882.5 ;
      RECT  39470.0 31677.5 39335.0 31742.5 ;
      RECT  40175.0 32097.5 40040.0 32162.5 ;
      RECT  40880.0 31957.5 40745.0 32022.5 ;
      RECT  41585.0 31817.5 41450.0 31882.5 ;
      RECT  42290.0 31677.5 42155.0 31742.5 ;
      RECT  42995.0 32097.5 42860.0 32162.5 ;
      RECT  43700.0 31957.5 43565.0 32022.5 ;
      RECT  44405.0 31817.5 44270.0 31882.5 ;
      RECT  45110.0 31677.5 44975.0 31742.5 ;
      RECT  45815.0 32097.5 45680.0 32162.5 ;
      RECT  46520.0 31957.5 46385.0 32022.5 ;
      RECT  47225.0 31817.5 47090.0 31882.5 ;
      RECT  47930.0 31677.5 47795.0 31742.5 ;
      RECT  48635.0 32097.5 48500.0 32162.5 ;
      RECT  49340.0 31957.5 49205.0 32022.5 ;
      RECT  50045.0 31817.5 49910.0 31882.5 ;
      RECT  50750.0 31677.5 50615.0 31742.5 ;
      RECT  51455.0 32097.5 51320.0 32162.5 ;
      RECT  52160.0 31957.5 52025.0 32022.5 ;
      RECT  52865.0 31817.5 52730.0 31882.5 ;
      RECT  53570.0 31677.5 53435.0 31742.5 ;
      RECT  54275.0 32097.5 54140.0 32162.5 ;
      RECT  54980.0 31957.5 54845.0 32022.5 ;
      RECT  55685.0 31817.5 55550.0 31882.5 ;
      RECT  56390.0 31677.5 56255.0 31742.5 ;
      RECT  57095.0 32097.5 56960.0 32162.5 ;
      RECT  57800.0 31957.5 57665.0 32022.5 ;
      RECT  58505.0 31817.5 58370.0 31882.5 ;
      RECT  59210.0 31677.5 59075.0 31742.5 ;
      RECT  59915.0 32097.5 59780.0 32162.5 ;
      RECT  60620.0 31957.5 60485.0 32022.5 ;
      RECT  61325.0 31817.5 61190.0 31882.5 ;
      RECT  62030.0 31677.5 61895.0 31742.5 ;
      RECT  62735.0 32097.5 62600.0 32162.5 ;
      RECT  63440.0 31957.5 63305.0 32022.5 ;
      RECT  64145.0 31817.5 64010.0 31882.5 ;
      RECT  64850.0 31677.5 64715.0 31742.5 ;
      RECT  65555.0 32097.5 65420.0 32162.5 ;
      RECT  66260.0 31957.5 66125.0 32022.5 ;
      RECT  66965.0 31817.5 66830.0 31882.5 ;
      RECT  67670.0 31677.5 67535.0 31742.5 ;
      RECT  68375.0 32097.5 68240.0 32162.5 ;
      RECT  69080.0 31957.5 68945.0 32022.5 ;
      RECT  69785.0 31817.5 69650.0 31882.5 ;
      RECT  70490.0 31677.5 70355.0 31742.5 ;
      RECT  71195.0 32097.5 71060.0 32162.5 ;
      RECT  71900.0 31957.5 71765.0 32022.5 ;
      RECT  72605.0 31817.5 72470.0 31882.5 ;
      RECT  73310.0 31677.5 73175.0 31742.5 ;
      RECT  74015.0 32097.5 73880.0 32162.5 ;
      RECT  74720.0 31957.5 74585.0 32022.5 ;
      RECT  75425.0 31817.5 75290.0 31882.5 ;
      RECT  76130.0 31677.5 75995.0 31742.5 ;
      RECT  76835.0 32097.5 76700.0 32162.5 ;
      RECT  77540.0 31957.5 77405.0 32022.5 ;
      RECT  78245.0 31817.5 78110.0 31882.5 ;
      RECT  78950.0 31677.5 78815.0 31742.5 ;
      RECT  79655.0 32097.5 79520.0 32162.5 ;
      RECT  80360.0 31957.5 80225.0 32022.5 ;
      RECT  81065.0 31817.5 80930.0 31882.5 ;
      RECT  81770.0 31677.5 81635.0 31742.5 ;
      RECT  82475.0 32097.5 82340.0 32162.5 ;
      RECT  83180.0 31957.5 83045.0 32022.5 ;
      RECT  83885.0 31817.5 83750.0 31882.5 ;
      RECT  84590.0 31677.5 84455.0 31742.5 ;
      RECT  85295.0 32097.5 85160.0 32162.5 ;
      RECT  86000.0 31957.5 85865.0 32022.5 ;
      RECT  86705.0 31817.5 86570.0 31882.5 ;
      RECT  87410.0 31677.5 87275.0 31742.5 ;
      RECT  88115.0 32097.5 87980.0 32162.5 ;
      RECT  88820.0 31957.5 88685.0 32022.5 ;
      RECT  89525.0 31817.5 89390.0 31882.5 ;
      RECT  90230.0 31677.5 90095.0 31742.5 ;
      RECT  90935.0 32097.5 90800.0 32162.5 ;
      RECT  91640.0 31957.5 91505.0 32022.5 ;
      RECT  92345.0 31817.5 92210.0 31882.5 ;
      RECT  93050.0 31677.5 92915.0 31742.5 ;
      RECT  93755.0 32097.5 93620.0 32162.5 ;
      RECT  94460.0 31957.5 94325.0 32022.5 ;
      RECT  95165.0 31817.5 95030.0 31882.5 ;
      RECT  95870.0 31677.5 95735.0 31742.5 ;
      RECT  96575.0 32097.5 96440.0 32162.5 ;
      RECT  97280.0 31957.5 97145.0 32022.5 ;
      RECT  97985.0 31817.5 97850.0 31882.5 ;
      RECT  98690.0 31677.5 98555.0 31742.5 ;
      RECT  99395.0 32097.5 99260.0 32162.5 ;
      RECT  100100.0 31957.5 99965.0 32022.5 ;
      RECT  100805.0 31817.5 100670.0 31882.5 ;
      RECT  101510.0 31677.5 101375.0 31742.5 ;
      RECT  102215.0 32097.5 102080.0 32162.5 ;
      RECT  102920.0 31957.5 102785.0 32022.5 ;
      RECT  103625.0 31817.5 103490.0 31882.5 ;
      RECT  104330.0 31677.5 104195.0 31742.5 ;
      RECT  105035.0 32097.5 104900.0 32162.5 ;
      RECT  105740.0 31957.5 105605.0 32022.5 ;
      RECT  106445.0 31817.5 106310.0 31882.5 ;
      RECT  107150.0 31677.5 107015.0 31742.5 ;
      RECT  17480.0 31537.5 17345.0 31602.5 ;
      RECT  17680.0 31397.5 17545.0 31462.5 ;
      RECT  18185.0 31537.5 18050.0 31602.5 ;
      RECT  18385.0 31397.5 18250.0 31462.5 ;
      RECT  18890.0 31537.5 18755.0 31602.5 ;
      RECT  19090.0 31397.5 18955.0 31462.5 ;
      RECT  19595.0 31537.5 19460.0 31602.5 ;
      RECT  19795.0 31397.5 19660.0 31462.5 ;
      RECT  20300.0 31537.5 20165.0 31602.5 ;
      RECT  20500.0 31397.5 20365.0 31462.5 ;
      RECT  21005.0 31537.5 20870.0 31602.5 ;
      RECT  21205.0 31397.5 21070.0 31462.5 ;
      RECT  21710.0 31537.5 21575.0 31602.5 ;
      RECT  21910.0 31397.5 21775.0 31462.5 ;
      RECT  22415.0 31537.5 22280.0 31602.5 ;
      RECT  22615.0 31397.5 22480.0 31462.5 ;
      RECT  23120.0 31537.5 22985.0 31602.5 ;
      RECT  23320.0 31397.5 23185.0 31462.5 ;
      RECT  23825.0 31537.5 23690.0 31602.5 ;
      RECT  24025.0 31397.5 23890.0 31462.5 ;
      RECT  24530.0 31537.5 24395.0 31602.5 ;
      RECT  24730.0 31397.5 24595.0 31462.5 ;
      RECT  25235.0 31537.5 25100.0 31602.5 ;
      RECT  25435.0 31397.5 25300.0 31462.5 ;
      RECT  25940.0 31537.5 25805.0 31602.5 ;
      RECT  26140.0 31397.5 26005.0 31462.5 ;
      RECT  26645.0 31537.5 26510.0 31602.5 ;
      RECT  26845.0 31397.5 26710.0 31462.5 ;
      RECT  27350.0 31537.5 27215.0 31602.5 ;
      RECT  27550.0 31397.5 27415.0 31462.5 ;
      RECT  28055.0 31537.5 27920.0 31602.5 ;
      RECT  28255.0 31397.5 28120.0 31462.5 ;
      RECT  28760.0 31537.5 28625.0 31602.5 ;
      RECT  28960.0 31397.5 28825.0 31462.5 ;
      RECT  29465.0 31537.5 29330.0 31602.5 ;
      RECT  29665.0 31397.5 29530.0 31462.5 ;
      RECT  30170.0 31537.5 30035.0 31602.5 ;
      RECT  30370.0 31397.5 30235.0 31462.5 ;
      RECT  30875.0 31537.5 30740.0 31602.5 ;
      RECT  31075.0 31397.5 30940.0 31462.5 ;
      RECT  31580.0 31537.5 31445.0 31602.5 ;
      RECT  31780.0 31397.5 31645.0 31462.5 ;
      RECT  32285.0 31537.5 32150.0 31602.5 ;
      RECT  32485.0 31397.5 32350.0 31462.5 ;
      RECT  32990.0 31537.5 32855.0 31602.5 ;
      RECT  33190.0 31397.5 33055.0 31462.5 ;
      RECT  33695.0 31537.5 33560.0 31602.5 ;
      RECT  33895.0 31397.5 33760.0 31462.5 ;
      RECT  34400.0 31537.5 34265.0 31602.5 ;
      RECT  34600.0 31397.5 34465.0 31462.5 ;
      RECT  35105.0 31537.5 34970.0 31602.5 ;
      RECT  35305.0 31397.5 35170.0 31462.5 ;
      RECT  35810.0 31537.5 35675.0 31602.5 ;
      RECT  36010.0 31397.5 35875.0 31462.5 ;
      RECT  36515.0 31537.5 36380.0 31602.5 ;
      RECT  36715.0 31397.5 36580.0 31462.5 ;
      RECT  37220.0 31537.5 37085.0 31602.5 ;
      RECT  37420.0 31397.5 37285.0 31462.5 ;
      RECT  37925.0 31537.5 37790.0 31602.5 ;
      RECT  38125.0 31397.5 37990.0 31462.5 ;
      RECT  38630.0 31537.5 38495.0 31602.5 ;
      RECT  38830.0 31397.5 38695.0 31462.5 ;
      RECT  39335.0 31537.5 39200.0 31602.5 ;
      RECT  39535.0 31397.5 39400.0 31462.5 ;
      RECT  40040.0 31537.5 39905.0 31602.5 ;
      RECT  40240.0 31397.5 40105.0 31462.5 ;
      RECT  40745.0 31537.5 40610.0 31602.5 ;
      RECT  40945.0 31397.5 40810.0 31462.5 ;
      RECT  41450.0 31537.5 41315.0 31602.5 ;
      RECT  41650.0 31397.5 41515.0 31462.5 ;
      RECT  42155.0 31537.5 42020.0 31602.5 ;
      RECT  42355.0 31397.5 42220.0 31462.5 ;
      RECT  42860.0 31537.5 42725.0 31602.5 ;
      RECT  43060.0 31397.5 42925.0 31462.5 ;
      RECT  43565.0 31537.5 43430.0 31602.5 ;
      RECT  43765.0 31397.5 43630.0 31462.5 ;
      RECT  44270.0 31537.5 44135.0 31602.5 ;
      RECT  44470.0 31397.5 44335.0 31462.5 ;
      RECT  44975.0 31537.5 44840.0 31602.5 ;
      RECT  45175.0 31397.5 45040.0 31462.5 ;
      RECT  45680.0 31537.5 45545.0 31602.5 ;
      RECT  45880.0 31397.5 45745.0 31462.5 ;
      RECT  46385.0 31537.5 46250.0 31602.5 ;
      RECT  46585.0 31397.5 46450.0 31462.5 ;
      RECT  47090.0 31537.5 46955.0 31602.5 ;
      RECT  47290.0 31397.5 47155.0 31462.5 ;
      RECT  47795.0 31537.5 47660.0 31602.5 ;
      RECT  47995.0 31397.5 47860.0 31462.5 ;
      RECT  48500.0 31537.5 48365.0 31602.5 ;
      RECT  48700.0 31397.5 48565.0 31462.5 ;
      RECT  49205.0 31537.5 49070.0 31602.5 ;
      RECT  49405.0 31397.5 49270.0 31462.5 ;
      RECT  49910.0 31537.5 49775.0 31602.5 ;
      RECT  50110.0 31397.5 49975.0 31462.5 ;
      RECT  50615.0 31537.5 50480.0 31602.5 ;
      RECT  50815.0 31397.5 50680.0 31462.5 ;
      RECT  51320.0 31537.5 51185.0 31602.5 ;
      RECT  51520.0 31397.5 51385.0 31462.5 ;
      RECT  52025.0 31537.5 51890.0 31602.5 ;
      RECT  52225.0 31397.5 52090.0 31462.5 ;
      RECT  52730.0 31537.5 52595.0 31602.5 ;
      RECT  52930.0 31397.5 52795.0 31462.5 ;
      RECT  53435.0 31537.5 53300.0 31602.5 ;
      RECT  53635.0 31397.5 53500.0 31462.5 ;
      RECT  54140.0 31537.5 54005.0 31602.5 ;
      RECT  54340.0 31397.5 54205.0 31462.5 ;
      RECT  54845.0 31537.5 54710.0 31602.5 ;
      RECT  55045.0 31397.5 54910.0 31462.5 ;
      RECT  55550.0 31537.5 55415.0 31602.5 ;
      RECT  55750.0 31397.5 55615.0 31462.5 ;
      RECT  56255.0 31537.5 56120.0 31602.5 ;
      RECT  56455.0 31397.5 56320.0 31462.5 ;
      RECT  56960.0 31537.5 56825.0 31602.5 ;
      RECT  57160.0 31397.5 57025.0 31462.5 ;
      RECT  57665.0 31537.5 57530.0 31602.5 ;
      RECT  57865.0 31397.5 57730.0 31462.5 ;
      RECT  58370.0 31537.5 58235.0 31602.5 ;
      RECT  58570.0 31397.5 58435.0 31462.5 ;
      RECT  59075.0 31537.5 58940.0 31602.5 ;
      RECT  59275.0 31397.5 59140.0 31462.5 ;
      RECT  59780.0 31537.5 59645.0 31602.5 ;
      RECT  59980.0 31397.5 59845.0 31462.5 ;
      RECT  60485.0 31537.5 60350.0 31602.5 ;
      RECT  60685.0 31397.5 60550.0 31462.5 ;
      RECT  61190.0 31537.5 61055.0 31602.5 ;
      RECT  61390.0 31397.5 61255.0 31462.5 ;
      RECT  61895.0 31537.5 61760.0 31602.5 ;
      RECT  62095.0 31397.5 61960.0 31462.5 ;
      RECT  62600.0 31537.5 62465.0 31602.5 ;
      RECT  62800.0 31397.5 62665.0 31462.5 ;
      RECT  63305.0 31537.5 63170.0 31602.5 ;
      RECT  63505.0 31397.5 63370.0 31462.5 ;
      RECT  64010.0 31537.5 63875.0 31602.5 ;
      RECT  64210.0 31397.5 64075.0 31462.5 ;
      RECT  64715.0 31537.5 64580.0 31602.5 ;
      RECT  64915.0 31397.5 64780.0 31462.5 ;
      RECT  65420.0 31537.5 65285.0 31602.5 ;
      RECT  65620.0 31397.5 65485.0 31462.5 ;
      RECT  66125.0 31537.5 65990.0 31602.5 ;
      RECT  66325.0 31397.5 66190.0 31462.5 ;
      RECT  66830.0 31537.5 66695.0 31602.5 ;
      RECT  67030.0 31397.5 66895.0 31462.5 ;
      RECT  67535.0 31537.5 67400.0 31602.5 ;
      RECT  67735.0 31397.5 67600.0 31462.5 ;
      RECT  68240.0 31537.5 68105.0 31602.5 ;
      RECT  68440.0 31397.5 68305.0 31462.5 ;
      RECT  68945.0 31537.5 68810.0 31602.5 ;
      RECT  69145.0 31397.5 69010.0 31462.5 ;
      RECT  69650.0 31537.5 69515.0 31602.5 ;
      RECT  69850.0 31397.5 69715.0 31462.5 ;
      RECT  70355.0 31537.5 70220.0 31602.5 ;
      RECT  70555.0 31397.5 70420.0 31462.5 ;
      RECT  71060.0 31537.5 70925.0 31602.5 ;
      RECT  71260.0 31397.5 71125.0 31462.5 ;
      RECT  71765.0 31537.5 71630.0 31602.5 ;
      RECT  71965.0 31397.5 71830.0 31462.5 ;
      RECT  72470.0 31537.5 72335.0 31602.5 ;
      RECT  72670.0 31397.5 72535.0 31462.5 ;
      RECT  73175.0 31537.5 73040.0 31602.5 ;
      RECT  73375.0 31397.5 73240.0 31462.5 ;
      RECT  73880.0 31537.5 73745.0 31602.5 ;
      RECT  74080.0 31397.5 73945.0 31462.5 ;
      RECT  74585.0 31537.5 74450.0 31602.5 ;
      RECT  74785.0 31397.5 74650.0 31462.5 ;
      RECT  75290.0 31537.5 75155.0 31602.5 ;
      RECT  75490.0 31397.5 75355.0 31462.5 ;
      RECT  75995.0 31537.5 75860.0 31602.5 ;
      RECT  76195.0 31397.5 76060.0 31462.5 ;
      RECT  76700.0 31537.5 76565.0 31602.5 ;
      RECT  76900.0 31397.5 76765.0 31462.5 ;
      RECT  77405.0 31537.5 77270.0 31602.5 ;
      RECT  77605.0 31397.5 77470.0 31462.5 ;
      RECT  78110.0 31537.5 77975.0 31602.5 ;
      RECT  78310.0 31397.5 78175.0 31462.5 ;
      RECT  78815.0 31537.5 78680.0 31602.5 ;
      RECT  79015.0 31397.5 78880.0 31462.5 ;
      RECT  79520.0 31537.5 79385.0 31602.5 ;
      RECT  79720.0 31397.5 79585.0 31462.5 ;
      RECT  80225.0 31537.5 80090.0 31602.5 ;
      RECT  80425.0 31397.5 80290.0 31462.5 ;
      RECT  80930.0 31537.5 80795.0 31602.5 ;
      RECT  81130.0 31397.5 80995.0 31462.5 ;
      RECT  81635.0 31537.5 81500.0 31602.5 ;
      RECT  81835.0 31397.5 81700.0 31462.5 ;
      RECT  82340.0 31537.5 82205.0 31602.5 ;
      RECT  82540.0 31397.5 82405.0 31462.5 ;
      RECT  83045.0 31537.5 82910.0 31602.5 ;
      RECT  83245.0 31397.5 83110.0 31462.5 ;
      RECT  83750.0 31537.5 83615.0 31602.5 ;
      RECT  83950.0 31397.5 83815.0 31462.5 ;
      RECT  84455.0 31537.5 84320.0 31602.5 ;
      RECT  84655.0 31397.5 84520.0 31462.5 ;
      RECT  85160.0 31537.5 85025.0 31602.5 ;
      RECT  85360.0 31397.5 85225.0 31462.5 ;
      RECT  85865.0 31537.5 85730.0 31602.5 ;
      RECT  86065.0 31397.5 85930.0 31462.5 ;
      RECT  86570.0 31537.5 86435.0 31602.5 ;
      RECT  86770.0 31397.5 86635.0 31462.5 ;
      RECT  87275.0 31537.5 87140.0 31602.5 ;
      RECT  87475.0 31397.5 87340.0 31462.5 ;
      RECT  87980.0 31537.5 87845.0 31602.5 ;
      RECT  88180.0 31397.5 88045.0 31462.5 ;
      RECT  88685.0 31537.5 88550.0 31602.5 ;
      RECT  88885.0 31397.5 88750.0 31462.5 ;
      RECT  89390.0 31537.5 89255.0 31602.5 ;
      RECT  89590.0 31397.5 89455.0 31462.5 ;
      RECT  90095.0 31537.5 89960.0 31602.5 ;
      RECT  90295.0 31397.5 90160.0 31462.5 ;
      RECT  90800.0 31537.5 90665.0 31602.5 ;
      RECT  91000.0 31397.5 90865.0 31462.5 ;
      RECT  91505.0 31537.5 91370.0 31602.5 ;
      RECT  91705.0 31397.5 91570.0 31462.5 ;
      RECT  92210.0 31537.5 92075.0 31602.5 ;
      RECT  92410.0 31397.5 92275.0 31462.5 ;
      RECT  92915.0 31537.5 92780.0 31602.5 ;
      RECT  93115.0 31397.5 92980.0 31462.5 ;
      RECT  93620.0 31537.5 93485.0 31602.5 ;
      RECT  93820.0 31397.5 93685.0 31462.5 ;
      RECT  94325.0 31537.5 94190.0 31602.5 ;
      RECT  94525.0 31397.5 94390.0 31462.5 ;
      RECT  95030.0 31537.5 94895.0 31602.5 ;
      RECT  95230.0 31397.5 95095.0 31462.5 ;
      RECT  95735.0 31537.5 95600.0 31602.5 ;
      RECT  95935.0 31397.5 95800.0 31462.5 ;
      RECT  96440.0 31537.5 96305.0 31602.5 ;
      RECT  96640.0 31397.5 96505.0 31462.5 ;
      RECT  97145.0 31537.5 97010.0 31602.5 ;
      RECT  97345.0 31397.5 97210.0 31462.5 ;
      RECT  97850.0 31537.5 97715.0 31602.5 ;
      RECT  98050.0 31397.5 97915.0 31462.5 ;
      RECT  98555.0 31537.5 98420.0 31602.5 ;
      RECT  98755.0 31397.5 98620.0 31462.5 ;
      RECT  99260.0 31537.5 99125.0 31602.5 ;
      RECT  99460.0 31397.5 99325.0 31462.5 ;
      RECT  99965.0 31537.5 99830.0 31602.5 ;
      RECT  100165.0 31397.5 100030.0 31462.5 ;
      RECT  100670.0 31537.5 100535.0 31602.5 ;
      RECT  100870.0 31397.5 100735.0 31462.5 ;
      RECT  101375.0 31537.5 101240.0 31602.5 ;
      RECT  101575.0 31397.5 101440.0 31462.5 ;
      RECT  102080.0 31537.5 101945.0 31602.5 ;
      RECT  102280.0 31397.5 102145.0 31462.5 ;
      RECT  102785.0 31537.5 102650.0 31602.5 ;
      RECT  102985.0 31397.5 102850.0 31462.5 ;
      RECT  103490.0 31537.5 103355.0 31602.5 ;
      RECT  103690.0 31397.5 103555.0 31462.5 ;
      RECT  104195.0 31537.5 104060.0 31602.5 ;
      RECT  104395.0 31397.5 104260.0 31462.5 ;
      RECT  104900.0 31537.5 104765.0 31602.5 ;
      RECT  105100.0 31397.5 104965.0 31462.5 ;
      RECT  105605.0 31537.5 105470.0 31602.5 ;
      RECT  105805.0 31397.5 105670.0 31462.5 ;
      RECT  106310.0 31537.5 106175.0 31602.5 ;
      RECT  106510.0 31397.5 106375.0 31462.5 ;
      RECT  107015.0 31537.5 106880.0 31602.5 ;
      RECT  107215.0 31397.5 107080.0 31462.5 ;
      RECT  17195.0 32095.0 107435.0 32165.0 ;
      RECT  17195.0 31955.0 107435.0 32025.0 ;
      RECT  17195.0 31815.0 107435.0 31885.0 ;
      RECT  17195.0 31675.0 107435.0 31745.0 ;
      RECT  9102.5 630.0 9167.5 695.0 ;
      RECT  9102.5 1152.5 9167.5 1217.5 ;
      RECT  8865.0 630.0 9135.0 695.0 ;
      RECT  9102.5 662.5 9167.5 1185.0 ;
      RECT  9135.0 1152.5 9380.0 1217.5 ;
      RECT  7995.0 630.0 8635.0 695.0 ;
      RECT  9102.5 2065.0 9167.5 2130.0 ;
      RECT  9102.5 2497.5 9167.5 2562.5 ;
      RECT  8865.0 2065.0 9135.0 2130.0 ;
      RECT  9102.5 2097.5 9167.5 2530.0 ;
      RECT  9135.0 2497.5 9655.0 2562.5 ;
      RECT  8270.0 2065.0 8635.0 2130.0 ;
      RECT  7995.0 2827.5 9930.0 2892.5 ;
      RECT  8270.0 4172.5 10205.0 4237.5 ;
      RECT  9380.0 642.5 10505.0 707.5 ;
      RECT  9655.0 427.5 10762.5 492.5 ;
      RECT  9930.0 2052.5 10505.0 2117.5 ;
      RECT  9655.0 2267.5 10762.5 2332.5 ;
      RECT  9380.0 3332.5 10505.0 3397.5 ;
      RECT  10205.0 3117.5 10762.5 3182.5 ;
      RECT  9930.0 4742.5 10505.0 4807.5 ;
      RECT  10205.0 4957.5 10762.5 5022.5 ;
      RECT  11210.0 642.5 11275.0 707.5 ;
      RECT  11210.0 630.0 11275.0 695.0 ;
      RECT  10992.5 642.5 11242.5 707.5 ;
      RECT  11210.0 662.5 11275.0 675.0 ;
      RECT  11242.5 630.0 11490.0 695.0 ;
      RECT  11210.0 2052.5 11275.0 2117.5 ;
      RECT  11210.0 2065.0 11275.0 2130.0 ;
      RECT  10992.5 2052.5 11242.5 2117.5 ;
      RECT  11210.0 2085.0 11275.0 2097.5 ;
      RECT  11242.5 2065.0 11490.0 2130.0 ;
      RECT  11210.0 3332.5 11275.0 3397.5 ;
      RECT  11210.0 3320.0 11275.0 3385.0 ;
      RECT  10992.5 3332.5 11242.5 3397.5 ;
      RECT  11210.0 3352.5 11275.0 3365.0 ;
      RECT  11242.5 3320.0 11490.0 3385.0 ;
      RECT  11210.0 4742.5 11275.0 4807.5 ;
      RECT  11210.0 4755.0 11275.0 4820.0 ;
      RECT  10992.5 4742.5 11242.5 4807.5 ;
      RECT  11210.0 4775.0 11275.0 4787.5 ;
      RECT  11242.5 4755.0 11490.0 4820.0 ;
      RECT  8937.5 1195.0 9002.5 1380.0 ;
      RECT  8937.5 35.0 9002.5 220.0 ;
      RECT  8577.5 152.5 8642.5 2.5 ;
      RECT  8577.5 1037.5 8642.5 1412.5 ;
      RECT  8767.5 152.5 8832.5 1037.5 ;
      RECT  8577.5 1037.5 8642.5 1172.5 ;
      RECT  8767.5 1037.5 8832.5 1172.5 ;
      RECT  8767.5 1037.5 8832.5 1172.5 ;
      RECT  8577.5 1037.5 8642.5 1172.5 ;
      RECT  8577.5 152.5 8642.5 287.5 ;
      RECT  8767.5 152.5 8832.5 287.5 ;
      RECT  8767.5 152.5 8832.5 287.5 ;
      RECT  8577.5 152.5 8642.5 287.5 ;
      RECT  8937.5 1127.5 9002.5 1262.5 ;
      RECT  8937.5 152.5 9002.5 287.5 ;
      RECT  8635.0 595.0 8700.0 730.0 ;
      RECT  8635.0 595.0 8700.0 730.0 ;
      RECT  8800.0 630.0 8865.0 695.0 ;
      RECT  8510.0 1347.5 9070.0 1412.5 ;
      RECT  8510.0 2.5 9070.0 67.5 ;
      RECT  8937.5 1565.0 9002.5 1380.0 ;
      RECT  8937.5 2725.0 9002.5 2540.0 ;
      RECT  8577.5 2607.5 8642.5 2757.5 ;
      RECT  8577.5 1722.5 8642.5 1347.5 ;
      RECT  8767.5 2607.5 8832.5 1722.5 ;
      RECT  8577.5 1722.5 8642.5 1587.5 ;
      RECT  8767.5 1722.5 8832.5 1587.5 ;
      RECT  8767.5 1722.5 8832.5 1587.5 ;
      RECT  8577.5 1722.5 8642.5 1587.5 ;
      RECT  8577.5 2607.5 8642.5 2472.5 ;
      RECT  8767.5 2607.5 8832.5 2472.5 ;
      RECT  8767.5 2607.5 8832.5 2472.5 ;
      RECT  8577.5 2607.5 8642.5 2472.5 ;
      RECT  8937.5 1632.5 9002.5 1497.5 ;
      RECT  8937.5 2607.5 9002.5 2472.5 ;
      RECT  8635.0 2165.0 8700.0 2030.0 ;
      RECT  8635.0 2165.0 8700.0 2030.0 ;
      RECT  8800.0 2130.0 8865.0 2065.0 ;
      RECT  8510.0 1412.5 9070.0 1347.5 ;
      RECT  8510.0 2757.5 9070.0 2692.5 ;
      RECT  11792.5 1195.0 11857.5 1380.0 ;
      RECT  11792.5 35.0 11857.5 220.0 ;
      RECT  11432.5 152.5 11497.5 2.5 ;
      RECT  11432.5 1037.5 11497.5 1412.5 ;
      RECT  11622.5 152.5 11687.5 1037.5 ;
      RECT  11432.5 1037.5 11497.5 1172.5 ;
      RECT  11622.5 1037.5 11687.5 1172.5 ;
      RECT  11622.5 1037.5 11687.5 1172.5 ;
      RECT  11432.5 1037.5 11497.5 1172.5 ;
      RECT  11432.5 152.5 11497.5 287.5 ;
      RECT  11622.5 152.5 11687.5 287.5 ;
      RECT  11622.5 152.5 11687.5 287.5 ;
      RECT  11432.5 152.5 11497.5 287.5 ;
      RECT  11792.5 1127.5 11857.5 1262.5 ;
      RECT  11792.5 152.5 11857.5 287.5 ;
      RECT  11490.0 595.0 11555.0 730.0 ;
      RECT  11490.0 595.0 11555.0 730.0 ;
      RECT  11655.0 630.0 11720.0 695.0 ;
      RECT  11365.0 1347.5 11925.0 1412.5 ;
      RECT  11365.0 2.5 11925.0 67.5 ;
      RECT  11792.5 1565.0 11857.5 1380.0 ;
      RECT  11792.5 2725.0 11857.5 2540.0 ;
      RECT  11432.5 2607.5 11497.5 2757.5 ;
      RECT  11432.5 1722.5 11497.5 1347.5 ;
      RECT  11622.5 2607.5 11687.5 1722.5 ;
      RECT  11432.5 1722.5 11497.5 1587.5 ;
      RECT  11622.5 1722.5 11687.5 1587.5 ;
      RECT  11622.5 1722.5 11687.5 1587.5 ;
      RECT  11432.5 1722.5 11497.5 1587.5 ;
      RECT  11432.5 2607.5 11497.5 2472.5 ;
      RECT  11622.5 2607.5 11687.5 2472.5 ;
      RECT  11622.5 2607.5 11687.5 2472.5 ;
      RECT  11432.5 2607.5 11497.5 2472.5 ;
      RECT  11792.5 1632.5 11857.5 1497.5 ;
      RECT  11792.5 2607.5 11857.5 2472.5 ;
      RECT  11490.0 2165.0 11555.0 2030.0 ;
      RECT  11490.0 2165.0 11555.0 2030.0 ;
      RECT  11655.0 2130.0 11720.0 2065.0 ;
      RECT  11365.0 1412.5 11925.0 1347.5 ;
      RECT  11365.0 2757.5 11925.0 2692.5 ;
      RECT  11792.5 3885.0 11857.5 4070.0 ;
      RECT  11792.5 2725.0 11857.5 2910.0 ;
      RECT  11432.5 2842.5 11497.5 2692.5 ;
      RECT  11432.5 3727.5 11497.5 4102.5 ;
      RECT  11622.5 2842.5 11687.5 3727.5 ;
      RECT  11432.5 3727.5 11497.5 3862.5 ;
      RECT  11622.5 3727.5 11687.5 3862.5 ;
      RECT  11622.5 3727.5 11687.5 3862.5 ;
      RECT  11432.5 3727.5 11497.5 3862.5 ;
      RECT  11432.5 2842.5 11497.5 2977.5 ;
      RECT  11622.5 2842.5 11687.5 2977.5 ;
      RECT  11622.5 2842.5 11687.5 2977.5 ;
      RECT  11432.5 2842.5 11497.5 2977.5 ;
      RECT  11792.5 3817.5 11857.5 3952.5 ;
      RECT  11792.5 2842.5 11857.5 2977.5 ;
      RECT  11490.0 3285.0 11555.0 3420.0 ;
      RECT  11490.0 3285.0 11555.0 3420.0 ;
      RECT  11655.0 3320.0 11720.0 3385.0 ;
      RECT  11365.0 4037.5 11925.0 4102.5 ;
      RECT  11365.0 2692.5 11925.0 2757.5 ;
      RECT  11792.5 4255.0 11857.5 4070.0 ;
      RECT  11792.5 5415.0 11857.5 5230.0 ;
      RECT  11432.5 5297.5 11497.5 5447.5 ;
      RECT  11432.5 4412.5 11497.5 4037.5 ;
      RECT  11622.5 5297.5 11687.5 4412.5 ;
      RECT  11432.5 4412.5 11497.5 4277.5 ;
      RECT  11622.5 4412.5 11687.5 4277.5 ;
      RECT  11622.5 4412.5 11687.5 4277.5 ;
      RECT  11432.5 4412.5 11497.5 4277.5 ;
      RECT  11432.5 5297.5 11497.5 5162.5 ;
      RECT  11622.5 5297.5 11687.5 5162.5 ;
      RECT  11622.5 5297.5 11687.5 5162.5 ;
      RECT  11432.5 5297.5 11497.5 5162.5 ;
      RECT  11792.5 4322.5 11857.5 4187.5 ;
      RECT  11792.5 5297.5 11857.5 5162.5 ;
      RECT  11490.0 4855.0 11555.0 4720.0 ;
      RECT  11490.0 4855.0 11555.0 4720.0 ;
      RECT  11655.0 4820.0 11720.0 4755.0 ;
      RECT  11365.0 4102.5 11925.0 4037.5 ;
      RECT  11365.0 5447.5 11925.0 5382.5 ;
      RECT  10512.5 197.5 10577.5 2.5 ;
      RECT  10512.5 1037.5 10577.5 1412.5 ;
      RECT  10892.5 1037.5 10957.5 1412.5 ;
      RECT  11062.5 1195.0 11127.5 1380.0 ;
      RECT  11062.5 35.0 11127.5 220.0 ;
      RECT  10512.5 1037.5 10577.5 1172.5 ;
      RECT  10702.5 1037.5 10767.5 1172.5 ;
      RECT  10702.5 1037.5 10767.5 1172.5 ;
      RECT  10512.5 1037.5 10577.5 1172.5 ;
      RECT  10702.5 1037.5 10767.5 1172.5 ;
      RECT  10892.5 1037.5 10957.5 1172.5 ;
      RECT  10892.5 1037.5 10957.5 1172.5 ;
      RECT  10702.5 1037.5 10767.5 1172.5 ;
      RECT  10512.5 197.5 10577.5 332.5 ;
      RECT  10702.5 197.5 10767.5 332.5 ;
      RECT  10702.5 197.5 10767.5 332.5 ;
      RECT  10512.5 197.5 10577.5 332.5 ;
      RECT  10702.5 197.5 10767.5 332.5 ;
      RECT  10892.5 197.5 10957.5 332.5 ;
      RECT  10892.5 197.5 10957.5 332.5 ;
      RECT  10702.5 197.5 10767.5 332.5 ;
      RECT  11062.5 1127.5 11127.5 1262.5 ;
      RECT  11062.5 152.5 11127.5 287.5 ;
      RECT  10897.5 427.5 10762.5 492.5 ;
      RECT  10640.0 642.5 10505.0 707.5 ;
      RECT  10702.5 1037.5 10767.5 1172.5 ;
      RECT  10892.5 197.5 10957.5 332.5 ;
      RECT  10992.5 642.5 10857.5 707.5 ;
      RECT  10505.0 642.5 10640.0 707.5 ;
      RECT  10762.5 427.5 10897.5 492.5 ;
      RECT  10857.5 642.5 10992.5 707.5 ;
      RECT  10445.0 1347.5 11365.0 1412.5 ;
      RECT  10445.0 2.5 11365.0 67.5 ;
      RECT  10512.5 2562.5 10577.5 2757.5 ;
      RECT  10512.5 1722.5 10577.5 1347.5 ;
      RECT  10892.5 1722.5 10957.5 1347.5 ;
      RECT  11062.5 1565.0 11127.5 1380.0 ;
      RECT  11062.5 2725.0 11127.5 2540.0 ;
      RECT  10512.5 1722.5 10577.5 1587.5 ;
      RECT  10702.5 1722.5 10767.5 1587.5 ;
      RECT  10702.5 1722.5 10767.5 1587.5 ;
      RECT  10512.5 1722.5 10577.5 1587.5 ;
      RECT  10702.5 1722.5 10767.5 1587.5 ;
      RECT  10892.5 1722.5 10957.5 1587.5 ;
      RECT  10892.5 1722.5 10957.5 1587.5 ;
      RECT  10702.5 1722.5 10767.5 1587.5 ;
      RECT  10512.5 2562.5 10577.5 2427.5 ;
      RECT  10702.5 2562.5 10767.5 2427.5 ;
      RECT  10702.5 2562.5 10767.5 2427.5 ;
      RECT  10512.5 2562.5 10577.5 2427.5 ;
      RECT  10702.5 2562.5 10767.5 2427.5 ;
      RECT  10892.5 2562.5 10957.5 2427.5 ;
      RECT  10892.5 2562.5 10957.5 2427.5 ;
      RECT  10702.5 2562.5 10767.5 2427.5 ;
      RECT  11062.5 1632.5 11127.5 1497.5 ;
      RECT  11062.5 2607.5 11127.5 2472.5 ;
      RECT  10897.5 2332.5 10762.5 2267.5 ;
      RECT  10640.0 2117.5 10505.0 2052.5 ;
      RECT  10702.5 1722.5 10767.5 1587.5 ;
      RECT  10892.5 2562.5 10957.5 2427.5 ;
      RECT  10992.5 2117.5 10857.5 2052.5 ;
      RECT  10505.0 2117.5 10640.0 2052.5 ;
      RECT  10762.5 2332.5 10897.5 2267.5 ;
      RECT  10857.5 2117.5 10992.5 2052.5 ;
      RECT  10445.0 1412.5 11365.0 1347.5 ;
      RECT  10445.0 2757.5 11365.0 2692.5 ;
      RECT  10512.5 2887.5 10577.5 2692.5 ;
      RECT  10512.5 3727.5 10577.5 4102.5 ;
      RECT  10892.5 3727.5 10957.5 4102.5 ;
      RECT  11062.5 3885.0 11127.5 4070.0 ;
      RECT  11062.5 2725.0 11127.5 2910.0 ;
      RECT  10512.5 3727.5 10577.5 3862.5 ;
      RECT  10702.5 3727.5 10767.5 3862.5 ;
      RECT  10702.5 3727.5 10767.5 3862.5 ;
      RECT  10512.5 3727.5 10577.5 3862.5 ;
      RECT  10702.5 3727.5 10767.5 3862.5 ;
      RECT  10892.5 3727.5 10957.5 3862.5 ;
      RECT  10892.5 3727.5 10957.5 3862.5 ;
      RECT  10702.5 3727.5 10767.5 3862.5 ;
      RECT  10512.5 2887.5 10577.5 3022.5 ;
      RECT  10702.5 2887.5 10767.5 3022.5 ;
      RECT  10702.5 2887.5 10767.5 3022.5 ;
      RECT  10512.5 2887.5 10577.5 3022.5 ;
      RECT  10702.5 2887.5 10767.5 3022.5 ;
      RECT  10892.5 2887.5 10957.5 3022.5 ;
      RECT  10892.5 2887.5 10957.5 3022.5 ;
      RECT  10702.5 2887.5 10767.5 3022.5 ;
      RECT  11062.5 3817.5 11127.5 3952.5 ;
      RECT  11062.5 2842.5 11127.5 2977.5 ;
      RECT  10897.5 3117.5 10762.5 3182.5 ;
      RECT  10640.0 3332.5 10505.0 3397.5 ;
      RECT  10702.5 3727.5 10767.5 3862.5 ;
      RECT  10892.5 2887.5 10957.5 3022.5 ;
      RECT  10992.5 3332.5 10857.5 3397.5 ;
      RECT  10505.0 3332.5 10640.0 3397.5 ;
      RECT  10762.5 3117.5 10897.5 3182.5 ;
      RECT  10857.5 3332.5 10992.5 3397.5 ;
      RECT  10445.0 4037.5 11365.0 4102.5 ;
      RECT  10445.0 2692.5 11365.0 2757.5 ;
      RECT  10512.5 5252.5 10577.5 5447.5 ;
      RECT  10512.5 4412.5 10577.5 4037.5 ;
      RECT  10892.5 4412.5 10957.5 4037.5 ;
      RECT  11062.5 4255.0 11127.5 4070.0 ;
      RECT  11062.5 5415.0 11127.5 5230.0 ;
      RECT  10512.5 4412.5 10577.5 4277.5 ;
      RECT  10702.5 4412.5 10767.5 4277.5 ;
      RECT  10702.5 4412.5 10767.5 4277.5 ;
      RECT  10512.5 4412.5 10577.5 4277.5 ;
      RECT  10702.5 4412.5 10767.5 4277.5 ;
      RECT  10892.5 4412.5 10957.5 4277.5 ;
      RECT  10892.5 4412.5 10957.5 4277.5 ;
      RECT  10702.5 4412.5 10767.5 4277.5 ;
      RECT  10512.5 5252.5 10577.5 5117.5 ;
      RECT  10702.5 5252.5 10767.5 5117.5 ;
      RECT  10702.5 5252.5 10767.5 5117.5 ;
      RECT  10512.5 5252.5 10577.5 5117.5 ;
      RECT  10702.5 5252.5 10767.5 5117.5 ;
      RECT  10892.5 5252.5 10957.5 5117.5 ;
      RECT  10892.5 5252.5 10957.5 5117.5 ;
      RECT  10702.5 5252.5 10767.5 5117.5 ;
      RECT  11062.5 4322.5 11127.5 4187.5 ;
      RECT  11062.5 5297.5 11127.5 5162.5 ;
      RECT  10897.5 5022.5 10762.5 4957.5 ;
      RECT  10640.0 4807.5 10505.0 4742.5 ;
      RECT  10702.5 4412.5 10767.5 4277.5 ;
      RECT  10892.5 5252.5 10957.5 5117.5 ;
      RECT  10992.5 4807.5 10857.5 4742.5 ;
      RECT  10505.0 4807.5 10640.0 4742.5 ;
      RECT  10762.5 5022.5 10897.5 4957.5 ;
      RECT  10857.5 4807.5 10992.5 4742.5 ;
      RECT  10445.0 4102.5 11365.0 4037.5 ;
      RECT  10445.0 5447.5 11365.0 5382.5 ;
      RECT  9447.5 1152.5 9312.5 1217.5 ;
      RECT  8062.5 630.0 7927.5 695.0 ;
      RECT  9722.5 2497.5 9587.5 2562.5 ;
      RECT  8337.5 2065.0 8202.5 2130.0 ;
      RECT  8062.5 2827.5 7927.5 2892.5 ;
      RECT  9997.5 2827.5 9862.5 2892.5 ;
      RECT  8337.5 4172.5 8202.5 4237.5 ;
      RECT  10272.5 4172.5 10137.5 4237.5 ;
      RECT  9447.5 642.5 9312.5 707.5 ;
      RECT  9722.5 427.5 9587.5 492.5 ;
      RECT  9997.5 2052.5 9862.5 2117.5 ;
      RECT  9722.5 2267.5 9587.5 2332.5 ;
      RECT  9447.5 3332.5 9312.5 3397.5 ;
      RECT  10272.5 3117.5 10137.5 3182.5 ;
      RECT  9997.5 4742.5 9862.5 4807.5 ;
      RECT  10272.5 4957.5 10137.5 5022.5 ;
      RECT  11720.0 630.0 11925.0 695.0 ;
      RECT  11720.0 2065.0 11925.0 2130.0 ;
      RECT  11720.0 3320.0 11925.0 3385.0 ;
      RECT  11720.0 4755.0 11925.0 4820.0 ;
      RECT  7960.0 1347.5 11925.0 1412.5 ;
      RECT  7960.0 4037.5 11925.0 4102.5 ;
      RECT  7960.0 2.5 11925.0 67.5 ;
      RECT  7960.0 2692.5 11925.0 2757.5 ;
      RECT  7960.0 5382.5 11925.0 5447.5 ;
      RECT  17195.0 26370.0 17900.0 31255.0 ;
      RECT  20015.0 26370.0 20720.0 31255.0 ;
      RECT  22835.0 26370.0 23540.0 31255.0 ;
      RECT  25655.0 26370.0 26360.0 31255.0 ;
      RECT  28475.0 26370.0 29180.0 31255.0 ;
      RECT  31295.0 26370.0 32000.0 31255.0 ;
      RECT  34115.0 26370.0 34820.0 31255.0 ;
      RECT  36935.0 26370.0 37640.0 31255.0 ;
      RECT  39755.0 26370.0 40460.0 31255.0 ;
      RECT  42575.0 26370.0 43280.0 31255.0 ;
      RECT  45395.0 26370.0 46100.0 31255.0 ;
      RECT  48215.0 26370.0 48920.0 31255.0 ;
      RECT  51035.0 26370.0 51740.0 31255.0 ;
      RECT  53855.0 26370.0 54560.0 31255.0 ;
      RECT  56675.0 26370.0 57380.0 31255.0 ;
      RECT  59495.0 26370.0 60200.0 31255.0 ;
      RECT  62315.0 26370.0 63020.0 31255.0 ;
      RECT  65135.0 26370.0 65840.0 31255.0 ;
      RECT  67955.0 26370.0 68660.0 31255.0 ;
      RECT  70775.0 26370.0 71480.0 31255.0 ;
      RECT  73595.0 26370.0 74300.0 31255.0 ;
      RECT  76415.0 26370.0 77120.0 31255.0 ;
      RECT  79235.0 26370.0 79940.0 31255.0 ;
      RECT  82055.0 26370.0 82760.0 31255.0 ;
      RECT  84875.0 26370.0 85580.0 31255.0 ;
      RECT  87695.0 26370.0 88400.0 31255.0 ;
      RECT  90515.0 26370.0 91220.0 31255.0 ;
      RECT  93335.0 26370.0 94040.0 31255.0 ;
      RECT  96155.0 26370.0 96860.0 31255.0 ;
      RECT  98975.0 26370.0 99680.0 31255.0 ;
      RECT  101795.0 26370.0 102500.0 31255.0 ;
      RECT  104615.0 26370.0 105320.0 31255.0 ;
      RECT  17195.0 26487.5 107435.0 26552.5 ;
      RECT  17195.0 31060.0 107435.0 31125.0 ;
      RECT  17195.0 26617.5 107435.0 26682.5 ;
      RECT  17195.0 22195.0 17900.0 26370.0 ;
      RECT  20015.0 22195.0 20720.0 26370.0 ;
      RECT  22835.0 22195.0 23540.0 26370.0 ;
      RECT  25655.0 22195.0 26360.0 26370.0 ;
      RECT  28475.0 22195.0 29180.0 26370.0 ;
      RECT  31295.0 22195.0 32000.0 26370.0 ;
      RECT  34115.0 22195.0 34820.0 26370.0 ;
      RECT  36935.0 22195.0 37640.0 26370.0 ;
      RECT  39755.0 22195.0 40460.0 26370.0 ;
      RECT  42575.0 22195.0 43280.0 26370.0 ;
      RECT  45395.0 22195.0 46100.0 26370.0 ;
      RECT  48215.0 22195.0 48920.0 26370.0 ;
      RECT  51035.0 22195.0 51740.0 26370.0 ;
      RECT  53855.0 22195.0 54560.0 26370.0 ;
      RECT  56675.0 22195.0 57380.0 26370.0 ;
      RECT  59495.0 22195.0 60200.0 26370.0 ;
      RECT  62315.0 22195.0 63020.0 26370.0 ;
      RECT  65135.0 22195.0 65840.0 26370.0 ;
      RECT  67955.0 22195.0 68660.0 26370.0 ;
      RECT  70775.0 22195.0 71480.0 26370.0 ;
      RECT  73595.0 22195.0 74300.0 26370.0 ;
      RECT  76415.0 22195.0 77120.0 26370.0 ;
      RECT  79235.0 22195.0 79940.0 26370.0 ;
      RECT  82055.0 22195.0 82760.0 26370.0 ;
      RECT  84875.0 22195.0 85580.0 26370.0 ;
      RECT  87695.0 22195.0 88400.0 26370.0 ;
      RECT  90515.0 22195.0 91220.0 26370.0 ;
      RECT  93335.0 22195.0 94040.0 26370.0 ;
      RECT  96155.0 22195.0 96860.0 26370.0 ;
      RECT  98975.0 22195.0 99680.0 26370.0 ;
      RECT  101795.0 22195.0 102500.0 26370.0 ;
      RECT  104615.0 22195.0 105320.0 26370.0 ;
      RECT  17195.0 22462.5 107435.0 22527.5 ;
      RECT  17195.0 22592.5 107435.0 22657.5 ;
      RECT  17195.0 23395.0 107435.0 23460.0 ;
      RECT  17195.0 15755.0 17900.0 22195.0 ;
      RECT  20015.0 15755.0 20720.0 22195.0 ;
      RECT  22835.0 15755.0 23540.0 22195.0 ;
      RECT  25655.0 15755.0 26360.0 22195.0 ;
      RECT  28475.0 15755.0 29180.0 22195.0 ;
      RECT  31295.0 15755.0 32000.0 22195.0 ;
      RECT  34115.0 15755.0 34820.0 22195.0 ;
      RECT  36935.0 15755.0 37640.0 22195.0 ;
      RECT  39755.0 15755.0 40460.0 22195.0 ;
      RECT  42575.0 15755.0 43280.0 22195.0 ;
      RECT  45395.0 15755.0 46100.0 22195.0 ;
      RECT  48215.0 15755.0 48920.0 22195.0 ;
      RECT  51035.0 15755.0 51740.0 22195.0 ;
      RECT  53855.0 15755.0 54560.0 22195.0 ;
      RECT  56675.0 15755.0 57380.0 22195.0 ;
      RECT  59495.0 15755.0 60200.0 22195.0 ;
      RECT  62315.0 15755.0 63020.0 22195.0 ;
      RECT  65135.0 15755.0 65840.0 22195.0 ;
      RECT  67955.0 15755.0 68660.0 22195.0 ;
      RECT  70775.0 15755.0 71480.0 22195.0 ;
      RECT  73595.0 15755.0 74300.0 22195.0 ;
      RECT  76415.0 15755.0 77120.0 22195.0 ;
      RECT  79235.0 15755.0 79940.0 22195.0 ;
      RECT  82055.0 15755.0 82760.0 22195.0 ;
      RECT  84875.0 15755.0 85580.0 22195.0 ;
      RECT  87695.0 15755.0 88400.0 22195.0 ;
      RECT  90515.0 15755.0 91220.0 22195.0 ;
      RECT  93335.0 15755.0 94040.0 22195.0 ;
      RECT  96155.0 15755.0 96860.0 22195.0 ;
      RECT  98975.0 15755.0 99680.0 22195.0 ;
      RECT  101795.0 15755.0 102500.0 22195.0 ;
      RECT  104615.0 15755.0 105320.0 22195.0 ;
      RECT  17195.0 15960.0 107435.0 16025.0 ;
      RECT  17195.0 18965.0 107435.0 19030.0 ;
      RECT  17195.0 21925.0 107435.0 21990.0 ;
      RECT  17195.0 16975.0 107435.0 17040.0 ;
      RECT  17195.0 19935.0 107435.0 20000.0 ;
      RECT  17195.0 16120.0 107435.0 16185.0 ;
      RECT  17195.0 15755.0 17900.0 12780.0 ;
      RECT  20015.0 15755.0 20720.0 12780.0 ;
      RECT  22835.0 15755.0 23540.0 12780.0 ;
      RECT  25655.0 15755.0 26360.0 12780.0 ;
      RECT  28475.0 15755.0 29180.0 12780.0 ;
      RECT  31295.0 15755.0 32000.0 12780.0 ;
      RECT  34115.0 15755.0 34820.0 12780.0 ;
      RECT  36935.0 15755.0 37640.0 12780.0 ;
      RECT  39755.0 15755.0 40460.0 12780.0 ;
      RECT  42575.0 15755.0 43280.0 12780.0 ;
      RECT  45395.0 15755.0 46100.0 12780.0 ;
      RECT  48215.0 15755.0 48920.0 12780.0 ;
      RECT  51035.0 15755.0 51740.0 12780.0 ;
      RECT  53855.0 15755.0 54560.0 12780.0 ;
      RECT  56675.0 15755.0 57380.0 12780.0 ;
      RECT  59495.0 15755.0 60200.0 12780.0 ;
      RECT  62315.0 15755.0 63020.0 12780.0 ;
      RECT  65135.0 15755.0 65840.0 12780.0 ;
      RECT  67955.0 15755.0 68660.0 12780.0 ;
      RECT  70775.0 15755.0 71480.0 12780.0 ;
      RECT  73595.0 15755.0 74300.0 12780.0 ;
      RECT  76415.0 15755.0 77120.0 12780.0 ;
      RECT  79235.0 15755.0 79940.0 12780.0 ;
      RECT  82055.0 15755.0 82760.0 12780.0 ;
      RECT  84875.0 15755.0 85580.0 12780.0 ;
      RECT  87695.0 15755.0 88400.0 12780.0 ;
      RECT  90515.0 15755.0 91220.0 12780.0 ;
      RECT  93335.0 15755.0 94040.0 12780.0 ;
      RECT  96155.0 15755.0 96860.0 12780.0 ;
      RECT  98975.0 15755.0 99680.0 12780.0 ;
      RECT  101795.0 15755.0 102500.0 12780.0 ;
      RECT  104615.0 15755.0 105320.0 12780.0 ;
      RECT  17195.0 15387.5 105320.0 15322.5 ;
      RECT  17195.0 13840.0 105320.0 13775.0 ;
      RECT  17195.0 13970.0 105320.0 13905.0 ;
      RECT  17195.0 15257.5 105320.0 15192.5 ;
      RECT  8342.5 34755.0 8407.5 34820.0 ;
      RECT  8342.5 34695.0 8407.5 34760.0 ;
      RECT  8157.5 34755.0 8375.0 34820.0 ;
      RECT  8342.5 34727.5 8407.5 34787.5 ;
      RECT  8375.0 34695.0 8590.0 34760.0 ;
      RECT  8342.5 36070.0 8407.5 36135.0 ;
      RECT  8342.5 36130.0 8407.5 36195.0 ;
      RECT  8157.5 36070.0 8375.0 36135.0 ;
      RECT  8342.5 36102.5 8407.5 36162.5 ;
      RECT  8375.0 36130.0 8590.0 36195.0 ;
      RECT  8342.5 37445.0 8407.5 37510.0 ;
      RECT  8342.5 37385.0 8407.5 37450.0 ;
      RECT  8157.5 37445.0 8375.0 37510.0 ;
      RECT  8342.5 37417.5 8407.5 37477.5 ;
      RECT  8375.0 37385.0 8590.0 37450.0 ;
      RECT  8342.5 38760.0 8407.5 38825.0 ;
      RECT  8342.5 38820.0 8407.5 38885.0 ;
      RECT  8157.5 38760.0 8375.0 38825.0 ;
      RECT  8342.5 38792.5 8407.5 38852.5 ;
      RECT  8375.0 38820.0 8590.0 38885.0 ;
      RECT  8342.5 40135.0 8407.5 40200.0 ;
      RECT  8342.5 40075.0 8407.5 40140.0 ;
      RECT  8157.5 40135.0 8375.0 40200.0 ;
      RECT  8342.5 40107.5 8407.5 40167.5 ;
      RECT  8375.0 40075.0 8590.0 40140.0 ;
      RECT  8342.5 41450.0 8407.5 41515.0 ;
      RECT  8342.5 41510.0 8407.5 41575.0 ;
      RECT  8157.5 41450.0 8375.0 41515.0 ;
      RECT  8342.5 41482.5 8407.5 41542.5 ;
      RECT  8375.0 41510.0 8590.0 41575.0 ;
      RECT  8342.5 42825.0 8407.5 42890.0 ;
      RECT  8342.5 42765.0 8407.5 42830.0 ;
      RECT  8157.5 42825.0 8375.0 42890.0 ;
      RECT  8342.5 42797.5 8407.5 42857.5 ;
      RECT  8375.0 42765.0 8590.0 42830.0 ;
      RECT  8342.5 44140.0 8407.5 44205.0 ;
      RECT  8342.5 44200.0 8407.5 44265.0 ;
      RECT  8157.5 44140.0 8375.0 44205.0 ;
      RECT  8342.5 44172.5 8407.5 44232.5 ;
      RECT  8375.0 44200.0 8590.0 44265.0 ;
      RECT  8342.5 45515.0 8407.5 45580.0 ;
      RECT  8342.5 45455.0 8407.5 45520.0 ;
      RECT  8157.5 45515.0 8375.0 45580.0 ;
      RECT  8342.5 45487.5 8407.5 45547.5 ;
      RECT  8375.0 45455.0 8590.0 45520.0 ;
      RECT  8342.5 46830.0 8407.5 46895.0 ;
      RECT  8342.5 46890.0 8407.5 46955.0 ;
      RECT  8157.5 46830.0 8375.0 46895.0 ;
      RECT  8342.5 46862.5 8407.5 46922.5 ;
      RECT  8375.0 46890.0 8590.0 46955.0 ;
      RECT  8342.5 48205.0 8407.5 48270.0 ;
      RECT  8342.5 48145.0 8407.5 48210.0 ;
      RECT  8157.5 48205.0 8375.0 48270.0 ;
      RECT  8342.5 48177.5 8407.5 48237.5 ;
      RECT  8375.0 48145.0 8590.0 48210.0 ;
      RECT  8342.5 49520.0 8407.5 49585.0 ;
      RECT  8342.5 49580.0 8407.5 49645.0 ;
      RECT  8157.5 49520.0 8375.0 49585.0 ;
      RECT  8342.5 49552.5 8407.5 49612.5 ;
      RECT  8375.0 49580.0 8590.0 49645.0 ;
      RECT  8342.5 50895.0 8407.5 50960.0 ;
      RECT  8342.5 50835.0 8407.5 50900.0 ;
      RECT  8157.5 50895.0 8375.0 50960.0 ;
      RECT  8342.5 50867.5 8407.5 50927.5 ;
      RECT  8375.0 50835.0 8590.0 50900.0 ;
      RECT  8342.5 52210.0 8407.5 52275.0 ;
      RECT  8342.5 52270.0 8407.5 52335.0 ;
      RECT  8157.5 52210.0 8375.0 52275.0 ;
      RECT  8342.5 52242.5 8407.5 52302.5 ;
      RECT  8375.0 52270.0 8590.0 52335.0 ;
      RECT  8342.5 53585.0 8407.5 53650.0 ;
      RECT  8342.5 53525.0 8407.5 53590.0 ;
      RECT  8157.5 53585.0 8375.0 53650.0 ;
      RECT  8342.5 53557.5 8407.5 53617.5 ;
      RECT  8375.0 53525.0 8590.0 53590.0 ;
      RECT  8342.5 54900.0 8407.5 54965.0 ;
      RECT  8342.5 54960.0 8407.5 55025.0 ;
      RECT  8157.5 54900.0 8375.0 54965.0 ;
      RECT  8342.5 54932.5 8407.5 54992.5 ;
      RECT  8375.0 54960.0 8590.0 55025.0 ;
      RECT  8342.5 56275.0 8407.5 56340.0 ;
      RECT  8342.5 56215.0 8407.5 56280.0 ;
      RECT  8157.5 56275.0 8375.0 56340.0 ;
      RECT  8342.5 56247.5 8407.5 56307.5 ;
      RECT  8375.0 56215.0 8590.0 56280.0 ;
      RECT  8342.5 57590.0 8407.5 57655.0 ;
      RECT  8342.5 57650.0 8407.5 57715.0 ;
      RECT  8157.5 57590.0 8375.0 57655.0 ;
      RECT  8342.5 57622.5 8407.5 57682.5 ;
      RECT  8375.0 57650.0 8590.0 57715.0 ;
      RECT  8342.5 58965.0 8407.5 59030.0 ;
      RECT  8342.5 58905.0 8407.5 58970.0 ;
      RECT  8157.5 58965.0 8375.0 59030.0 ;
      RECT  8342.5 58937.5 8407.5 58997.5 ;
      RECT  8375.0 58905.0 8590.0 58970.0 ;
      RECT  8342.5 60280.0 8407.5 60345.0 ;
      RECT  8342.5 60340.0 8407.5 60405.0 ;
      RECT  8157.5 60280.0 8375.0 60345.0 ;
      RECT  8342.5 60312.5 8407.5 60372.5 ;
      RECT  8375.0 60340.0 8590.0 60405.0 ;
      RECT  8342.5 61655.0 8407.5 61720.0 ;
      RECT  8342.5 61595.0 8407.5 61660.0 ;
      RECT  8157.5 61655.0 8375.0 61720.0 ;
      RECT  8342.5 61627.5 8407.5 61687.5 ;
      RECT  8375.0 61595.0 8590.0 61660.0 ;
      RECT  8342.5 62970.0 8407.5 63035.0 ;
      RECT  8342.5 63030.0 8407.5 63095.0 ;
      RECT  8157.5 62970.0 8375.0 63035.0 ;
      RECT  8342.5 63002.5 8407.5 63062.5 ;
      RECT  8375.0 63030.0 8590.0 63095.0 ;
      RECT  8342.5 64345.0 8407.5 64410.0 ;
      RECT  8342.5 64285.0 8407.5 64350.0 ;
      RECT  8157.5 64345.0 8375.0 64410.0 ;
      RECT  8342.5 64317.5 8407.5 64377.5 ;
      RECT  8375.0 64285.0 8590.0 64350.0 ;
      RECT  8342.5 65660.0 8407.5 65725.0 ;
      RECT  8342.5 65720.0 8407.5 65785.0 ;
      RECT  8157.5 65660.0 8375.0 65725.0 ;
      RECT  8342.5 65692.5 8407.5 65752.5 ;
      RECT  8375.0 65720.0 8590.0 65785.0 ;
      RECT  8342.5 67035.0 8407.5 67100.0 ;
      RECT  8342.5 66975.0 8407.5 67040.0 ;
      RECT  8157.5 67035.0 8375.0 67100.0 ;
      RECT  8342.5 67007.5 8407.5 67067.5 ;
      RECT  8375.0 66975.0 8590.0 67040.0 ;
      RECT  8342.5 68350.0 8407.5 68415.0 ;
      RECT  8342.5 68410.0 8407.5 68475.0 ;
      RECT  8157.5 68350.0 8375.0 68415.0 ;
      RECT  8342.5 68382.5 8407.5 68442.5 ;
      RECT  8375.0 68410.0 8590.0 68475.0 ;
      RECT  8342.5 69725.0 8407.5 69790.0 ;
      RECT  8342.5 69665.0 8407.5 69730.0 ;
      RECT  8157.5 69725.0 8375.0 69790.0 ;
      RECT  8342.5 69697.5 8407.5 69757.5 ;
      RECT  8375.0 69665.0 8590.0 69730.0 ;
      RECT  8342.5 71040.0 8407.5 71105.0 ;
      RECT  8342.5 71100.0 8407.5 71165.0 ;
      RECT  8157.5 71040.0 8375.0 71105.0 ;
      RECT  8342.5 71072.5 8407.5 71132.5 ;
      RECT  8375.0 71100.0 8590.0 71165.0 ;
      RECT  8342.5 72415.0 8407.5 72480.0 ;
      RECT  8342.5 72355.0 8407.5 72420.0 ;
      RECT  8157.5 72415.0 8375.0 72480.0 ;
      RECT  8342.5 72387.5 8407.5 72447.5 ;
      RECT  8375.0 72355.0 8590.0 72420.0 ;
      RECT  8342.5 73730.0 8407.5 73795.0 ;
      RECT  8342.5 73790.0 8407.5 73855.0 ;
      RECT  8157.5 73730.0 8375.0 73795.0 ;
      RECT  8342.5 73762.5 8407.5 73822.5 ;
      RECT  8375.0 73790.0 8590.0 73855.0 ;
      RECT  8342.5 75105.0 8407.5 75170.0 ;
      RECT  8342.5 75045.0 8407.5 75110.0 ;
      RECT  8157.5 75105.0 8375.0 75170.0 ;
      RECT  8342.5 75077.5 8407.5 75137.5 ;
      RECT  8375.0 75045.0 8590.0 75110.0 ;
      RECT  8342.5 76420.0 8407.5 76485.0 ;
      RECT  8342.5 76480.0 8407.5 76545.0 ;
      RECT  8157.5 76420.0 8375.0 76485.0 ;
      RECT  8342.5 76452.5 8407.5 76512.5 ;
      RECT  8375.0 76480.0 8590.0 76545.0 ;
      RECT  8342.5 77795.0 8407.5 77860.0 ;
      RECT  8342.5 77735.0 8407.5 77800.0 ;
      RECT  8157.5 77795.0 8375.0 77860.0 ;
      RECT  8342.5 77767.5 8407.5 77827.5 ;
      RECT  8375.0 77735.0 8590.0 77800.0 ;
      RECT  8342.5 79110.0 8407.5 79175.0 ;
      RECT  8342.5 79170.0 8407.5 79235.0 ;
      RECT  8157.5 79110.0 8375.0 79175.0 ;
      RECT  8342.5 79142.5 8407.5 79202.5 ;
      RECT  8375.0 79170.0 8590.0 79235.0 ;
      RECT  8342.5 80485.0 8407.5 80550.0 ;
      RECT  8342.5 80425.0 8407.5 80490.0 ;
      RECT  8157.5 80485.0 8375.0 80550.0 ;
      RECT  8342.5 80457.5 8407.5 80517.5 ;
      RECT  8375.0 80425.0 8590.0 80490.0 ;
      RECT  8342.5 81800.0 8407.5 81865.0 ;
      RECT  8342.5 81860.0 8407.5 81925.0 ;
      RECT  8157.5 81800.0 8375.0 81865.0 ;
      RECT  8342.5 81832.5 8407.5 81892.5 ;
      RECT  8375.0 81860.0 8590.0 81925.0 ;
      RECT  8342.5 83175.0 8407.5 83240.0 ;
      RECT  8342.5 83115.0 8407.5 83180.0 ;
      RECT  8157.5 83175.0 8375.0 83240.0 ;
      RECT  8342.5 83147.5 8407.5 83207.5 ;
      RECT  8375.0 83115.0 8590.0 83180.0 ;
      RECT  8342.5 84490.0 8407.5 84555.0 ;
      RECT  8342.5 84550.0 8407.5 84615.0 ;
      RECT  8157.5 84490.0 8375.0 84555.0 ;
      RECT  8342.5 84522.5 8407.5 84582.5 ;
      RECT  8375.0 84550.0 8590.0 84615.0 ;
      RECT  8342.5 85865.0 8407.5 85930.0 ;
      RECT  8342.5 85805.0 8407.5 85870.0 ;
      RECT  8157.5 85865.0 8375.0 85930.0 ;
      RECT  8342.5 85837.5 8407.5 85897.5 ;
      RECT  8375.0 85805.0 8590.0 85870.0 ;
      RECT  8342.5 87180.0 8407.5 87245.0 ;
      RECT  8342.5 87240.0 8407.5 87305.0 ;
      RECT  8157.5 87180.0 8375.0 87245.0 ;
      RECT  8342.5 87212.5 8407.5 87272.5 ;
      RECT  8375.0 87240.0 8590.0 87305.0 ;
      RECT  8342.5 88555.0 8407.5 88620.0 ;
      RECT  8342.5 88495.0 8407.5 88560.0 ;
      RECT  8157.5 88555.0 8375.0 88620.0 ;
      RECT  8342.5 88527.5 8407.5 88587.5 ;
      RECT  8375.0 88495.0 8590.0 88560.0 ;
      RECT  8342.5 89870.0 8407.5 89935.0 ;
      RECT  8342.5 89930.0 8407.5 89995.0 ;
      RECT  8157.5 89870.0 8375.0 89935.0 ;
      RECT  8342.5 89902.5 8407.5 89962.5 ;
      RECT  8375.0 89930.0 8590.0 89995.0 ;
      RECT  8342.5 91245.0 8407.5 91310.0 ;
      RECT  8342.5 91185.0 8407.5 91250.0 ;
      RECT  8157.5 91245.0 8375.0 91310.0 ;
      RECT  8342.5 91217.5 8407.5 91277.5 ;
      RECT  8375.0 91185.0 8590.0 91250.0 ;
      RECT  8342.5 92560.0 8407.5 92625.0 ;
      RECT  8342.5 92620.0 8407.5 92685.0 ;
      RECT  8157.5 92560.0 8375.0 92625.0 ;
      RECT  8342.5 92592.5 8407.5 92652.5 ;
      RECT  8375.0 92620.0 8590.0 92685.0 ;
      RECT  8342.5 93935.0 8407.5 94000.0 ;
      RECT  8342.5 93875.0 8407.5 93940.0 ;
      RECT  8157.5 93935.0 8375.0 94000.0 ;
      RECT  8342.5 93907.5 8407.5 93967.5 ;
      RECT  8375.0 93875.0 8590.0 93940.0 ;
      RECT  8342.5 95250.0 8407.5 95315.0 ;
      RECT  8342.5 95310.0 8407.5 95375.0 ;
      RECT  8157.5 95250.0 8375.0 95315.0 ;
      RECT  8342.5 95282.5 8407.5 95342.5 ;
      RECT  8375.0 95310.0 8590.0 95375.0 ;
      RECT  8342.5 96625.0 8407.5 96690.0 ;
      RECT  8342.5 96565.0 8407.5 96630.0 ;
      RECT  8157.5 96625.0 8375.0 96690.0 ;
      RECT  8342.5 96597.5 8407.5 96657.5 ;
      RECT  8375.0 96565.0 8590.0 96630.0 ;
      RECT  8342.5 97940.0 8407.5 98005.0 ;
      RECT  8342.5 98000.0 8407.5 98065.0 ;
      RECT  8157.5 97940.0 8375.0 98005.0 ;
      RECT  8342.5 97972.5 8407.5 98032.5 ;
      RECT  8375.0 98000.0 8590.0 98065.0 ;
      RECT  8342.5 99315.0 8407.5 99380.0 ;
      RECT  8342.5 99255.0 8407.5 99320.0 ;
      RECT  8157.5 99315.0 8375.0 99380.0 ;
      RECT  8342.5 99287.5 8407.5 99347.5 ;
      RECT  8375.0 99255.0 8590.0 99320.0 ;
      RECT  8342.5 100630.0 8407.5 100695.0 ;
      RECT  8342.5 100690.0 8407.5 100755.0 ;
      RECT  8157.5 100630.0 8375.0 100695.0 ;
      RECT  8342.5 100662.5 8407.5 100722.5 ;
      RECT  8375.0 100690.0 8590.0 100755.0 ;
      RECT  8342.5 102005.0 8407.5 102070.0 ;
      RECT  8342.5 101945.0 8407.5 102010.0 ;
      RECT  8157.5 102005.0 8375.0 102070.0 ;
      RECT  8342.5 101977.5 8407.5 102037.5 ;
      RECT  8375.0 101945.0 8590.0 102010.0 ;
      RECT  8342.5 103320.0 8407.5 103385.0 ;
      RECT  8342.5 103380.0 8407.5 103445.0 ;
      RECT  8157.5 103320.0 8375.0 103385.0 ;
      RECT  8342.5 103352.5 8407.5 103412.5 ;
      RECT  8375.0 103380.0 8590.0 103445.0 ;
      RECT  8342.5 104695.0 8407.5 104760.0 ;
      RECT  8342.5 104635.0 8407.5 104700.0 ;
      RECT  8157.5 104695.0 8375.0 104760.0 ;
      RECT  8342.5 104667.5 8407.5 104727.5 ;
      RECT  8375.0 104635.0 8590.0 104700.0 ;
      RECT  8342.5 106010.0 8407.5 106075.0 ;
      RECT  8342.5 106070.0 8407.5 106135.0 ;
      RECT  8157.5 106010.0 8375.0 106075.0 ;
      RECT  8342.5 106042.5 8407.5 106102.5 ;
      RECT  8375.0 106070.0 8590.0 106135.0 ;
      RECT  8342.5 107385.0 8407.5 107450.0 ;
      RECT  8342.5 107325.0 8407.5 107390.0 ;
      RECT  8157.5 107385.0 8375.0 107450.0 ;
      RECT  8342.5 107357.5 8407.5 107417.5 ;
      RECT  8375.0 107325.0 8590.0 107390.0 ;
      RECT  8342.5 108700.0 8407.5 108765.0 ;
      RECT  8342.5 108760.0 8407.5 108825.0 ;
      RECT  8157.5 108700.0 8375.0 108765.0 ;
      RECT  8342.5 108732.5 8407.5 108792.5 ;
      RECT  8375.0 108760.0 8590.0 108825.0 ;
      RECT  8342.5 110075.0 8407.5 110140.0 ;
      RECT  8342.5 110015.0 8407.5 110080.0 ;
      RECT  8157.5 110075.0 8375.0 110140.0 ;
      RECT  8342.5 110047.5 8407.5 110107.5 ;
      RECT  8375.0 110015.0 8590.0 110080.0 ;
      RECT  8342.5 111390.0 8407.5 111455.0 ;
      RECT  8342.5 111450.0 8407.5 111515.0 ;
      RECT  8157.5 111390.0 8375.0 111455.0 ;
      RECT  8342.5 111422.5 8407.5 111482.5 ;
      RECT  8375.0 111450.0 8590.0 111515.0 ;
      RECT  8342.5 112765.0 8407.5 112830.0 ;
      RECT  8342.5 112705.0 8407.5 112770.0 ;
      RECT  8157.5 112765.0 8375.0 112830.0 ;
      RECT  8342.5 112737.5 8407.5 112797.5 ;
      RECT  8375.0 112705.0 8590.0 112770.0 ;
      RECT  8342.5 114080.0 8407.5 114145.0 ;
      RECT  8342.5 114140.0 8407.5 114205.0 ;
      RECT  8157.5 114080.0 8375.0 114145.0 ;
      RECT  8342.5 114112.5 8407.5 114172.5 ;
      RECT  8375.0 114140.0 8590.0 114205.0 ;
      RECT  8342.5 115455.0 8407.5 115520.0 ;
      RECT  8342.5 115395.0 8407.5 115460.0 ;
      RECT  8157.5 115455.0 8375.0 115520.0 ;
      RECT  8342.5 115427.5 8407.5 115487.5 ;
      RECT  8375.0 115395.0 8590.0 115460.0 ;
      RECT  8342.5 116770.0 8407.5 116835.0 ;
      RECT  8342.5 116830.0 8407.5 116895.0 ;
      RECT  8157.5 116770.0 8375.0 116835.0 ;
      RECT  8342.5 116802.5 8407.5 116862.5 ;
      RECT  8375.0 116830.0 8590.0 116895.0 ;
      RECT  8342.5 118145.0 8407.5 118210.0 ;
      RECT  8342.5 118085.0 8407.5 118150.0 ;
      RECT  8157.5 118145.0 8375.0 118210.0 ;
      RECT  8342.5 118117.5 8407.5 118177.5 ;
      RECT  8375.0 118085.0 8590.0 118150.0 ;
      RECT  8342.5 119460.0 8407.5 119525.0 ;
      RECT  8342.5 119520.0 8407.5 119585.0 ;
      RECT  8157.5 119460.0 8375.0 119525.0 ;
      RECT  8342.5 119492.5 8407.5 119552.5 ;
      RECT  8375.0 119520.0 8590.0 119585.0 ;
      RECT  8342.5 120835.0 8407.5 120900.0 ;
      RECT  8342.5 120775.0 8407.5 120840.0 ;
      RECT  8157.5 120835.0 8375.0 120900.0 ;
      RECT  8342.5 120807.5 8407.5 120867.5 ;
      RECT  8375.0 120775.0 8590.0 120840.0 ;
      RECT  8342.5 122150.0 8407.5 122215.0 ;
      RECT  8342.5 122210.0 8407.5 122275.0 ;
      RECT  8157.5 122150.0 8375.0 122215.0 ;
      RECT  8342.5 122182.5 8407.5 122242.5 ;
      RECT  8375.0 122210.0 8590.0 122275.0 ;
      RECT  8342.5 123525.0 8407.5 123590.0 ;
      RECT  8342.5 123465.0 8407.5 123530.0 ;
      RECT  8157.5 123525.0 8375.0 123590.0 ;
      RECT  8342.5 123497.5 8407.5 123557.5 ;
      RECT  8375.0 123465.0 8590.0 123530.0 ;
      RECT  8342.5 124840.0 8407.5 124905.0 ;
      RECT  8342.5 124900.0 8407.5 124965.0 ;
      RECT  8157.5 124840.0 8375.0 124905.0 ;
      RECT  8342.5 124872.5 8407.5 124932.5 ;
      RECT  8375.0 124900.0 8590.0 124965.0 ;
      RECT  8342.5 126215.0 8407.5 126280.0 ;
      RECT  8342.5 126155.0 8407.5 126220.0 ;
      RECT  8157.5 126215.0 8375.0 126280.0 ;
      RECT  8342.5 126187.5 8407.5 126247.5 ;
      RECT  8375.0 126155.0 8590.0 126220.0 ;
      RECT  8342.5 127530.0 8407.5 127595.0 ;
      RECT  8342.5 127590.0 8407.5 127655.0 ;
      RECT  8157.5 127530.0 8375.0 127595.0 ;
      RECT  8342.5 127562.5 8407.5 127622.5 ;
      RECT  8375.0 127590.0 8590.0 127655.0 ;
      RECT  8342.5 128905.0 8407.5 128970.0 ;
      RECT  8342.5 128845.0 8407.5 128910.0 ;
      RECT  8157.5 128905.0 8375.0 128970.0 ;
      RECT  8342.5 128877.5 8407.5 128937.5 ;
      RECT  8375.0 128845.0 8590.0 128910.0 ;
      RECT  8342.5 130220.0 8407.5 130285.0 ;
      RECT  8342.5 130280.0 8407.5 130345.0 ;
      RECT  8157.5 130220.0 8375.0 130285.0 ;
      RECT  8342.5 130252.5 8407.5 130312.5 ;
      RECT  8375.0 130280.0 8590.0 130345.0 ;
      RECT  8342.5 131595.0 8407.5 131660.0 ;
      RECT  8342.5 131535.0 8407.5 131600.0 ;
      RECT  8157.5 131595.0 8375.0 131660.0 ;
      RECT  8342.5 131567.5 8407.5 131627.5 ;
      RECT  8375.0 131535.0 8590.0 131600.0 ;
      RECT  8342.5 132910.0 8407.5 132975.0 ;
      RECT  8342.5 132970.0 8407.5 133035.0 ;
      RECT  8157.5 132910.0 8375.0 132975.0 ;
      RECT  8342.5 132942.5 8407.5 133002.5 ;
      RECT  8375.0 132970.0 8590.0 133035.0 ;
      RECT  8342.5 134285.0 8407.5 134350.0 ;
      RECT  8342.5 134225.0 8407.5 134290.0 ;
      RECT  8157.5 134285.0 8375.0 134350.0 ;
      RECT  8342.5 134257.5 8407.5 134317.5 ;
      RECT  8375.0 134225.0 8590.0 134290.0 ;
      RECT  8342.5 135600.0 8407.5 135665.0 ;
      RECT  8342.5 135660.0 8407.5 135725.0 ;
      RECT  8157.5 135600.0 8375.0 135665.0 ;
      RECT  8342.5 135632.5 8407.5 135692.5 ;
      RECT  8375.0 135660.0 8590.0 135725.0 ;
      RECT  8342.5 136975.0 8407.5 137040.0 ;
      RECT  8342.5 136915.0 8407.5 136980.0 ;
      RECT  8157.5 136975.0 8375.0 137040.0 ;
      RECT  8342.5 136947.5 8407.5 137007.5 ;
      RECT  8375.0 136915.0 8590.0 136980.0 ;
      RECT  8342.5 138290.0 8407.5 138355.0 ;
      RECT  8342.5 138350.0 8407.5 138415.0 ;
      RECT  8157.5 138290.0 8375.0 138355.0 ;
      RECT  8342.5 138322.5 8407.5 138382.5 ;
      RECT  8375.0 138350.0 8590.0 138415.0 ;
      RECT  8342.5 139665.0 8407.5 139730.0 ;
      RECT  8342.5 139605.0 8407.5 139670.0 ;
      RECT  8157.5 139665.0 8375.0 139730.0 ;
      RECT  8342.5 139637.5 8407.5 139697.5 ;
      RECT  8375.0 139605.0 8590.0 139670.0 ;
      RECT  8342.5 140980.0 8407.5 141045.0 ;
      RECT  8342.5 141040.0 8407.5 141105.0 ;
      RECT  8157.5 140980.0 8375.0 141045.0 ;
      RECT  8342.5 141012.5 8407.5 141072.5 ;
      RECT  8375.0 141040.0 8590.0 141105.0 ;
      RECT  8342.5 142355.0 8407.5 142420.0 ;
      RECT  8342.5 142295.0 8407.5 142360.0 ;
      RECT  8157.5 142355.0 8375.0 142420.0 ;
      RECT  8342.5 142327.5 8407.5 142387.5 ;
      RECT  8375.0 142295.0 8590.0 142360.0 ;
      RECT  8342.5 143670.0 8407.5 143735.0 ;
      RECT  8342.5 143730.0 8407.5 143795.0 ;
      RECT  8157.5 143670.0 8375.0 143735.0 ;
      RECT  8342.5 143702.5 8407.5 143762.5 ;
      RECT  8375.0 143730.0 8590.0 143795.0 ;
      RECT  8342.5 145045.0 8407.5 145110.0 ;
      RECT  8342.5 144985.0 8407.5 145050.0 ;
      RECT  8157.5 145045.0 8375.0 145110.0 ;
      RECT  8342.5 145017.5 8407.5 145077.5 ;
      RECT  8375.0 144985.0 8590.0 145050.0 ;
      RECT  8342.5 146360.0 8407.5 146425.0 ;
      RECT  8342.5 146420.0 8407.5 146485.0 ;
      RECT  8157.5 146360.0 8375.0 146425.0 ;
      RECT  8342.5 146392.5 8407.5 146452.5 ;
      RECT  8375.0 146420.0 8590.0 146485.0 ;
      RECT  8342.5 147735.0 8407.5 147800.0 ;
      RECT  8342.5 147675.0 8407.5 147740.0 ;
      RECT  8157.5 147735.0 8375.0 147800.0 ;
      RECT  8342.5 147707.5 8407.5 147767.5 ;
      RECT  8375.0 147675.0 8590.0 147740.0 ;
      RECT  8342.5 149050.0 8407.5 149115.0 ;
      RECT  8342.5 149110.0 8407.5 149175.0 ;
      RECT  8157.5 149050.0 8375.0 149115.0 ;
      RECT  8342.5 149082.5 8407.5 149142.5 ;
      RECT  8375.0 149110.0 8590.0 149175.0 ;
      RECT  8342.5 150425.0 8407.5 150490.0 ;
      RECT  8342.5 150365.0 8407.5 150430.0 ;
      RECT  8157.5 150425.0 8375.0 150490.0 ;
      RECT  8342.5 150397.5 8407.5 150457.5 ;
      RECT  8375.0 150365.0 8590.0 150430.0 ;
      RECT  8342.5 151740.0 8407.5 151805.0 ;
      RECT  8342.5 151800.0 8407.5 151865.0 ;
      RECT  8157.5 151740.0 8375.0 151805.0 ;
      RECT  8342.5 151772.5 8407.5 151832.5 ;
      RECT  8375.0 151800.0 8590.0 151865.0 ;
      RECT  8342.5 153115.0 8407.5 153180.0 ;
      RECT  8342.5 153055.0 8407.5 153120.0 ;
      RECT  8157.5 153115.0 8375.0 153180.0 ;
      RECT  8342.5 153087.5 8407.5 153147.5 ;
      RECT  8375.0 153055.0 8590.0 153120.0 ;
      RECT  8342.5 154430.0 8407.5 154495.0 ;
      RECT  8342.5 154490.0 8407.5 154555.0 ;
      RECT  8157.5 154430.0 8375.0 154495.0 ;
      RECT  8342.5 154462.5 8407.5 154522.5 ;
      RECT  8375.0 154490.0 8590.0 154555.0 ;
      RECT  8342.5 155805.0 8407.5 155870.0 ;
      RECT  8342.5 155745.0 8407.5 155810.0 ;
      RECT  8157.5 155805.0 8375.0 155870.0 ;
      RECT  8342.5 155777.5 8407.5 155837.5 ;
      RECT  8375.0 155745.0 8590.0 155810.0 ;
      RECT  8342.5 157120.0 8407.5 157185.0 ;
      RECT  8342.5 157180.0 8407.5 157245.0 ;
      RECT  8157.5 157120.0 8375.0 157185.0 ;
      RECT  8342.5 157152.5 8407.5 157212.5 ;
      RECT  8375.0 157180.0 8590.0 157245.0 ;
      RECT  8342.5 158495.0 8407.5 158560.0 ;
      RECT  8342.5 158435.0 8407.5 158500.0 ;
      RECT  8157.5 158495.0 8375.0 158560.0 ;
      RECT  8342.5 158467.5 8407.5 158527.5 ;
      RECT  8375.0 158435.0 8590.0 158500.0 ;
      RECT  8342.5 159810.0 8407.5 159875.0 ;
      RECT  8342.5 159870.0 8407.5 159935.0 ;
      RECT  8157.5 159810.0 8375.0 159875.0 ;
      RECT  8342.5 159842.5 8407.5 159902.5 ;
      RECT  8375.0 159870.0 8590.0 159935.0 ;
      RECT  8342.5 161185.0 8407.5 161250.0 ;
      RECT  8342.5 161125.0 8407.5 161190.0 ;
      RECT  8157.5 161185.0 8375.0 161250.0 ;
      RECT  8342.5 161157.5 8407.5 161217.5 ;
      RECT  8375.0 161125.0 8590.0 161190.0 ;
      RECT  8342.5 162500.0 8407.5 162565.0 ;
      RECT  8342.5 162560.0 8407.5 162625.0 ;
      RECT  8157.5 162500.0 8375.0 162565.0 ;
      RECT  8342.5 162532.5 8407.5 162592.5 ;
      RECT  8375.0 162560.0 8590.0 162625.0 ;
      RECT  8342.5 163875.0 8407.5 163940.0 ;
      RECT  8342.5 163815.0 8407.5 163880.0 ;
      RECT  8157.5 163875.0 8375.0 163940.0 ;
      RECT  8342.5 163847.5 8407.5 163907.5 ;
      RECT  8375.0 163815.0 8590.0 163880.0 ;
      RECT  8342.5 165190.0 8407.5 165255.0 ;
      RECT  8342.5 165250.0 8407.5 165315.0 ;
      RECT  8157.5 165190.0 8375.0 165255.0 ;
      RECT  8342.5 165222.5 8407.5 165282.5 ;
      RECT  8375.0 165250.0 8590.0 165315.0 ;
      RECT  8342.5 166565.0 8407.5 166630.0 ;
      RECT  8342.5 166505.0 8407.5 166570.0 ;
      RECT  8157.5 166565.0 8375.0 166630.0 ;
      RECT  8342.5 166537.5 8407.5 166597.5 ;
      RECT  8375.0 166505.0 8590.0 166570.0 ;
      RECT  8342.5 167880.0 8407.5 167945.0 ;
      RECT  8342.5 167940.0 8407.5 168005.0 ;
      RECT  8157.5 167880.0 8375.0 167945.0 ;
      RECT  8342.5 167912.5 8407.5 167972.5 ;
      RECT  8375.0 167940.0 8590.0 168005.0 ;
      RECT  8342.5 169255.0 8407.5 169320.0 ;
      RECT  8342.5 169195.0 8407.5 169260.0 ;
      RECT  8157.5 169255.0 8375.0 169320.0 ;
      RECT  8342.5 169227.5 8407.5 169287.5 ;
      RECT  8375.0 169195.0 8590.0 169260.0 ;
      RECT  8342.5 170570.0 8407.5 170635.0 ;
      RECT  8342.5 170630.0 8407.5 170695.0 ;
      RECT  8157.5 170570.0 8375.0 170635.0 ;
      RECT  8342.5 170602.5 8407.5 170662.5 ;
      RECT  8375.0 170630.0 8590.0 170695.0 ;
      RECT  8342.5 171945.0 8407.5 172010.0 ;
      RECT  8342.5 171885.0 8407.5 171950.0 ;
      RECT  8157.5 171945.0 8375.0 172010.0 ;
      RECT  8342.5 171917.5 8407.5 171977.5 ;
      RECT  8375.0 171885.0 8590.0 171950.0 ;
      RECT  8342.5 173260.0 8407.5 173325.0 ;
      RECT  8342.5 173320.0 8407.5 173385.0 ;
      RECT  8157.5 173260.0 8375.0 173325.0 ;
      RECT  8342.5 173292.5 8407.5 173352.5 ;
      RECT  8375.0 173320.0 8590.0 173385.0 ;
      RECT  8342.5 174635.0 8407.5 174700.0 ;
      RECT  8342.5 174575.0 8407.5 174640.0 ;
      RECT  8157.5 174635.0 8375.0 174700.0 ;
      RECT  8342.5 174607.5 8407.5 174667.5 ;
      RECT  8375.0 174575.0 8590.0 174640.0 ;
      RECT  8342.5 175950.0 8407.5 176015.0 ;
      RECT  8342.5 176010.0 8407.5 176075.0 ;
      RECT  8157.5 175950.0 8375.0 176015.0 ;
      RECT  8342.5 175982.5 8407.5 176042.5 ;
      RECT  8375.0 176010.0 8590.0 176075.0 ;
      RECT  8342.5 177325.0 8407.5 177390.0 ;
      RECT  8342.5 177265.0 8407.5 177330.0 ;
      RECT  8157.5 177325.0 8375.0 177390.0 ;
      RECT  8342.5 177297.5 8407.5 177357.5 ;
      RECT  8375.0 177265.0 8590.0 177330.0 ;
      RECT  8342.5 178640.0 8407.5 178705.0 ;
      RECT  8342.5 178700.0 8407.5 178765.0 ;
      RECT  8157.5 178640.0 8375.0 178705.0 ;
      RECT  8342.5 178672.5 8407.5 178732.5 ;
      RECT  8375.0 178700.0 8590.0 178765.0 ;
      RECT  8342.5 180015.0 8407.5 180080.0 ;
      RECT  8342.5 179955.0 8407.5 180020.0 ;
      RECT  8157.5 180015.0 8375.0 180080.0 ;
      RECT  8342.5 179987.5 8407.5 180047.5 ;
      RECT  8375.0 179955.0 8590.0 180020.0 ;
      RECT  8342.5 181330.0 8407.5 181395.0 ;
      RECT  8342.5 181390.0 8407.5 181455.0 ;
      RECT  8157.5 181330.0 8375.0 181395.0 ;
      RECT  8342.5 181362.5 8407.5 181422.5 ;
      RECT  8375.0 181390.0 8590.0 181455.0 ;
      RECT  8342.5 182705.0 8407.5 182770.0 ;
      RECT  8342.5 182645.0 8407.5 182710.0 ;
      RECT  8157.5 182705.0 8375.0 182770.0 ;
      RECT  8342.5 182677.5 8407.5 182737.5 ;
      RECT  8375.0 182645.0 8590.0 182710.0 ;
      RECT  8342.5 184020.0 8407.5 184085.0 ;
      RECT  8342.5 184080.0 8407.5 184145.0 ;
      RECT  8157.5 184020.0 8375.0 184085.0 ;
      RECT  8342.5 184052.5 8407.5 184112.5 ;
      RECT  8375.0 184080.0 8590.0 184145.0 ;
      RECT  8342.5 185395.0 8407.5 185460.0 ;
      RECT  8342.5 185335.0 8407.5 185400.0 ;
      RECT  8157.5 185395.0 8375.0 185460.0 ;
      RECT  8342.5 185367.5 8407.5 185427.5 ;
      RECT  8375.0 185335.0 8590.0 185400.0 ;
      RECT  8342.5 186710.0 8407.5 186775.0 ;
      RECT  8342.5 186770.0 8407.5 186835.0 ;
      RECT  8157.5 186710.0 8375.0 186775.0 ;
      RECT  8342.5 186742.5 8407.5 186802.5 ;
      RECT  8375.0 186770.0 8590.0 186835.0 ;
      RECT  8342.5 188085.0 8407.5 188150.0 ;
      RECT  8342.5 188025.0 8407.5 188090.0 ;
      RECT  8157.5 188085.0 8375.0 188150.0 ;
      RECT  8342.5 188057.5 8407.5 188117.5 ;
      RECT  8375.0 188025.0 8590.0 188090.0 ;
      RECT  8342.5 189400.0 8407.5 189465.0 ;
      RECT  8342.5 189460.0 8407.5 189525.0 ;
      RECT  8157.5 189400.0 8375.0 189465.0 ;
      RECT  8342.5 189432.5 8407.5 189492.5 ;
      RECT  8375.0 189460.0 8590.0 189525.0 ;
      RECT  8342.5 190775.0 8407.5 190840.0 ;
      RECT  8342.5 190715.0 8407.5 190780.0 ;
      RECT  8157.5 190775.0 8375.0 190840.0 ;
      RECT  8342.5 190747.5 8407.5 190807.5 ;
      RECT  8375.0 190715.0 8590.0 190780.0 ;
      RECT  8342.5 192090.0 8407.5 192155.0 ;
      RECT  8342.5 192150.0 8407.5 192215.0 ;
      RECT  8157.5 192090.0 8375.0 192155.0 ;
      RECT  8342.5 192122.5 8407.5 192182.5 ;
      RECT  8375.0 192150.0 8590.0 192215.0 ;
      RECT  8342.5 193465.0 8407.5 193530.0 ;
      RECT  8342.5 193405.0 8407.5 193470.0 ;
      RECT  8157.5 193465.0 8375.0 193530.0 ;
      RECT  8342.5 193437.5 8407.5 193497.5 ;
      RECT  8375.0 193405.0 8590.0 193470.0 ;
      RECT  8342.5 194780.0 8407.5 194845.0 ;
      RECT  8342.5 194840.0 8407.5 194905.0 ;
      RECT  8157.5 194780.0 8375.0 194845.0 ;
      RECT  8342.5 194812.5 8407.5 194872.5 ;
      RECT  8375.0 194840.0 8590.0 194905.0 ;
      RECT  8342.5 196155.0 8407.5 196220.0 ;
      RECT  8342.5 196095.0 8407.5 196160.0 ;
      RECT  8157.5 196155.0 8375.0 196220.0 ;
      RECT  8342.5 196127.5 8407.5 196187.5 ;
      RECT  8375.0 196095.0 8590.0 196160.0 ;
      RECT  8342.5 197470.0 8407.5 197535.0 ;
      RECT  8342.5 197530.0 8407.5 197595.0 ;
      RECT  8157.5 197470.0 8375.0 197535.0 ;
      RECT  8342.5 197502.5 8407.5 197562.5 ;
      RECT  8375.0 197530.0 8590.0 197595.0 ;
      RECT  8342.5 198845.0 8407.5 198910.0 ;
      RECT  8342.5 198785.0 8407.5 198850.0 ;
      RECT  8157.5 198845.0 8375.0 198910.0 ;
      RECT  8342.5 198817.5 8407.5 198877.5 ;
      RECT  8375.0 198785.0 8590.0 198850.0 ;
      RECT  8342.5 200160.0 8407.5 200225.0 ;
      RECT  8342.5 200220.0 8407.5 200285.0 ;
      RECT  8157.5 200160.0 8375.0 200225.0 ;
      RECT  8342.5 200192.5 8407.5 200252.5 ;
      RECT  8375.0 200220.0 8590.0 200285.0 ;
      RECT  8342.5 201535.0 8407.5 201600.0 ;
      RECT  8342.5 201475.0 8407.5 201540.0 ;
      RECT  8157.5 201535.0 8375.0 201600.0 ;
      RECT  8342.5 201507.5 8407.5 201567.5 ;
      RECT  8375.0 201475.0 8590.0 201540.0 ;
      RECT  8342.5 202850.0 8407.5 202915.0 ;
      RECT  8342.5 202910.0 8407.5 202975.0 ;
      RECT  8157.5 202850.0 8375.0 202915.0 ;
      RECT  8342.5 202882.5 8407.5 202942.5 ;
      RECT  8375.0 202910.0 8590.0 202975.0 ;
      RECT  8342.5 204225.0 8407.5 204290.0 ;
      RECT  8342.5 204165.0 8407.5 204230.0 ;
      RECT  8157.5 204225.0 8375.0 204290.0 ;
      RECT  8342.5 204197.5 8407.5 204257.5 ;
      RECT  8375.0 204165.0 8590.0 204230.0 ;
      RECT  8342.5 205540.0 8407.5 205605.0 ;
      RECT  8342.5 205600.0 8407.5 205665.0 ;
      RECT  8157.5 205540.0 8375.0 205605.0 ;
      RECT  8342.5 205572.5 8407.5 205632.5 ;
      RECT  8375.0 205600.0 8590.0 205665.0 ;
      RECT  4690.0 13175.0 7455.0 13240.0 ;
      RECT  4865.0 14610.0 7455.0 14675.0 ;
      RECT  5040.0 15865.0 7455.0 15930.0 ;
      RECT  5215.0 17300.0 7455.0 17365.0 ;
      RECT  5390.0 18555.0 7455.0 18620.0 ;
      RECT  5565.0 19990.0 7455.0 20055.0 ;
      RECT  5740.0 21245.0 7455.0 21310.0 ;
      RECT  5915.0 22680.0 7455.0 22745.0 ;
      RECT  6090.0 23935.0 7455.0 24000.0 ;
      RECT  6265.0 25370.0 7455.0 25435.0 ;
      RECT  6440.0 26625.0 7455.0 26690.0 ;
      RECT  6615.0 28060.0 7455.0 28125.0 ;
      RECT  6790.0 29315.0 7455.0 29380.0 ;
      RECT  6965.0 30750.0 7455.0 30815.0 ;
      RECT  7140.0 32005.0 7455.0 32070.0 ;
      RECT  7315.0 33440.0 7455.0 33505.0 ;
      RECT  4690.0 34755.0 7582.5 34820.0 ;
      RECT  5390.0 34615.0 7772.5 34680.0 ;
      RECT  6090.0 34475.0 7962.5 34540.0 ;
      RECT  4690.0 36070.0 7582.5 36135.0 ;
      RECT  5390.0 36210.0 7772.5 36275.0 ;
      RECT  6265.0 36350.0 7962.5 36415.0 ;
      RECT  4690.0 37445.0 7582.5 37510.0 ;
      RECT  5390.0 37305.0 7772.5 37370.0 ;
      RECT  6440.0 37165.0 7962.5 37230.0 ;
      RECT  4690.0 38760.0 7582.5 38825.0 ;
      RECT  5390.0 38900.0 7772.5 38965.0 ;
      RECT  6615.0 39040.0 7962.5 39105.0 ;
      RECT  4690.0 40135.0 7582.5 40200.0 ;
      RECT  5390.0 39995.0 7772.5 40060.0 ;
      RECT  6790.0 39855.0 7962.5 39920.0 ;
      RECT  4690.0 41450.0 7582.5 41515.0 ;
      RECT  5390.0 41590.0 7772.5 41655.0 ;
      RECT  6965.0 41730.0 7962.5 41795.0 ;
      RECT  4690.0 42825.0 7582.5 42890.0 ;
      RECT  5390.0 42685.0 7772.5 42750.0 ;
      RECT  7140.0 42545.0 7962.5 42610.0 ;
      RECT  4690.0 44140.0 7582.5 44205.0 ;
      RECT  5390.0 44280.0 7772.5 44345.0 ;
      RECT  7315.0 44420.0 7962.5 44485.0 ;
      RECT  4690.0 45515.0 7582.5 45580.0 ;
      RECT  5565.0 45375.0 7772.5 45440.0 ;
      RECT  6090.0 45235.0 7962.5 45300.0 ;
      RECT  4690.0 46830.0 7582.5 46895.0 ;
      RECT  5565.0 46970.0 7772.5 47035.0 ;
      RECT  6265.0 47110.0 7962.5 47175.0 ;
      RECT  4690.0 48205.0 7582.5 48270.0 ;
      RECT  5565.0 48065.0 7772.5 48130.0 ;
      RECT  6440.0 47925.0 7962.5 47990.0 ;
      RECT  4690.0 49520.0 7582.5 49585.0 ;
      RECT  5565.0 49660.0 7772.5 49725.0 ;
      RECT  6615.0 49800.0 7962.5 49865.0 ;
      RECT  4690.0 50895.0 7582.5 50960.0 ;
      RECT  5565.0 50755.0 7772.5 50820.0 ;
      RECT  6790.0 50615.0 7962.5 50680.0 ;
      RECT  4690.0 52210.0 7582.5 52275.0 ;
      RECT  5565.0 52350.0 7772.5 52415.0 ;
      RECT  6965.0 52490.0 7962.5 52555.0 ;
      RECT  4690.0 53585.0 7582.5 53650.0 ;
      RECT  5565.0 53445.0 7772.5 53510.0 ;
      RECT  7140.0 53305.0 7962.5 53370.0 ;
      RECT  4690.0 54900.0 7582.5 54965.0 ;
      RECT  5565.0 55040.0 7772.5 55105.0 ;
      RECT  7315.0 55180.0 7962.5 55245.0 ;
      RECT  4690.0 56275.0 7582.5 56340.0 ;
      RECT  5740.0 56135.0 7772.5 56200.0 ;
      RECT  6090.0 55995.0 7962.5 56060.0 ;
      RECT  4690.0 57590.0 7582.5 57655.0 ;
      RECT  5740.0 57730.0 7772.5 57795.0 ;
      RECT  6265.0 57870.0 7962.5 57935.0 ;
      RECT  4690.0 58965.0 7582.5 59030.0 ;
      RECT  5740.0 58825.0 7772.5 58890.0 ;
      RECT  6440.0 58685.0 7962.5 58750.0 ;
      RECT  4690.0 60280.0 7582.5 60345.0 ;
      RECT  5740.0 60420.0 7772.5 60485.0 ;
      RECT  6615.0 60560.0 7962.5 60625.0 ;
      RECT  4690.0 61655.0 7582.5 61720.0 ;
      RECT  5740.0 61515.0 7772.5 61580.0 ;
      RECT  6790.0 61375.0 7962.5 61440.0 ;
      RECT  4690.0 62970.0 7582.5 63035.0 ;
      RECT  5740.0 63110.0 7772.5 63175.0 ;
      RECT  6965.0 63250.0 7962.5 63315.0 ;
      RECT  4690.0 64345.0 7582.5 64410.0 ;
      RECT  5740.0 64205.0 7772.5 64270.0 ;
      RECT  7140.0 64065.0 7962.5 64130.0 ;
      RECT  4690.0 65660.0 7582.5 65725.0 ;
      RECT  5740.0 65800.0 7772.5 65865.0 ;
      RECT  7315.0 65940.0 7962.5 66005.0 ;
      RECT  4690.0 67035.0 7582.5 67100.0 ;
      RECT  5915.0 66895.0 7772.5 66960.0 ;
      RECT  6090.0 66755.0 7962.5 66820.0 ;
      RECT  4690.0 68350.0 7582.5 68415.0 ;
      RECT  5915.0 68490.0 7772.5 68555.0 ;
      RECT  6265.0 68630.0 7962.5 68695.0 ;
      RECT  4690.0 69725.0 7582.5 69790.0 ;
      RECT  5915.0 69585.0 7772.5 69650.0 ;
      RECT  6440.0 69445.0 7962.5 69510.0 ;
      RECT  4690.0 71040.0 7582.5 71105.0 ;
      RECT  5915.0 71180.0 7772.5 71245.0 ;
      RECT  6615.0 71320.0 7962.5 71385.0 ;
      RECT  4690.0 72415.0 7582.5 72480.0 ;
      RECT  5915.0 72275.0 7772.5 72340.0 ;
      RECT  6790.0 72135.0 7962.5 72200.0 ;
      RECT  4690.0 73730.0 7582.5 73795.0 ;
      RECT  5915.0 73870.0 7772.5 73935.0 ;
      RECT  6965.0 74010.0 7962.5 74075.0 ;
      RECT  4690.0 75105.0 7582.5 75170.0 ;
      RECT  5915.0 74965.0 7772.5 75030.0 ;
      RECT  7140.0 74825.0 7962.5 74890.0 ;
      RECT  4690.0 76420.0 7582.5 76485.0 ;
      RECT  5915.0 76560.0 7772.5 76625.0 ;
      RECT  7315.0 76700.0 7962.5 76765.0 ;
      RECT  4865.0 77795.0 7582.5 77860.0 ;
      RECT  5390.0 77655.0 7772.5 77720.0 ;
      RECT  6090.0 77515.0 7962.5 77580.0 ;
      RECT  4865.0 79110.0 7582.5 79175.0 ;
      RECT  5390.0 79250.0 7772.5 79315.0 ;
      RECT  6265.0 79390.0 7962.5 79455.0 ;
      RECT  4865.0 80485.0 7582.5 80550.0 ;
      RECT  5390.0 80345.0 7772.5 80410.0 ;
      RECT  6440.0 80205.0 7962.5 80270.0 ;
      RECT  4865.0 81800.0 7582.5 81865.0 ;
      RECT  5390.0 81940.0 7772.5 82005.0 ;
      RECT  6615.0 82080.0 7962.5 82145.0 ;
      RECT  4865.0 83175.0 7582.5 83240.0 ;
      RECT  5390.0 83035.0 7772.5 83100.0 ;
      RECT  6790.0 82895.0 7962.5 82960.0 ;
      RECT  4865.0 84490.0 7582.5 84555.0 ;
      RECT  5390.0 84630.0 7772.5 84695.0 ;
      RECT  6965.0 84770.0 7962.5 84835.0 ;
      RECT  4865.0 85865.0 7582.5 85930.0 ;
      RECT  5390.0 85725.0 7772.5 85790.0 ;
      RECT  7140.0 85585.0 7962.5 85650.0 ;
      RECT  4865.0 87180.0 7582.5 87245.0 ;
      RECT  5390.0 87320.0 7772.5 87385.0 ;
      RECT  7315.0 87460.0 7962.5 87525.0 ;
      RECT  4865.0 88555.0 7582.5 88620.0 ;
      RECT  5565.0 88415.0 7772.5 88480.0 ;
      RECT  6090.0 88275.0 7962.5 88340.0 ;
      RECT  4865.0 89870.0 7582.5 89935.0 ;
      RECT  5565.0 90010.0 7772.5 90075.0 ;
      RECT  6265.0 90150.0 7962.5 90215.0 ;
      RECT  4865.0 91245.0 7582.5 91310.0 ;
      RECT  5565.0 91105.0 7772.5 91170.0 ;
      RECT  6440.0 90965.0 7962.5 91030.0 ;
      RECT  4865.0 92560.0 7582.5 92625.0 ;
      RECT  5565.0 92700.0 7772.5 92765.0 ;
      RECT  6615.0 92840.0 7962.5 92905.0 ;
      RECT  4865.0 93935.0 7582.5 94000.0 ;
      RECT  5565.0 93795.0 7772.5 93860.0 ;
      RECT  6790.0 93655.0 7962.5 93720.0 ;
      RECT  4865.0 95250.0 7582.5 95315.0 ;
      RECT  5565.0 95390.0 7772.5 95455.0 ;
      RECT  6965.0 95530.0 7962.5 95595.0 ;
      RECT  4865.0 96625.0 7582.5 96690.0 ;
      RECT  5565.0 96485.0 7772.5 96550.0 ;
      RECT  7140.0 96345.0 7962.5 96410.0 ;
      RECT  4865.0 97940.0 7582.5 98005.0 ;
      RECT  5565.0 98080.0 7772.5 98145.0 ;
      RECT  7315.0 98220.0 7962.5 98285.0 ;
      RECT  4865.0 99315.0 7582.5 99380.0 ;
      RECT  5740.0 99175.0 7772.5 99240.0 ;
      RECT  6090.0 99035.0 7962.5 99100.0 ;
      RECT  4865.0 100630.0 7582.5 100695.0 ;
      RECT  5740.0 100770.0 7772.5 100835.0 ;
      RECT  6265.0 100910.0 7962.5 100975.0 ;
      RECT  4865.0 102005.0 7582.5 102070.0 ;
      RECT  5740.0 101865.0 7772.5 101930.0 ;
      RECT  6440.0 101725.0 7962.5 101790.0 ;
      RECT  4865.0 103320.0 7582.5 103385.0 ;
      RECT  5740.0 103460.0 7772.5 103525.0 ;
      RECT  6615.0 103600.0 7962.5 103665.0 ;
      RECT  4865.0 104695.0 7582.5 104760.0 ;
      RECT  5740.0 104555.0 7772.5 104620.0 ;
      RECT  6790.0 104415.0 7962.5 104480.0 ;
      RECT  4865.0 106010.0 7582.5 106075.0 ;
      RECT  5740.0 106150.0 7772.5 106215.0 ;
      RECT  6965.0 106290.0 7962.5 106355.0 ;
      RECT  4865.0 107385.0 7582.5 107450.0 ;
      RECT  5740.0 107245.0 7772.5 107310.0 ;
      RECT  7140.0 107105.0 7962.5 107170.0 ;
      RECT  4865.0 108700.0 7582.5 108765.0 ;
      RECT  5740.0 108840.0 7772.5 108905.0 ;
      RECT  7315.0 108980.0 7962.5 109045.0 ;
      RECT  4865.0 110075.0 7582.5 110140.0 ;
      RECT  5915.0 109935.0 7772.5 110000.0 ;
      RECT  6090.0 109795.0 7962.5 109860.0 ;
      RECT  4865.0 111390.0 7582.5 111455.0 ;
      RECT  5915.0 111530.0 7772.5 111595.0 ;
      RECT  6265.0 111670.0 7962.5 111735.0 ;
      RECT  4865.0 112765.0 7582.5 112830.0 ;
      RECT  5915.0 112625.0 7772.5 112690.0 ;
      RECT  6440.0 112485.0 7962.5 112550.0 ;
      RECT  4865.0 114080.0 7582.5 114145.0 ;
      RECT  5915.0 114220.0 7772.5 114285.0 ;
      RECT  6615.0 114360.0 7962.5 114425.0 ;
      RECT  4865.0 115455.0 7582.5 115520.0 ;
      RECT  5915.0 115315.0 7772.5 115380.0 ;
      RECT  6790.0 115175.0 7962.5 115240.0 ;
      RECT  4865.0 116770.0 7582.5 116835.0 ;
      RECT  5915.0 116910.0 7772.5 116975.0 ;
      RECT  6965.0 117050.0 7962.5 117115.0 ;
      RECT  4865.0 118145.0 7582.5 118210.0 ;
      RECT  5915.0 118005.0 7772.5 118070.0 ;
      RECT  7140.0 117865.0 7962.5 117930.0 ;
      RECT  4865.0 119460.0 7582.5 119525.0 ;
      RECT  5915.0 119600.0 7772.5 119665.0 ;
      RECT  7315.0 119740.0 7962.5 119805.0 ;
      RECT  5040.0 120835.0 7582.5 120900.0 ;
      RECT  5390.0 120695.0 7772.5 120760.0 ;
      RECT  6090.0 120555.0 7962.5 120620.0 ;
      RECT  5040.0 122150.0 7582.5 122215.0 ;
      RECT  5390.0 122290.0 7772.5 122355.0 ;
      RECT  6265.0 122430.0 7962.5 122495.0 ;
      RECT  5040.0 123525.0 7582.5 123590.0 ;
      RECT  5390.0 123385.0 7772.5 123450.0 ;
      RECT  6440.0 123245.0 7962.5 123310.0 ;
      RECT  5040.0 124840.0 7582.5 124905.0 ;
      RECT  5390.0 124980.0 7772.5 125045.0 ;
      RECT  6615.0 125120.0 7962.5 125185.0 ;
      RECT  5040.0 126215.0 7582.5 126280.0 ;
      RECT  5390.0 126075.0 7772.5 126140.0 ;
      RECT  6790.0 125935.0 7962.5 126000.0 ;
      RECT  5040.0 127530.0 7582.5 127595.0 ;
      RECT  5390.0 127670.0 7772.5 127735.0 ;
      RECT  6965.0 127810.0 7962.5 127875.0 ;
      RECT  5040.0 128905.0 7582.5 128970.0 ;
      RECT  5390.0 128765.0 7772.5 128830.0 ;
      RECT  7140.0 128625.0 7962.5 128690.0 ;
      RECT  5040.0 130220.0 7582.5 130285.0 ;
      RECT  5390.0 130360.0 7772.5 130425.0 ;
      RECT  7315.0 130500.0 7962.5 130565.0 ;
      RECT  5040.0 131595.0 7582.5 131660.0 ;
      RECT  5565.0 131455.0 7772.5 131520.0 ;
      RECT  6090.0 131315.0 7962.5 131380.0 ;
      RECT  5040.0 132910.0 7582.5 132975.0 ;
      RECT  5565.0 133050.0 7772.5 133115.0 ;
      RECT  6265.0 133190.0 7962.5 133255.0 ;
      RECT  5040.0 134285.0 7582.5 134350.0 ;
      RECT  5565.0 134145.0 7772.5 134210.0 ;
      RECT  6440.0 134005.0 7962.5 134070.0 ;
      RECT  5040.0 135600.0 7582.5 135665.0 ;
      RECT  5565.0 135740.0 7772.5 135805.0 ;
      RECT  6615.0 135880.0 7962.5 135945.0 ;
      RECT  5040.0 136975.0 7582.5 137040.0 ;
      RECT  5565.0 136835.0 7772.5 136900.0 ;
      RECT  6790.0 136695.0 7962.5 136760.0 ;
      RECT  5040.0 138290.0 7582.5 138355.0 ;
      RECT  5565.0 138430.0 7772.5 138495.0 ;
      RECT  6965.0 138570.0 7962.5 138635.0 ;
      RECT  5040.0 139665.0 7582.5 139730.0 ;
      RECT  5565.0 139525.0 7772.5 139590.0 ;
      RECT  7140.0 139385.0 7962.5 139450.0 ;
      RECT  5040.0 140980.0 7582.5 141045.0 ;
      RECT  5565.0 141120.0 7772.5 141185.0 ;
      RECT  7315.0 141260.0 7962.5 141325.0 ;
      RECT  5040.0 142355.0 7582.5 142420.0 ;
      RECT  5740.0 142215.0 7772.5 142280.0 ;
      RECT  6090.0 142075.0 7962.5 142140.0 ;
      RECT  5040.0 143670.0 7582.5 143735.0 ;
      RECT  5740.0 143810.0 7772.5 143875.0 ;
      RECT  6265.0 143950.0 7962.5 144015.0 ;
      RECT  5040.0 145045.0 7582.5 145110.0 ;
      RECT  5740.0 144905.0 7772.5 144970.0 ;
      RECT  6440.0 144765.0 7962.5 144830.0 ;
      RECT  5040.0 146360.0 7582.5 146425.0 ;
      RECT  5740.0 146500.0 7772.5 146565.0 ;
      RECT  6615.0 146640.0 7962.5 146705.0 ;
      RECT  5040.0 147735.0 7582.5 147800.0 ;
      RECT  5740.0 147595.0 7772.5 147660.0 ;
      RECT  6790.0 147455.0 7962.5 147520.0 ;
      RECT  5040.0 149050.0 7582.5 149115.0 ;
      RECT  5740.0 149190.0 7772.5 149255.0 ;
      RECT  6965.0 149330.0 7962.5 149395.0 ;
      RECT  5040.0 150425.0 7582.5 150490.0 ;
      RECT  5740.0 150285.0 7772.5 150350.0 ;
      RECT  7140.0 150145.0 7962.5 150210.0 ;
      RECT  5040.0 151740.0 7582.5 151805.0 ;
      RECT  5740.0 151880.0 7772.5 151945.0 ;
      RECT  7315.0 152020.0 7962.5 152085.0 ;
      RECT  5040.0 153115.0 7582.5 153180.0 ;
      RECT  5915.0 152975.0 7772.5 153040.0 ;
      RECT  6090.0 152835.0 7962.5 152900.0 ;
      RECT  5040.0 154430.0 7582.5 154495.0 ;
      RECT  5915.0 154570.0 7772.5 154635.0 ;
      RECT  6265.0 154710.0 7962.5 154775.0 ;
      RECT  5040.0 155805.0 7582.5 155870.0 ;
      RECT  5915.0 155665.0 7772.5 155730.0 ;
      RECT  6440.0 155525.0 7962.5 155590.0 ;
      RECT  5040.0 157120.0 7582.5 157185.0 ;
      RECT  5915.0 157260.0 7772.5 157325.0 ;
      RECT  6615.0 157400.0 7962.5 157465.0 ;
      RECT  5040.0 158495.0 7582.5 158560.0 ;
      RECT  5915.0 158355.0 7772.5 158420.0 ;
      RECT  6790.0 158215.0 7962.5 158280.0 ;
      RECT  5040.0 159810.0 7582.5 159875.0 ;
      RECT  5915.0 159950.0 7772.5 160015.0 ;
      RECT  6965.0 160090.0 7962.5 160155.0 ;
      RECT  5040.0 161185.0 7582.5 161250.0 ;
      RECT  5915.0 161045.0 7772.5 161110.0 ;
      RECT  7140.0 160905.0 7962.5 160970.0 ;
      RECT  5040.0 162500.0 7582.5 162565.0 ;
      RECT  5915.0 162640.0 7772.5 162705.0 ;
      RECT  7315.0 162780.0 7962.5 162845.0 ;
      RECT  5215.0 163875.0 7582.5 163940.0 ;
      RECT  5390.0 163735.0 7772.5 163800.0 ;
      RECT  6090.0 163595.0 7962.5 163660.0 ;
      RECT  5215.0 165190.0 7582.5 165255.0 ;
      RECT  5390.0 165330.0 7772.5 165395.0 ;
      RECT  6265.0 165470.0 7962.5 165535.0 ;
      RECT  5215.0 166565.0 7582.5 166630.0 ;
      RECT  5390.0 166425.0 7772.5 166490.0 ;
      RECT  6440.0 166285.0 7962.5 166350.0 ;
      RECT  5215.0 167880.0 7582.5 167945.0 ;
      RECT  5390.0 168020.0 7772.5 168085.0 ;
      RECT  6615.0 168160.0 7962.5 168225.0 ;
      RECT  5215.0 169255.0 7582.5 169320.0 ;
      RECT  5390.0 169115.0 7772.5 169180.0 ;
      RECT  6790.0 168975.0 7962.5 169040.0 ;
      RECT  5215.0 170570.0 7582.5 170635.0 ;
      RECT  5390.0 170710.0 7772.5 170775.0 ;
      RECT  6965.0 170850.0 7962.5 170915.0 ;
      RECT  5215.0 171945.0 7582.5 172010.0 ;
      RECT  5390.0 171805.0 7772.5 171870.0 ;
      RECT  7140.0 171665.0 7962.5 171730.0 ;
      RECT  5215.0 173260.0 7582.5 173325.0 ;
      RECT  5390.0 173400.0 7772.5 173465.0 ;
      RECT  7315.0 173540.0 7962.5 173605.0 ;
      RECT  5215.0 174635.0 7582.5 174700.0 ;
      RECT  5565.0 174495.0 7772.5 174560.0 ;
      RECT  6090.0 174355.0 7962.5 174420.0 ;
      RECT  5215.0 175950.0 7582.5 176015.0 ;
      RECT  5565.0 176090.0 7772.5 176155.0 ;
      RECT  6265.0 176230.0 7962.5 176295.0 ;
      RECT  5215.0 177325.0 7582.5 177390.0 ;
      RECT  5565.0 177185.0 7772.5 177250.0 ;
      RECT  6440.0 177045.0 7962.5 177110.0 ;
      RECT  5215.0 178640.0 7582.5 178705.0 ;
      RECT  5565.0 178780.0 7772.5 178845.0 ;
      RECT  6615.0 178920.0 7962.5 178985.0 ;
      RECT  5215.0 180015.0 7582.5 180080.0 ;
      RECT  5565.0 179875.0 7772.5 179940.0 ;
      RECT  6790.0 179735.0 7962.5 179800.0 ;
      RECT  5215.0 181330.0 7582.5 181395.0 ;
      RECT  5565.0 181470.0 7772.5 181535.0 ;
      RECT  6965.0 181610.0 7962.5 181675.0 ;
      RECT  5215.0 182705.0 7582.5 182770.0 ;
      RECT  5565.0 182565.0 7772.5 182630.0 ;
      RECT  7140.0 182425.0 7962.5 182490.0 ;
      RECT  5215.0 184020.0 7582.5 184085.0 ;
      RECT  5565.0 184160.0 7772.5 184225.0 ;
      RECT  7315.0 184300.0 7962.5 184365.0 ;
      RECT  5215.0 185395.0 7582.5 185460.0 ;
      RECT  5740.0 185255.0 7772.5 185320.0 ;
      RECT  6090.0 185115.0 7962.5 185180.0 ;
      RECT  5215.0 186710.0 7582.5 186775.0 ;
      RECT  5740.0 186850.0 7772.5 186915.0 ;
      RECT  6265.0 186990.0 7962.5 187055.0 ;
      RECT  5215.0 188085.0 7582.5 188150.0 ;
      RECT  5740.0 187945.0 7772.5 188010.0 ;
      RECT  6440.0 187805.0 7962.5 187870.0 ;
      RECT  5215.0 189400.0 7582.5 189465.0 ;
      RECT  5740.0 189540.0 7772.5 189605.0 ;
      RECT  6615.0 189680.0 7962.5 189745.0 ;
      RECT  5215.0 190775.0 7582.5 190840.0 ;
      RECT  5740.0 190635.0 7772.5 190700.0 ;
      RECT  6790.0 190495.0 7962.5 190560.0 ;
      RECT  5215.0 192090.0 7582.5 192155.0 ;
      RECT  5740.0 192230.0 7772.5 192295.0 ;
      RECT  6965.0 192370.0 7962.5 192435.0 ;
      RECT  5215.0 193465.0 7582.5 193530.0 ;
      RECT  5740.0 193325.0 7772.5 193390.0 ;
      RECT  7140.0 193185.0 7962.5 193250.0 ;
      RECT  5215.0 194780.0 7582.5 194845.0 ;
      RECT  5740.0 194920.0 7772.5 194985.0 ;
      RECT  7315.0 195060.0 7962.5 195125.0 ;
      RECT  5215.0 196155.0 7582.5 196220.0 ;
      RECT  5915.0 196015.0 7772.5 196080.0 ;
      RECT  6090.0 195875.0 7962.5 195940.0 ;
      RECT  5215.0 197470.0 7582.5 197535.0 ;
      RECT  5915.0 197610.0 7772.5 197675.0 ;
      RECT  6265.0 197750.0 7962.5 197815.0 ;
      RECT  5215.0 198845.0 7582.5 198910.0 ;
      RECT  5915.0 198705.0 7772.5 198770.0 ;
      RECT  6440.0 198565.0 7962.5 198630.0 ;
      RECT  5215.0 200160.0 7582.5 200225.0 ;
      RECT  5915.0 200300.0 7772.5 200365.0 ;
      RECT  6615.0 200440.0 7962.5 200505.0 ;
      RECT  5215.0 201535.0 7582.5 201600.0 ;
      RECT  5915.0 201395.0 7772.5 201460.0 ;
      RECT  6790.0 201255.0 7962.5 201320.0 ;
      RECT  5215.0 202850.0 7582.5 202915.0 ;
      RECT  5915.0 202990.0 7772.5 203055.0 ;
      RECT  6965.0 203130.0 7962.5 203195.0 ;
      RECT  5215.0 204225.0 7582.5 204290.0 ;
      RECT  5915.0 204085.0 7772.5 204150.0 ;
      RECT  7140.0 203945.0 7962.5 204010.0 ;
      RECT  5215.0 205540.0 7582.5 205605.0 ;
      RECT  5915.0 205680.0 7772.5 205745.0 ;
      RECT  7315.0 205820.0 7962.5 205885.0 ;
      RECT  10277.5 13175.0 10212.5 13240.0 ;
      RECT  10277.5 13697.5 10212.5 13762.5 ;
      RECT  10515.0 13175.0 10245.0 13240.0 ;
      RECT  10277.5 13207.5 10212.5 13730.0 ;
      RECT  10245.0 13697.5 10000.0 13762.5 ;
      RECT  11385.0 13175.0 10745.0 13240.0 ;
      RECT  10277.5 14610.0 10212.5 14675.0 ;
      RECT  10277.5 15042.5 10212.5 15107.5 ;
      RECT  10515.0 14610.0 10245.0 14675.0 ;
      RECT  10277.5 14642.5 10212.5 15075.0 ;
      RECT  10245.0 15042.5 9725.0 15107.5 ;
      RECT  11110.0 14610.0 10745.0 14675.0 ;
      RECT  11385.0 15372.5 9450.0 15437.5 ;
      RECT  11110.0 16717.5 9175.0 16782.5 ;
      RECT  10000.0 13187.5 8875.0 13252.5 ;
      RECT  9725.0 12972.5 8617.5 13037.5 ;
      RECT  9450.0 14597.5 8875.0 14662.5 ;
      RECT  9725.0 14812.5 8617.5 14877.5 ;
      RECT  10000.0 15877.5 8875.0 15942.5 ;
      RECT  9175.0 15662.5 8617.5 15727.5 ;
      RECT  9450.0 17287.5 8875.0 17352.5 ;
      RECT  9175.0 17502.5 8617.5 17567.5 ;
      RECT  8170.0 13187.5 8105.0 13252.5 ;
      RECT  8170.0 13175.0 8105.0 13240.0 ;
      RECT  8387.5 13187.5 8137.5 13252.5 ;
      RECT  8170.0 13207.5 8105.0 13220.0 ;
      RECT  8137.5 13175.0 7890.0 13240.0 ;
      RECT  8170.0 14597.5 8105.0 14662.5 ;
      RECT  8170.0 14610.0 8105.0 14675.0 ;
      RECT  8387.5 14597.5 8137.5 14662.5 ;
      RECT  8170.0 14630.0 8105.0 14642.5 ;
      RECT  8137.5 14610.0 7890.0 14675.0 ;
      RECT  8170.0 15877.5 8105.0 15942.5 ;
      RECT  8170.0 15865.0 8105.0 15930.0 ;
      RECT  8387.5 15877.5 8137.5 15942.5 ;
      RECT  8170.0 15897.5 8105.0 15910.0 ;
      RECT  8137.5 15865.0 7890.0 15930.0 ;
      RECT  8170.0 17287.5 8105.0 17352.5 ;
      RECT  8170.0 17300.0 8105.0 17365.0 ;
      RECT  8387.5 17287.5 8137.5 17352.5 ;
      RECT  8170.0 17320.0 8105.0 17332.5 ;
      RECT  8137.5 17300.0 7890.0 17365.0 ;
      RECT  10442.5 13740.0 10377.5 13925.0 ;
      RECT  10442.5 12580.0 10377.5 12765.0 ;
      RECT  10802.5 12697.5 10737.5 12547.5 ;
      RECT  10802.5 13582.5 10737.5 13957.5 ;
      RECT  10612.5 12697.5 10547.5 13582.5 ;
      RECT  10802.5 13582.5 10737.5 13717.5 ;
      RECT  10612.5 13582.5 10547.5 13717.5 ;
      RECT  10612.5 13582.5 10547.5 13717.5 ;
      RECT  10802.5 13582.5 10737.5 13717.5 ;
      RECT  10802.5 12697.5 10737.5 12832.5 ;
      RECT  10612.5 12697.5 10547.5 12832.5 ;
      RECT  10612.5 12697.5 10547.5 12832.5 ;
      RECT  10802.5 12697.5 10737.5 12832.5 ;
      RECT  10442.5 13672.5 10377.5 13807.5 ;
      RECT  10442.5 12697.5 10377.5 12832.5 ;
      RECT  10745.0 13140.0 10680.0 13275.0 ;
      RECT  10745.0 13140.0 10680.0 13275.0 ;
      RECT  10580.0 13175.0 10515.0 13240.0 ;
      RECT  10870.0 13892.5 10310.0 13957.5 ;
      RECT  10870.0 12547.5 10310.0 12612.5 ;
      RECT  10442.5 14110.0 10377.5 13925.0 ;
      RECT  10442.5 15270.0 10377.5 15085.0 ;
      RECT  10802.5 15152.5 10737.5 15302.5 ;
      RECT  10802.5 14267.5 10737.5 13892.5 ;
      RECT  10612.5 15152.5 10547.5 14267.5 ;
      RECT  10802.5 14267.5 10737.5 14132.5 ;
      RECT  10612.5 14267.5 10547.5 14132.5 ;
      RECT  10612.5 14267.5 10547.5 14132.5 ;
      RECT  10802.5 14267.5 10737.5 14132.5 ;
      RECT  10802.5 15152.5 10737.5 15017.5 ;
      RECT  10612.5 15152.5 10547.5 15017.5 ;
      RECT  10612.5 15152.5 10547.5 15017.5 ;
      RECT  10802.5 15152.5 10737.5 15017.5 ;
      RECT  10442.5 14177.5 10377.5 14042.5 ;
      RECT  10442.5 15152.5 10377.5 15017.5 ;
      RECT  10745.0 14710.0 10680.0 14575.0 ;
      RECT  10745.0 14710.0 10680.0 14575.0 ;
      RECT  10580.0 14675.0 10515.0 14610.0 ;
      RECT  10870.0 13957.5 10310.0 13892.5 ;
      RECT  10870.0 15302.5 10310.0 15237.5 ;
      RECT  7587.5 13740.0 7522.5 13925.0 ;
      RECT  7587.5 12580.0 7522.5 12765.0 ;
      RECT  7947.5 12697.5 7882.5 12547.5 ;
      RECT  7947.5 13582.5 7882.5 13957.5 ;
      RECT  7757.5 12697.5 7692.5 13582.5 ;
      RECT  7947.5 13582.5 7882.5 13717.5 ;
      RECT  7757.5 13582.5 7692.5 13717.5 ;
      RECT  7757.5 13582.5 7692.5 13717.5 ;
      RECT  7947.5 13582.5 7882.5 13717.5 ;
      RECT  7947.5 12697.5 7882.5 12832.5 ;
      RECT  7757.5 12697.5 7692.5 12832.5 ;
      RECT  7757.5 12697.5 7692.5 12832.5 ;
      RECT  7947.5 12697.5 7882.5 12832.5 ;
      RECT  7587.5 13672.5 7522.5 13807.5 ;
      RECT  7587.5 12697.5 7522.5 12832.5 ;
      RECT  7890.0 13140.0 7825.0 13275.0 ;
      RECT  7890.0 13140.0 7825.0 13275.0 ;
      RECT  7725.0 13175.0 7660.0 13240.0 ;
      RECT  8015.0 13892.5 7455.0 13957.5 ;
      RECT  8015.0 12547.5 7455.0 12612.5 ;
      RECT  7587.5 14110.0 7522.5 13925.0 ;
      RECT  7587.5 15270.0 7522.5 15085.0 ;
      RECT  7947.5 15152.5 7882.5 15302.5 ;
      RECT  7947.5 14267.5 7882.5 13892.5 ;
      RECT  7757.5 15152.5 7692.5 14267.5 ;
      RECT  7947.5 14267.5 7882.5 14132.5 ;
      RECT  7757.5 14267.5 7692.5 14132.5 ;
      RECT  7757.5 14267.5 7692.5 14132.5 ;
      RECT  7947.5 14267.5 7882.5 14132.5 ;
      RECT  7947.5 15152.5 7882.5 15017.5 ;
      RECT  7757.5 15152.5 7692.5 15017.5 ;
      RECT  7757.5 15152.5 7692.5 15017.5 ;
      RECT  7947.5 15152.5 7882.5 15017.5 ;
      RECT  7587.5 14177.5 7522.5 14042.5 ;
      RECT  7587.5 15152.5 7522.5 15017.5 ;
      RECT  7890.0 14710.0 7825.0 14575.0 ;
      RECT  7890.0 14710.0 7825.0 14575.0 ;
      RECT  7725.0 14675.0 7660.0 14610.0 ;
      RECT  8015.0 13957.5 7455.0 13892.5 ;
      RECT  8015.0 15302.5 7455.0 15237.5 ;
      RECT  7587.5 16430.0 7522.5 16615.0 ;
      RECT  7587.5 15270.0 7522.5 15455.0 ;
      RECT  7947.5 15387.5 7882.5 15237.5 ;
      RECT  7947.5 16272.5 7882.5 16647.5 ;
      RECT  7757.5 15387.5 7692.5 16272.5 ;
      RECT  7947.5 16272.5 7882.5 16407.5 ;
      RECT  7757.5 16272.5 7692.5 16407.5 ;
      RECT  7757.5 16272.5 7692.5 16407.5 ;
      RECT  7947.5 16272.5 7882.5 16407.5 ;
      RECT  7947.5 15387.5 7882.5 15522.5 ;
      RECT  7757.5 15387.5 7692.5 15522.5 ;
      RECT  7757.5 15387.5 7692.5 15522.5 ;
      RECT  7947.5 15387.5 7882.5 15522.5 ;
      RECT  7587.5 16362.5 7522.5 16497.5 ;
      RECT  7587.5 15387.5 7522.5 15522.5 ;
      RECT  7890.0 15830.0 7825.0 15965.0 ;
      RECT  7890.0 15830.0 7825.0 15965.0 ;
      RECT  7725.0 15865.0 7660.0 15930.0 ;
      RECT  8015.0 16582.5 7455.0 16647.5 ;
      RECT  8015.0 15237.5 7455.0 15302.5 ;
      RECT  7587.5 16800.0 7522.5 16615.0 ;
      RECT  7587.5 17960.0 7522.5 17775.0 ;
      RECT  7947.5 17842.5 7882.5 17992.5 ;
      RECT  7947.5 16957.5 7882.5 16582.5 ;
      RECT  7757.5 17842.5 7692.5 16957.5 ;
      RECT  7947.5 16957.5 7882.5 16822.5 ;
      RECT  7757.5 16957.5 7692.5 16822.5 ;
      RECT  7757.5 16957.5 7692.5 16822.5 ;
      RECT  7947.5 16957.5 7882.5 16822.5 ;
      RECT  7947.5 17842.5 7882.5 17707.5 ;
      RECT  7757.5 17842.5 7692.5 17707.5 ;
      RECT  7757.5 17842.5 7692.5 17707.5 ;
      RECT  7947.5 17842.5 7882.5 17707.5 ;
      RECT  7587.5 16867.5 7522.5 16732.5 ;
      RECT  7587.5 17842.5 7522.5 17707.5 ;
      RECT  7890.0 17400.0 7825.0 17265.0 ;
      RECT  7890.0 17400.0 7825.0 17265.0 ;
      RECT  7725.0 17365.0 7660.0 17300.0 ;
      RECT  8015.0 16647.5 7455.0 16582.5 ;
      RECT  8015.0 17992.5 7455.0 17927.5 ;
      RECT  8867.5 12742.5 8802.5 12547.5 ;
      RECT  8867.5 13582.5 8802.5 13957.5 ;
      RECT  8487.5 13582.5 8422.5 13957.5 ;
      RECT  8317.5 13740.0 8252.5 13925.0 ;
      RECT  8317.5 12580.0 8252.5 12765.0 ;
      RECT  8867.5 13582.5 8802.5 13717.5 ;
      RECT  8677.5 13582.5 8612.5 13717.5 ;
      RECT  8677.5 13582.5 8612.5 13717.5 ;
      RECT  8867.5 13582.5 8802.5 13717.5 ;
      RECT  8677.5 13582.5 8612.5 13717.5 ;
      RECT  8487.5 13582.5 8422.5 13717.5 ;
      RECT  8487.5 13582.5 8422.5 13717.5 ;
      RECT  8677.5 13582.5 8612.5 13717.5 ;
      RECT  8867.5 12742.5 8802.5 12877.5 ;
      RECT  8677.5 12742.5 8612.5 12877.5 ;
      RECT  8677.5 12742.5 8612.5 12877.5 ;
      RECT  8867.5 12742.5 8802.5 12877.5 ;
      RECT  8677.5 12742.5 8612.5 12877.5 ;
      RECT  8487.5 12742.5 8422.5 12877.5 ;
      RECT  8487.5 12742.5 8422.5 12877.5 ;
      RECT  8677.5 12742.5 8612.5 12877.5 ;
      RECT  8317.5 13672.5 8252.5 13807.5 ;
      RECT  8317.5 12697.5 8252.5 12832.5 ;
      RECT  8482.5 12972.5 8617.5 13037.5 ;
      RECT  8740.0 13187.5 8875.0 13252.5 ;
      RECT  8677.5 13582.5 8612.5 13717.5 ;
      RECT  8487.5 12742.5 8422.5 12877.5 ;
      RECT  8387.5 13187.5 8522.5 13252.5 ;
      RECT  8875.0 13187.5 8740.0 13252.5 ;
      RECT  8617.5 12972.5 8482.5 13037.5 ;
      RECT  8522.5 13187.5 8387.5 13252.5 ;
      RECT  8935.0 13892.5 8015.0 13957.5 ;
      RECT  8935.0 12547.5 8015.0 12612.5 ;
      RECT  8867.5 15107.5 8802.5 15302.5 ;
      RECT  8867.5 14267.5 8802.5 13892.5 ;
      RECT  8487.5 14267.5 8422.5 13892.5 ;
      RECT  8317.5 14110.0 8252.5 13925.0 ;
      RECT  8317.5 15270.0 8252.5 15085.0 ;
      RECT  8867.5 14267.5 8802.5 14132.5 ;
      RECT  8677.5 14267.5 8612.5 14132.5 ;
      RECT  8677.5 14267.5 8612.5 14132.5 ;
      RECT  8867.5 14267.5 8802.5 14132.5 ;
      RECT  8677.5 14267.5 8612.5 14132.5 ;
      RECT  8487.5 14267.5 8422.5 14132.5 ;
      RECT  8487.5 14267.5 8422.5 14132.5 ;
      RECT  8677.5 14267.5 8612.5 14132.5 ;
      RECT  8867.5 15107.5 8802.5 14972.5 ;
      RECT  8677.5 15107.5 8612.5 14972.5 ;
      RECT  8677.5 15107.5 8612.5 14972.5 ;
      RECT  8867.5 15107.5 8802.5 14972.5 ;
      RECT  8677.5 15107.5 8612.5 14972.5 ;
      RECT  8487.5 15107.5 8422.5 14972.5 ;
      RECT  8487.5 15107.5 8422.5 14972.5 ;
      RECT  8677.5 15107.5 8612.5 14972.5 ;
      RECT  8317.5 14177.5 8252.5 14042.5 ;
      RECT  8317.5 15152.5 8252.5 15017.5 ;
      RECT  8482.5 14877.5 8617.5 14812.5 ;
      RECT  8740.0 14662.5 8875.0 14597.5 ;
      RECT  8677.5 14267.5 8612.5 14132.5 ;
      RECT  8487.5 15107.5 8422.5 14972.5 ;
      RECT  8387.5 14662.5 8522.5 14597.5 ;
      RECT  8875.0 14662.5 8740.0 14597.5 ;
      RECT  8617.5 14877.5 8482.5 14812.5 ;
      RECT  8522.5 14662.5 8387.5 14597.5 ;
      RECT  8935.0 13957.5 8015.0 13892.5 ;
      RECT  8935.0 15302.5 8015.0 15237.5 ;
      RECT  8867.5 15432.5 8802.5 15237.5 ;
      RECT  8867.5 16272.5 8802.5 16647.5 ;
      RECT  8487.5 16272.5 8422.5 16647.5 ;
      RECT  8317.5 16430.0 8252.5 16615.0 ;
      RECT  8317.5 15270.0 8252.5 15455.0 ;
      RECT  8867.5 16272.5 8802.5 16407.5 ;
      RECT  8677.5 16272.5 8612.5 16407.5 ;
      RECT  8677.5 16272.5 8612.5 16407.5 ;
      RECT  8867.5 16272.5 8802.5 16407.5 ;
      RECT  8677.5 16272.5 8612.5 16407.5 ;
      RECT  8487.5 16272.5 8422.5 16407.5 ;
      RECT  8487.5 16272.5 8422.5 16407.5 ;
      RECT  8677.5 16272.5 8612.5 16407.5 ;
      RECT  8867.5 15432.5 8802.5 15567.5 ;
      RECT  8677.5 15432.5 8612.5 15567.5 ;
      RECT  8677.5 15432.5 8612.5 15567.5 ;
      RECT  8867.5 15432.5 8802.5 15567.5 ;
      RECT  8677.5 15432.5 8612.5 15567.5 ;
      RECT  8487.5 15432.5 8422.5 15567.5 ;
      RECT  8487.5 15432.5 8422.5 15567.5 ;
      RECT  8677.5 15432.5 8612.5 15567.5 ;
      RECT  8317.5 16362.5 8252.5 16497.5 ;
      RECT  8317.5 15387.5 8252.5 15522.5 ;
      RECT  8482.5 15662.5 8617.5 15727.5 ;
      RECT  8740.0 15877.5 8875.0 15942.5 ;
      RECT  8677.5 16272.5 8612.5 16407.5 ;
      RECT  8487.5 15432.5 8422.5 15567.5 ;
      RECT  8387.5 15877.5 8522.5 15942.5 ;
      RECT  8875.0 15877.5 8740.0 15942.5 ;
      RECT  8617.5 15662.5 8482.5 15727.5 ;
      RECT  8522.5 15877.5 8387.5 15942.5 ;
      RECT  8935.0 16582.5 8015.0 16647.5 ;
      RECT  8935.0 15237.5 8015.0 15302.5 ;
      RECT  8867.5 17797.5 8802.5 17992.5 ;
      RECT  8867.5 16957.5 8802.5 16582.5 ;
      RECT  8487.5 16957.5 8422.5 16582.5 ;
      RECT  8317.5 16800.0 8252.5 16615.0 ;
      RECT  8317.5 17960.0 8252.5 17775.0 ;
      RECT  8867.5 16957.5 8802.5 16822.5 ;
      RECT  8677.5 16957.5 8612.5 16822.5 ;
      RECT  8677.5 16957.5 8612.5 16822.5 ;
      RECT  8867.5 16957.5 8802.5 16822.5 ;
      RECT  8677.5 16957.5 8612.5 16822.5 ;
      RECT  8487.5 16957.5 8422.5 16822.5 ;
      RECT  8487.5 16957.5 8422.5 16822.5 ;
      RECT  8677.5 16957.5 8612.5 16822.5 ;
      RECT  8867.5 17797.5 8802.5 17662.5 ;
      RECT  8677.5 17797.5 8612.5 17662.5 ;
      RECT  8677.5 17797.5 8612.5 17662.5 ;
      RECT  8867.5 17797.5 8802.5 17662.5 ;
      RECT  8677.5 17797.5 8612.5 17662.5 ;
      RECT  8487.5 17797.5 8422.5 17662.5 ;
      RECT  8487.5 17797.5 8422.5 17662.5 ;
      RECT  8677.5 17797.5 8612.5 17662.5 ;
      RECT  8317.5 16867.5 8252.5 16732.5 ;
      RECT  8317.5 17842.5 8252.5 17707.5 ;
      RECT  8482.5 17567.5 8617.5 17502.5 ;
      RECT  8740.0 17352.5 8875.0 17287.5 ;
      RECT  8677.5 16957.5 8612.5 16822.5 ;
      RECT  8487.5 17797.5 8422.5 17662.5 ;
      RECT  8387.5 17352.5 8522.5 17287.5 ;
      RECT  8875.0 17352.5 8740.0 17287.5 ;
      RECT  8617.5 17567.5 8482.5 17502.5 ;
      RECT  8522.5 17352.5 8387.5 17287.5 ;
      RECT  8935.0 16647.5 8015.0 16582.5 ;
      RECT  8935.0 17992.5 8015.0 17927.5 ;
      RECT  9932.5 13697.5 10067.5 13762.5 ;
      RECT  11317.5 13175.0 11452.5 13240.0 ;
      RECT  9657.5 15042.5 9792.5 15107.5 ;
      RECT  11042.5 14610.0 11177.5 14675.0 ;
      RECT  11317.5 15372.5 11452.5 15437.5 ;
      RECT  9382.5 15372.5 9517.5 15437.5 ;
      RECT  11042.5 16717.5 11177.5 16782.5 ;
      RECT  9107.5 16717.5 9242.5 16782.5 ;
      RECT  9932.5 13187.5 10067.5 13252.5 ;
      RECT  9657.5 12972.5 9792.5 13037.5 ;
      RECT  9382.5 14597.5 9517.5 14662.5 ;
      RECT  9657.5 14812.5 9792.5 14877.5 ;
      RECT  9932.5 15877.5 10067.5 15942.5 ;
      RECT  9107.5 15662.5 9242.5 15727.5 ;
      RECT  9382.5 17287.5 9517.5 17352.5 ;
      RECT  9107.5 17502.5 9242.5 17567.5 ;
      RECT  7660.0 13175.0 7455.0 13240.0 ;
      RECT  7660.0 14610.0 7455.0 14675.0 ;
      RECT  7660.0 15865.0 7455.0 15930.0 ;
      RECT  7660.0 17300.0 7455.0 17365.0 ;
      RECT  11420.0 13892.5 7455.0 13957.5 ;
      RECT  11420.0 16582.5 7455.0 16647.5 ;
      RECT  11420.0 12547.5 7455.0 12612.5 ;
      RECT  11420.0 15237.5 7455.0 15302.5 ;
      RECT  11420.0 17927.5 7455.0 17992.5 ;
      RECT  10277.5 18555.0 10212.5 18620.0 ;
      RECT  10277.5 19077.5 10212.5 19142.5 ;
      RECT  10515.0 18555.0 10245.0 18620.0 ;
      RECT  10277.5 18587.5 10212.5 19110.0 ;
      RECT  10245.0 19077.5 10000.0 19142.5 ;
      RECT  11385.0 18555.0 10745.0 18620.0 ;
      RECT  10277.5 19990.0 10212.5 20055.0 ;
      RECT  10277.5 20422.5 10212.5 20487.5 ;
      RECT  10515.0 19990.0 10245.0 20055.0 ;
      RECT  10277.5 20022.5 10212.5 20455.0 ;
      RECT  10245.0 20422.5 9725.0 20487.5 ;
      RECT  11110.0 19990.0 10745.0 20055.0 ;
      RECT  11385.0 20752.5 9450.0 20817.5 ;
      RECT  11110.0 22097.5 9175.0 22162.5 ;
      RECT  10000.0 18567.5 8875.0 18632.5 ;
      RECT  9725.0 18352.5 8617.5 18417.5 ;
      RECT  9450.0 19977.5 8875.0 20042.5 ;
      RECT  9725.0 20192.5 8617.5 20257.5 ;
      RECT  10000.0 21257.5 8875.0 21322.5 ;
      RECT  9175.0 21042.5 8617.5 21107.5 ;
      RECT  9450.0 22667.5 8875.0 22732.5 ;
      RECT  9175.0 22882.5 8617.5 22947.5 ;
      RECT  8170.0 18567.5 8105.0 18632.5 ;
      RECT  8170.0 18555.0 8105.0 18620.0 ;
      RECT  8387.5 18567.5 8137.5 18632.5 ;
      RECT  8170.0 18587.5 8105.0 18600.0 ;
      RECT  8137.5 18555.0 7890.0 18620.0 ;
      RECT  8170.0 19977.5 8105.0 20042.5 ;
      RECT  8170.0 19990.0 8105.0 20055.0 ;
      RECT  8387.5 19977.5 8137.5 20042.5 ;
      RECT  8170.0 20010.0 8105.0 20022.5 ;
      RECT  8137.5 19990.0 7890.0 20055.0 ;
      RECT  8170.0 21257.5 8105.0 21322.5 ;
      RECT  8170.0 21245.0 8105.0 21310.0 ;
      RECT  8387.5 21257.5 8137.5 21322.5 ;
      RECT  8170.0 21277.5 8105.0 21290.0 ;
      RECT  8137.5 21245.0 7890.0 21310.0 ;
      RECT  8170.0 22667.5 8105.0 22732.5 ;
      RECT  8170.0 22680.0 8105.0 22745.0 ;
      RECT  8387.5 22667.5 8137.5 22732.5 ;
      RECT  8170.0 22700.0 8105.0 22712.5 ;
      RECT  8137.5 22680.0 7890.0 22745.0 ;
      RECT  10442.5 19120.0 10377.5 19305.0 ;
      RECT  10442.5 17960.0 10377.5 18145.0 ;
      RECT  10802.5 18077.5 10737.5 17927.5 ;
      RECT  10802.5 18962.5 10737.5 19337.5 ;
      RECT  10612.5 18077.5 10547.5 18962.5 ;
      RECT  10802.5 18962.5 10737.5 19097.5 ;
      RECT  10612.5 18962.5 10547.5 19097.5 ;
      RECT  10612.5 18962.5 10547.5 19097.5 ;
      RECT  10802.5 18962.5 10737.5 19097.5 ;
      RECT  10802.5 18077.5 10737.5 18212.5 ;
      RECT  10612.5 18077.5 10547.5 18212.5 ;
      RECT  10612.5 18077.5 10547.5 18212.5 ;
      RECT  10802.5 18077.5 10737.5 18212.5 ;
      RECT  10442.5 19052.5 10377.5 19187.5 ;
      RECT  10442.5 18077.5 10377.5 18212.5 ;
      RECT  10745.0 18520.0 10680.0 18655.0 ;
      RECT  10745.0 18520.0 10680.0 18655.0 ;
      RECT  10580.0 18555.0 10515.0 18620.0 ;
      RECT  10870.0 19272.5 10310.0 19337.5 ;
      RECT  10870.0 17927.5 10310.0 17992.5 ;
      RECT  10442.5 19490.0 10377.5 19305.0 ;
      RECT  10442.5 20650.0 10377.5 20465.0 ;
      RECT  10802.5 20532.5 10737.5 20682.5 ;
      RECT  10802.5 19647.5 10737.5 19272.5 ;
      RECT  10612.5 20532.5 10547.5 19647.5 ;
      RECT  10802.5 19647.5 10737.5 19512.5 ;
      RECT  10612.5 19647.5 10547.5 19512.5 ;
      RECT  10612.5 19647.5 10547.5 19512.5 ;
      RECT  10802.5 19647.5 10737.5 19512.5 ;
      RECT  10802.5 20532.5 10737.5 20397.5 ;
      RECT  10612.5 20532.5 10547.5 20397.5 ;
      RECT  10612.5 20532.5 10547.5 20397.5 ;
      RECT  10802.5 20532.5 10737.5 20397.5 ;
      RECT  10442.5 19557.5 10377.5 19422.5 ;
      RECT  10442.5 20532.5 10377.5 20397.5 ;
      RECT  10745.0 20090.0 10680.0 19955.0 ;
      RECT  10745.0 20090.0 10680.0 19955.0 ;
      RECT  10580.0 20055.0 10515.0 19990.0 ;
      RECT  10870.0 19337.5 10310.0 19272.5 ;
      RECT  10870.0 20682.5 10310.0 20617.5 ;
      RECT  7587.5 19120.0 7522.5 19305.0 ;
      RECT  7587.5 17960.0 7522.5 18145.0 ;
      RECT  7947.5 18077.5 7882.5 17927.5 ;
      RECT  7947.5 18962.5 7882.5 19337.5 ;
      RECT  7757.5 18077.5 7692.5 18962.5 ;
      RECT  7947.5 18962.5 7882.5 19097.5 ;
      RECT  7757.5 18962.5 7692.5 19097.5 ;
      RECT  7757.5 18962.5 7692.5 19097.5 ;
      RECT  7947.5 18962.5 7882.5 19097.5 ;
      RECT  7947.5 18077.5 7882.5 18212.5 ;
      RECT  7757.5 18077.5 7692.5 18212.5 ;
      RECT  7757.5 18077.5 7692.5 18212.5 ;
      RECT  7947.5 18077.5 7882.5 18212.5 ;
      RECT  7587.5 19052.5 7522.5 19187.5 ;
      RECT  7587.5 18077.5 7522.5 18212.5 ;
      RECT  7890.0 18520.0 7825.0 18655.0 ;
      RECT  7890.0 18520.0 7825.0 18655.0 ;
      RECT  7725.0 18555.0 7660.0 18620.0 ;
      RECT  8015.0 19272.5 7455.0 19337.5 ;
      RECT  8015.0 17927.5 7455.0 17992.5 ;
      RECT  7587.5 19490.0 7522.5 19305.0 ;
      RECT  7587.5 20650.0 7522.5 20465.0 ;
      RECT  7947.5 20532.5 7882.5 20682.5 ;
      RECT  7947.5 19647.5 7882.5 19272.5 ;
      RECT  7757.5 20532.5 7692.5 19647.5 ;
      RECT  7947.5 19647.5 7882.5 19512.5 ;
      RECT  7757.5 19647.5 7692.5 19512.5 ;
      RECT  7757.5 19647.5 7692.5 19512.5 ;
      RECT  7947.5 19647.5 7882.5 19512.5 ;
      RECT  7947.5 20532.5 7882.5 20397.5 ;
      RECT  7757.5 20532.5 7692.5 20397.5 ;
      RECT  7757.5 20532.5 7692.5 20397.5 ;
      RECT  7947.5 20532.5 7882.5 20397.5 ;
      RECT  7587.5 19557.5 7522.5 19422.5 ;
      RECT  7587.5 20532.5 7522.5 20397.5 ;
      RECT  7890.0 20090.0 7825.0 19955.0 ;
      RECT  7890.0 20090.0 7825.0 19955.0 ;
      RECT  7725.0 20055.0 7660.0 19990.0 ;
      RECT  8015.0 19337.5 7455.0 19272.5 ;
      RECT  8015.0 20682.5 7455.0 20617.5 ;
      RECT  7587.5 21810.0 7522.5 21995.0 ;
      RECT  7587.5 20650.0 7522.5 20835.0 ;
      RECT  7947.5 20767.5 7882.5 20617.5 ;
      RECT  7947.5 21652.5 7882.5 22027.5 ;
      RECT  7757.5 20767.5 7692.5 21652.5 ;
      RECT  7947.5 21652.5 7882.5 21787.5 ;
      RECT  7757.5 21652.5 7692.5 21787.5 ;
      RECT  7757.5 21652.5 7692.5 21787.5 ;
      RECT  7947.5 21652.5 7882.5 21787.5 ;
      RECT  7947.5 20767.5 7882.5 20902.5 ;
      RECT  7757.5 20767.5 7692.5 20902.5 ;
      RECT  7757.5 20767.5 7692.5 20902.5 ;
      RECT  7947.5 20767.5 7882.5 20902.5 ;
      RECT  7587.5 21742.5 7522.5 21877.5 ;
      RECT  7587.5 20767.5 7522.5 20902.5 ;
      RECT  7890.0 21210.0 7825.0 21345.0 ;
      RECT  7890.0 21210.0 7825.0 21345.0 ;
      RECT  7725.0 21245.0 7660.0 21310.0 ;
      RECT  8015.0 21962.5 7455.0 22027.5 ;
      RECT  8015.0 20617.5 7455.0 20682.5 ;
      RECT  7587.5 22180.0 7522.5 21995.0 ;
      RECT  7587.5 23340.0 7522.5 23155.0 ;
      RECT  7947.5 23222.5 7882.5 23372.5 ;
      RECT  7947.5 22337.5 7882.5 21962.5 ;
      RECT  7757.5 23222.5 7692.5 22337.5 ;
      RECT  7947.5 22337.5 7882.5 22202.5 ;
      RECT  7757.5 22337.5 7692.5 22202.5 ;
      RECT  7757.5 22337.5 7692.5 22202.5 ;
      RECT  7947.5 22337.5 7882.5 22202.5 ;
      RECT  7947.5 23222.5 7882.5 23087.5 ;
      RECT  7757.5 23222.5 7692.5 23087.5 ;
      RECT  7757.5 23222.5 7692.5 23087.5 ;
      RECT  7947.5 23222.5 7882.5 23087.5 ;
      RECT  7587.5 22247.5 7522.5 22112.5 ;
      RECT  7587.5 23222.5 7522.5 23087.5 ;
      RECT  7890.0 22780.0 7825.0 22645.0 ;
      RECT  7890.0 22780.0 7825.0 22645.0 ;
      RECT  7725.0 22745.0 7660.0 22680.0 ;
      RECT  8015.0 22027.5 7455.0 21962.5 ;
      RECT  8015.0 23372.5 7455.0 23307.5 ;
      RECT  8867.5 18122.5 8802.5 17927.5 ;
      RECT  8867.5 18962.5 8802.5 19337.5 ;
      RECT  8487.5 18962.5 8422.5 19337.5 ;
      RECT  8317.5 19120.0 8252.5 19305.0 ;
      RECT  8317.5 17960.0 8252.5 18145.0 ;
      RECT  8867.5 18962.5 8802.5 19097.5 ;
      RECT  8677.5 18962.5 8612.5 19097.5 ;
      RECT  8677.5 18962.5 8612.5 19097.5 ;
      RECT  8867.5 18962.5 8802.5 19097.5 ;
      RECT  8677.5 18962.5 8612.5 19097.5 ;
      RECT  8487.5 18962.5 8422.5 19097.5 ;
      RECT  8487.5 18962.5 8422.5 19097.5 ;
      RECT  8677.5 18962.5 8612.5 19097.5 ;
      RECT  8867.5 18122.5 8802.5 18257.5 ;
      RECT  8677.5 18122.5 8612.5 18257.5 ;
      RECT  8677.5 18122.5 8612.5 18257.5 ;
      RECT  8867.5 18122.5 8802.5 18257.5 ;
      RECT  8677.5 18122.5 8612.5 18257.5 ;
      RECT  8487.5 18122.5 8422.5 18257.5 ;
      RECT  8487.5 18122.5 8422.5 18257.5 ;
      RECT  8677.5 18122.5 8612.5 18257.5 ;
      RECT  8317.5 19052.5 8252.5 19187.5 ;
      RECT  8317.5 18077.5 8252.5 18212.5 ;
      RECT  8482.5 18352.5 8617.5 18417.5 ;
      RECT  8740.0 18567.5 8875.0 18632.5 ;
      RECT  8677.5 18962.5 8612.5 19097.5 ;
      RECT  8487.5 18122.5 8422.5 18257.5 ;
      RECT  8387.5 18567.5 8522.5 18632.5 ;
      RECT  8875.0 18567.5 8740.0 18632.5 ;
      RECT  8617.5 18352.5 8482.5 18417.5 ;
      RECT  8522.5 18567.5 8387.5 18632.5 ;
      RECT  8935.0 19272.5 8015.0 19337.5 ;
      RECT  8935.0 17927.5 8015.0 17992.5 ;
      RECT  8867.5 20487.5 8802.5 20682.5 ;
      RECT  8867.5 19647.5 8802.5 19272.5 ;
      RECT  8487.5 19647.5 8422.5 19272.5 ;
      RECT  8317.5 19490.0 8252.5 19305.0 ;
      RECT  8317.5 20650.0 8252.5 20465.0 ;
      RECT  8867.5 19647.5 8802.5 19512.5 ;
      RECT  8677.5 19647.5 8612.5 19512.5 ;
      RECT  8677.5 19647.5 8612.5 19512.5 ;
      RECT  8867.5 19647.5 8802.5 19512.5 ;
      RECT  8677.5 19647.5 8612.5 19512.5 ;
      RECT  8487.5 19647.5 8422.5 19512.5 ;
      RECT  8487.5 19647.5 8422.5 19512.5 ;
      RECT  8677.5 19647.5 8612.5 19512.5 ;
      RECT  8867.5 20487.5 8802.5 20352.5 ;
      RECT  8677.5 20487.5 8612.5 20352.5 ;
      RECT  8677.5 20487.5 8612.5 20352.5 ;
      RECT  8867.5 20487.5 8802.5 20352.5 ;
      RECT  8677.5 20487.5 8612.5 20352.5 ;
      RECT  8487.5 20487.5 8422.5 20352.5 ;
      RECT  8487.5 20487.5 8422.5 20352.5 ;
      RECT  8677.5 20487.5 8612.5 20352.5 ;
      RECT  8317.5 19557.5 8252.5 19422.5 ;
      RECT  8317.5 20532.5 8252.5 20397.5 ;
      RECT  8482.5 20257.5 8617.5 20192.5 ;
      RECT  8740.0 20042.5 8875.0 19977.5 ;
      RECT  8677.5 19647.5 8612.5 19512.5 ;
      RECT  8487.5 20487.5 8422.5 20352.5 ;
      RECT  8387.5 20042.5 8522.5 19977.5 ;
      RECT  8875.0 20042.5 8740.0 19977.5 ;
      RECT  8617.5 20257.5 8482.5 20192.5 ;
      RECT  8522.5 20042.5 8387.5 19977.5 ;
      RECT  8935.0 19337.5 8015.0 19272.5 ;
      RECT  8935.0 20682.5 8015.0 20617.5 ;
      RECT  8867.5 20812.5 8802.5 20617.5 ;
      RECT  8867.5 21652.5 8802.5 22027.5 ;
      RECT  8487.5 21652.5 8422.5 22027.5 ;
      RECT  8317.5 21810.0 8252.5 21995.0 ;
      RECT  8317.5 20650.0 8252.5 20835.0 ;
      RECT  8867.5 21652.5 8802.5 21787.5 ;
      RECT  8677.5 21652.5 8612.5 21787.5 ;
      RECT  8677.5 21652.5 8612.5 21787.5 ;
      RECT  8867.5 21652.5 8802.5 21787.5 ;
      RECT  8677.5 21652.5 8612.5 21787.5 ;
      RECT  8487.5 21652.5 8422.5 21787.5 ;
      RECT  8487.5 21652.5 8422.5 21787.5 ;
      RECT  8677.5 21652.5 8612.5 21787.5 ;
      RECT  8867.5 20812.5 8802.5 20947.5 ;
      RECT  8677.5 20812.5 8612.5 20947.5 ;
      RECT  8677.5 20812.5 8612.5 20947.5 ;
      RECT  8867.5 20812.5 8802.5 20947.5 ;
      RECT  8677.5 20812.5 8612.5 20947.5 ;
      RECT  8487.5 20812.5 8422.5 20947.5 ;
      RECT  8487.5 20812.5 8422.5 20947.5 ;
      RECT  8677.5 20812.5 8612.5 20947.5 ;
      RECT  8317.5 21742.5 8252.5 21877.5 ;
      RECT  8317.5 20767.5 8252.5 20902.5 ;
      RECT  8482.5 21042.5 8617.5 21107.5 ;
      RECT  8740.0 21257.5 8875.0 21322.5 ;
      RECT  8677.5 21652.5 8612.5 21787.5 ;
      RECT  8487.5 20812.5 8422.5 20947.5 ;
      RECT  8387.5 21257.5 8522.5 21322.5 ;
      RECT  8875.0 21257.5 8740.0 21322.5 ;
      RECT  8617.5 21042.5 8482.5 21107.5 ;
      RECT  8522.5 21257.5 8387.5 21322.5 ;
      RECT  8935.0 21962.5 8015.0 22027.5 ;
      RECT  8935.0 20617.5 8015.0 20682.5 ;
      RECT  8867.5 23177.5 8802.5 23372.5 ;
      RECT  8867.5 22337.5 8802.5 21962.5 ;
      RECT  8487.5 22337.5 8422.5 21962.5 ;
      RECT  8317.5 22180.0 8252.5 21995.0 ;
      RECT  8317.5 23340.0 8252.5 23155.0 ;
      RECT  8867.5 22337.5 8802.5 22202.5 ;
      RECT  8677.5 22337.5 8612.5 22202.5 ;
      RECT  8677.5 22337.5 8612.5 22202.5 ;
      RECT  8867.5 22337.5 8802.5 22202.5 ;
      RECT  8677.5 22337.5 8612.5 22202.5 ;
      RECT  8487.5 22337.5 8422.5 22202.5 ;
      RECT  8487.5 22337.5 8422.5 22202.5 ;
      RECT  8677.5 22337.5 8612.5 22202.5 ;
      RECT  8867.5 23177.5 8802.5 23042.5 ;
      RECT  8677.5 23177.5 8612.5 23042.5 ;
      RECT  8677.5 23177.5 8612.5 23042.5 ;
      RECT  8867.5 23177.5 8802.5 23042.5 ;
      RECT  8677.5 23177.5 8612.5 23042.5 ;
      RECT  8487.5 23177.5 8422.5 23042.5 ;
      RECT  8487.5 23177.5 8422.5 23042.5 ;
      RECT  8677.5 23177.5 8612.5 23042.5 ;
      RECT  8317.5 22247.5 8252.5 22112.5 ;
      RECT  8317.5 23222.5 8252.5 23087.5 ;
      RECT  8482.5 22947.5 8617.5 22882.5 ;
      RECT  8740.0 22732.5 8875.0 22667.5 ;
      RECT  8677.5 22337.5 8612.5 22202.5 ;
      RECT  8487.5 23177.5 8422.5 23042.5 ;
      RECT  8387.5 22732.5 8522.5 22667.5 ;
      RECT  8875.0 22732.5 8740.0 22667.5 ;
      RECT  8617.5 22947.5 8482.5 22882.5 ;
      RECT  8522.5 22732.5 8387.5 22667.5 ;
      RECT  8935.0 22027.5 8015.0 21962.5 ;
      RECT  8935.0 23372.5 8015.0 23307.5 ;
      RECT  9932.5 19077.5 10067.5 19142.5 ;
      RECT  11317.5 18555.0 11452.5 18620.0 ;
      RECT  9657.5 20422.5 9792.5 20487.5 ;
      RECT  11042.5 19990.0 11177.5 20055.0 ;
      RECT  11317.5 20752.5 11452.5 20817.5 ;
      RECT  9382.5 20752.5 9517.5 20817.5 ;
      RECT  11042.5 22097.5 11177.5 22162.5 ;
      RECT  9107.5 22097.5 9242.5 22162.5 ;
      RECT  9932.5 18567.5 10067.5 18632.5 ;
      RECT  9657.5 18352.5 9792.5 18417.5 ;
      RECT  9382.5 19977.5 9517.5 20042.5 ;
      RECT  9657.5 20192.5 9792.5 20257.5 ;
      RECT  9932.5 21257.5 10067.5 21322.5 ;
      RECT  9107.5 21042.5 9242.5 21107.5 ;
      RECT  9382.5 22667.5 9517.5 22732.5 ;
      RECT  9107.5 22882.5 9242.5 22947.5 ;
      RECT  7660.0 18555.0 7455.0 18620.0 ;
      RECT  7660.0 19990.0 7455.0 20055.0 ;
      RECT  7660.0 21245.0 7455.0 21310.0 ;
      RECT  7660.0 22680.0 7455.0 22745.0 ;
      RECT  11420.0 19272.5 7455.0 19337.5 ;
      RECT  11420.0 21962.5 7455.0 22027.5 ;
      RECT  11420.0 17927.5 7455.0 17992.5 ;
      RECT  11420.0 20617.5 7455.0 20682.5 ;
      RECT  11420.0 23307.5 7455.0 23372.5 ;
      RECT  10917.5 23935.0 10852.5 24000.0 ;
      RECT  10917.5 24457.5 10852.5 24522.5 ;
      RECT  11155.0 23935.0 10885.0 24000.0 ;
      RECT  10917.5 23967.5 10852.5 24490.0 ;
      RECT  10885.0 24457.5 10640.0 24522.5 ;
      RECT  12300.0 23935.0 11385.0 24000.0 ;
      RECT  10917.5 25370.0 10852.5 25435.0 ;
      RECT  10917.5 25802.5 10852.5 25867.5 ;
      RECT  11155.0 25370.0 10885.0 25435.0 ;
      RECT  10917.5 25402.5 10852.5 25835.0 ;
      RECT  10885.0 25802.5 10365.0 25867.5 ;
      RECT  12025.0 25370.0 11385.0 25435.0 ;
      RECT  10917.5 26625.0 10852.5 26690.0 ;
      RECT  10917.5 27147.5 10852.5 27212.5 ;
      RECT  11155.0 26625.0 10885.0 26690.0 ;
      RECT  10917.5 26657.5 10852.5 27180.0 ;
      RECT  10885.0 27147.5 10090.0 27212.5 ;
      RECT  11750.0 26625.0 11385.0 26690.0 ;
      RECT  12300.0 27477.5 9815.0 27542.5 ;
      RECT  12025.0 28822.5 9540.0 28887.5 ;
      RECT  11750.0 30167.5 9265.0 30232.5 ;
      RECT  10640.0 23995.0 8897.5 24060.0 ;
      RECT  10365.0 23855.0 8707.5 23920.0 ;
      RECT  10090.0 23715.0 8517.5 23780.0 ;
      RECT  9815.0 25310.0 8897.5 25375.0 ;
      RECT  10365.0 25450.0 8707.5 25515.0 ;
      RECT  10090.0 25590.0 8517.5 25655.0 ;
      RECT  10640.0 26685.0 8897.5 26750.0 ;
      RECT  9540.0 26545.0 8707.5 26610.0 ;
      RECT  10090.0 26405.0 8517.5 26470.0 ;
      RECT  9815.0 28000.0 8897.5 28065.0 ;
      RECT  9540.0 28140.0 8707.5 28205.0 ;
      RECT  10090.0 28280.0 8517.5 28345.0 ;
      RECT  10640.0 29375.0 8897.5 29440.0 ;
      RECT  10365.0 29235.0 8707.5 29300.0 ;
      RECT  9265.0 29095.0 8517.5 29160.0 ;
      RECT  9815.0 30690.0 8897.5 30755.0 ;
      RECT  10365.0 30830.0 8707.5 30895.0 ;
      RECT  9265.0 30970.0 8517.5 31035.0 ;
      RECT  10640.0 32065.0 8897.5 32130.0 ;
      RECT  9540.0 31925.0 8707.5 31990.0 ;
      RECT  9265.0 31785.0 8517.5 31850.0 ;
      RECT  9815.0 33380.0 8897.5 33445.0 ;
      RECT  9540.0 33520.0 8707.5 33585.0 ;
      RECT  9265.0 33660.0 8517.5 33725.0 ;
      RECT  8137.5 23995.0 8072.5 24060.0 ;
      RECT  8137.5 23935.0 8072.5 24000.0 ;
      RECT  8322.5 23995.0 8105.0 24060.0 ;
      RECT  8137.5 23967.5 8072.5 24027.5 ;
      RECT  8105.0 23935.0 7890.0 24000.0 ;
      RECT  8137.5 25310.0 8072.5 25375.0 ;
      RECT  8137.5 25370.0 8072.5 25435.0 ;
      RECT  8322.5 25310.0 8105.0 25375.0 ;
      RECT  8137.5 25342.5 8072.5 25402.5 ;
      RECT  8105.0 25370.0 7890.0 25435.0 ;
      RECT  8137.5 26685.0 8072.5 26750.0 ;
      RECT  8137.5 26625.0 8072.5 26690.0 ;
      RECT  8322.5 26685.0 8105.0 26750.0 ;
      RECT  8137.5 26657.5 8072.5 26717.5 ;
      RECT  8105.0 26625.0 7890.0 26690.0 ;
      RECT  8137.5 28000.0 8072.5 28065.0 ;
      RECT  8137.5 28060.0 8072.5 28125.0 ;
      RECT  8322.5 28000.0 8105.0 28065.0 ;
      RECT  8137.5 28032.5 8072.5 28092.5 ;
      RECT  8105.0 28060.0 7890.0 28125.0 ;
      RECT  8137.5 29375.0 8072.5 29440.0 ;
      RECT  8137.5 29315.0 8072.5 29380.0 ;
      RECT  8322.5 29375.0 8105.0 29440.0 ;
      RECT  8137.5 29347.5 8072.5 29407.5 ;
      RECT  8105.0 29315.0 7890.0 29380.0 ;
      RECT  8137.5 30690.0 8072.5 30755.0 ;
      RECT  8137.5 30750.0 8072.5 30815.0 ;
      RECT  8322.5 30690.0 8105.0 30755.0 ;
      RECT  8137.5 30722.5 8072.5 30782.5 ;
      RECT  8105.0 30750.0 7890.0 30815.0 ;
      RECT  8137.5 32065.0 8072.5 32130.0 ;
      RECT  8137.5 32005.0 8072.5 32070.0 ;
      RECT  8322.5 32065.0 8105.0 32130.0 ;
      RECT  8137.5 32037.5 8072.5 32097.5 ;
      RECT  8105.0 32005.0 7890.0 32070.0 ;
      RECT  8137.5 33380.0 8072.5 33445.0 ;
      RECT  8137.5 33440.0 8072.5 33505.0 ;
      RECT  8322.5 33380.0 8105.0 33445.0 ;
      RECT  8137.5 33412.5 8072.5 33472.5 ;
      RECT  8105.0 33440.0 7890.0 33505.0 ;
      RECT  11082.5 24500.0 11017.5 24685.0 ;
      RECT  11082.5 23340.0 11017.5 23525.0 ;
      RECT  11442.5 23457.5 11377.5 23307.5 ;
      RECT  11442.5 24342.5 11377.5 24717.5 ;
      RECT  11252.5 23457.5 11187.5 24342.5 ;
      RECT  11442.5 24342.5 11377.5 24477.5 ;
      RECT  11252.5 24342.5 11187.5 24477.5 ;
      RECT  11252.5 24342.5 11187.5 24477.5 ;
      RECT  11442.5 24342.5 11377.5 24477.5 ;
      RECT  11442.5 23457.5 11377.5 23592.5 ;
      RECT  11252.5 23457.5 11187.5 23592.5 ;
      RECT  11252.5 23457.5 11187.5 23592.5 ;
      RECT  11442.5 23457.5 11377.5 23592.5 ;
      RECT  11082.5 24432.5 11017.5 24567.5 ;
      RECT  11082.5 23457.5 11017.5 23592.5 ;
      RECT  11385.0 23900.0 11320.0 24035.0 ;
      RECT  11385.0 23900.0 11320.0 24035.0 ;
      RECT  11220.0 23935.0 11155.0 24000.0 ;
      RECT  11510.0 24652.5 10950.0 24717.5 ;
      RECT  11510.0 23307.5 10950.0 23372.5 ;
      RECT  11082.5 24870.0 11017.5 24685.0 ;
      RECT  11082.5 26030.0 11017.5 25845.0 ;
      RECT  11442.5 25912.5 11377.5 26062.5 ;
      RECT  11442.5 25027.5 11377.5 24652.5 ;
      RECT  11252.5 25912.5 11187.5 25027.5 ;
      RECT  11442.5 25027.5 11377.5 24892.5 ;
      RECT  11252.5 25027.5 11187.5 24892.5 ;
      RECT  11252.5 25027.5 11187.5 24892.5 ;
      RECT  11442.5 25027.5 11377.5 24892.5 ;
      RECT  11442.5 25912.5 11377.5 25777.5 ;
      RECT  11252.5 25912.5 11187.5 25777.5 ;
      RECT  11252.5 25912.5 11187.5 25777.5 ;
      RECT  11442.5 25912.5 11377.5 25777.5 ;
      RECT  11082.5 24937.5 11017.5 24802.5 ;
      RECT  11082.5 25912.5 11017.5 25777.5 ;
      RECT  11385.0 25470.0 11320.0 25335.0 ;
      RECT  11385.0 25470.0 11320.0 25335.0 ;
      RECT  11220.0 25435.0 11155.0 25370.0 ;
      RECT  11510.0 24717.5 10950.0 24652.5 ;
      RECT  11510.0 26062.5 10950.0 25997.5 ;
      RECT  11082.5 27190.0 11017.5 27375.0 ;
      RECT  11082.5 26030.0 11017.5 26215.0 ;
      RECT  11442.5 26147.5 11377.5 25997.5 ;
      RECT  11442.5 27032.5 11377.5 27407.5 ;
      RECT  11252.5 26147.5 11187.5 27032.5 ;
      RECT  11442.5 27032.5 11377.5 27167.5 ;
      RECT  11252.5 27032.5 11187.5 27167.5 ;
      RECT  11252.5 27032.5 11187.5 27167.5 ;
      RECT  11442.5 27032.5 11377.5 27167.5 ;
      RECT  11442.5 26147.5 11377.5 26282.5 ;
      RECT  11252.5 26147.5 11187.5 26282.5 ;
      RECT  11252.5 26147.5 11187.5 26282.5 ;
      RECT  11442.5 26147.5 11377.5 26282.5 ;
      RECT  11082.5 27122.5 11017.5 27257.5 ;
      RECT  11082.5 26147.5 11017.5 26282.5 ;
      RECT  11385.0 26590.0 11320.0 26725.0 ;
      RECT  11385.0 26590.0 11320.0 26725.0 ;
      RECT  11220.0 26625.0 11155.0 26690.0 ;
      RECT  11510.0 27342.5 10950.0 27407.5 ;
      RECT  11510.0 25997.5 10950.0 26062.5 ;
      RECT  7587.5 24500.0 7522.5 24685.0 ;
      RECT  7587.5 23340.0 7522.5 23525.0 ;
      RECT  7947.5 23457.5 7882.5 23307.5 ;
      RECT  7947.5 24342.5 7882.5 24717.5 ;
      RECT  7757.5 23457.5 7692.5 24342.5 ;
      RECT  7947.5 24342.5 7882.5 24477.5 ;
      RECT  7757.5 24342.5 7692.5 24477.5 ;
      RECT  7757.5 24342.5 7692.5 24477.5 ;
      RECT  7947.5 24342.5 7882.5 24477.5 ;
      RECT  7947.5 23457.5 7882.5 23592.5 ;
      RECT  7757.5 23457.5 7692.5 23592.5 ;
      RECT  7757.5 23457.5 7692.5 23592.5 ;
      RECT  7947.5 23457.5 7882.5 23592.5 ;
      RECT  7587.5 24432.5 7522.5 24567.5 ;
      RECT  7587.5 23457.5 7522.5 23592.5 ;
      RECT  7890.0 23900.0 7825.0 24035.0 ;
      RECT  7890.0 23900.0 7825.0 24035.0 ;
      RECT  7725.0 23935.0 7660.0 24000.0 ;
      RECT  8015.0 24652.5 7455.0 24717.5 ;
      RECT  8015.0 23307.5 7455.0 23372.5 ;
      RECT  7587.5 24870.0 7522.5 24685.0 ;
      RECT  7587.5 26030.0 7522.5 25845.0 ;
      RECT  7947.5 25912.5 7882.5 26062.5 ;
      RECT  7947.5 25027.5 7882.5 24652.5 ;
      RECT  7757.5 25912.5 7692.5 25027.5 ;
      RECT  7947.5 25027.5 7882.5 24892.5 ;
      RECT  7757.5 25027.5 7692.5 24892.5 ;
      RECT  7757.5 25027.5 7692.5 24892.5 ;
      RECT  7947.5 25027.5 7882.5 24892.5 ;
      RECT  7947.5 25912.5 7882.5 25777.5 ;
      RECT  7757.5 25912.5 7692.5 25777.5 ;
      RECT  7757.5 25912.5 7692.5 25777.5 ;
      RECT  7947.5 25912.5 7882.5 25777.5 ;
      RECT  7587.5 24937.5 7522.5 24802.5 ;
      RECT  7587.5 25912.5 7522.5 25777.5 ;
      RECT  7890.0 25470.0 7825.0 25335.0 ;
      RECT  7890.0 25470.0 7825.0 25335.0 ;
      RECT  7725.0 25435.0 7660.0 25370.0 ;
      RECT  8015.0 24717.5 7455.0 24652.5 ;
      RECT  8015.0 26062.5 7455.0 25997.5 ;
      RECT  7587.5 27190.0 7522.5 27375.0 ;
      RECT  7587.5 26030.0 7522.5 26215.0 ;
      RECT  7947.5 26147.5 7882.5 25997.5 ;
      RECT  7947.5 27032.5 7882.5 27407.5 ;
      RECT  7757.5 26147.5 7692.5 27032.5 ;
      RECT  7947.5 27032.5 7882.5 27167.5 ;
      RECT  7757.5 27032.5 7692.5 27167.5 ;
      RECT  7757.5 27032.5 7692.5 27167.5 ;
      RECT  7947.5 27032.5 7882.5 27167.5 ;
      RECT  7947.5 26147.5 7882.5 26282.5 ;
      RECT  7757.5 26147.5 7692.5 26282.5 ;
      RECT  7757.5 26147.5 7692.5 26282.5 ;
      RECT  7947.5 26147.5 7882.5 26282.5 ;
      RECT  7587.5 27122.5 7522.5 27257.5 ;
      RECT  7587.5 26147.5 7522.5 26282.5 ;
      RECT  7890.0 26590.0 7825.0 26725.0 ;
      RECT  7890.0 26590.0 7825.0 26725.0 ;
      RECT  7725.0 26625.0 7660.0 26690.0 ;
      RECT  8015.0 27342.5 7455.0 27407.5 ;
      RECT  8015.0 25997.5 7455.0 26062.5 ;
      RECT  7587.5 27560.0 7522.5 27375.0 ;
      RECT  7587.5 28720.0 7522.5 28535.0 ;
      RECT  7947.5 28602.5 7882.5 28752.5 ;
      RECT  7947.5 27717.5 7882.5 27342.5 ;
      RECT  7757.5 28602.5 7692.5 27717.5 ;
      RECT  7947.5 27717.5 7882.5 27582.5 ;
      RECT  7757.5 27717.5 7692.5 27582.5 ;
      RECT  7757.5 27717.5 7692.5 27582.5 ;
      RECT  7947.5 27717.5 7882.5 27582.5 ;
      RECT  7947.5 28602.5 7882.5 28467.5 ;
      RECT  7757.5 28602.5 7692.5 28467.5 ;
      RECT  7757.5 28602.5 7692.5 28467.5 ;
      RECT  7947.5 28602.5 7882.5 28467.5 ;
      RECT  7587.5 27627.5 7522.5 27492.5 ;
      RECT  7587.5 28602.5 7522.5 28467.5 ;
      RECT  7890.0 28160.0 7825.0 28025.0 ;
      RECT  7890.0 28160.0 7825.0 28025.0 ;
      RECT  7725.0 28125.0 7660.0 28060.0 ;
      RECT  8015.0 27407.5 7455.0 27342.5 ;
      RECT  8015.0 28752.5 7455.0 28687.5 ;
      RECT  7587.5 29880.0 7522.5 30065.0 ;
      RECT  7587.5 28720.0 7522.5 28905.0 ;
      RECT  7947.5 28837.5 7882.5 28687.5 ;
      RECT  7947.5 29722.5 7882.5 30097.5 ;
      RECT  7757.5 28837.5 7692.5 29722.5 ;
      RECT  7947.5 29722.5 7882.5 29857.5 ;
      RECT  7757.5 29722.5 7692.5 29857.5 ;
      RECT  7757.5 29722.5 7692.5 29857.5 ;
      RECT  7947.5 29722.5 7882.5 29857.5 ;
      RECT  7947.5 28837.5 7882.5 28972.5 ;
      RECT  7757.5 28837.5 7692.5 28972.5 ;
      RECT  7757.5 28837.5 7692.5 28972.5 ;
      RECT  7947.5 28837.5 7882.5 28972.5 ;
      RECT  7587.5 29812.5 7522.5 29947.5 ;
      RECT  7587.5 28837.5 7522.5 28972.5 ;
      RECT  7890.0 29280.0 7825.0 29415.0 ;
      RECT  7890.0 29280.0 7825.0 29415.0 ;
      RECT  7725.0 29315.0 7660.0 29380.0 ;
      RECT  8015.0 30032.5 7455.0 30097.5 ;
      RECT  8015.0 28687.5 7455.0 28752.5 ;
      RECT  7587.5 30250.0 7522.5 30065.0 ;
      RECT  7587.5 31410.0 7522.5 31225.0 ;
      RECT  7947.5 31292.5 7882.5 31442.5 ;
      RECT  7947.5 30407.5 7882.5 30032.5 ;
      RECT  7757.5 31292.5 7692.5 30407.5 ;
      RECT  7947.5 30407.5 7882.5 30272.5 ;
      RECT  7757.5 30407.5 7692.5 30272.5 ;
      RECT  7757.5 30407.5 7692.5 30272.5 ;
      RECT  7947.5 30407.5 7882.5 30272.5 ;
      RECT  7947.5 31292.5 7882.5 31157.5 ;
      RECT  7757.5 31292.5 7692.5 31157.5 ;
      RECT  7757.5 31292.5 7692.5 31157.5 ;
      RECT  7947.5 31292.5 7882.5 31157.5 ;
      RECT  7587.5 30317.5 7522.5 30182.5 ;
      RECT  7587.5 31292.5 7522.5 31157.5 ;
      RECT  7890.0 30850.0 7825.0 30715.0 ;
      RECT  7890.0 30850.0 7825.0 30715.0 ;
      RECT  7725.0 30815.0 7660.0 30750.0 ;
      RECT  8015.0 30097.5 7455.0 30032.5 ;
      RECT  8015.0 31442.5 7455.0 31377.5 ;
      RECT  7587.5 32570.0 7522.5 32755.0 ;
      RECT  7587.5 31410.0 7522.5 31595.0 ;
      RECT  7947.5 31527.5 7882.5 31377.5 ;
      RECT  7947.5 32412.5 7882.5 32787.5 ;
      RECT  7757.5 31527.5 7692.5 32412.5 ;
      RECT  7947.5 32412.5 7882.5 32547.5 ;
      RECT  7757.5 32412.5 7692.5 32547.5 ;
      RECT  7757.5 32412.5 7692.5 32547.5 ;
      RECT  7947.5 32412.5 7882.5 32547.5 ;
      RECT  7947.5 31527.5 7882.5 31662.5 ;
      RECT  7757.5 31527.5 7692.5 31662.5 ;
      RECT  7757.5 31527.5 7692.5 31662.5 ;
      RECT  7947.5 31527.5 7882.5 31662.5 ;
      RECT  7587.5 32502.5 7522.5 32637.5 ;
      RECT  7587.5 31527.5 7522.5 31662.5 ;
      RECT  7890.0 31970.0 7825.0 32105.0 ;
      RECT  7890.0 31970.0 7825.0 32105.0 ;
      RECT  7725.0 32005.0 7660.0 32070.0 ;
      RECT  8015.0 32722.5 7455.0 32787.5 ;
      RECT  8015.0 31377.5 7455.0 31442.5 ;
      RECT  7587.5 32940.0 7522.5 32755.0 ;
      RECT  7587.5 34100.0 7522.5 33915.0 ;
      RECT  7947.5 33982.5 7882.5 34132.5 ;
      RECT  7947.5 33097.5 7882.5 32722.5 ;
      RECT  7757.5 33982.5 7692.5 33097.5 ;
      RECT  7947.5 33097.5 7882.5 32962.5 ;
      RECT  7757.5 33097.5 7692.5 32962.5 ;
      RECT  7757.5 33097.5 7692.5 32962.5 ;
      RECT  7947.5 33097.5 7882.5 32962.5 ;
      RECT  7947.5 33982.5 7882.5 33847.5 ;
      RECT  7757.5 33982.5 7692.5 33847.5 ;
      RECT  7757.5 33982.5 7692.5 33847.5 ;
      RECT  7947.5 33982.5 7882.5 33847.5 ;
      RECT  7587.5 33007.5 7522.5 32872.5 ;
      RECT  7587.5 33982.5 7522.5 33847.5 ;
      RECT  7890.0 33540.0 7825.0 33405.0 ;
      RECT  7890.0 33540.0 7825.0 33405.0 ;
      RECT  7725.0 33505.0 7660.0 33440.0 ;
      RECT  8015.0 32787.5 7455.0 32722.5 ;
      RECT  8015.0 34132.5 7455.0 34067.5 ;
      RECT  8957.5 23502.5 8892.5 23307.5 ;
      RECT  8957.5 24342.5 8892.5 24717.5 ;
      RECT  8577.5 24342.5 8512.5 24717.5 ;
      RECT  8217.5 24500.0 8152.5 24685.0 ;
      RECT  8217.5 23340.0 8152.5 23525.0 ;
      RECT  8957.5 24342.5 8892.5 24477.5 ;
      RECT  8767.5 24342.5 8702.5 24477.5 ;
      RECT  8767.5 24342.5 8702.5 24477.5 ;
      RECT  8957.5 24342.5 8892.5 24477.5 ;
      RECT  8767.5 24342.5 8702.5 24477.5 ;
      RECT  8577.5 24342.5 8512.5 24477.5 ;
      RECT  8577.5 24342.5 8512.5 24477.5 ;
      RECT  8767.5 24342.5 8702.5 24477.5 ;
      RECT  8577.5 24342.5 8512.5 24477.5 ;
      RECT  8387.5 24342.5 8322.5 24477.5 ;
      RECT  8387.5 24342.5 8322.5 24477.5 ;
      RECT  8577.5 24342.5 8512.5 24477.5 ;
      RECT  8957.5 23502.5 8892.5 23637.5 ;
      RECT  8767.5 23502.5 8702.5 23637.5 ;
      RECT  8767.5 23502.5 8702.5 23637.5 ;
      RECT  8957.5 23502.5 8892.5 23637.5 ;
      RECT  8767.5 23502.5 8702.5 23637.5 ;
      RECT  8577.5 23502.5 8512.5 23637.5 ;
      RECT  8577.5 23502.5 8512.5 23637.5 ;
      RECT  8767.5 23502.5 8702.5 23637.5 ;
      RECT  8577.5 23502.5 8512.5 23637.5 ;
      RECT  8387.5 23502.5 8322.5 23637.5 ;
      RECT  8387.5 23502.5 8322.5 23637.5 ;
      RECT  8577.5 23502.5 8512.5 23637.5 ;
      RECT  8217.5 24432.5 8152.5 24567.5 ;
      RECT  8217.5 23457.5 8152.5 23592.5 ;
      RECT  8382.5 23715.0 8517.5 23780.0 ;
      RECT  8572.5 23855.0 8707.5 23920.0 ;
      RECT  8762.5 23995.0 8897.5 24060.0 ;
      RECT  8767.5 24342.5 8702.5 24477.5 ;
      RECT  8387.5 24342.5 8322.5 24477.5 ;
      RECT  8387.5 23502.5 8322.5 23637.5 ;
      RECT  8387.5 23960.0 8322.5 24095.0 ;
      RECT  8897.5 23995.0 8762.5 24060.0 ;
      RECT  8707.5 23855.0 8572.5 23920.0 ;
      RECT  8517.5 23715.0 8382.5 23780.0 ;
      RECT  8387.5 23960.0 8322.5 24095.0 ;
      RECT  9025.0 24652.5 8015.0 24717.5 ;
      RECT  9025.0 23307.5 8015.0 23372.5 ;
      RECT  8957.5 25867.5 8892.5 26062.5 ;
      RECT  8957.5 25027.5 8892.5 24652.5 ;
      RECT  8577.5 25027.5 8512.5 24652.5 ;
      RECT  8217.5 24870.0 8152.5 24685.0 ;
      RECT  8217.5 26030.0 8152.5 25845.0 ;
      RECT  8957.5 25027.5 8892.5 24892.5 ;
      RECT  8767.5 25027.5 8702.5 24892.5 ;
      RECT  8767.5 25027.5 8702.5 24892.5 ;
      RECT  8957.5 25027.5 8892.5 24892.5 ;
      RECT  8767.5 25027.5 8702.5 24892.5 ;
      RECT  8577.5 25027.5 8512.5 24892.5 ;
      RECT  8577.5 25027.5 8512.5 24892.5 ;
      RECT  8767.5 25027.5 8702.5 24892.5 ;
      RECT  8577.5 25027.5 8512.5 24892.5 ;
      RECT  8387.5 25027.5 8322.5 24892.5 ;
      RECT  8387.5 25027.5 8322.5 24892.5 ;
      RECT  8577.5 25027.5 8512.5 24892.5 ;
      RECT  8957.5 25867.5 8892.5 25732.5 ;
      RECT  8767.5 25867.5 8702.5 25732.5 ;
      RECT  8767.5 25867.5 8702.5 25732.5 ;
      RECT  8957.5 25867.5 8892.5 25732.5 ;
      RECT  8767.5 25867.5 8702.5 25732.5 ;
      RECT  8577.5 25867.5 8512.5 25732.5 ;
      RECT  8577.5 25867.5 8512.5 25732.5 ;
      RECT  8767.5 25867.5 8702.5 25732.5 ;
      RECT  8577.5 25867.5 8512.5 25732.5 ;
      RECT  8387.5 25867.5 8322.5 25732.5 ;
      RECT  8387.5 25867.5 8322.5 25732.5 ;
      RECT  8577.5 25867.5 8512.5 25732.5 ;
      RECT  8217.5 24937.5 8152.5 24802.5 ;
      RECT  8217.5 25912.5 8152.5 25777.5 ;
      RECT  8382.5 25655.0 8517.5 25590.0 ;
      RECT  8572.5 25515.0 8707.5 25450.0 ;
      RECT  8762.5 25375.0 8897.5 25310.0 ;
      RECT  8767.5 25027.5 8702.5 24892.5 ;
      RECT  8387.5 25027.5 8322.5 24892.5 ;
      RECT  8387.5 25867.5 8322.5 25732.5 ;
      RECT  8387.5 25410.0 8322.5 25275.0 ;
      RECT  8897.5 25375.0 8762.5 25310.0 ;
      RECT  8707.5 25515.0 8572.5 25450.0 ;
      RECT  8517.5 25655.0 8382.5 25590.0 ;
      RECT  8387.5 25410.0 8322.5 25275.0 ;
      RECT  9025.0 24717.5 8015.0 24652.5 ;
      RECT  9025.0 26062.5 8015.0 25997.5 ;
      RECT  8957.5 26192.5 8892.5 25997.5 ;
      RECT  8957.5 27032.5 8892.5 27407.5 ;
      RECT  8577.5 27032.5 8512.5 27407.5 ;
      RECT  8217.5 27190.0 8152.5 27375.0 ;
      RECT  8217.5 26030.0 8152.5 26215.0 ;
      RECT  8957.5 27032.5 8892.5 27167.5 ;
      RECT  8767.5 27032.5 8702.5 27167.5 ;
      RECT  8767.5 27032.5 8702.5 27167.5 ;
      RECT  8957.5 27032.5 8892.5 27167.5 ;
      RECT  8767.5 27032.5 8702.5 27167.5 ;
      RECT  8577.5 27032.5 8512.5 27167.5 ;
      RECT  8577.5 27032.5 8512.5 27167.5 ;
      RECT  8767.5 27032.5 8702.5 27167.5 ;
      RECT  8577.5 27032.5 8512.5 27167.5 ;
      RECT  8387.5 27032.5 8322.5 27167.5 ;
      RECT  8387.5 27032.5 8322.5 27167.5 ;
      RECT  8577.5 27032.5 8512.5 27167.5 ;
      RECT  8957.5 26192.5 8892.5 26327.5 ;
      RECT  8767.5 26192.5 8702.5 26327.5 ;
      RECT  8767.5 26192.5 8702.5 26327.5 ;
      RECT  8957.5 26192.5 8892.5 26327.5 ;
      RECT  8767.5 26192.5 8702.5 26327.5 ;
      RECT  8577.5 26192.5 8512.5 26327.5 ;
      RECT  8577.5 26192.5 8512.5 26327.5 ;
      RECT  8767.5 26192.5 8702.5 26327.5 ;
      RECT  8577.5 26192.5 8512.5 26327.5 ;
      RECT  8387.5 26192.5 8322.5 26327.5 ;
      RECT  8387.5 26192.5 8322.5 26327.5 ;
      RECT  8577.5 26192.5 8512.5 26327.5 ;
      RECT  8217.5 27122.5 8152.5 27257.5 ;
      RECT  8217.5 26147.5 8152.5 26282.5 ;
      RECT  8382.5 26405.0 8517.5 26470.0 ;
      RECT  8572.5 26545.0 8707.5 26610.0 ;
      RECT  8762.5 26685.0 8897.5 26750.0 ;
      RECT  8767.5 27032.5 8702.5 27167.5 ;
      RECT  8387.5 27032.5 8322.5 27167.5 ;
      RECT  8387.5 26192.5 8322.5 26327.5 ;
      RECT  8387.5 26650.0 8322.5 26785.0 ;
      RECT  8897.5 26685.0 8762.5 26750.0 ;
      RECT  8707.5 26545.0 8572.5 26610.0 ;
      RECT  8517.5 26405.0 8382.5 26470.0 ;
      RECT  8387.5 26650.0 8322.5 26785.0 ;
      RECT  9025.0 27342.5 8015.0 27407.5 ;
      RECT  9025.0 25997.5 8015.0 26062.5 ;
      RECT  8957.5 28557.5 8892.5 28752.5 ;
      RECT  8957.5 27717.5 8892.5 27342.5 ;
      RECT  8577.5 27717.5 8512.5 27342.5 ;
      RECT  8217.5 27560.0 8152.5 27375.0 ;
      RECT  8217.5 28720.0 8152.5 28535.0 ;
      RECT  8957.5 27717.5 8892.5 27582.5 ;
      RECT  8767.5 27717.5 8702.5 27582.5 ;
      RECT  8767.5 27717.5 8702.5 27582.5 ;
      RECT  8957.5 27717.5 8892.5 27582.5 ;
      RECT  8767.5 27717.5 8702.5 27582.5 ;
      RECT  8577.5 27717.5 8512.5 27582.5 ;
      RECT  8577.5 27717.5 8512.5 27582.5 ;
      RECT  8767.5 27717.5 8702.5 27582.5 ;
      RECT  8577.5 27717.5 8512.5 27582.5 ;
      RECT  8387.5 27717.5 8322.5 27582.5 ;
      RECT  8387.5 27717.5 8322.5 27582.5 ;
      RECT  8577.5 27717.5 8512.5 27582.5 ;
      RECT  8957.5 28557.5 8892.5 28422.5 ;
      RECT  8767.5 28557.5 8702.5 28422.5 ;
      RECT  8767.5 28557.5 8702.5 28422.5 ;
      RECT  8957.5 28557.5 8892.5 28422.5 ;
      RECT  8767.5 28557.5 8702.5 28422.5 ;
      RECT  8577.5 28557.5 8512.5 28422.5 ;
      RECT  8577.5 28557.5 8512.5 28422.5 ;
      RECT  8767.5 28557.5 8702.5 28422.5 ;
      RECT  8577.5 28557.5 8512.5 28422.5 ;
      RECT  8387.5 28557.5 8322.5 28422.5 ;
      RECT  8387.5 28557.5 8322.5 28422.5 ;
      RECT  8577.5 28557.5 8512.5 28422.5 ;
      RECT  8217.5 27627.5 8152.5 27492.5 ;
      RECT  8217.5 28602.5 8152.5 28467.5 ;
      RECT  8382.5 28345.0 8517.5 28280.0 ;
      RECT  8572.5 28205.0 8707.5 28140.0 ;
      RECT  8762.5 28065.0 8897.5 28000.0 ;
      RECT  8767.5 27717.5 8702.5 27582.5 ;
      RECT  8387.5 27717.5 8322.5 27582.5 ;
      RECT  8387.5 28557.5 8322.5 28422.5 ;
      RECT  8387.5 28100.0 8322.5 27965.0 ;
      RECT  8897.5 28065.0 8762.5 28000.0 ;
      RECT  8707.5 28205.0 8572.5 28140.0 ;
      RECT  8517.5 28345.0 8382.5 28280.0 ;
      RECT  8387.5 28100.0 8322.5 27965.0 ;
      RECT  9025.0 27407.5 8015.0 27342.5 ;
      RECT  9025.0 28752.5 8015.0 28687.5 ;
      RECT  8957.5 28882.5 8892.5 28687.5 ;
      RECT  8957.5 29722.5 8892.5 30097.5 ;
      RECT  8577.5 29722.5 8512.5 30097.5 ;
      RECT  8217.5 29880.0 8152.5 30065.0 ;
      RECT  8217.5 28720.0 8152.5 28905.0 ;
      RECT  8957.5 29722.5 8892.5 29857.5 ;
      RECT  8767.5 29722.5 8702.5 29857.5 ;
      RECT  8767.5 29722.5 8702.5 29857.5 ;
      RECT  8957.5 29722.5 8892.5 29857.5 ;
      RECT  8767.5 29722.5 8702.5 29857.5 ;
      RECT  8577.5 29722.5 8512.5 29857.5 ;
      RECT  8577.5 29722.5 8512.5 29857.5 ;
      RECT  8767.5 29722.5 8702.5 29857.5 ;
      RECT  8577.5 29722.5 8512.5 29857.5 ;
      RECT  8387.5 29722.5 8322.5 29857.5 ;
      RECT  8387.5 29722.5 8322.5 29857.5 ;
      RECT  8577.5 29722.5 8512.5 29857.5 ;
      RECT  8957.5 28882.5 8892.5 29017.5 ;
      RECT  8767.5 28882.5 8702.5 29017.5 ;
      RECT  8767.5 28882.5 8702.5 29017.5 ;
      RECT  8957.5 28882.5 8892.5 29017.5 ;
      RECT  8767.5 28882.5 8702.5 29017.5 ;
      RECT  8577.5 28882.5 8512.5 29017.5 ;
      RECT  8577.5 28882.5 8512.5 29017.5 ;
      RECT  8767.5 28882.5 8702.5 29017.5 ;
      RECT  8577.5 28882.5 8512.5 29017.5 ;
      RECT  8387.5 28882.5 8322.5 29017.5 ;
      RECT  8387.5 28882.5 8322.5 29017.5 ;
      RECT  8577.5 28882.5 8512.5 29017.5 ;
      RECT  8217.5 29812.5 8152.5 29947.5 ;
      RECT  8217.5 28837.5 8152.5 28972.5 ;
      RECT  8382.5 29095.0 8517.5 29160.0 ;
      RECT  8572.5 29235.0 8707.5 29300.0 ;
      RECT  8762.5 29375.0 8897.5 29440.0 ;
      RECT  8767.5 29722.5 8702.5 29857.5 ;
      RECT  8387.5 29722.5 8322.5 29857.5 ;
      RECT  8387.5 28882.5 8322.5 29017.5 ;
      RECT  8387.5 29340.0 8322.5 29475.0 ;
      RECT  8897.5 29375.0 8762.5 29440.0 ;
      RECT  8707.5 29235.0 8572.5 29300.0 ;
      RECT  8517.5 29095.0 8382.5 29160.0 ;
      RECT  8387.5 29340.0 8322.5 29475.0 ;
      RECT  9025.0 30032.5 8015.0 30097.5 ;
      RECT  9025.0 28687.5 8015.0 28752.5 ;
      RECT  8957.5 31247.5 8892.5 31442.5 ;
      RECT  8957.5 30407.5 8892.5 30032.5 ;
      RECT  8577.5 30407.5 8512.5 30032.5 ;
      RECT  8217.5 30250.0 8152.5 30065.0 ;
      RECT  8217.5 31410.0 8152.5 31225.0 ;
      RECT  8957.5 30407.5 8892.5 30272.5 ;
      RECT  8767.5 30407.5 8702.5 30272.5 ;
      RECT  8767.5 30407.5 8702.5 30272.5 ;
      RECT  8957.5 30407.5 8892.5 30272.5 ;
      RECT  8767.5 30407.5 8702.5 30272.5 ;
      RECT  8577.5 30407.5 8512.5 30272.5 ;
      RECT  8577.5 30407.5 8512.5 30272.5 ;
      RECT  8767.5 30407.5 8702.5 30272.5 ;
      RECT  8577.5 30407.5 8512.5 30272.5 ;
      RECT  8387.5 30407.5 8322.5 30272.5 ;
      RECT  8387.5 30407.5 8322.5 30272.5 ;
      RECT  8577.5 30407.5 8512.5 30272.5 ;
      RECT  8957.5 31247.5 8892.5 31112.5 ;
      RECT  8767.5 31247.5 8702.5 31112.5 ;
      RECT  8767.5 31247.5 8702.5 31112.5 ;
      RECT  8957.5 31247.5 8892.5 31112.5 ;
      RECT  8767.5 31247.5 8702.5 31112.5 ;
      RECT  8577.5 31247.5 8512.5 31112.5 ;
      RECT  8577.5 31247.5 8512.5 31112.5 ;
      RECT  8767.5 31247.5 8702.5 31112.5 ;
      RECT  8577.5 31247.5 8512.5 31112.5 ;
      RECT  8387.5 31247.5 8322.5 31112.5 ;
      RECT  8387.5 31247.5 8322.5 31112.5 ;
      RECT  8577.5 31247.5 8512.5 31112.5 ;
      RECT  8217.5 30317.5 8152.5 30182.5 ;
      RECT  8217.5 31292.5 8152.5 31157.5 ;
      RECT  8382.5 31035.0 8517.5 30970.0 ;
      RECT  8572.5 30895.0 8707.5 30830.0 ;
      RECT  8762.5 30755.0 8897.5 30690.0 ;
      RECT  8767.5 30407.5 8702.5 30272.5 ;
      RECT  8387.5 30407.5 8322.5 30272.5 ;
      RECT  8387.5 31247.5 8322.5 31112.5 ;
      RECT  8387.5 30790.0 8322.5 30655.0 ;
      RECT  8897.5 30755.0 8762.5 30690.0 ;
      RECT  8707.5 30895.0 8572.5 30830.0 ;
      RECT  8517.5 31035.0 8382.5 30970.0 ;
      RECT  8387.5 30790.0 8322.5 30655.0 ;
      RECT  9025.0 30097.5 8015.0 30032.5 ;
      RECT  9025.0 31442.5 8015.0 31377.5 ;
      RECT  8957.5 31572.5 8892.5 31377.5 ;
      RECT  8957.5 32412.5 8892.5 32787.5 ;
      RECT  8577.5 32412.5 8512.5 32787.5 ;
      RECT  8217.5 32570.0 8152.5 32755.0 ;
      RECT  8217.5 31410.0 8152.5 31595.0 ;
      RECT  8957.5 32412.5 8892.5 32547.5 ;
      RECT  8767.5 32412.5 8702.5 32547.5 ;
      RECT  8767.5 32412.5 8702.5 32547.5 ;
      RECT  8957.5 32412.5 8892.5 32547.5 ;
      RECT  8767.5 32412.5 8702.5 32547.5 ;
      RECT  8577.5 32412.5 8512.5 32547.5 ;
      RECT  8577.5 32412.5 8512.5 32547.5 ;
      RECT  8767.5 32412.5 8702.5 32547.5 ;
      RECT  8577.5 32412.5 8512.5 32547.5 ;
      RECT  8387.5 32412.5 8322.5 32547.5 ;
      RECT  8387.5 32412.5 8322.5 32547.5 ;
      RECT  8577.5 32412.5 8512.5 32547.5 ;
      RECT  8957.5 31572.5 8892.5 31707.5 ;
      RECT  8767.5 31572.5 8702.5 31707.5 ;
      RECT  8767.5 31572.5 8702.5 31707.5 ;
      RECT  8957.5 31572.5 8892.5 31707.5 ;
      RECT  8767.5 31572.5 8702.5 31707.5 ;
      RECT  8577.5 31572.5 8512.5 31707.5 ;
      RECT  8577.5 31572.5 8512.5 31707.5 ;
      RECT  8767.5 31572.5 8702.5 31707.5 ;
      RECT  8577.5 31572.5 8512.5 31707.5 ;
      RECT  8387.5 31572.5 8322.5 31707.5 ;
      RECT  8387.5 31572.5 8322.5 31707.5 ;
      RECT  8577.5 31572.5 8512.5 31707.5 ;
      RECT  8217.5 32502.5 8152.5 32637.5 ;
      RECT  8217.5 31527.5 8152.5 31662.5 ;
      RECT  8382.5 31785.0 8517.5 31850.0 ;
      RECT  8572.5 31925.0 8707.5 31990.0 ;
      RECT  8762.5 32065.0 8897.5 32130.0 ;
      RECT  8767.5 32412.5 8702.5 32547.5 ;
      RECT  8387.5 32412.5 8322.5 32547.5 ;
      RECT  8387.5 31572.5 8322.5 31707.5 ;
      RECT  8387.5 32030.0 8322.5 32165.0 ;
      RECT  8897.5 32065.0 8762.5 32130.0 ;
      RECT  8707.5 31925.0 8572.5 31990.0 ;
      RECT  8517.5 31785.0 8382.5 31850.0 ;
      RECT  8387.5 32030.0 8322.5 32165.0 ;
      RECT  9025.0 32722.5 8015.0 32787.5 ;
      RECT  9025.0 31377.5 8015.0 31442.5 ;
      RECT  8957.5 33937.5 8892.5 34132.5 ;
      RECT  8957.5 33097.5 8892.5 32722.5 ;
      RECT  8577.5 33097.5 8512.5 32722.5 ;
      RECT  8217.5 32940.0 8152.5 32755.0 ;
      RECT  8217.5 34100.0 8152.5 33915.0 ;
      RECT  8957.5 33097.5 8892.5 32962.5 ;
      RECT  8767.5 33097.5 8702.5 32962.5 ;
      RECT  8767.5 33097.5 8702.5 32962.5 ;
      RECT  8957.5 33097.5 8892.5 32962.5 ;
      RECT  8767.5 33097.5 8702.5 32962.5 ;
      RECT  8577.5 33097.5 8512.5 32962.5 ;
      RECT  8577.5 33097.5 8512.5 32962.5 ;
      RECT  8767.5 33097.5 8702.5 32962.5 ;
      RECT  8577.5 33097.5 8512.5 32962.5 ;
      RECT  8387.5 33097.5 8322.5 32962.5 ;
      RECT  8387.5 33097.5 8322.5 32962.5 ;
      RECT  8577.5 33097.5 8512.5 32962.5 ;
      RECT  8957.5 33937.5 8892.5 33802.5 ;
      RECT  8767.5 33937.5 8702.5 33802.5 ;
      RECT  8767.5 33937.5 8702.5 33802.5 ;
      RECT  8957.5 33937.5 8892.5 33802.5 ;
      RECT  8767.5 33937.5 8702.5 33802.5 ;
      RECT  8577.5 33937.5 8512.5 33802.5 ;
      RECT  8577.5 33937.5 8512.5 33802.5 ;
      RECT  8767.5 33937.5 8702.5 33802.5 ;
      RECT  8577.5 33937.5 8512.5 33802.5 ;
      RECT  8387.5 33937.5 8322.5 33802.5 ;
      RECT  8387.5 33937.5 8322.5 33802.5 ;
      RECT  8577.5 33937.5 8512.5 33802.5 ;
      RECT  8217.5 33007.5 8152.5 32872.5 ;
      RECT  8217.5 33982.5 8152.5 33847.5 ;
      RECT  8382.5 33725.0 8517.5 33660.0 ;
      RECT  8572.5 33585.0 8707.5 33520.0 ;
      RECT  8762.5 33445.0 8897.5 33380.0 ;
      RECT  8767.5 33097.5 8702.5 32962.5 ;
      RECT  8387.5 33097.5 8322.5 32962.5 ;
      RECT  8387.5 33937.5 8322.5 33802.5 ;
      RECT  8387.5 33480.0 8322.5 33345.0 ;
      RECT  8897.5 33445.0 8762.5 33380.0 ;
      RECT  8707.5 33585.0 8572.5 33520.0 ;
      RECT  8517.5 33725.0 8382.5 33660.0 ;
      RECT  8387.5 33480.0 8322.5 33345.0 ;
      RECT  9025.0 32787.5 8015.0 32722.5 ;
      RECT  9025.0 34132.5 8015.0 34067.5 ;
      RECT  10572.5 24457.5 10707.5 24522.5 ;
      RECT  12232.5 23935.0 12367.5 24000.0 ;
      RECT  10297.5 25802.5 10432.5 25867.5 ;
      RECT  11957.5 25370.0 12092.5 25435.0 ;
      RECT  10022.5 27147.5 10157.5 27212.5 ;
      RECT  11682.5 26625.0 11817.5 26690.0 ;
      RECT  12232.5 27477.5 12367.5 27542.5 ;
      RECT  9747.5 27477.5 9882.5 27542.5 ;
      RECT  11957.5 28822.5 12092.5 28887.5 ;
      RECT  9472.5 28822.5 9607.5 28887.5 ;
      RECT  11682.5 30167.5 11817.5 30232.5 ;
      RECT  9197.5 30167.5 9332.5 30232.5 ;
      RECT  10572.5 23995.0 10707.5 24060.0 ;
      RECT  10297.5 23855.0 10432.5 23920.0 ;
      RECT  10022.5 23715.0 10157.5 23780.0 ;
      RECT  9747.5 25310.0 9882.5 25375.0 ;
      RECT  10297.5 25450.0 10432.5 25515.0 ;
      RECT  10022.5 25590.0 10157.5 25655.0 ;
      RECT  10572.5 26685.0 10707.5 26750.0 ;
      RECT  9472.5 26545.0 9607.5 26610.0 ;
      RECT  10022.5 26405.0 10157.5 26470.0 ;
      RECT  9747.5 28000.0 9882.5 28065.0 ;
      RECT  9472.5 28140.0 9607.5 28205.0 ;
      RECT  10022.5 28280.0 10157.5 28345.0 ;
      RECT  10572.5 29375.0 10707.5 29440.0 ;
      RECT  10297.5 29235.0 10432.5 29300.0 ;
      RECT  9197.5 29095.0 9332.5 29160.0 ;
      RECT  9747.5 30690.0 9882.5 30755.0 ;
      RECT  10297.5 30830.0 10432.5 30895.0 ;
      RECT  9197.5 30970.0 9332.5 31035.0 ;
      RECT  10572.5 32065.0 10707.5 32130.0 ;
      RECT  9472.5 31925.0 9607.5 31990.0 ;
      RECT  9197.5 31785.0 9332.5 31850.0 ;
      RECT  9747.5 33380.0 9882.5 33445.0 ;
      RECT  9472.5 33520.0 9607.5 33585.0 ;
      RECT  9197.5 33660.0 9332.5 33725.0 ;
      RECT  7660.0 23935.0 7455.0 24000.0 ;
      RECT  7660.0 25370.0 7455.0 25435.0 ;
      RECT  7660.0 26625.0 7455.0 26690.0 ;
      RECT  7660.0 28060.0 7455.0 28125.0 ;
      RECT  7660.0 29315.0 7455.0 29380.0 ;
      RECT  7660.0 30750.0 7455.0 30815.0 ;
      RECT  7660.0 32005.0 7455.0 32070.0 ;
      RECT  7660.0 33440.0 7455.0 33505.0 ;
      RECT  12335.0 24652.5 7455.0 24717.5 ;
      RECT  12335.0 27342.5 7455.0 27407.5 ;
      RECT  12335.0 30032.5 7455.0 30097.5 ;
      RECT  12335.0 32722.5 7455.0 32787.5 ;
      RECT  12335.0 23307.5 7455.0 23372.5 ;
      RECT  12335.0 25997.5 7455.0 26062.5 ;
      RECT  12335.0 28687.5 7455.0 28752.5 ;
      RECT  12335.0 31377.5 7455.0 31442.5 ;
      RECT  12335.0 34067.5 7455.0 34132.5 ;
      RECT  7522.5 34262.5 7587.5 34067.5 ;
      RECT  7522.5 35102.5 7587.5 35477.5 ;
      RECT  7902.5 35102.5 7967.5 35477.5 ;
      RECT  8262.5 35260.0 8327.5 35445.0 ;
      RECT  8262.5 34100.0 8327.5 34285.0 ;
      RECT  7522.5 35102.5 7587.5 35237.5 ;
      RECT  7712.5 35102.5 7777.5 35237.5 ;
      RECT  7712.5 35102.5 7777.5 35237.5 ;
      RECT  7522.5 35102.5 7587.5 35237.5 ;
      RECT  7712.5 35102.5 7777.5 35237.5 ;
      RECT  7902.5 35102.5 7967.5 35237.5 ;
      RECT  7902.5 35102.5 7967.5 35237.5 ;
      RECT  7712.5 35102.5 7777.5 35237.5 ;
      RECT  7902.5 35102.5 7967.5 35237.5 ;
      RECT  8092.5 35102.5 8157.5 35237.5 ;
      RECT  8092.5 35102.5 8157.5 35237.5 ;
      RECT  7902.5 35102.5 7967.5 35237.5 ;
      RECT  7522.5 34262.5 7587.5 34397.5 ;
      RECT  7712.5 34262.5 7777.5 34397.5 ;
      RECT  7712.5 34262.5 7777.5 34397.5 ;
      RECT  7522.5 34262.5 7587.5 34397.5 ;
      RECT  7712.5 34262.5 7777.5 34397.5 ;
      RECT  7902.5 34262.5 7967.5 34397.5 ;
      RECT  7902.5 34262.5 7967.5 34397.5 ;
      RECT  7712.5 34262.5 7777.5 34397.5 ;
      RECT  7902.5 34262.5 7967.5 34397.5 ;
      RECT  8092.5 34262.5 8157.5 34397.5 ;
      RECT  8092.5 34262.5 8157.5 34397.5 ;
      RECT  7902.5 34262.5 7967.5 34397.5 ;
      RECT  8262.5 35192.5 8327.5 35327.5 ;
      RECT  8262.5 34217.5 8327.5 34352.5 ;
      RECT  8097.5 34475.0 7962.5 34540.0 ;
      RECT  7907.5 34615.0 7772.5 34680.0 ;
      RECT  7717.5 34755.0 7582.5 34820.0 ;
      RECT  7712.5 35102.5 7777.5 35237.5 ;
      RECT  8092.5 35102.5 8157.5 35237.5 ;
      RECT  8092.5 34262.5 8157.5 34397.5 ;
      RECT  8092.5 34720.0 8157.5 34855.0 ;
      RECT  7582.5 34755.0 7717.5 34820.0 ;
      RECT  7772.5 34615.0 7907.5 34680.0 ;
      RECT  7962.5 34475.0 8097.5 34540.0 ;
      RECT  8092.5 34720.0 8157.5 34855.0 ;
      RECT  7455.0 35412.5 8465.0 35477.5 ;
      RECT  7455.0 34067.5 8465.0 34132.5 ;
      RECT  7522.5 36627.5 7587.5 36822.5 ;
      RECT  7522.5 35787.5 7587.5 35412.5 ;
      RECT  7902.5 35787.5 7967.5 35412.5 ;
      RECT  8262.5 35630.0 8327.5 35445.0 ;
      RECT  8262.5 36790.0 8327.5 36605.0 ;
      RECT  7522.5 35787.5 7587.5 35652.5 ;
      RECT  7712.5 35787.5 7777.5 35652.5 ;
      RECT  7712.5 35787.5 7777.5 35652.5 ;
      RECT  7522.5 35787.5 7587.5 35652.5 ;
      RECT  7712.5 35787.5 7777.5 35652.5 ;
      RECT  7902.5 35787.5 7967.5 35652.5 ;
      RECT  7902.5 35787.5 7967.5 35652.5 ;
      RECT  7712.5 35787.5 7777.5 35652.5 ;
      RECT  7902.5 35787.5 7967.5 35652.5 ;
      RECT  8092.5 35787.5 8157.5 35652.5 ;
      RECT  8092.5 35787.5 8157.5 35652.5 ;
      RECT  7902.5 35787.5 7967.5 35652.5 ;
      RECT  7522.5 36627.5 7587.5 36492.5 ;
      RECT  7712.5 36627.5 7777.5 36492.5 ;
      RECT  7712.5 36627.5 7777.5 36492.5 ;
      RECT  7522.5 36627.5 7587.5 36492.5 ;
      RECT  7712.5 36627.5 7777.5 36492.5 ;
      RECT  7902.5 36627.5 7967.5 36492.5 ;
      RECT  7902.5 36627.5 7967.5 36492.5 ;
      RECT  7712.5 36627.5 7777.5 36492.5 ;
      RECT  7902.5 36627.5 7967.5 36492.5 ;
      RECT  8092.5 36627.5 8157.5 36492.5 ;
      RECT  8092.5 36627.5 8157.5 36492.5 ;
      RECT  7902.5 36627.5 7967.5 36492.5 ;
      RECT  8262.5 35697.5 8327.5 35562.5 ;
      RECT  8262.5 36672.5 8327.5 36537.5 ;
      RECT  8097.5 36415.0 7962.5 36350.0 ;
      RECT  7907.5 36275.0 7772.5 36210.0 ;
      RECT  7717.5 36135.0 7582.5 36070.0 ;
      RECT  7712.5 35787.5 7777.5 35652.5 ;
      RECT  8092.5 35787.5 8157.5 35652.5 ;
      RECT  8092.5 36627.5 8157.5 36492.5 ;
      RECT  8092.5 36170.0 8157.5 36035.0 ;
      RECT  7582.5 36135.0 7717.5 36070.0 ;
      RECT  7772.5 36275.0 7907.5 36210.0 ;
      RECT  7962.5 36415.0 8097.5 36350.0 ;
      RECT  8092.5 36170.0 8157.5 36035.0 ;
      RECT  7455.0 35477.5 8465.0 35412.5 ;
      RECT  7455.0 36822.5 8465.0 36757.5 ;
      RECT  7522.5 36952.5 7587.5 36757.5 ;
      RECT  7522.5 37792.5 7587.5 38167.5 ;
      RECT  7902.5 37792.5 7967.5 38167.5 ;
      RECT  8262.5 37950.0 8327.5 38135.0 ;
      RECT  8262.5 36790.0 8327.5 36975.0 ;
      RECT  7522.5 37792.5 7587.5 37927.5 ;
      RECT  7712.5 37792.5 7777.5 37927.5 ;
      RECT  7712.5 37792.5 7777.5 37927.5 ;
      RECT  7522.5 37792.5 7587.5 37927.5 ;
      RECT  7712.5 37792.5 7777.5 37927.5 ;
      RECT  7902.5 37792.5 7967.5 37927.5 ;
      RECT  7902.5 37792.5 7967.5 37927.5 ;
      RECT  7712.5 37792.5 7777.5 37927.5 ;
      RECT  7902.5 37792.5 7967.5 37927.5 ;
      RECT  8092.5 37792.5 8157.5 37927.5 ;
      RECT  8092.5 37792.5 8157.5 37927.5 ;
      RECT  7902.5 37792.5 7967.5 37927.5 ;
      RECT  7522.5 36952.5 7587.5 37087.5 ;
      RECT  7712.5 36952.5 7777.5 37087.5 ;
      RECT  7712.5 36952.5 7777.5 37087.5 ;
      RECT  7522.5 36952.5 7587.5 37087.5 ;
      RECT  7712.5 36952.5 7777.5 37087.5 ;
      RECT  7902.5 36952.5 7967.5 37087.5 ;
      RECT  7902.5 36952.5 7967.5 37087.5 ;
      RECT  7712.5 36952.5 7777.5 37087.5 ;
      RECT  7902.5 36952.5 7967.5 37087.5 ;
      RECT  8092.5 36952.5 8157.5 37087.5 ;
      RECT  8092.5 36952.5 8157.5 37087.5 ;
      RECT  7902.5 36952.5 7967.5 37087.5 ;
      RECT  8262.5 37882.5 8327.5 38017.5 ;
      RECT  8262.5 36907.5 8327.5 37042.5 ;
      RECT  8097.5 37165.0 7962.5 37230.0 ;
      RECT  7907.5 37305.0 7772.5 37370.0 ;
      RECT  7717.5 37445.0 7582.5 37510.0 ;
      RECT  7712.5 37792.5 7777.5 37927.5 ;
      RECT  8092.5 37792.5 8157.5 37927.5 ;
      RECT  8092.5 36952.5 8157.5 37087.5 ;
      RECT  8092.5 37410.0 8157.5 37545.0 ;
      RECT  7582.5 37445.0 7717.5 37510.0 ;
      RECT  7772.5 37305.0 7907.5 37370.0 ;
      RECT  7962.5 37165.0 8097.5 37230.0 ;
      RECT  8092.5 37410.0 8157.5 37545.0 ;
      RECT  7455.0 38102.5 8465.0 38167.5 ;
      RECT  7455.0 36757.5 8465.0 36822.5 ;
      RECT  7522.5 39317.5 7587.5 39512.5 ;
      RECT  7522.5 38477.5 7587.5 38102.5 ;
      RECT  7902.5 38477.5 7967.5 38102.5 ;
      RECT  8262.5 38320.0 8327.5 38135.0 ;
      RECT  8262.5 39480.0 8327.5 39295.0 ;
      RECT  7522.5 38477.5 7587.5 38342.5 ;
      RECT  7712.5 38477.5 7777.5 38342.5 ;
      RECT  7712.5 38477.5 7777.5 38342.5 ;
      RECT  7522.5 38477.5 7587.5 38342.5 ;
      RECT  7712.5 38477.5 7777.5 38342.5 ;
      RECT  7902.5 38477.5 7967.5 38342.5 ;
      RECT  7902.5 38477.5 7967.5 38342.5 ;
      RECT  7712.5 38477.5 7777.5 38342.5 ;
      RECT  7902.5 38477.5 7967.5 38342.5 ;
      RECT  8092.5 38477.5 8157.5 38342.5 ;
      RECT  8092.5 38477.5 8157.5 38342.5 ;
      RECT  7902.5 38477.5 7967.5 38342.5 ;
      RECT  7522.5 39317.5 7587.5 39182.5 ;
      RECT  7712.5 39317.5 7777.5 39182.5 ;
      RECT  7712.5 39317.5 7777.5 39182.5 ;
      RECT  7522.5 39317.5 7587.5 39182.5 ;
      RECT  7712.5 39317.5 7777.5 39182.5 ;
      RECT  7902.5 39317.5 7967.5 39182.5 ;
      RECT  7902.5 39317.5 7967.5 39182.5 ;
      RECT  7712.5 39317.5 7777.5 39182.5 ;
      RECT  7902.5 39317.5 7967.5 39182.5 ;
      RECT  8092.5 39317.5 8157.5 39182.5 ;
      RECT  8092.5 39317.5 8157.5 39182.5 ;
      RECT  7902.5 39317.5 7967.5 39182.5 ;
      RECT  8262.5 38387.5 8327.5 38252.5 ;
      RECT  8262.5 39362.5 8327.5 39227.5 ;
      RECT  8097.5 39105.0 7962.5 39040.0 ;
      RECT  7907.5 38965.0 7772.5 38900.0 ;
      RECT  7717.5 38825.0 7582.5 38760.0 ;
      RECT  7712.5 38477.5 7777.5 38342.5 ;
      RECT  8092.5 38477.5 8157.5 38342.5 ;
      RECT  8092.5 39317.5 8157.5 39182.5 ;
      RECT  8092.5 38860.0 8157.5 38725.0 ;
      RECT  7582.5 38825.0 7717.5 38760.0 ;
      RECT  7772.5 38965.0 7907.5 38900.0 ;
      RECT  7962.5 39105.0 8097.5 39040.0 ;
      RECT  8092.5 38860.0 8157.5 38725.0 ;
      RECT  7455.0 38167.5 8465.0 38102.5 ;
      RECT  7455.0 39512.5 8465.0 39447.5 ;
      RECT  7522.5 39642.5 7587.5 39447.5 ;
      RECT  7522.5 40482.5 7587.5 40857.5 ;
      RECT  7902.5 40482.5 7967.5 40857.5 ;
      RECT  8262.5 40640.0 8327.5 40825.0 ;
      RECT  8262.5 39480.0 8327.5 39665.0 ;
      RECT  7522.5 40482.5 7587.5 40617.5 ;
      RECT  7712.5 40482.5 7777.5 40617.5 ;
      RECT  7712.5 40482.5 7777.5 40617.5 ;
      RECT  7522.5 40482.5 7587.5 40617.5 ;
      RECT  7712.5 40482.5 7777.5 40617.5 ;
      RECT  7902.5 40482.5 7967.5 40617.5 ;
      RECT  7902.5 40482.5 7967.5 40617.5 ;
      RECT  7712.5 40482.5 7777.5 40617.5 ;
      RECT  7902.5 40482.5 7967.5 40617.5 ;
      RECT  8092.5 40482.5 8157.5 40617.5 ;
      RECT  8092.5 40482.5 8157.5 40617.5 ;
      RECT  7902.5 40482.5 7967.5 40617.5 ;
      RECT  7522.5 39642.5 7587.5 39777.5 ;
      RECT  7712.5 39642.5 7777.5 39777.5 ;
      RECT  7712.5 39642.5 7777.5 39777.5 ;
      RECT  7522.5 39642.5 7587.5 39777.5 ;
      RECT  7712.5 39642.5 7777.5 39777.5 ;
      RECT  7902.5 39642.5 7967.5 39777.5 ;
      RECT  7902.5 39642.5 7967.5 39777.5 ;
      RECT  7712.5 39642.5 7777.5 39777.5 ;
      RECT  7902.5 39642.5 7967.5 39777.5 ;
      RECT  8092.5 39642.5 8157.5 39777.5 ;
      RECT  8092.5 39642.5 8157.5 39777.5 ;
      RECT  7902.5 39642.5 7967.5 39777.5 ;
      RECT  8262.5 40572.5 8327.5 40707.5 ;
      RECT  8262.5 39597.5 8327.5 39732.5 ;
      RECT  8097.5 39855.0 7962.5 39920.0 ;
      RECT  7907.5 39995.0 7772.5 40060.0 ;
      RECT  7717.5 40135.0 7582.5 40200.0 ;
      RECT  7712.5 40482.5 7777.5 40617.5 ;
      RECT  8092.5 40482.5 8157.5 40617.5 ;
      RECT  8092.5 39642.5 8157.5 39777.5 ;
      RECT  8092.5 40100.0 8157.5 40235.0 ;
      RECT  7582.5 40135.0 7717.5 40200.0 ;
      RECT  7772.5 39995.0 7907.5 40060.0 ;
      RECT  7962.5 39855.0 8097.5 39920.0 ;
      RECT  8092.5 40100.0 8157.5 40235.0 ;
      RECT  7455.0 40792.5 8465.0 40857.5 ;
      RECT  7455.0 39447.5 8465.0 39512.5 ;
      RECT  7522.5 42007.5 7587.5 42202.5 ;
      RECT  7522.5 41167.5 7587.5 40792.5 ;
      RECT  7902.5 41167.5 7967.5 40792.5 ;
      RECT  8262.5 41010.0 8327.5 40825.0 ;
      RECT  8262.5 42170.0 8327.5 41985.0 ;
      RECT  7522.5 41167.5 7587.5 41032.5 ;
      RECT  7712.5 41167.5 7777.5 41032.5 ;
      RECT  7712.5 41167.5 7777.5 41032.5 ;
      RECT  7522.5 41167.5 7587.5 41032.5 ;
      RECT  7712.5 41167.5 7777.5 41032.5 ;
      RECT  7902.5 41167.5 7967.5 41032.5 ;
      RECT  7902.5 41167.5 7967.5 41032.5 ;
      RECT  7712.5 41167.5 7777.5 41032.5 ;
      RECT  7902.5 41167.5 7967.5 41032.5 ;
      RECT  8092.5 41167.5 8157.5 41032.5 ;
      RECT  8092.5 41167.5 8157.5 41032.5 ;
      RECT  7902.5 41167.5 7967.5 41032.5 ;
      RECT  7522.5 42007.5 7587.5 41872.5 ;
      RECT  7712.5 42007.5 7777.5 41872.5 ;
      RECT  7712.5 42007.5 7777.5 41872.5 ;
      RECT  7522.5 42007.5 7587.5 41872.5 ;
      RECT  7712.5 42007.5 7777.5 41872.5 ;
      RECT  7902.5 42007.5 7967.5 41872.5 ;
      RECT  7902.5 42007.5 7967.5 41872.5 ;
      RECT  7712.5 42007.5 7777.5 41872.5 ;
      RECT  7902.5 42007.5 7967.5 41872.5 ;
      RECT  8092.5 42007.5 8157.5 41872.5 ;
      RECT  8092.5 42007.5 8157.5 41872.5 ;
      RECT  7902.5 42007.5 7967.5 41872.5 ;
      RECT  8262.5 41077.5 8327.5 40942.5 ;
      RECT  8262.5 42052.5 8327.5 41917.5 ;
      RECT  8097.5 41795.0 7962.5 41730.0 ;
      RECT  7907.5 41655.0 7772.5 41590.0 ;
      RECT  7717.5 41515.0 7582.5 41450.0 ;
      RECT  7712.5 41167.5 7777.5 41032.5 ;
      RECT  8092.5 41167.5 8157.5 41032.5 ;
      RECT  8092.5 42007.5 8157.5 41872.5 ;
      RECT  8092.5 41550.0 8157.5 41415.0 ;
      RECT  7582.5 41515.0 7717.5 41450.0 ;
      RECT  7772.5 41655.0 7907.5 41590.0 ;
      RECT  7962.5 41795.0 8097.5 41730.0 ;
      RECT  8092.5 41550.0 8157.5 41415.0 ;
      RECT  7455.0 40857.5 8465.0 40792.5 ;
      RECT  7455.0 42202.5 8465.0 42137.5 ;
      RECT  7522.5 42332.5 7587.5 42137.5 ;
      RECT  7522.5 43172.5 7587.5 43547.5 ;
      RECT  7902.5 43172.5 7967.5 43547.5 ;
      RECT  8262.5 43330.0 8327.5 43515.0 ;
      RECT  8262.5 42170.0 8327.5 42355.0 ;
      RECT  7522.5 43172.5 7587.5 43307.5 ;
      RECT  7712.5 43172.5 7777.5 43307.5 ;
      RECT  7712.5 43172.5 7777.5 43307.5 ;
      RECT  7522.5 43172.5 7587.5 43307.5 ;
      RECT  7712.5 43172.5 7777.5 43307.5 ;
      RECT  7902.5 43172.5 7967.5 43307.5 ;
      RECT  7902.5 43172.5 7967.5 43307.5 ;
      RECT  7712.5 43172.5 7777.5 43307.5 ;
      RECT  7902.5 43172.5 7967.5 43307.5 ;
      RECT  8092.5 43172.5 8157.5 43307.5 ;
      RECT  8092.5 43172.5 8157.5 43307.5 ;
      RECT  7902.5 43172.5 7967.5 43307.5 ;
      RECT  7522.5 42332.5 7587.5 42467.5 ;
      RECT  7712.5 42332.5 7777.5 42467.5 ;
      RECT  7712.5 42332.5 7777.5 42467.5 ;
      RECT  7522.5 42332.5 7587.5 42467.5 ;
      RECT  7712.5 42332.5 7777.5 42467.5 ;
      RECT  7902.5 42332.5 7967.5 42467.5 ;
      RECT  7902.5 42332.5 7967.5 42467.5 ;
      RECT  7712.5 42332.5 7777.5 42467.5 ;
      RECT  7902.5 42332.5 7967.5 42467.5 ;
      RECT  8092.5 42332.5 8157.5 42467.5 ;
      RECT  8092.5 42332.5 8157.5 42467.5 ;
      RECT  7902.5 42332.5 7967.5 42467.5 ;
      RECT  8262.5 43262.5 8327.5 43397.5 ;
      RECT  8262.5 42287.5 8327.5 42422.5 ;
      RECT  8097.5 42545.0 7962.5 42610.0 ;
      RECT  7907.5 42685.0 7772.5 42750.0 ;
      RECT  7717.5 42825.0 7582.5 42890.0 ;
      RECT  7712.5 43172.5 7777.5 43307.5 ;
      RECT  8092.5 43172.5 8157.5 43307.5 ;
      RECT  8092.5 42332.5 8157.5 42467.5 ;
      RECT  8092.5 42790.0 8157.5 42925.0 ;
      RECT  7582.5 42825.0 7717.5 42890.0 ;
      RECT  7772.5 42685.0 7907.5 42750.0 ;
      RECT  7962.5 42545.0 8097.5 42610.0 ;
      RECT  8092.5 42790.0 8157.5 42925.0 ;
      RECT  7455.0 43482.5 8465.0 43547.5 ;
      RECT  7455.0 42137.5 8465.0 42202.5 ;
      RECT  7522.5 44697.5 7587.5 44892.5 ;
      RECT  7522.5 43857.5 7587.5 43482.5 ;
      RECT  7902.5 43857.5 7967.5 43482.5 ;
      RECT  8262.5 43700.0 8327.5 43515.0 ;
      RECT  8262.5 44860.0 8327.5 44675.0 ;
      RECT  7522.5 43857.5 7587.5 43722.5 ;
      RECT  7712.5 43857.5 7777.5 43722.5 ;
      RECT  7712.5 43857.5 7777.5 43722.5 ;
      RECT  7522.5 43857.5 7587.5 43722.5 ;
      RECT  7712.5 43857.5 7777.5 43722.5 ;
      RECT  7902.5 43857.5 7967.5 43722.5 ;
      RECT  7902.5 43857.5 7967.5 43722.5 ;
      RECT  7712.5 43857.5 7777.5 43722.5 ;
      RECT  7902.5 43857.5 7967.5 43722.5 ;
      RECT  8092.5 43857.5 8157.5 43722.5 ;
      RECT  8092.5 43857.5 8157.5 43722.5 ;
      RECT  7902.5 43857.5 7967.5 43722.5 ;
      RECT  7522.5 44697.5 7587.5 44562.5 ;
      RECT  7712.5 44697.5 7777.5 44562.5 ;
      RECT  7712.5 44697.5 7777.5 44562.5 ;
      RECT  7522.5 44697.5 7587.5 44562.5 ;
      RECT  7712.5 44697.5 7777.5 44562.5 ;
      RECT  7902.5 44697.5 7967.5 44562.5 ;
      RECT  7902.5 44697.5 7967.5 44562.5 ;
      RECT  7712.5 44697.5 7777.5 44562.5 ;
      RECT  7902.5 44697.5 7967.5 44562.5 ;
      RECT  8092.5 44697.5 8157.5 44562.5 ;
      RECT  8092.5 44697.5 8157.5 44562.5 ;
      RECT  7902.5 44697.5 7967.5 44562.5 ;
      RECT  8262.5 43767.5 8327.5 43632.5 ;
      RECT  8262.5 44742.5 8327.5 44607.5 ;
      RECT  8097.5 44485.0 7962.5 44420.0 ;
      RECT  7907.5 44345.0 7772.5 44280.0 ;
      RECT  7717.5 44205.0 7582.5 44140.0 ;
      RECT  7712.5 43857.5 7777.5 43722.5 ;
      RECT  8092.5 43857.5 8157.5 43722.5 ;
      RECT  8092.5 44697.5 8157.5 44562.5 ;
      RECT  8092.5 44240.0 8157.5 44105.0 ;
      RECT  7582.5 44205.0 7717.5 44140.0 ;
      RECT  7772.5 44345.0 7907.5 44280.0 ;
      RECT  7962.5 44485.0 8097.5 44420.0 ;
      RECT  8092.5 44240.0 8157.5 44105.0 ;
      RECT  7455.0 43547.5 8465.0 43482.5 ;
      RECT  7455.0 44892.5 8465.0 44827.5 ;
      RECT  7522.5 45022.5 7587.5 44827.5 ;
      RECT  7522.5 45862.5 7587.5 46237.5 ;
      RECT  7902.5 45862.5 7967.5 46237.5 ;
      RECT  8262.5 46020.0 8327.5 46205.0 ;
      RECT  8262.5 44860.0 8327.5 45045.0 ;
      RECT  7522.5 45862.5 7587.5 45997.5 ;
      RECT  7712.5 45862.5 7777.5 45997.5 ;
      RECT  7712.5 45862.5 7777.5 45997.5 ;
      RECT  7522.5 45862.5 7587.5 45997.5 ;
      RECT  7712.5 45862.5 7777.5 45997.5 ;
      RECT  7902.5 45862.5 7967.5 45997.5 ;
      RECT  7902.5 45862.5 7967.5 45997.5 ;
      RECT  7712.5 45862.5 7777.5 45997.5 ;
      RECT  7902.5 45862.5 7967.5 45997.5 ;
      RECT  8092.5 45862.5 8157.5 45997.5 ;
      RECT  8092.5 45862.5 8157.5 45997.5 ;
      RECT  7902.5 45862.5 7967.5 45997.5 ;
      RECT  7522.5 45022.5 7587.5 45157.5 ;
      RECT  7712.5 45022.5 7777.5 45157.5 ;
      RECT  7712.5 45022.5 7777.5 45157.5 ;
      RECT  7522.5 45022.5 7587.5 45157.5 ;
      RECT  7712.5 45022.5 7777.5 45157.5 ;
      RECT  7902.5 45022.5 7967.5 45157.5 ;
      RECT  7902.5 45022.5 7967.5 45157.5 ;
      RECT  7712.5 45022.5 7777.5 45157.5 ;
      RECT  7902.5 45022.5 7967.5 45157.5 ;
      RECT  8092.5 45022.5 8157.5 45157.5 ;
      RECT  8092.5 45022.5 8157.5 45157.5 ;
      RECT  7902.5 45022.5 7967.5 45157.5 ;
      RECT  8262.5 45952.5 8327.5 46087.5 ;
      RECT  8262.5 44977.5 8327.5 45112.5 ;
      RECT  8097.5 45235.0 7962.5 45300.0 ;
      RECT  7907.5 45375.0 7772.5 45440.0 ;
      RECT  7717.5 45515.0 7582.5 45580.0 ;
      RECT  7712.5 45862.5 7777.5 45997.5 ;
      RECT  8092.5 45862.5 8157.5 45997.5 ;
      RECT  8092.5 45022.5 8157.5 45157.5 ;
      RECT  8092.5 45480.0 8157.5 45615.0 ;
      RECT  7582.5 45515.0 7717.5 45580.0 ;
      RECT  7772.5 45375.0 7907.5 45440.0 ;
      RECT  7962.5 45235.0 8097.5 45300.0 ;
      RECT  8092.5 45480.0 8157.5 45615.0 ;
      RECT  7455.0 46172.5 8465.0 46237.5 ;
      RECT  7455.0 44827.5 8465.0 44892.5 ;
      RECT  7522.5 47387.5 7587.5 47582.5 ;
      RECT  7522.5 46547.5 7587.5 46172.5 ;
      RECT  7902.5 46547.5 7967.5 46172.5 ;
      RECT  8262.5 46390.0 8327.5 46205.0 ;
      RECT  8262.5 47550.0 8327.5 47365.0 ;
      RECT  7522.5 46547.5 7587.5 46412.5 ;
      RECT  7712.5 46547.5 7777.5 46412.5 ;
      RECT  7712.5 46547.5 7777.5 46412.5 ;
      RECT  7522.5 46547.5 7587.5 46412.5 ;
      RECT  7712.5 46547.5 7777.5 46412.5 ;
      RECT  7902.5 46547.5 7967.5 46412.5 ;
      RECT  7902.5 46547.5 7967.5 46412.5 ;
      RECT  7712.5 46547.5 7777.5 46412.5 ;
      RECT  7902.5 46547.5 7967.5 46412.5 ;
      RECT  8092.5 46547.5 8157.5 46412.5 ;
      RECT  8092.5 46547.5 8157.5 46412.5 ;
      RECT  7902.5 46547.5 7967.5 46412.5 ;
      RECT  7522.5 47387.5 7587.5 47252.5 ;
      RECT  7712.5 47387.5 7777.5 47252.5 ;
      RECT  7712.5 47387.5 7777.5 47252.5 ;
      RECT  7522.5 47387.5 7587.5 47252.5 ;
      RECT  7712.5 47387.5 7777.5 47252.5 ;
      RECT  7902.5 47387.5 7967.5 47252.5 ;
      RECT  7902.5 47387.5 7967.5 47252.5 ;
      RECT  7712.5 47387.5 7777.5 47252.5 ;
      RECT  7902.5 47387.5 7967.5 47252.5 ;
      RECT  8092.5 47387.5 8157.5 47252.5 ;
      RECT  8092.5 47387.5 8157.5 47252.5 ;
      RECT  7902.5 47387.5 7967.5 47252.5 ;
      RECT  8262.5 46457.5 8327.5 46322.5 ;
      RECT  8262.5 47432.5 8327.5 47297.5 ;
      RECT  8097.5 47175.0 7962.5 47110.0 ;
      RECT  7907.5 47035.0 7772.5 46970.0 ;
      RECT  7717.5 46895.0 7582.5 46830.0 ;
      RECT  7712.5 46547.5 7777.5 46412.5 ;
      RECT  8092.5 46547.5 8157.5 46412.5 ;
      RECT  8092.5 47387.5 8157.5 47252.5 ;
      RECT  8092.5 46930.0 8157.5 46795.0 ;
      RECT  7582.5 46895.0 7717.5 46830.0 ;
      RECT  7772.5 47035.0 7907.5 46970.0 ;
      RECT  7962.5 47175.0 8097.5 47110.0 ;
      RECT  8092.5 46930.0 8157.5 46795.0 ;
      RECT  7455.0 46237.5 8465.0 46172.5 ;
      RECT  7455.0 47582.5 8465.0 47517.5 ;
      RECT  7522.5 47712.5 7587.5 47517.5 ;
      RECT  7522.5 48552.5 7587.5 48927.5 ;
      RECT  7902.5 48552.5 7967.5 48927.5 ;
      RECT  8262.5 48710.0 8327.5 48895.0 ;
      RECT  8262.5 47550.0 8327.5 47735.0 ;
      RECT  7522.5 48552.5 7587.5 48687.5 ;
      RECT  7712.5 48552.5 7777.5 48687.5 ;
      RECT  7712.5 48552.5 7777.5 48687.5 ;
      RECT  7522.5 48552.5 7587.5 48687.5 ;
      RECT  7712.5 48552.5 7777.5 48687.5 ;
      RECT  7902.5 48552.5 7967.5 48687.5 ;
      RECT  7902.5 48552.5 7967.5 48687.5 ;
      RECT  7712.5 48552.5 7777.5 48687.5 ;
      RECT  7902.5 48552.5 7967.5 48687.5 ;
      RECT  8092.5 48552.5 8157.5 48687.5 ;
      RECT  8092.5 48552.5 8157.5 48687.5 ;
      RECT  7902.5 48552.5 7967.5 48687.5 ;
      RECT  7522.5 47712.5 7587.5 47847.5 ;
      RECT  7712.5 47712.5 7777.5 47847.5 ;
      RECT  7712.5 47712.5 7777.5 47847.5 ;
      RECT  7522.5 47712.5 7587.5 47847.5 ;
      RECT  7712.5 47712.5 7777.5 47847.5 ;
      RECT  7902.5 47712.5 7967.5 47847.5 ;
      RECT  7902.5 47712.5 7967.5 47847.5 ;
      RECT  7712.5 47712.5 7777.5 47847.5 ;
      RECT  7902.5 47712.5 7967.5 47847.5 ;
      RECT  8092.5 47712.5 8157.5 47847.5 ;
      RECT  8092.5 47712.5 8157.5 47847.5 ;
      RECT  7902.5 47712.5 7967.5 47847.5 ;
      RECT  8262.5 48642.5 8327.5 48777.5 ;
      RECT  8262.5 47667.5 8327.5 47802.5 ;
      RECT  8097.5 47925.0 7962.5 47990.0 ;
      RECT  7907.5 48065.0 7772.5 48130.0 ;
      RECT  7717.5 48205.0 7582.5 48270.0 ;
      RECT  7712.5 48552.5 7777.5 48687.5 ;
      RECT  8092.5 48552.5 8157.5 48687.5 ;
      RECT  8092.5 47712.5 8157.5 47847.5 ;
      RECT  8092.5 48170.0 8157.5 48305.0 ;
      RECT  7582.5 48205.0 7717.5 48270.0 ;
      RECT  7772.5 48065.0 7907.5 48130.0 ;
      RECT  7962.5 47925.0 8097.5 47990.0 ;
      RECT  8092.5 48170.0 8157.5 48305.0 ;
      RECT  7455.0 48862.5 8465.0 48927.5 ;
      RECT  7455.0 47517.5 8465.0 47582.5 ;
      RECT  7522.5 50077.5 7587.5 50272.5 ;
      RECT  7522.5 49237.5 7587.5 48862.5 ;
      RECT  7902.5 49237.5 7967.5 48862.5 ;
      RECT  8262.5 49080.0 8327.5 48895.0 ;
      RECT  8262.5 50240.0 8327.5 50055.0 ;
      RECT  7522.5 49237.5 7587.5 49102.5 ;
      RECT  7712.5 49237.5 7777.5 49102.5 ;
      RECT  7712.5 49237.5 7777.5 49102.5 ;
      RECT  7522.5 49237.5 7587.5 49102.5 ;
      RECT  7712.5 49237.5 7777.5 49102.5 ;
      RECT  7902.5 49237.5 7967.5 49102.5 ;
      RECT  7902.5 49237.5 7967.5 49102.5 ;
      RECT  7712.5 49237.5 7777.5 49102.5 ;
      RECT  7902.5 49237.5 7967.5 49102.5 ;
      RECT  8092.5 49237.5 8157.5 49102.5 ;
      RECT  8092.5 49237.5 8157.5 49102.5 ;
      RECT  7902.5 49237.5 7967.5 49102.5 ;
      RECT  7522.5 50077.5 7587.5 49942.5 ;
      RECT  7712.5 50077.5 7777.5 49942.5 ;
      RECT  7712.5 50077.5 7777.5 49942.5 ;
      RECT  7522.5 50077.5 7587.5 49942.5 ;
      RECT  7712.5 50077.5 7777.5 49942.5 ;
      RECT  7902.5 50077.5 7967.5 49942.5 ;
      RECT  7902.5 50077.5 7967.5 49942.5 ;
      RECT  7712.5 50077.5 7777.5 49942.5 ;
      RECT  7902.5 50077.5 7967.5 49942.5 ;
      RECT  8092.5 50077.5 8157.5 49942.5 ;
      RECT  8092.5 50077.5 8157.5 49942.5 ;
      RECT  7902.5 50077.5 7967.5 49942.5 ;
      RECT  8262.5 49147.5 8327.5 49012.5 ;
      RECT  8262.5 50122.5 8327.5 49987.5 ;
      RECT  8097.5 49865.0 7962.5 49800.0 ;
      RECT  7907.5 49725.0 7772.5 49660.0 ;
      RECT  7717.5 49585.0 7582.5 49520.0 ;
      RECT  7712.5 49237.5 7777.5 49102.5 ;
      RECT  8092.5 49237.5 8157.5 49102.5 ;
      RECT  8092.5 50077.5 8157.5 49942.5 ;
      RECT  8092.5 49620.0 8157.5 49485.0 ;
      RECT  7582.5 49585.0 7717.5 49520.0 ;
      RECT  7772.5 49725.0 7907.5 49660.0 ;
      RECT  7962.5 49865.0 8097.5 49800.0 ;
      RECT  8092.5 49620.0 8157.5 49485.0 ;
      RECT  7455.0 48927.5 8465.0 48862.5 ;
      RECT  7455.0 50272.5 8465.0 50207.5 ;
      RECT  7522.5 50402.5 7587.5 50207.5 ;
      RECT  7522.5 51242.5 7587.5 51617.5 ;
      RECT  7902.5 51242.5 7967.5 51617.5 ;
      RECT  8262.5 51400.0 8327.5 51585.0 ;
      RECT  8262.5 50240.0 8327.5 50425.0 ;
      RECT  7522.5 51242.5 7587.5 51377.5 ;
      RECT  7712.5 51242.5 7777.5 51377.5 ;
      RECT  7712.5 51242.5 7777.5 51377.5 ;
      RECT  7522.5 51242.5 7587.5 51377.5 ;
      RECT  7712.5 51242.5 7777.5 51377.5 ;
      RECT  7902.5 51242.5 7967.5 51377.5 ;
      RECT  7902.5 51242.5 7967.5 51377.5 ;
      RECT  7712.5 51242.5 7777.5 51377.5 ;
      RECT  7902.5 51242.5 7967.5 51377.5 ;
      RECT  8092.5 51242.5 8157.5 51377.5 ;
      RECT  8092.5 51242.5 8157.5 51377.5 ;
      RECT  7902.5 51242.5 7967.5 51377.5 ;
      RECT  7522.5 50402.5 7587.5 50537.5 ;
      RECT  7712.5 50402.5 7777.5 50537.5 ;
      RECT  7712.5 50402.5 7777.5 50537.5 ;
      RECT  7522.5 50402.5 7587.5 50537.5 ;
      RECT  7712.5 50402.5 7777.5 50537.5 ;
      RECT  7902.5 50402.5 7967.5 50537.5 ;
      RECT  7902.5 50402.5 7967.5 50537.5 ;
      RECT  7712.5 50402.5 7777.5 50537.5 ;
      RECT  7902.5 50402.5 7967.5 50537.5 ;
      RECT  8092.5 50402.5 8157.5 50537.5 ;
      RECT  8092.5 50402.5 8157.5 50537.5 ;
      RECT  7902.5 50402.5 7967.5 50537.5 ;
      RECT  8262.5 51332.5 8327.5 51467.5 ;
      RECT  8262.5 50357.5 8327.5 50492.5 ;
      RECT  8097.5 50615.0 7962.5 50680.0 ;
      RECT  7907.5 50755.0 7772.5 50820.0 ;
      RECT  7717.5 50895.0 7582.5 50960.0 ;
      RECT  7712.5 51242.5 7777.5 51377.5 ;
      RECT  8092.5 51242.5 8157.5 51377.5 ;
      RECT  8092.5 50402.5 8157.5 50537.5 ;
      RECT  8092.5 50860.0 8157.5 50995.0 ;
      RECT  7582.5 50895.0 7717.5 50960.0 ;
      RECT  7772.5 50755.0 7907.5 50820.0 ;
      RECT  7962.5 50615.0 8097.5 50680.0 ;
      RECT  8092.5 50860.0 8157.5 50995.0 ;
      RECT  7455.0 51552.5 8465.0 51617.5 ;
      RECT  7455.0 50207.5 8465.0 50272.5 ;
      RECT  7522.5 52767.5 7587.5 52962.5 ;
      RECT  7522.5 51927.5 7587.5 51552.5 ;
      RECT  7902.5 51927.5 7967.5 51552.5 ;
      RECT  8262.5 51770.0 8327.5 51585.0 ;
      RECT  8262.5 52930.0 8327.5 52745.0 ;
      RECT  7522.5 51927.5 7587.5 51792.5 ;
      RECT  7712.5 51927.5 7777.5 51792.5 ;
      RECT  7712.5 51927.5 7777.5 51792.5 ;
      RECT  7522.5 51927.5 7587.5 51792.5 ;
      RECT  7712.5 51927.5 7777.5 51792.5 ;
      RECT  7902.5 51927.5 7967.5 51792.5 ;
      RECT  7902.5 51927.5 7967.5 51792.5 ;
      RECT  7712.5 51927.5 7777.5 51792.5 ;
      RECT  7902.5 51927.5 7967.5 51792.5 ;
      RECT  8092.5 51927.5 8157.5 51792.5 ;
      RECT  8092.5 51927.5 8157.5 51792.5 ;
      RECT  7902.5 51927.5 7967.5 51792.5 ;
      RECT  7522.5 52767.5 7587.5 52632.5 ;
      RECT  7712.5 52767.5 7777.5 52632.5 ;
      RECT  7712.5 52767.5 7777.5 52632.5 ;
      RECT  7522.5 52767.5 7587.5 52632.5 ;
      RECT  7712.5 52767.5 7777.5 52632.5 ;
      RECT  7902.5 52767.5 7967.5 52632.5 ;
      RECT  7902.5 52767.5 7967.5 52632.5 ;
      RECT  7712.5 52767.5 7777.5 52632.5 ;
      RECT  7902.5 52767.5 7967.5 52632.5 ;
      RECT  8092.5 52767.5 8157.5 52632.5 ;
      RECT  8092.5 52767.5 8157.5 52632.5 ;
      RECT  7902.5 52767.5 7967.5 52632.5 ;
      RECT  8262.5 51837.5 8327.5 51702.5 ;
      RECT  8262.5 52812.5 8327.5 52677.5 ;
      RECT  8097.5 52555.0 7962.5 52490.0 ;
      RECT  7907.5 52415.0 7772.5 52350.0 ;
      RECT  7717.5 52275.0 7582.5 52210.0 ;
      RECT  7712.5 51927.5 7777.5 51792.5 ;
      RECT  8092.5 51927.5 8157.5 51792.5 ;
      RECT  8092.5 52767.5 8157.5 52632.5 ;
      RECT  8092.5 52310.0 8157.5 52175.0 ;
      RECT  7582.5 52275.0 7717.5 52210.0 ;
      RECT  7772.5 52415.0 7907.5 52350.0 ;
      RECT  7962.5 52555.0 8097.5 52490.0 ;
      RECT  8092.5 52310.0 8157.5 52175.0 ;
      RECT  7455.0 51617.5 8465.0 51552.5 ;
      RECT  7455.0 52962.5 8465.0 52897.5 ;
      RECT  7522.5 53092.5 7587.5 52897.5 ;
      RECT  7522.5 53932.5 7587.5 54307.5 ;
      RECT  7902.5 53932.5 7967.5 54307.5 ;
      RECT  8262.5 54090.0 8327.5 54275.0 ;
      RECT  8262.5 52930.0 8327.5 53115.0 ;
      RECT  7522.5 53932.5 7587.5 54067.5 ;
      RECT  7712.5 53932.5 7777.5 54067.5 ;
      RECT  7712.5 53932.5 7777.5 54067.5 ;
      RECT  7522.5 53932.5 7587.5 54067.5 ;
      RECT  7712.5 53932.5 7777.5 54067.5 ;
      RECT  7902.5 53932.5 7967.5 54067.5 ;
      RECT  7902.5 53932.5 7967.5 54067.5 ;
      RECT  7712.5 53932.5 7777.5 54067.5 ;
      RECT  7902.5 53932.5 7967.5 54067.5 ;
      RECT  8092.5 53932.5 8157.5 54067.5 ;
      RECT  8092.5 53932.5 8157.5 54067.5 ;
      RECT  7902.5 53932.5 7967.5 54067.5 ;
      RECT  7522.5 53092.5 7587.5 53227.5 ;
      RECT  7712.5 53092.5 7777.5 53227.5 ;
      RECT  7712.5 53092.5 7777.5 53227.5 ;
      RECT  7522.5 53092.5 7587.5 53227.5 ;
      RECT  7712.5 53092.5 7777.5 53227.5 ;
      RECT  7902.5 53092.5 7967.5 53227.5 ;
      RECT  7902.5 53092.5 7967.5 53227.5 ;
      RECT  7712.5 53092.5 7777.5 53227.5 ;
      RECT  7902.5 53092.5 7967.5 53227.5 ;
      RECT  8092.5 53092.5 8157.5 53227.5 ;
      RECT  8092.5 53092.5 8157.5 53227.5 ;
      RECT  7902.5 53092.5 7967.5 53227.5 ;
      RECT  8262.5 54022.5 8327.5 54157.5 ;
      RECT  8262.5 53047.5 8327.5 53182.5 ;
      RECT  8097.5 53305.0 7962.5 53370.0 ;
      RECT  7907.5 53445.0 7772.5 53510.0 ;
      RECT  7717.5 53585.0 7582.5 53650.0 ;
      RECT  7712.5 53932.5 7777.5 54067.5 ;
      RECT  8092.5 53932.5 8157.5 54067.5 ;
      RECT  8092.5 53092.5 8157.5 53227.5 ;
      RECT  8092.5 53550.0 8157.5 53685.0 ;
      RECT  7582.5 53585.0 7717.5 53650.0 ;
      RECT  7772.5 53445.0 7907.5 53510.0 ;
      RECT  7962.5 53305.0 8097.5 53370.0 ;
      RECT  8092.5 53550.0 8157.5 53685.0 ;
      RECT  7455.0 54242.5 8465.0 54307.5 ;
      RECT  7455.0 52897.5 8465.0 52962.5 ;
      RECT  7522.5 55457.5 7587.5 55652.5 ;
      RECT  7522.5 54617.5 7587.5 54242.5 ;
      RECT  7902.5 54617.5 7967.5 54242.5 ;
      RECT  8262.5 54460.0 8327.5 54275.0 ;
      RECT  8262.5 55620.0 8327.5 55435.0 ;
      RECT  7522.5 54617.5 7587.5 54482.5 ;
      RECT  7712.5 54617.5 7777.5 54482.5 ;
      RECT  7712.5 54617.5 7777.5 54482.5 ;
      RECT  7522.5 54617.5 7587.5 54482.5 ;
      RECT  7712.5 54617.5 7777.5 54482.5 ;
      RECT  7902.5 54617.5 7967.5 54482.5 ;
      RECT  7902.5 54617.5 7967.5 54482.5 ;
      RECT  7712.5 54617.5 7777.5 54482.5 ;
      RECT  7902.5 54617.5 7967.5 54482.5 ;
      RECT  8092.5 54617.5 8157.5 54482.5 ;
      RECT  8092.5 54617.5 8157.5 54482.5 ;
      RECT  7902.5 54617.5 7967.5 54482.5 ;
      RECT  7522.5 55457.5 7587.5 55322.5 ;
      RECT  7712.5 55457.5 7777.5 55322.5 ;
      RECT  7712.5 55457.5 7777.5 55322.5 ;
      RECT  7522.5 55457.5 7587.5 55322.5 ;
      RECT  7712.5 55457.5 7777.5 55322.5 ;
      RECT  7902.5 55457.5 7967.5 55322.5 ;
      RECT  7902.5 55457.5 7967.5 55322.5 ;
      RECT  7712.5 55457.5 7777.5 55322.5 ;
      RECT  7902.5 55457.5 7967.5 55322.5 ;
      RECT  8092.5 55457.5 8157.5 55322.5 ;
      RECT  8092.5 55457.5 8157.5 55322.5 ;
      RECT  7902.5 55457.5 7967.5 55322.5 ;
      RECT  8262.5 54527.5 8327.5 54392.5 ;
      RECT  8262.5 55502.5 8327.5 55367.5 ;
      RECT  8097.5 55245.0 7962.5 55180.0 ;
      RECT  7907.5 55105.0 7772.5 55040.0 ;
      RECT  7717.5 54965.0 7582.5 54900.0 ;
      RECT  7712.5 54617.5 7777.5 54482.5 ;
      RECT  8092.5 54617.5 8157.5 54482.5 ;
      RECT  8092.5 55457.5 8157.5 55322.5 ;
      RECT  8092.5 55000.0 8157.5 54865.0 ;
      RECT  7582.5 54965.0 7717.5 54900.0 ;
      RECT  7772.5 55105.0 7907.5 55040.0 ;
      RECT  7962.5 55245.0 8097.5 55180.0 ;
      RECT  8092.5 55000.0 8157.5 54865.0 ;
      RECT  7455.0 54307.5 8465.0 54242.5 ;
      RECT  7455.0 55652.5 8465.0 55587.5 ;
      RECT  7522.5 55782.5 7587.5 55587.5 ;
      RECT  7522.5 56622.5 7587.5 56997.5 ;
      RECT  7902.5 56622.5 7967.5 56997.5 ;
      RECT  8262.5 56780.0 8327.5 56965.0 ;
      RECT  8262.5 55620.0 8327.5 55805.0 ;
      RECT  7522.5 56622.5 7587.5 56757.5 ;
      RECT  7712.5 56622.5 7777.5 56757.5 ;
      RECT  7712.5 56622.5 7777.5 56757.5 ;
      RECT  7522.5 56622.5 7587.5 56757.5 ;
      RECT  7712.5 56622.5 7777.5 56757.5 ;
      RECT  7902.5 56622.5 7967.5 56757.5 ;
      RECT  7902.5 56622.5 7967.5 56757.5 ;
      RECT  7712.5 56622.5 7777.5 56757.5 ;
      RECT  7902.5 56622.5 7967.5 56757.5 ;
      RECT  8092.5 56622.5 8157.5 56757.5 ;
      RECT  8092.5 56622.5 8157.5 56757.5 ;
      RECT  7902.5 56622.5 7967.5 56757.5 ;
      RECT  7522.5 55782.5 7587.5 55917.5 ;
      RECT  7712.5 55782.5 7777.5 55917.5 ;
      RECT  7712.5 55782.5 7777.5 55917.5 ;
      RECT  7522.5 55782.5 7587.5 55917.5 ;
      RECT  7712.5 55782.5 7777.5 55917.5 ;
      RECT  7902.5 55782.5 7967.5 55917.5 ;
      RECT  7902.5 55782.5 7967.5 55917.5 ;
      RECT  7712.5 55782.5 7777.5 55917.5 ;
      RECT  7902.5 55782.5 7967.5 55917.5 ;
      RECT  8092.5 55782.5 8157.5 55917.5 ;
      RECT  8092.5 55782.5 8157.5 55917.5 ;
      RECT  7902.5 55782.5 7967.5 55917.5 ;
      RECT  8262.5 56712.5 8327.5 56847.5 ;
      RECT  8262.5 55737.5 8327.5 55872.5 ;
      RECT  8097.5 55995.0 7962.5 56060.0 ;
      RECT  7907.5 56135.0 7772.5 56200.0 ;
      RECT  7717.5 56275.0 7582.5 56340.0 ;
      RECT  7712.5 56622.5 7777.5 56757.5 ;
      RECT  8092.5 56622.5 8157.5 56757.5 ;
      RECT  8092.5 55782.5 8157.5 55917.5 ;
      RECT  8092.5 56240.0 8157.5 56375.0 ;
      RECT  7582.5 56275.0 7717.5 56340.0 ;
      RECT  7772.5 56135.0 7907.5 56200.0 ;
      RECT  7962.5 55995.0 8097.5 56060.0 ;
      RECT  8092.5 56240.0 8157.5 56375.0 ;
      RECT  7455.0 56932.5 8465.0 56997.5 ;
      RECT  7455.0 55587.5 8465.0 55652.5 ;
      RECT  7522.5 58147.5 7587.5 58342.5 ;
      RECT  7522.5 57307.5 7587.5 56932.5 ;
      RECT  7902.5 57307.5 7967.5 56932.5 ;
      RECT  8262.5 57150.0 8327.5 56965.0 ;
      RECT  8262.5 58310.0 8327.5 58125.0 ;
      RECT  7522.5 57307.5 7587.5 57172.5 ;
      RECT  7712.5 57307.5 7777.5 57172.5 ;
      RECT  7712.5 57307.5 7777.5 57172.5 ;
      RECT  7522.5 57307.5 7587.5 57172.5 ;
      RECT  7712.5 57307.5 7777.5 57172.5 ;
      RECT  7902.5 57307.5 7967.5 57172.5 ;
      RECT  7902.5 57307.5 7967.5 57172.5 ;
      RECT  7712.5 57307.5 7777.5 57172.5 ;
      RECT  7902.5 57307.5 7967.5 57172.5 ;
      RECT  8092.5 57307.5 8157.5 57172.5 ;
      RECT  8092.5 57307.5 8157.5 57172.5 ;
      RECT  7902.5 57307.5 7967.5 57172.5 ;
      RECT  7522.5 58147.5 7587.5 58012.5 ;
      RECT  7712.5 58147.5 7777.5 58012.5 ;
      RECT  7712.5 58147.5 7777.5 58012.5 ;
      RECT  7522.5 58147.5 7587.5 58012.5 ;
      RECT  7712.5 58147.5 7777.5 58012.5 ;
      RECT  7902.5 58147.5 7967.5 58012.5 ;
      RECT  7902.5 58147.5 7967.5 58012.5 ;
      RECT  7712.5 58147.5 7777.5 58012.5 ;
      RECT  7902.5 58147.5 7967.5 58012.5 ;
      RECT  8092.5 58147.5 8157.5 58012.5 ;
      RECT  8092.5 58147.5 8157.5 58012.5 ;
      RECT  7902.5 58147.5 7967.5 58012.5 ;
      RECT  8262.5 57217.5 8327.5 57082.5 ;
      RECT  8262.5 58192.5 8327.5 58057.5 ;
      RECT  8097.5 57935.0 7962.5 57870.0 ;
      RECT  7907.5 57795.0 7772.5 57730.0 ;
      RECT  7717.5 57655.0 7582.5 57590.0 ;
      RECT  7712.5 57307.5 7777.5 57172.5 ;
      RECT  8092.5 57307.5 8157.5 57172.5 ;
      RECT  8092.5 58147.5 8157.5 58012.5 ;
      RECT  8092.5 57690.0 8157.5 57555.0 ;
      RECT  7582.5 57655.0 7717.5 57590.0 ;
      RECT  7772.5 57795.0 7907.5 57730.0 ;
      RECT  7962.5 57935.0 8097.5 57870.0 ;
      RECT  8092.5 57690.0 8157.5 57555.0 ;
      RECT  7455.0 56997.5 8465.0 56932.5 ;
      RECT  7455.0 58342.5 8465.0 58277.5 ;
      RECT  7522.5 58472.5 7587.5 58277.5 ;
      RECT  7522.5 59312.5 7587.5 59687.5 ;
      RECT  7902.5 59312.5 7967.5 59687.5 ;
      RECT  8262.5 59470.0 8327.5 59655.0 ;
      RECT  8262.5 58310.0 8327.5 58495.0 ;
      RECT  7522.5 59312.5 7587.5 59447.5 ;
      RECT  7712.5 59312.5 7777.5 59447.5 ;
      RECT  7712.5 59312.5 7777.5 59447.5 ;
      RECT  7522.5 59312.5 7587.5 59447.5 ;
      RECT  7712.5 59312.5 7777.5 59447.5 ;
      RECT  7902.5 59312.5 7967.5 59447.5 ;
      RECT  7902.5 59312.5 7967.5 59447.5 ;
      RECT  7712.5 59312.5 7777.5 59447.5 ;
      RECT  7902.5 59312.5 7967.5 59447.5 ;
      RECT  8092.5 59312.5 8157.5 59447.5 ;
      RECT  8092.5 59312.5 8157.5 59447.5 ;
      RECT  7902.5 59312.5 7967.5 59447.5 ;
      RECT  7522.5 58472.5 7587.5 58607.5 ;
      RECT  7712.5 58472.5 7777.5 58607.5 ;
      RECT  7712.5 58472.5 7777.5 58607.5 ;
      RECT  7522.5 58472.5 7587.5 58607.5 ;
      RECT  7712.5 58472.5 7777.5 58607.5 ;
      RECT  7902.5 58472.5 7967.5 58607.5 ;
      RECT  7902.5 58472.5 7967.5 58607.5 ;
      RECT  7712.5 58472.5 7777.5 58607.5 ;
      RECT  7902.5 58472.5 7967.5 58607.5 ;
      RECT  8092.5 58472.5 8157.5 58607.5 ;
      RECT  8092.5 58472.5 8157.5 58607.5 ;
      RECT  7902.5 58472.5 7967.5 58607.5 ;
      RECT  8262.5 59402.5 8327.5 59537.5 ;
      RECT  8262.5 58427.5 8327.5 58562.5 ;
      RECT  8097.5 58685.0 7962.5 58750.0 ;
      RECT  7907.5 58825.0 7772.5 58890.0 ;
      RECT  7717.5 58965.0 7582.5 59030.0 ;
      RECT  7712.5 59312.5 7777.5 59447.5 ;
      RECT  8092.5 59312.5 8157.5 59447.5 ;
      RECT  8092.5 58472.5 8157.5 58607.5 ;
      RECT  8092.5 58930.0 8157.5 59065.0 ;
      RECT  7582.5 58965.0 7717.5 59030.0 ;
      RECT  7772.5 58825.0 7907.5 58890.0 ;
      RECT  7962.5 58685.0 8097.5 58750.0 ;
      RECT  8092.5 58930.0 8157.5 59065.0 ;
      RECT  7455.0 59622.5 8465.0 59687.5 ;
      RECT  7455.0 58277.5 8465.0 58342.5 ;
      RECT  7522.5 60837.5 7587.5 61032.5 ;
      RECT  7522.5 59997.5 7587.5 59622.5 ;
      RECT  7902.5 59997.5 7967.5 59622.5 ;
      RECT  8262.5 59840.0 8327.5 59655.0 ;
      RECT  8262.5 61000.0 8327.5 60815.0 ;
      RECT  7522.5 59997.5 7587.5 59862.5 ;
      RECT  7712.5 59997.5 7777.5 59862.5 ;
      RECT  7712.5 59997.5 7777.5 59862.5 ;
      RECT  7522.5 59997.5 7587.5 59862.5 ;
      RECT  7712.5 59997.5 7777.5 59862.5 ;
      RECT  7902.5 59997.5 7967.5 59862.5 ;
      RECT  7902.5 59997.5 7967.5 59862.5 ;
      RECT  7712.5 59997.5 7777.5 59862.5 ;
      RECT  7902.5 59997.5 7967.5 59862.5 ;
      RECT  8092.5 59997.5 8157.5 59862.5 ;
      RECT  8092.5 59997.5 8157.5 59862.5 ;
      RECT  7902.5 59997.5 7967.5 59862.5 ;
      RECT  7522.5 60837.5 7587.5 60702.5 ;
      RECT  7712.5 60837.5 7777.5 60702.5 ;
      RECT  7712.5 60837.5 7777.5 60702.5 ;
      RECT  7522.5 60837.5 7587.5 60702.5 ;
      RECT  7712.5 60837.5 7777.5 60702.5 ;
      RECT  7902.5 60837.5 7967.5 60702.5 ;
      RECT  7902.5 60837.5 7967.5 60702.5 ;
      RECT  7712.5 60837.5 7777.5 60702.5 ;
      RECT  7902.5 60837.5 7967.5 60702.5 ;
      RECT  8092.5 60837.5 8157.5 60702.5 ;
      RECT  8092.5 60837.5 8157.5 60702.5 ;
      RECT  7902.5 60837.5 7967.5 60702.5 ;
      RECT  8262.5 59907.5 8327.5 59772.5 ;
      RECT  8262.5 60882.5 8327.5 60747.5 ;
      RECT  8097.5 60625.0 7962.5 60560.0 ;
      RECT  7907.5 60485.0 7772.5 60420.0 ;
      RECT  7717.5 60345.0 7582.5 60280.0 ;
      RECT  7712.5 59997.5 7777.5 59862.5 ;
      RECT  8092.5 59997.5 8157.5 59862.5 ;
      RECT  8092.5 60837.5 8157.5 60702.5 ;
      RECT  8092.5 60380.0 8157.5 60245.0 ;
      RECT  7582.5 60345.0 7717.5 60280.0 ;
      RECT  7772.5 60485.0 7907.5 60420.0 ;
      RECT  7962.5 60625.0 8097.5 60560.0 ;
      RECT  8092.5 60380.0 8157.5 60245.0 ;
      RECT  7455.0 59687.5 8465.0 59622.5 ;
      RECT  7455.0 61032.5 8465.0 60967.5 ;
      RECT  7522.5 61162.5 7587.5 60967.5 ;
      RECT  7522.5 62002.5 7587.5 62377.5 ;
      RECT  7902.5 62002.5 7967.5 62377.5 ;
      RECT  8262.5 62160.0 8327.5 62345.0 ;
      RECT  8262.5 61000.0 8327.5 61185.0 ;
      RECT  7522.5 62002.5 7587.5 62137.5 ;
      RECT  7712.5 62002.5 7777.5 62137.5 ;
      RECT  7712.5 62002.5 7777.5 62137.5 ;
      RECT  7522.5 62002.5 7587.5 62137.5 ;
      RECT  7712.5 62002.5 7777.5 62137.5 ;
      RECT  7902.5 62002.5 7967.5 62137.5 ;
      RECT  7902.5 62002.5 7967.5 62137.5 ;
      RECT  7712.5 62002.5 7777.5 62137.5 ;
      RECT  7902.5 62002.5 7967.5 62137.5 ;
      RECT  8092.5 62002.5 8157.5 62137.5 ;
      RECT  8092.5 62002.5 8157.5 62137.5 ;
      RECT  7902.5 62002.5 7967.5 62137.5 ;
      RECT  7522.5 61162.5 7587.5 61297.5 ;
      RECT  7712.5 61162.5 7777.5 61297.5 ;
      RECT  7712.5 61162.5 7777.5 61297.5 ;
      RECT  7522.5 61162.5 7587.5 61297.5 ;
      RECT  7712.5 61162.5 7777.5 61297.5 ;
      RECT  7902.5 61162.5 7967.5 61297.5 ;
      RECT  7902.5 61162.5 7967.5 61297.5 ;
      RECT  7712.5 61162.5 7777.5 61297.5 ;
      RECT  7902.5 61162.5 7967.5 61297.5 ;
      RECT  8092.5 61162.5 8157.5 61297.5 ;
      RECT  8092.5 61162.5 8157.5 61297.5 ;
      RECT  7902.5 61162.5 7967.5 61297.5 ;
      RECT  8262.5 62092.5 8327.5 62227.5 ;
      RECT  8262.5 61117.5 8327.5 61252.5 ;
      RECT  8097.5 61375.0 7962.5 61440.0 ;
      RECT  7907.5 61515.0 7772.5 61580.0 ;
      RECT  7717.5 61655.0 7582.5 61720.0 ;
      RECT  7712.5 62002.5 7777.5 62137.5 ;
      RECT  8092.5 62002.5 8157.5 62137.5 ;
      RECT  8092.5 61162.5 8157.5 61297.5 ;
      RECT  8092.5 61620.0 8157.5 61755.0 ;
      RECT  7582.5 61655.0 7717.5 61720.0 ;
      RECT  7772.5 61515.0 7907.5 61580.0 ;
      RECT  7962.5 61375.0 8097.5 61440.0 ;
      RECT  8092.5 61620.0 8157.5 61755.0 ;
      RECT  7455.0 62312.5 8465.0 62377.5 ;
      RECT  7455.0 60967.5 8465.0 61032.5 ;
      RECT  7522.5 63527.5 7587.5 63722.5 ;
      RECT  7522.5 62687.5 7587.5 62312.5 ;
      RECT  7902.5 62687.5 7967.5 62312.5 ;
      RECT  8262.5 62530.0 8327.5 62345.0 ;
      RECT  8262.5 63690.0 8327.5 63505.0 ;
      RECT  7522.5 62687.5 7587.5 62552.5 ;
      RECT  7712.5 62687.5 7777.5 62552.5 ;
      RECT  7712.5 62687.5 7777.5 62552.5 ;
      RECT  7522.5 62687.5 7587.5 62552.5 ;
      RECT  7712.5 62687.5 7777.5 62552.5 ;
      RECT  7902.5 62687.5 7967.5 62552.5 ;
      RECT  7902.5 62687.5 7967.5 62552.5 ;
      RECT  7712.5 62687.5 7777.5 62552.5 ;
      RECT  7902.5 62687.5 7967.5 62552.5 ;
      RECT  8092.5 62687.5 8157.5 62552.5 ;
      RECT  8092.5 62687.5 8157.5 62552.5 ;
      RECT  7902.5 62687.5 7967.5 62552.5 ;
      RECT  7522.5 63527.5 7587.5 63392.5 ;
      RECT  7712.5 63527.5 7777.5 63392.5 ;
      RECT  7712.5 63527.5 7777.5 63392.5 ;
      RECT  7522.5 63527.5 7587.5 63392.5 ;
      RECT  7712.5 63527.5 7777.5 63392.5 ;
      RECT  7902.5 63527.5 7967.5 63392.5 ;
      RECT  7902.5 63527.5 7967.5 63392.5 ;
      RECT  7712.5 63527.5 7777.5 63392.5 ;
      RECT  7902.5 63527.5 7967.5 63392.5 ;
      RECT  8092.5 63527.5 8157.5 63392.5 ;
      RECT  8092.5 63527.5 8157.5 63392.5 ;
      RECT  7902.5 63527.5 7967.5 63392.5 ;
      RECT  8262.5 62597.5 8327.5 62462.5 ;
      RECT  8262.5 63572.5 8327.5 63437.5 ;
      RECT  8097.5 63315.0 7962.5 63250.0 ;
      RECT  7907.5 63175.0 7772.5 63110.0 ;
      RECT  7717.5 63035.0 7582.5 62970.0 ;
      RECT  7712.5 62687.5 7777.5 62552.5 ;
      RECT  8092.5 62687.5 8157.5 62552.5 ;
      RECT  8092.5 63527.5 8157.5 63392.5 ;
      RECT  8092.5 63070.0 8157.5 62935.0 ;
      RECT  7582.5 63035.0 7717.5 62970.0 ;
      RECT  7772.5 63175.0 7907.5 63110.0 ;
      RECT  7962.5 63315.0 8097.5 63250.0 ;
      RECT  8092.5 63070.0 8157.5 62935.0 ;
      RECT  7455.0 62377.5 8465.0 62312.5 ;
      RECT  7455.0 63722.5 8465.0 63657.5 ;
      RECT  7522.5 63852.5 7587.5 63657.5 ;
      RECT  7522.5 64692.5 7587.5 65067.5 ;
      RECT  7902.5 64692.5 7967.5 65067.5 ;
      RECT  8262.5 64850.0 8327.5 65035.0 ;
      RECT  8262.5 63690.0 8327.5 63875.0 ;
      RECT  7522.5 64692.5 7587.5 64827.5 ;
      RECT  7712.5 64692.5 7777.5 64827.5 ;
      RECT  7712.5 64692.5 7777.5 64827.5 ;
      RECT  7522.5 64692.5 7587.5 64827.5 ;
      RECT  7712.5 64692.5 7777.5 64827.5 ;
      RECT  7902.5 64692.5 7967.5 64827.5 ;
      RECT  7902.5 64692.5 7967.5 64827.5 ;
      RECT  7712.5 64692.5 7777.5 64827.5 ;
      RECT  7902.5 64692.5 7967.5 64827.5 ;
      RECT  8092.5 64692.5 8157.5 64827.5 ;
      RECT  8092.5 64692.5 8157.5 64827.5 ;
      RECT  7902.5 64692.5 7967.5 64827.5 ;
      RECT  7522.5 63852.5 7587.5 63987.5 ;
      RECT  7712.5 63852.5 7777.5 63987.5 ;
      RECT  7712.5 63852.5 7777.5 63987.5 ;
      RECT  7522.5 63852.5 7587.5 63987.5 ;
      RECT  7712.5 63852.5 7777.5 63987.5 ;
      RECT  7902.5 63852.5 7967.5 63987.5 ;
      RECT  7902.5 63852.5 7967.5 63987.5 ;
      RECT  7712.5 63852.5 7777.5 63987.5 ;
      RECT  7902.5 63852.5 7967.5 63987.5 ;
      RECT  8092.5 63852.5 8157.5 63987.5 ;
      RECT  8092.5 63852.5 8157.5 63987.5 ;
      RECT  7902.5 63852.5 7967.5 63987.5 ;
      RECT  8262.5 64782.5 8327.5 64917.5 ;
      RECT  8262.5 63807.5 8327.5 63942.5 ;
      RECT  8097.5 64065.0 7962.5 64130.0 ;
      RECT  7907.5 64205.0 7772.5 64270.0 ;
      RECT  7717.5 64345.0 7582.5 64410.0 ;
      RECT  7712.5 64692.5 7777.5 64827.5 ;
      RECT  8092.5 64692.5 8157.5 64827.5 ;
      RECT  8092.5 63852.5 8157.5 63987.5 ;
      RECT  8092.5 64310.0 8157.5 64445.0 ;
      RECT  7582.5 64345.0 7717.5 64410.0 ;
      RECT  7772.5 64205.0 7907.5 64270.0 ;
      RECT  7962.5 64065.0 8097.5 64130.0 ;
      RECT  8092.5 64310.0 8157.5 64445.0 ;
      RECT  7455.0 65002.5 8465.0 65067.5 ;
      RECT  7455.0 63657.5 8465.0 63722.5 ;
      RECT  7522.5 66217.5 7587.5 66412.5 ;
      RECT  7522.5 65377.5 7587.5 65002.5 ;
      RECT  7902.5 65377.5 7967.5 65002.5 ;
      RECT  8262.5 65220.0 8327.5 65035.0 ;
      RECT  8262.5 66380.0 8327.5 66195.0 ;
      RECT  7522.5 65377.5 7587.5 65242.5 ;
      RECT  7712.5 65377.5 7777.5 65242.5 ;
      RECT  7712.5 65377.5 7777.5 65242.5 ;
      RECT  7522.5 65377.5 7587.5 65242.5 ;
      RECT  7712.5 65377.5 7777.5 65242.5 ;
      RECT  7902.5 65377.5 7967.5 65242.5 ;
      RECT  7902.5 65377.5 7967.5 65242.5 ;
      RECT  7712.5 65377.5 7777.5 65242.5 ;
      RECT  7902.5 65377.5 7967.5 65242.5 ;
      RECT  8092.5 65377.5 8157.5 65242.5 ;
      RECT  8092.5 65377.5 8157.5 65242.5 ;
      RECT  7902.5 65377.5 7967.5 65242.5 ;
      RECT  7522.5 66217.5 7587.5 66082.5 ;
      RECT  7712.5 66217.5 7777.5 66082.5 ;
      RECT  7712.5 66217.5 7777.5 66082.5 ;
      RECT  7522.5 66217.5 7587.5 66082.5 ;
      RECT  7712.5 66217.5 7777.5 66082.5 ;
      RECT  7902.5 66217.5 7967.5 66082.5 ;
      RECT  7902.5 66217.5 7967.5 66082.5 ;
      RECT  7712.5 66217.5 7777.5 66082.5 ;
      RECT  7902.5 66217.5 7967.5 66082.5 ;
      RECT  8092.5 66217.5 8157.5 66082.5 ;
      RECT  8092.5 66217.5 8157.5 66082.5 ;
      RECT  7902.5 66217.5 7967.5 66082.5 ;
      RECT  8262.5 65287.5 8327.5 65152.5 ;
      RECT  8262.5 66262.5 8327.5 66127.5 ;
      RECT  8097.5 66005.0 7962.5 65940.0 ;
      RECT  7907.5 65865.0 7772.5 65800.0 ;
      RECT  7717.5 65725.0 7582.5 65660.0 ;
      RECT  7712.5 65377.5 7777.5 65242.5 ;
      RECT  8092.5 65377.5 8157.5 65242.5 ;
      RECT  8092.5 66217.5 8157.5 66082.5 ;
      RECT  8092.5 65760.0 8157.5 65625.0 ;
      RECT  7582.5 65725.0 7717.5 65660.0 ;
      RECT  7772.5 65865.0 7907.5 65800.0 ;
      RECT  7962.5 66005.0 8097.5 65940.0 ;
      RECT  8092.5 65760.0 8157.5 65625.0 ;
      RECT  7455.0 65067.5 8465.0 65002.5 ;
      RECT  7455.0 66412.5 8465.0 66347.5 ;
      RECT  7522.5 66542.5 7587.5 66347.5 ;
      RECT  7522.5 67382.5 7587.5 67757.5 ;
      RECT  7902.5 67382.5 7967.5 67757.5 ;
      RECT  8262.5 67540.0 8327.5 67725.0 ;
      RECT  8262.5 66380.0 8327.5 66565.0 ;
      RECT  7522.5 67382.5 7587.5 67517.5 ;
      RECT  7712.5 67382.5 7777.5 67517.5 ;
      RECT  7712.5 67382.5 7777.5 67517.5 ;
      RECT  7522.5 67382.5 7587.5 67517.5 ;
      RECT  7712.5 67382.5 7777.5 67517.5 ;
      RECT  7902.5 67382.5 7967.5 67517.5 ;
      RECT  7902.5 67382.5 7967.5 67517.5 ;
      RECT  7712.5 67382.5 7777.5 67517.5 ;
      RECT  7902.5 67382.5 7967.5 67517.5 ;
      RECT  8092.5 67382.5 8157.5 67517.5 ;
      RECT  8092.5 67382.5 8157.5 67517.5 ;
      RECT  7902.5 67382.5 7967.5 67517.5 ;
      RECT  7522.5 66542.5 7587.5 66677.5 ;
      RECT  7712.5 66542.5 7777.5 66677.5 ;
      RECT  7712.5 66542.5 7777.5 66677.5 ;
      RECT  7522.5 66542.5 7587.5 66677.5 ;
      RECT  7712.5 66542.5 7777.5 66677.5 ;
      RECT  7902.5 66542.5 7967.5 66677.5 ;
      RECT  7902.5 66542.5 7967.5 66677.5 ;
      RECT  7712.5 66542.5 7777.5 66677.5 ;
      RECT  7902.5 66542.5 7967.5 66677.5 ;
      RECT  8092.5 66542.5 8157.5 66677.5 ;
      RECT  8092.5 66542.5 8157.5 66677.5 ;
      RECT  7902.5 66542.5 7967.5 66677.5 ;
      RECT  8262.5 67472.5 8327.5 67607.5 ;
      RECT  8262.5 66497.5 8327.5 66632.5 ;
      RECT  8097.5 66755.0 7962.5 66820.0 ;
      RECT  7907.5 66895.0 7772.5 66960.0 ;
      RECT  7717.5 67035.0 7582.5 67100.0 ;
      RECT  7712.5 67382.5 7777.5 67517.5 ;
      RECT  8092.5 67382.5 8157.5 67517.5 ;
      RECT  8092.5 66542.5 8157.5 66677.5 ;
      RECT  8092.5 67000.0 8157.5 67135.0 ;
      RECT  7582.5 67035.0 7717.5 67100.0 ;
      RECT  7772.5 66895.0 7907.5 66960.0 ;
      RECT  7962.5 66755.0 8097.5 66820.0 ;
      RECT  8092.5 67000.0 8157.5 67135.0 ;
      RECT  7455.0 67692.5 8465.0 67757.5 ;
      RECT  7455.0 66347.5 8465.0 66412.5 ;
      RECT  7522.5 68907.5 7587.5 69102.5 ;
      RECT  7522.5 68067.5 7587.5 67692.5 ;
      RECT  7902.5 68067.5 7967.5 67692.5 ;
      RECT  8262.5 67910.0 8327.5 67725.0 ;
      RECT  8262.5 69070.0 8327.5 68885.0 ;
      RECT  7522.5 68067.5 7587.5 67932.5 ;
      RECT  7712.5 68067.5 7777.5 67932.5 ;
      RECT  7712.5 68067.5 7777.5 67932.5 ;
      RECT  7522.5 68067.5 7587.5 67932.5 ;
      RECT  7712.5 68067.5 7777.5 67932.5 ;
      RECT  7902.5 68067.5 7967.5 67932.5 ;
      RECT  7902.5 68067.5 7967.5 67932.5 ;
      RECT  7712.5 68067.5 7777.5 67932.5 ;
      RECT  7902.5 68067.5 7967.5 67932.5 ;
      RECT  8092.5 68067.5 8157.5 67932.5 ;
      RECT  8092.5 68067.5 8157.5 67932.5 ;
      RECT  7902.5 68067.5 7967.5 67932.5 ;
      RECT  7522.5 68907.5 7587.5 68772.5 ;
      RECT  7712.5 68907.5 7777.5 68772.5 ;
      RECT  7712.5 68907.5 7777.5 68772.5 ;
      RECT  7522.5 68907.5 7587.5 68772.5 ;
      RECT  7712.5 68907.5 7777.5 68772.5 ;
      RECT  7902.5 68907.5 7967.5 68772.5 ;
      RECT  7902.5 68907.5 7967.5 68772.5 ;
      RECT  7712.5 68907.5 7777.5 68772.5 ;
      RECT  7902.5 68907.5 7967.5 68772.5 ;
      RECT  8092.5 68907.5 8157.5 68772.5 ;
      RECT  8092.5 68907.5 8157.5 68772.5 ;
      RECT  7902.5 68907.5 7967.5 68772.5 ;
      RECT  8262.5 67977.5 8327.5 67842.5 ;
      RECT  8262.5 68952.5 8327.5 68817.5 ;
      RECT  8097.5 68695.0 7962.5 68630.0 ;
      RECT  7907.5 68555.0 7772.5 68490.0 ;
      RECT  7717.5 68415.0 7582.5 68350.0 ;
      RECT  7712.5 68067.5 7777.5 67932.5 ;
      RECT  8092.5 68067.5 8157.5 67932.5 ;
      RECT  8092.5 68907.5 8157.5 68772.5 ;
      RECT  8092.5 68450.0 8157.5 68315.0 ;
      RECT  7582.5 68415.0 7717.5 68350.0 ;
      RECT  7772.5 68555.0 7907.5 68490.0 ;
      RECT  7962.5 68695.0 8097.5 68630.0 ;
      RECT  8092.5 68450.0 8157.5 68315.0 ;
      RECT  7455.0 67757.5 8465.0 67692.5 ;
      RECT  7455.0 69102.5 8465.0 69037.5 ;
      RECT  7522.5 69232.5 7587.5 69037.5 ;
      RECT  7522.5 70072.5 7587.5 70447.5 ;
      RECT  7902.5 70072.5 7967.5 70447.5 ;
      RECT  8262.5 70230.0 8327.5 70415.0 ;
      RECT  8262.5 69070.0 8327.5 69255.0 ;
      RECT  7522.5 70072.5 7587.5 70207.5 ;
      RECT  7712.5 70072.5 7777.5 70207.5 ;
      RECT  7712.5 70072.5 7777.5 70207.5 ;
      RECT  7522.5 70072.5 7587.5 70207.5 ;
      RECT  7712.5 70072.5 7777.5 70207.5 ;
      RECT  7902.5 70072.5 7967.5 70207.5 ;
      RECT  7902.5 70072.5 7967.5 70207.5 ;
      RECT  7712.5 70072.5 7777.5 70207.5 ;
      RECT  7902.5 70072.5 7967.5 70207.5 ;
      RECT  8092.5 70072.5 8157.5 70207.5 ;
      RECT  8092.5 70072.5 8157.5 70207.5 ;
      RECT  7902.5 70072.5 7967.5 70207.5 ;
      RECT  7522.5 69232.5 7587.5 69367.5 ;
      RECT  7712.5 69232.5 7777.5 69367.5 ;
      RECT  7712.5 69232.5 7777.5 69367.5 ;
      RECT  7522.5 69232.5 7587.5 69367.5 ;
      RECT  7712.5 69232.5 7777.5 69367.5 ;
      RECT  7902.5 69232.5 7967.5 69367.5 ;
      RECT  7902.5 69232.5 7967.5 69367.5 ;
      RECT  7712.5 69232.5 7777.5 69367.5 ;
      RECT  7902.5 69232.5 7967.5 69367.5 ;
      RECT  8092.5 69232.5 8157.5 69367.5 ;
      RECT  8092.5 69232.5 8157.5 69367.5 ;
      RECT  7902.5 69232.5 7967.5 69367.5 ;
      RECT  8262.5 70162.5 8327.5 70297.5 ;
      RECT  8262.5 69187.5 8327.5 69322.5 ;
      RECT  8097.5 69445.0 7962.5 69510.0 ;
      RECT  7907.5 69585.0 7772.5 69650.0 ;
      RECT  7717.5 69725.0 7582.5 69790.0 ;
      RECT  7712.5 70072.5 7777.5 70207.5 ;
      RECT  8092.5 70072.5 8157.5 70207.5 ;
      RECT  8092.5 69232.5 8157.5 69367.5 ;
      RECT  8092.5 69690.0 8157.5 69825.0 ;
      RECT  7582.5 69725.0 7717.5 69790.0 ;
      RECT  7772.5 69585.0 7907.5 69650.0 ;
      RECT  7962.5 69445.0 8097.5 69510.0 ;
      RECT  8092.5 69690.0 8157.5 69825.0 ;
      RECT  7455.0 70382.5 8465.0 70447.5 ;
      RECT  7455.0 69037.5 8465.0 69102.5 ;
      RECT  7522.5 71597.5 7587.5 71792.5 ;
      RECT  7522.5 70757.5 7587.5 70382.5 ;
      RECT  7902.5 70757.5 7967.5 70382.5 ;
      RECT  8262.5 70600.0 8327.5 70415.0 ;
      RECT  8262.5 71760.0 8327.5 71575.0 ;
      RECT  7522.5 70757.5 7587.5 70622.5 ;
      RECT  7712.5 70757.5 7777.5 70622.5 ;
      RECT  7712.5 70757.5 7777.5 70622.5 ;
      RECT  7522.5 70757.5 7587.5 70622.5 ;
      RECT  7712.5 70757.5 7777.5 70622.5 ;
      RECT  7902.5 70757.5 7967.5 70622.5 ;
      RECT  7902.5 70757.5 7967.5 70622.5 ;
      RECT  7712.5 70757.5 7777.5 70622.5 ;
      RECT  7902.5 70757.5 7967.5 70622.5 ;
      RECT  8092.5 70757.5 8157.5 70622.5 ;
      RECT  8092.5 70757.5 8157.5 70622.5 ;
      RECT  7902.5 70757.5 7967.5 70622.5 ;
      RECT  7522.5 71597.5 7587.5 71462.5 ;
      RECT  7712.5 71597.5 7777.5 71462.5 ;
      RECT  7712.5 71597.5 7777.5 71462.5 ;
      RECT  7522.5 71597.5 7587.5 71462.5 ;
      RECT  7712.5 71597.5 7777.5 71462.5 ;
      RECT  7902.5 71597.5 7967.5 71462.5 ;
      RECT  7902.5 71597.5 7967.5 71462.5 ;
      RECT  7712.5 71597.5 7777.5 71462.5 ;
      RECT  7902.5 71597.5 7967.5 71462.5 ;
      RECT  8092.5 71597.5 8157.5 71462.5 ;
      RECT  8092.5 71597.5 8157.5 71462.5 ;
      RECT  7902.5 71597.5 7967.5 71462.5 ;
      RECT  8262.5 70667.5 8327.5 70532.5 ;
      RECT  8262.5 71642.5 8327.5 71507.5 ;
      RECT  8097.5 71385.0 7962.5 71320.0 ;
      RECT  7907.5 71245.0 7772.5 71180.0 ;
      RECT  7717.5 71105.0 7582.5 71040.0 ;
      RECT  7712.5 70757.5 7777.5 70622.5 ;
      RECT  8092.5 70757.5 8157.5 70622.5 ;
      RECT  8092.5 71597.5 8157.5 71462.5 ;
      RECT  8092.5 71140.0 8157.5 71005.0 ;
      RECT  7582.5 71105.0 7717.5 71040.0 ;
      RECT  7772.5 71245.0 7907.5 71180.0 ;
      RECT  7962.5 71385.0 8097.5 71320.0 ;
      RECT  8092.5 71140.0 8157.5 71005.0 ;
      RECT  7455.0 70447.5 8465.0 70382.5 ;
      RECT  7455.0 71792.5 8465.0 71727.5 ;
      RECT  7522.5 71922.5 7587.5 71727.5 ;
      RECT  7522.5 72762.5 7587.5 73137.5 ;
      RECT  7902.5 72762.5 7967.5 73137.5 ;
      RECT  8262.5 72920.0 8327.5 73105.0 ;
      RECT  8262.5 71760.0 8327.5 71945.0 ;
      RECT  7522.5 72762.5 7587.5 72897.5 ;
      RECT  7712.5 72762.5 7777.5 72897.5 ;
      RECT  7712.5 72762.5 7777.5 72897.5 ;
      RECT  7522.5 72762.5 7587.5 72897.5 ;
      RECT  7712.5 72762.5 7777.5 72897.5 ;
      RECT  7902.5 72762.5 7967.5 72897.5 ;
      RECT  7902.5 72762.5 7967.5 72897.5 ;
      RECT  7712.5 72762.5 7777.5 72897.5 ;
      RECT  7902.5 72762.5 7967.5 72897.5 ;
      RECT  8092.5 72762.5 8157.5 72897.5 ;
      RECT  8092.5 72762.5 8157.5 72897.5 ;
      RECT  7902.5 72762.5 7967.5 72897.5 ;
      RECT  7522.5 71922.5 7587.5 72057.5 ;
      RECT  7712.5 71922.5 7777.5 72057.5 ;
      RECT  7712.5 71922.5 7777.5 72057.5 ;
      RECT  7522.5 71922.5 7587.5 72057.5 ;
      RECT  7712.5 71922.5 7777.5 72057.5 ;
      RECT  7902.5 71922.5 7967.5 72057.5 ;
      RECT  7902.5 71922.5 7967.5 72057.5 ;
      RECT  7712.5 71922.5 7777.5 72057.5 ;
      RECT  7902.5 71922.5 7967.5 72057.5 ;
      RECT  8092.5 71922.5 8157.5 72057.5 ;
      RECT  8092.5 71922.5 8157.5 72057.5 ;
      RECT  7902.5 71922.5 7967.5 72057.5 ;
      RECT  8262.5 72852.5 8327.5 72987.5 ;
      RECT  8262.5 71877.5 8327.5 72012.5 ;
      RECT  8097.5 72135.0 7962.5 72200.0 ;
      RECT  7907.5 72275.0 7772.5 72340.0 ;
      RECT  7717.5 72415.0 7582.5 72480.0 ;
      RECT  7712.5 72762.5 7777.5 72897.5 ;
      RECT  8092.5 72762.5 8157.5 72897.5 ;
      RECT  8092.5 71922.5 8157.5 72057.5 ;
      RECT  8092.5 72380.0 8157.5 72515.0 ;
      RECT  7582.5 72415.0 7717.5 72480.0 ;
      RECT  7772.5 72275.0 7907.5 72340.0 ;
      RECT  7962.5 72135.0 8097.5 72200.0 ;
      RECT  8092.5 72380.0 8157.5 72515.0 ;
      RECT  7455.0 73072.5 8465.0 73137.5 ;
      RECT  7455.0 71727.5 8465.0 71792.5 ;
      RECT  7522.5 74287.5 7587.5 74482.5 ;
      RECT  7522.5 73447.5 7587.5 73072.5 ;
      RECT  7902.5 73447.5 7967.5 73072.5 ;
      RECT  8262.5 73290.0 8327.5 73105.0 ;
      RECT  8262.5 74450.0 8327.5 74265.0 ;
      RECT  7522.5 73447.5 7587.5 73312.5 ;
      RECT  7712.5 73447.5 7777.5 73312.5 ;
      RECT  7712.5 73447.5 7777.5 73312.5 ;
      RECT  7522.5 73447.5 7587.5 73312.5 ;
      RECT  7712.5 73447.5 7777.5 73312.5 ;
      RECT  7902.5 73447.5 7967.5 73312.5 ;
      RECT  7902.5 73447.5 7967.5 73312.5 ;
      RECT  7712.5 73447.5 7777.5 73312.5 ;
      RECT  7902.5 73447.5 7967.5 73312.5 ;
      RECT  8092.5 73447.5 8157.5 73312.5 ;
      RECT  8092.5 73447.5 8157.5 73312.5 ;
      RECT  7902.5 73447.5 7967.5 73312.5 ;
      RECT  7522.5 74287.5 7587.5 74152.5 ;
      RECT  7712.5 74287.5 7777.5 74152.5 ;
      RECT  7712.5 74287.5 7777.5 74152.5 ;
      RECT  7522.5 74287.5 7587.5 74152.5 ;
      RECT  7712.5 74287.5 7777.5 74152.5 ;
      RECT  7902.5 74287.5 7967.5 74152.5 ;
      RECT  7902.5 74287.5 7967.5 74152.5 ;
      RECT  7712.5 74287.5 7777.5 74152.5 ;
      RECT  7902.5 74287.5 7967.5 74152.5 ;
      RECT  8092.5 74287.5 8157.5 74152.5 ;
      RECT  8092.5 74287.5 8157.5 74152.5 ;
      RECT  7902.5 74287.5 7967.5 74152.5 ;
      RECT  8262.5 73357.5 8327.5 73222.5 ;
      RECT  8262.5 74332.5 8327.5 74197.5 ;
      RECT  8097.5 74075.0 7962.5 74010.0 ;
      RECT  7907.5 73935.0 7772.5 73870.0 ;
      RECT  7717.5 73795.0 7582.5 73730.0 ;
      RECT  7712.5 73447.5 7777.5 73312.5 ;
      RECT  8092.5 73447.5 8157.5 73312.5 ;
      RECT  8092.5 74287.5 8157.5 74152.5 ;
      RECT  8092.5 73830.0 8157.5 73695.0 ;
      RECT  7582.5 73795.0 7717.5 73730.0 ;
      RECT  7772.5 73935.0 7907.5 73870.0 ;
      RECT  7962.5 74075.0 8097.5 74010.0 ;
      RECT  8092.5 73830.0 8157.5 73695.0 ;
      RECT  7455.0 73137.5 8465.0 73072.5 ;
      RECT  7455.0 74482.5 8465.0 74417.5 ;
      RECT  7522.5 74612.5 7587.5 74417.5 ;
      RECT  7522.5 75452.5 7587.5 75827.5 ;
      RECT  7902.5 75452.5 7967.5 75827.5 ;
      RECT  8262.5 75610.0 8327.5 75795.0 ;
      RECT  8262.5 74450.0 8327.5 74635.0 ;
      RECT  7522.5 75452.5 7587.5 75587.5 ;
      RECT  7712.5 75452.5 7777.5 75587.5 ;
      RECT  7712.5 75452.5 7777.5 75587.5 ;
      RECT  7522.5 75452.5 7587.5 75587.5 ;
      RECT  7712.5 75452.5 7777.5 75587.5 ;
      RECT  7902.5 75452.5 7967.5 75587.5 ;
      RECT  7902.5 75452.5 7967.5 75587.5 ;
      RECT  7712.5 75452.5 7777.5 75587.5 ;
      RECT  7902.5 75452.5 7967.5 75587.5 ;
      RECT  8092.5 75452.5 8157.5 75587.5 ;
      RECT  8092.5 75452.5 8157.5 75587.5 ;
      RECT  7902.5 75452.5 7967.5 75587.5 ;
      RECT  7522.5 74612.5 7587.5 74747.5 ;
      RECT  7712.5 74612.5 7777.5 74747.5 ;
      RECT  7712.5 74612.5 7777.5 74747.5 ;
      RECT  7522.5 74612.5 7587.5 74747.5 ;
      RECT  7712.5 74612.5 7777.5 74747.5 ;
      RECT  7902.5 74612.5 7967.5 74747.5 ;
      RECT  7902.5 74612.5 7967.5 74747.5 ;
      RECT  7712.5 74612.5 7777.5 74747.5 ;
      RECT  7902.5 74612.5 7967.5 74747.5 ;
      RECT  8092.5 74612.5 8157.5 74747.5 ;
      RECT  8092.5 74612.5 8157.5 74747.5 ;
      RECT  7902.5 74612.5 7967.5 74747.5 ;
      RECT  8262.5 75542.5 8327.5 75677.5 ;
      RECT  8262.5 74567.5 8327.5 74702.5 ;
      RECT  8097.5 74825.0 7962.5 74890.0 ;
      RECT  7907.5 74965.0 7772.5 75030.0 ;
      RECT  7717.5 75105.0 7582.5 75170.0 ;
      RECT  7712.5 75452.5 7777.5 75587.5 ;
      RECT  8092.5 75452.5 8157.5 75587.5 ;
      RECT  8092.5 74612.5 8157.5 74747.5 ;
      RECT  8092.5 75070.0 8157.5 75205.0 ;
      RECT  7582.5 75105.0 7717.5 75170.0 ;
      RECT  7772.5 74965.0 7907.5 75030.0 ;
      RECT  7962.5 74825.0 8097.5 74890.0 ;
      RECT  8092.5 75070.0 8157.5 75205.0 ;
      RECT  7455.0 75762.5 8465.0 75827.5 ;
      RECT  7455.0 74417.5 8465.0 74482.5 ;
      RECT  7522.5 76977.5 7587.5 77172.5 ;
      RECT  7522.5 76137.5 7587.5 75762.5 ;
      RECT  7902.5 76137.5 7967.5 75762.5 ;
      RECT  8262.5 75980.0 8327.5 75795.0 ;
      RECT  8262.5 77140.0 8327.5 76955.0 ;
      RECT  7522.5 76137.5 7587.5 76002.5 ;
      RECT  7712.5 76137.5 7777.5 76002.5 ;
      RECT  7712.5 76137.5 7777.5 76002.5 ;
      RECT  7522.5 76137.5 7587.5 76002.5 ;
      RECT  7712.5 76137.5 7777.5 76002.5 ;
      RECT  7902.5 76137.5 7967.5 76002.5 ;
      RECT  7902.5 76137.5 7967.5 76002.5 ;
      RECT  7712.5 76137.5 7777.5 76002.5 ;
      RECT  7902.5 76137.5 7967.5 76002.5 ;
      RECT  8092.5 76137.5 8157.5 76002.5 ;
      RECT  8092.5 76137.5 8157.5 76002.5 ;
      RECT  7902.5 76137.5 7967.5 76002.5 ;
      RECT  7522.5 76977.5 7587.5 76842.5 ;
      RECT  7712.5 76977.5 7777.5 76842.5 ;
      RECT  7712.5 76977.5 7777.5 76842.5 ;
      RECT  7522.5 76977.5 7587.5 76842.5 ;
      RECT  7712.5 76977.5 7777.5 76842.5 ;
      RECT  7902.5 76977.5 7967.5 76842.5 ;
      RECT  7902.5 76977.5 7967.5 76842.5 ;
      RECT  7712.5 76977.5 7777.5 76842.5 ;
      RECT  7902.5 76977.5 7967.5 76842.5 ;
      RECT  8092.5 76977.5 8157.5 76842.5 ;
      RECT  8092.5 76977.5 8157.5 76842.5 ;
      RECT  7902.5 76977.5 7967.5 76842.5 ;
      RECT  8262.5 76047.5 8327.5 75912.5 ;
      RECT  8262.5 77022.5 8327.5 76887.5 ;
      RECT  8097.5 76765.0 7962.5 76700.0 ;
      RECT  7907.5 76625.0 7772.5 76560.0 ;
      RECT  7717.5 76485.0 7582.5 76420.0 ;
      RECT  7712.5 76137.5 7777.5 76002.5 ;
      RECT  8092.5 76137.5 8157.5 76002.5 ;
      RECT  8092.5 76977.5 8157.5 76842.5 ;
      RECT  8092.5 76520.0 8157.5 76385.0 ;
      RECT  7582.5 76485.0 7717.5 76420.0 ;
      RECT  7772.5 76625.0 7907.5 76560.0 ;
      RECT  7962.5 76765.0 8097.5 76700.0 ;
      RECT  8092.5 76520.0 8157.5 76385.0 ;
      RECT  7455.0 75827.5 8465.0 75762.5 ;
      RECT  7455.0 77172.5 8465.0 77107.5 ;
      RECT  7522.5 77302.5 7587.5 77107.5 ;
      RECT  7522.5 78142.5 7587.5 78517.5 ;
      RECT  7902.5 78142.5 7967.5 78517.5 ;
      RECT  8262.5 78300.0 8327.5 78485.0 ;
      RECT  8262.5 77140.0 8327.5 77325.0 ;
      RECT  7522.5 78142.5 7587.5 78277.5 ;
      RECT  7712.5 78142.5 7777.5 78277.5 ;
      RECT  7712.5 78142.5 7777.5 78277.5 ;
      RECT  7522.5 78142.5 7587.5 78277.5 ;
      RECT  7712.5 78142.5 7777.5 78277.5 ;
      RECT  7902.5 78142.5 7967.5 78277.5 ;
      RECT  7902.5 78142.5 7967.5 78277.5 ;
      RECT  7712.5 78142.5 7777.5 78277.5 ;
      RECT  7902.5 78142.5 7967.5 78277.5 ;
      RECT  8092.5 78142.5 8157.5 78277.5 ;
      RECT  8092.5 78142.5 8157.5 78277.5 ;
      RECT  7902.5 78142.5 7967.5 78277.5 ;
      RECT  7522.5 77302.5 7587.5 77437.5 ;
      RECT  7712.5 77302.5 7777.5 77437.5 ;
      RECT  7712.5 77302.5 7777.5 77437.5 ;
      RECT  7522.5 77302.5 7587.5 77437.5 ;
      RECT  7712.5 77302.5 7777.5 77437.5 ;
      RECT  7902.5 77302.5 7967.5 77437.5 ;
      RECT  7902.5 77302.5 7967.5 77437.5 ;
      RECT  7712.5 77302.5 7777.5 77437.5 ;
      RECT  7902.5 77302.5 7967.5 77437.5 ;
      RECT  8092.5 77302.5 8157.5 77437.5 ;
      RECT  8092.5 77302.5 8157.5 77437.5 ;
      RECT  7902.5 77302.5 7967.5 77437.5 ;
      RECT  8262.5 78232.5 8327.5 78367.5 ;
      RECT  8262.5 77257.5 8327.5 77392.5 ;
      RECT  8097.5 77515.0 7962.5 77580.0 ;
      RECT  7907.5 77655.0 7772.5 77720.0 ;
      RECT  7717.5 77795.0 7582.5 77860.0 ;
      RECT  7712.5 78142.5 7777.5 78277.5 ;
      RECT  8092.5 78142.5 8157.5 78277.5 ;
      RECT  8092.5 77302.5 8157.5 77437.5 ;
      RECT  8092.5 77760.0 8157.5 77895.0 ;
      RECT  7582.5 77795.0 7717.5 77860.0 ;
      RECT  7772.5 77655.0 7907.5 77720.0 ;
      RECT  7962.5 77515.0 8097.5 77580.0 ;
      RECT  8092.5 77760.0 8157.5 77895.0 ;
      RECT  7455.0 78452.5 8465.0 78517.5 ;
      RECT  7455.0 77107.5 8465.0 77172.5 ;
      RECT  7522.5 79667.5 7587.5 79862.5 ;
      RECT  7522.5 78827.5 7587.5 78452.5 ;
      RECT  7902.5 78827.5 7967.5 78452.5 ;
      RECT  8262.5 78670.0 8327.5 78485.0 ;
      RECT  8262.5 79830.0 8327.5 79645.0 ;
      RECT  7522.5 78827.5 7587.5 78692.5 ;
      RECT  7712.5 78827.5 7777.5 78692.5 ;
      RECT  7712.5 78827.5 7777.5 78692.5 ;
      RECT  7522.5 78827.5 7587.5 78692.5 ;
      RECT  7712.5 78827.5 7777.5 78692.5 ;
      RECT  7902.5 78827.5 7967.5 78692.5 ;
      RECT  7902.5 78827.5 7967.5 78692.5 ;
      RECT  7712.5 78827.5 7777.5 78692.5 ;
      RECT  7902.5 78827.5 7967.5 78692.5 ;
      RECT  8092.5 78827.5 8157.5 78692.5 ;
      RECT  8092.5 78827.5 8157.5 78692.5 ;
      RECT  7902.5 78827.5 7967.5 78692.5 ;
      RECT  7522.5 79667.5 7587.5 79532.5 ;
      RECT  7712.5 79667.5 7777.5 79532.5 ;
      RECT  7712.5 79667.5 7777.5 79532.5 ;
      RECT  7522.5 79667.5 7587.5 79532.5 ;
      RECT  7712.5 79667.5 7777.5 79532.5 ;
      RECT  7902.5 79667.5 7967.5 79532.5 ;
      RECT  7902.5 79667.5 7967.5 79532.5 ;
      RECT  7712.5 79667.5 7777.5 79532.5 ;
      RECT  7902.5 79667.5 7967.5 79532.5 ;
      RECT  8092.5 79667.5 8157.5 79532.5 ;
      RECT  8092.5 79667.5 8157.5 79532.5 ;
      RECT  7902.5 79667.5 7967.5 79532.5 ;
      RECT  8262.5 78737.5 8327.5 78602.5 ;
      RECT  8262.5 79712.5 8327.5 79577.5 ;
      RECT  8097.5 79455.0 7962.5 79390.0 ;
      RECT  7907.5 79315.0 7772.5 79250.0 ;
      RECT  7717.5 79175.0 7582.5 79110.0 ;
      RECT  7712.5 78827.5 7777.5 78692.5 ;
      RECT  8092.5 78827.5 8157.5 78692.5 ;
      RECT  8092.5 79667.5 8157.5 79532.5 ;
      RECT  8092.5 79210.0 8157.5 79075.0 ;
      RECT  7582.5 79175.0 7717.5 79110.0 ;
      RECT  7772.5 79315.0 7907.5 79250.0 ;
      RECT  7962.5 79455.0 8097.5 79390.0 ;
      RECT  8092.5 79210.0 8157.5 79075.0 ;
      RECT  7455.0 78517.5 8465.0 78452.5 ;
      RECT  7455.0 79862.5 8465.0 79797.5 ;
      RECT  7522.5 79992.5 7587.5 79797.5 ;
      RECT  7522.5 80832.5 7587.5 81207.5 ;
      RECT  7902.5 80832.5 7967.5 81207.5 ;
      RECT  8262.5 80990.0 8327.5 81175.0 ;
      RECT  8262.5 79830.0 8327.5 80015.0 ;
      RECT  7522.5 80832.5 7587.5 80967.5 ;
      RECT  7712.5 80832.5 7777.5 80967.5 ;
      RECT  7712.5 80832.5 7777.5 80967.5 ;
      RECT  7522.5 80832.5 7587.5 80967.5 ;
      RECT  7712.5 80832.5 7777.5 80967.5 ;
      RECT  7902.5 80832.5 7967.5 80967.5 ;
      RECT  7902.5 80832.5 7967.5 80967.5 ;
      RECT  7712.5 80832.5 7777.5 80967.5 ;
      RECT  7902.5 80832.5 7967.5 80967.5 ;
      RECT  8092.5 80832.5 8157.5 80967.5 ;
      RECT  8092.5 80832.5 8157.5 80967.5 ;
      RECT  7902.5 80832.5 7967.5 80967.5 ;
      RECT  7522.5 79992.5 7587.5 80127.5 ;
      RECT  7712.5 79992.5 7777.5 80127.5 ;
      RECT  7712.5 79992.5 7777.5 80127.5 ;
      RECT  7522.5 79992.5 7587.5 80127.5 ;
      RECT  7712.5 79992.5 7777.5 80127.5 ;
      RECT  7902.5 79992.5 7967.5 80127.5 ;
      RECT  7902.5 79992.5 7967.5 80127.5 ;
      RECT  7712.5 79992.5 7777.5 80127.5 ;
      RECT  7902.5 79992.5 7967.5 80127.5 ;
      RECT  8092.5 79992.5 8157.5 80127.5 ;
      RECT  8092.5 79992.5 8157.5 80127.5 ;
      RECT  7902.5 79992.5 7967.5 80127.5 ;
      RECT  8262.5 80922.5 8327.5 81057.5 ;
      RECT  8262.5 79947.5 8327.5 80082.5 ;
      RECT  8097.5 80205.0 7962.5 80270.0 ;
      RECT  7907.5 80345.0 7772.5 80410.0 ;
      RECT  7717.5 80485.0 7582.5 80550.0 ;
      RECT  7712.5 80832.5 7777.5 80967.5 ;
      RECT  8092.5 80832.5 8157.5 80967.5 ;
      RECT  8092.5 79992.5 8157.5 80127.5 ;
      RECT  8092.5 80450.0 8157.5 80585.0 ;
      RECT  7582.5 80485.0 7717.5 80550.0 ;
      RECT  7772.5 80345.0 7907.5 80410.0 ;
      RECT  7962.5 80205.0 8097.5 80270.0 ;
      RECT  8092.5 80450.0 8157.5 80585.0 ;
      RECT  7455.0 81142.5 8465.0 81207.5 ;
      RECT  7455.0 79797.5 8465.0 79862.5 ;
      RECT  7522.5 82357.5 7587.5 82552.5 ;
      RECT  7522.5 81517.5 7587.5 81142.5 ;
      RECT  7902.5 81517.5 7967.5 81142.5 ;
      RECT  8262.5 81360.0 8327.5 81175.0 ;
      RECT  8262.5 82520.0 8327.5 82335.0 ;
      RECT  7522.5 81517.5 7587.5 81382.5 ;
      RECT  7712.5 81517.5 7777.5 81382.5 ;
      RECT  7712.5 81517.5 7777.5 81382.5 ;
      RECT  7522.5 81517.5 7587.5 81382.5 ;
      RECT  7712.5 81517.5 7777.5 81382.5 ;
      RECT  7902.5 81517.5 7967.5 81382.5 ;
      RECT  7902.5 81517.5 7967.5 81382.5 ;
      RECT  7712.5 81517.5 7777.5 81382.5 ;
      RECT  7902.5 81517.5 7967.5 81382.5 ;
      RECT  8092.5 81517.5 8157.5 81382.5 ;
      RECT  8092.5 81517.5 8157.5 81382.5 ;
      RECT  7902.5 81517.5 7967.5 81382.5 ;
      RECT  7522.5 82357.5 7587.5 82222.5 ;
      RECT  7712.5 82357.5 7777.5 82222.5 ;
      RECT  7712.5 82357.5 7777.5 82222.5 ;
      RECT  7522.5 82357.5 7587.5 82222.5 ;
      RECT  7712.5 82357.5 7777.5 82222.5 ;
      RECT  7902.5 82357.5 7967.5 82222.5 ;
      RECT  7902.5 82357.5 7967.5 82222.5 ;
      RECT  7712.5 82357.5 7777.5 82222.5 ;
      RECT  7902.5 82357.5 7967.5 82222.5 ;
      RECT  8092.5 82357.5 8157.5 82222.5 ;
      RECT  8092.5 82357.5 8157.5 82222.5 ;
      RECT  7902.5 82357.5 7967.5 82222.5 ;
      RECT  8262.5 81427.5 8327.5 81292.5 ;
      RECT  8262.5 82402.5 8327.5 82267.5 ;
      RECT  8097.5 82145.0 7962.5 82080.0 ;
      RECT  7907.5 82005.0 7772.5 81940.0 ;
      RECT  7717.5 81865.0 7582.5 81800.0 ;
      RECT  7712.5 81517.5 7777.5 81382.5 ;
      RECT  8092.5 81517.5 8157.5 81382.5 ;
      RECT  8092.5 82357.5 8157.5 82222.5 ;
      RECT  8092.5 81900.0 8157.5 81765.0 ;
      RECT  7582.5 81865.0 7717.5 81800.0 ;
      RECT  7772.5 82005.0 7907.5 81940.0 ;
      RECT  7962.5 82145.0 8097.5 82080.0 ;
      RECT  8092.5 81900.0 8157.5 81765.0 ;
      RECT  7455.0 81207.5 8465.0 81142.5 ;
      RECT  7455.0 82552.5 8465.0 82487.5 ;
      RECT  7522.5 82682.5 7587.5 82487.5 ;
      RECT  7522.5 83522.5 7587.5 83897.5 ;
      RECT  7902.5 83522.5 7967.5 83897.5 ;
      RECT  8262.5 83680.0 8327.5 83865.0 ;
      RECT  8262.5 82520.0 8327.5 82705.0 ;
      RECT  7522.5 83522.5 7587.5 83657.5 ;
      RECT  7712.5 83522.5 7777.5 83657.5 ;
      RECT  7712.5 83522.5 7777.5 83657.5 ;
      RECT  7522.5 83522.5 7587.5 83657.5 ;
      RECT  7712.5 83522.5 7777.5 83657.5 ;
      RECT  7902.5 83522.5 7967.5 83657.5 ;
      RECT  7902.5 83522.5 7967.5 83657.5 ;
      RECT  7712.5 83522.5 7777.5 83657.5 ;
      RECT  7902.5 83522.5 7967.5 83657.5 ;
      RECT  8092.5 83522.5 8157.5 83657.5 ;
      RECT  8092.5 83522.5 8157.5 83657.5 ;
      RECT  7902.5 83522.5 7967.5 83657.5 ;
      RECT  7522.5 82682.5 7587.5 82817.5 ;
      RECT  7712.5 82682.5 7777.5 82817.5 ;
      RECT  7712.5 82682.5 7777.5 82817.5 ;
      RECT  7522.5 82682.5 7587.5 82817.5 ;
      RECT  7712.5 82682.5 7777.5 82817.5 ;
      RECT  7902.5 82682.5 7967.5 82817.5 ;
      RECT  7902.5 82682.5 7967.5 82817.5 ;
      RECT  7712.5 82682.5 7777.5 82817.5 ;
      RECT  7902.5 82682.5 7967.5 82817.5 ;
      RECT  8092.5 82682.5 8157.5 82817.5 ;
      RECT  8092.5 82682.5 8157.5 82817.5 ;
      RECT  7902.5 82682.5 7967.5 82817.5 ;
      RECT  8262.5 83612.5 8327.5 83747.5 ;
      RECT  8262.5 82637.5 8327.5 82772.5 ;
      RECT  8097.5 82895.0 7962.5 82960.0 ;
      RECT  7907.5 83035.0 7772.5 83100.0 ;
      RECT  7717.5 83175.0 7582.5 83240.0 ;
      RECT  7712.5 83522.5 7777.5 83657.5 ;
      RECT  8092.5 83522.5 8157.5 83657.5 ;
      RECT  8092.5 82682.5 8157.5 82817.5 ;
      RECT  8092.5 83140.0 8157.5 83275.0 ;
      RECT  7582.5 83175.0 7717.5 83240.0 ;
      RECT  7772.5 83035.0 7907.5 83100.0 ;
      RECT  7962.5 82895.0 8097.5 82960.0 ;
      RECT  8092.5 83140.0 8157.5 83275.0 ;
      RECT  7455.0 83832.5 8465.0 83897.5 ;
      RECT  7455.0 82487.5 8465.0 82552.5 ;
      RECT  7522.5 85047.5 7587.5 85242.5 ;
      RECT  7522.5 84207.5 7587.5 83832.5 ;
      RECT  7902.5 84207.5 7967.5 83832.5 ;
      RECT  8262.5 84050.0 8327.5 83865.0 ;
      RECT  8262.5 85210.0 8327.5 85025.0 ;
      RECT  7522.5 84207.5 7587.5 84072.5 ;
      RECT  7712.5 84207.5 7777.5 84072.5 ;
      RECT  7712.5 84207.5 7777.5 84072.5 ;
      RECT  7522.5 84207.5 7587.5 84072.5 ;
      RECT  7712.5 84207.5 7777.5 84072.5 ;
      RECT  7902.5 84207.5 7967.5 84072.5 ;
      RECT  7902.5 84207.5 7967.5 84072.5 ;
      RECT  7712.5 84207.5 7777.5 84072.5 ;
      RECT  7902.5 84207.5 7967.5 84072.5 ;
      RECT  8092.5 84207.5 8157.5 84072.5 ;
      RECT  8092.5 84207.5 8157.5 84072.5 ;
      RECT  7902.5 84207.5 7967.5 84072.5 ;
      RECT  7522.5 85047.5 7587.5 84912.5 ;
      RECT  7712.5 85047.5 7777.5 84912.5 ;
      RECT  7712.5 85047.5 7777.5 84912.5 ;
      RECT  7522.5 85047.5 7587.5 84912.5 ;
      RECT  7712.5 85047.5 7777.5 84912.5 ;
      RECT  7902.5 85047.5 7967.5 84912.5 ;
      RECT  7902.5 85047.5 7967.5 84912.5 ;
      RECT  7712.5 85047.5 7777.5 84912.5 ;
      RECT  7902.5 85047.5 7967.5 84912.5 ;
      RECT  8092.5 85047.5 8157.5 84912.5 ;
      RECT  8092.5 85047.5 8157.5 84912.5 ;
      RECT  7902.5 85047.5 7967.5 84912.5 ;
      RECT  8262.5 84117.5 8327.5 83982.5 ;
      RECT  8262.5 85092.5 8327.5 84957.5 ;
      RECT  8097.5 84835.0 7962.5 84770.0 ;
      RECT  7907.5 84695.0 7772.5 84630.0 ;
      RECT  7717.5 84555.0 7582.5 84490.0 ;
      RECT  7712.5 84207.5 7777.5 84072.5 ;
      RECT  8092.5 84207.5 8157.5 84072.5 ;
      RECT  8092.5 85047.5 8157.5 84912.5 ;
      RECT  8092.5 84590.0 8157.5 84455.0 ;
      RECT  7582.5 84555.0 7717.5 84490.0 ;
      RECT  7772.5 84695.0 7907.5 84630.0 ;
      RECT  7962.5 84835.0 8097.5 84770.0 ;
      RECT  8092.5 84590.0 8157.5 84455.0 ;
      RECT  7455.0 83897.5 8465.0 83832.5 ;
      RECT  7455.0 85242.5 8465.0 85177.5 ;
      RECT  7522.5 85372.5 7587.5 85177.5 ;
      RECT  7522.5 86212.5 7587.5 86587.5 ;
      RECT  7902.5 86212.5 7967.5 86587.5 ;
      RECT  8262.5 86370.0 8327.5 86555.0 ;
      RECT  8262.5 85210.0 8327.5 85395.0 ;
      RECT  7522.5 86212.5 7587.5 86347.5 ;
      RECT  7712.5 86212.5 7777.5 86347.5 ;
      RECT  7712.5 86212.5 7777.5 86347.5 ;
      RECT  7522.5 86212.5 7587.5 86347.5 ;
      RECT  7712.5 86212.5 7777.5 86347.5 ;
      RECT  7902.5 86212.5 7967.5 86347.5 ;
      RECT  7902.5 86212.5 7967.5 86347.5 ;
      RECT  7712.5 86212.5 7777.5 86347.5 ;
      RECT  7902.5 86212.5 7967.5 86347.5 ;
      RECT  8092.5 86212.5 8157.5 86347.5 ;
      RECT  8092.5 86212.5 8157.5 86347.5 ;
      RECT  7902.5 86212.5 7967.5 86347.5 ;
      RECT  7522.5 85372.5 7587.5 85507.5 ;
      RECT  7712.5 85372.5 7777.5 85507.5 ;
      RECT  7712.5 85372.5 7777.5 85507.5 ;
      RECT  7522.5 85372.5 7587.5 85507.5 ;
      RECT  7712.5 85372.5 7777.5 85507.5 ;
      RECT  7902.5 85372.5 7967.5 85507.5 ;
      RECT  7902.5 85372.5 7967.5 85507.5 ;
      RECT  7712.5 85372.5 7777.5 85507.5 ;
      RECT  7902.5 85372.5 7967.5 85507.5 ;
      RECT  8092.5 85372.5 8157.5 85507.5 ;
      RECT  8092.5 85372.5 8157.5 85507.5 ;
      RECT  7902.5 85372.5 7967.5 85507.5 ;
      RECT  8262.5 86302.5 8327.5 86437.5 ;
      RECT  8262.5 85327.5 8327.5 85462.5 ;
      RECT  8097.5 85585.0 7962.5 85650.0 ;
      RECT  7907.5 85725.0 7772.5 85790.0 ;
      RECT  7717.5 85865.0 7582.5 85930.0 ;
      RECT  7712.5 86212.5 7777.5 86347.5 ;
      RECT  8092.5 86212.5 8157.5 86347.5 ;
      RECT  8092.5 85372.5 8157.5 85507.5 ;
      RECT  8092.5 85830.0 8157.5 85965.0 ;
      RECT  7582.5 85865.0 7717.5 85930.0 ;
      RECT  7772.5 85725.0 7907.5 85790.0 ;
      RECT  7962.5 85585.0 8097.5 85650.0 ;
      RECT  8092.5 85830.0 8157.5 85965.0 ;
      RECT  7455.0 86522.5 8465.0 86587.5 ;
      RECT  7455.0 85177.5 8465.0 85242.5 ;
      RECT  7522.5 87737.5 7587.5 87932.5 ;
      RECT  7522.5 86897.5 7587.5 86522.5 ;
      RECT  7902.5 86897.5 7967.5 86522.5 ;
      RECT  8262.5 86740.0 8327.5 86555.0 ;
      RECT  8262.5 87900.0 8327.5 87715.0 ;
      RECT  7522.5 86897.5 7587.5 86762.5 ;
      RECT  7712.5 86897.5 7777.5 86762.5 ;
      RECT  7712.5 86897.5 7777.5 86762.5 ;
      RECT  7522.5 86897.5 7587.5 86762.5 ;
      RECT  7712.5 86897.5 7777.5 86762.5 ;
      RECT  7902.5 86897.5 7967.5 86762.5 ;
      RECT  7902.5 86897.5 7967.5 86762.5 ;
      RECT  7712.5 86897.5 7777.5 86762.5 ;
      RECT  7902.5 86897.5 7967.5 86762.5 ;
      RECT  8092.5 86897.5 8157.5 86762.5 ;
      RECT  8092.5 86897.5 8157.5 86762.5 ;
      RECT  7902.5 86897.5 7967.5 86762.5 ;
      RECT  7522.5 87737.5 7587.5 87602.5 ;
      RECT  7712.5 87737.5 7777.5 87602.5 ;
      RECT  7712.5 87737.5 7777.5 87602.5 ;
      RECT  7522.5 87737.5 7587.5 87602.5 ;
      RECT  7712.5 87737.5 7777.5 87602.5 ;
      RECT  7902.5 87737.5 7967.5 87602.5 ;
      RECT  7902.5 87737.5 7967.5 87602.5 ;
      RECT  7712.5 87737.5 7777.5 87602.5 ;
      RECT  7902.5 87737.5 7967.5 87602.5 ;
      RECT  8092.5 87737.5 8157.5 87602.5 ;
      RECT  8092.5 87737.5 8157.5 87602.5 ;
      RECT  7902.5 87737.5 7967.5 87602.5 ;
      RECT  8262.5 86807.5 8327.5 86672.5 ;
      RECT  8262.5 87782.5 8327.5 87647.5 ;
      RECT  8097.5 87525.0 7962.5 87460.0 ;
      RECT  7907.5 87385.0 7772.5 87320.0 ;
      RECT  7717.5 87245.0 7582.5 87180.0 ;
      RECT  7712.5 86897.5 7777.5 86762.5 ;
      RECT  8092.5 86897.5 8157.5 86762.5 ;
      RECT  8092.5 87737.5 8157.5 87602.5 ;
      RECT  8092.5 87280.0 8157.5 87145.0 ;
      RECT  7582.5 87245.0 7717.5 87180.0 ;
      RECT  7772.5 87385.0 7907.5 87320.0 ;
      RECT  7962.5 87525.0 8097.5 87460.0 ;
      RECT  8092.5 87280.0 8157.5 87145.0 ;
      RECT  7455.0 86587.5 8465.0 86522.5 ;
      RECT  7455.0 87932.5 8465.0 87867.5 ;
      RECT  7522.5 88062.5 7587.5 87867.5 ;
      RECT  7522.5 88902.5 7587.5 89277.5 ;
      RECT  7902.5 88902.5 7967.5 89277.5 ;
      RECT  8262.5 89060.0 8327.5 89245.0 ;
      RECT  8262.5 87900.0 8327.5 88085.0 ;
      RECT  7522.5 88902.5 7587.5 89037.5 ;
      RECT  7712.5 88902.5 7777.5 89037.5 ;
      RECT  7712.5 88902.5 7777.5 89037.5 ;
      RECT  7522.5 88902.5 7587.5 89037.5 ;
      RECT  7712.5 88902.5 7777.5 89037.5 ;
      RECT  7902.5 88902.5 7967.5 89037.5 ;
      RECT  7902.5 88902.5 7967.5 89037.5 ;
      RECT  7712.5 88902.5 7777.5 89037.5 ;
      RECT  7902.5 88902.5 7967.5 89037.5 ;
      RECT  8092.5 88902.5 8157.5 89037.5 ;
      RECT  8092.5 88902.5 8157.5 89037.5 ;
      RECT  7902.5 88902.5 7967.5 89037.5 ;
      RECT  7522.5 88062.5 7587.5 88197.5 ;
      RECT  7712.5 88062.5 7777.5 88197.5 ;
      RECT  7712.5 88062.5 7777.5 88197.5 ;
      RECT  7522.5 88062.5 7587.5 88197.5 ;
      RECT  7712.5 88062.5 7777.5 88197.5 ;
      RECT  7902.5 88062.5 7967.5 88197.5 ;
      RECT  7902.5 88062.5 7967.5 88197.5 ;
      RECT  7712.5 88062.5 7777.5 88197.5 ;
      RECT  7902.5 88062.5 7967.5 88197.5 ;
      RECT  8092.5 88062.5 8157.5 88197.5 ;
      RECT  8092.5 88062.5 8157.5 88197.5 ;
      RECT  7902.5 88062.5 7967.5 88197.5 ;
      RECT  8262.5 88992.5 8327.5 89127.5 ;
      RECT  8262.5 88017.5 8327.5 88152.5 ;
      RECT  8097.5 88275.0 7962.5 88340.0 ;
      RECT  7907.5 88415.0 7772.5 88480.0 ;
      RECT  7717.5 88555.0 7582.5 88620.0 ;
      RECT  7712.5 88902.5 7777.5 89037.5 ;
      RECT  8092.5 88902.5 8157.5 89037.5 ;
      RECT  8092.5 88062.5 8157.5 88197.5 ;
      RECT  8092.5 88520.0 8157.5 88655.0 ;
      RECT  7582.5 88555.0 7717.5 88620.0 ;
      RECT  7772.5 88415.0 7907.5 88480.0 ;
      RECT  7962.5 88275.0 8097.5 88340.0 ;
      RECT  8092.5 88520.0 8157.5 88655.0 ;
      RECT  7455.0 89212.5 8465.0 89277.5 ;
      RECT  7455.0 87867.5 8465.0 87932.5 ;
      RECT  7522.5 90427.5 7587.5 90622.5 ;
      RECT  7522.5 89587.5 7587.5 89212.5 ;
      RECT  7902.5 89587.5 7967.5 89212.5 ;
      RECT  8262.5 89430.0 8327.5 89245.0 ;
      RECT  8262.5 90590.0 8327.5 90405.0 ;
      RECT  7522.5 89587.5 7587.5 89452.5 ;
      RECT  7712.5 89587.5 7777.5 89452.5 ;
      RECT  7712.5 89587.5 7777.5 89452.5 ;
      RECT  7522.5 89587.5 7587.5 89452.5 ;
      RECT  7712.5 89587.5 7777.5 89452.5 ;
      RECT  7902.5 89587.5 7967.5 89452.5 ;
      RECT  7902.5 89587.5 7967.5 89452.5 ;
      RECT  7712.5 89587.5 7777.5 89452.5 ;
      RECT  7902.5 89587.5 7967.5 89452.5 ;
      RECT  8092.5 89587.5 8157.5 89452.5 ;
      RECT  8092.5 89587.5 8157.5 89452.5 ;
      RECT  7902.5 89587.5 7967.5 89452.5 ;
      RECT  7522.5 90427.5 7587.5 90292.5 ;
      RECT  7712.5 90427.5 7777.5 90292.5 ;
      RECT  7712.5 90427.5 7777.5 90292.5 ;
      RECT  7522.5 90427.5 7587.5 90292.5 ;
      RECT  7712.5 90427.5 7777.5 90292.5 ;
      RECT  7902.5 90427.5 7967.5 90292.5 ;
      RECT  7902.5 90427.5 7967.5 90292.5 ;
      RECT  7712.5 90427.5 7777.5 90292.5 ;
      RECT  7902.5 90427.5 7967.5 90292.5 ;
      RECT  8092.5 90427.5 8157.5 90292.5 ;
      RECT  8092.5 90427.5 8157.5 90292.5 ;
      RECT  7902.5 90427.5 7967.5 90292.5 ;
      RECT  8262.5 89497.5 8327.5 89362.5 ;
      RECT  8262.5 90472.5 8327.5 90337.5 ;
      RECT  8097.5 90215.0 7962.5 90150.0 ;
      RECT  7907.5 90075.0 7772.5 90010.0 ;
      RECT  7717.5 89935.0 7582.5 89870.0 ;
      RECT  7712.5 89587.5 7777.5 89452.5 ;
      RECT  8092.5 89587.5 8157.5 89452.5 ;
      RECT  8092.5 90427.5 8157.5 90292.5 ;
      RECT  8092.5 89970.0 8157.5 89835.0 ;
      RECT  7582.5 89935.0 7717.5 89870.0 ;
      RECT  7772.5 90075.0 7907.5 90010.0 ;
      RECT  7962.5 90215.0 8097.5 90150.0 ;
      RECT  8092.5 89970.0 8157.5 89835.0 ;
      RECT  7455.0 89277.5 8465.0 89212.5 ;
      RECT  7455.0 90622.5 8465.0 90557.5 ;
      RECT  7522.5 90752.5 7587.5 90557.5 ;
      RECT  7522.5 91592.5 7587.5 91967.5 ;
      RECT  7902.5 91592.5 7967.5 91967.5 ;
      RECT  8262.5 91750.0 8327.5 91935.0 ;
      RECT  8262.5 90590.0 8327.5 90775.0 ;
      RECT  7522.5 91592.5 7587.5 91727.5 ;
      RECT  7712.5 91592.5 7777.5 91727.5 ;
      RECT  7712.5 91592.5 7777.5 91727.5 ;
      RECT  7522.5 91592.5 7587.5 91727.5 ;
      RECT  7712.5 91592.5 7777.5 91727.5 ;
      RECT  7902.5 91592.5 7967.5 91727.5 ;
      RECT  7902.5 91592.5 7967.5 91727.5 ;
      RECT  7712.5 91592.5 7777.5 91727.5 ;
      RECT  7902.5 91592.5 7967.5 91727.5 ;
      RECT  8092.5 91592.5 8157.5 91727.5 ;
      RECT  8092.5 91592.5 8157.5 91727.5 ;
      RECT  7902.5 91592.5 7967.5 91727.5 ;
      RECT  7522.5 90752.5 7587.5 90887.5 ;
      RECT  7712.5 90752.5 7777.5 90887.5 ;
      RECT  7712.5 90752.5 7777.5 90887.5 ;
      RECT  7522.5 90752.5 7587.5 90887.5 ;
      RECT  7712.5 90752.5 7777.5 90887.5 ;
      RECT  7902.5 90752.5 7967.5 90887.5 ;
      RECT  7902.5 90752.5 7967.5 90887.5 ;
      RECT  7712.5 90752.5 7777.5 90887.5 ;
      RECT  7902.5 90752.5 7967.5 90887.5 ;
      RECT  8092.5 90752.5 8157.5 90887.5 ;
      RECT  8092.5 90752.5 8157.5 90887.5 ;
      RECT  7902.5 90752.5 7967.5 90887.5 ;
      RECT  8262.5 91682.5 8327.5 91817.5 ;
      RECT  8262.5 90707.5 8327.5 90842.5 ;
      RECT  8097.5 90965.0 7962.5 91030.0 ;
      RECT  7907.5 91105.0 7772.5 91170.0 ;
      RECT  7717.5 91245.0 7582.5 91310.0 ;
      RECT  7712.5 91592.5 7777.5 91727.5 ;
      RECT  8092.5 91592.5 8157.5 91727.5 ;
      RECT  8092.5 90752.5 8157.5 90887.5 ;
      RECT  8092.5 91210.0 8157.5 91345.0 ;
      RECT  7582.5 91245.0 7717.5 91310.0 ;
      RECT  7772.5 91105.0 7907.5 91170.0 ;
      RECT  7962.5 90965.0 8097.5 91030.0 ;
      RECT  8092.5 91210.0 8157.5 91345.0 ;
      RECT  7455.0 91902.5 8465.0 91967.5 ;
      RECT  7455.0 90557.5 8465.0 90622.5 ;
      RECT  7522.5 93117.5 7587.5 93312.5 ;
      RECT  7522.5 92277.5 7587.5 91902.5 ;
      RECT  7902.5 92277.5 7967.5 91902.5 ;
      RECT  8262.5 92120.0 8327.5 91935.0 ;
      RECT  8262.5 93280.0 8327.5 93095.0 ;
      RECT  7522.5 92277.5 7587.5 92142.5 ;
      RECT  7712.5 92277.5 7777.5 92142.5 ;
      RECT  7712.5 92277.5 7777.5 92142.5 ;
      RECT  7522.5 92277.5 7587.5 92142.5 ;
      RECT  7712.5 92277.5 7777.5 92142.5 ;
      RECT  7902.5 92277.5 7967.5 92142.5 ;
      RECT  7902.5 92277.5 7967.5 92142.5 ;
      RECT  7712.5 92277.5 7777.5 92142.5 ;
      RECT  7902.5 92277.5 7967.5 92142.5 ;
      RECT  8092.5 92277.5 8157.5 92142.5 ;
      RECT  8092.5 92277.5 8157.5 92142.5 ;
      RECT  7902.5 92277.5 7967.5 92142.5 ;
      RECT  7522.5 93117.5 7587.5 92982.5 ;
      RECT  7712.5 93117.5 7777.5 92982.5 ;
      RECT  7712.5 93117.5 7777.5 92982.5 ;
      RECT  7522.5 93117.5 7587.5 92982.5 ;
      RECT  7712.5 93117.5 7777.5 92982.5 ;
      RECT  7902.5 93117.5 7967.5 92982.5 ;
      RECT  7902.5 93117.5 7967.5 92982.5 ;
      RECT  7712.5 93117.5 7777.5 92982.5 ;
      RECT  7902.5 93117.5 7967.5 92982.5 ;
      RECT  8092.5 93117.5 8157.5 92982.5 ;
      RECT  8092.5 93117.5 8157.5 92982.5 ;
      RECT  7902.5 93117.5 7967.5 92982.5 ;
      RECT  8262.5 92187.5 8327.5 92052.5 ;
      RECT  8262.5 93162.5 8327.5 93027.5 ;
      RECT  8097.5 92905.0 7962.5 92840.0 ;
      RECT  7907.5 92765.0 7772.5 92700.0 ;
      RECT  7717.5 92625.0 7582.5 92560.0 ;
      RECT  7712.5 92277.5 7777.5 92142.5 ;
      RECT  8092.5 92277.5 8157.5 92142.5 ;
      RECT  8092.5 93117.5 8157.5 92982.5 ;
      RECT  8092.5 92660.0 8157.5 92525.0 ;
      RECT  7582.5 92625.0 7717.5 92560.0 ;
      RECT  7772.5 92765.0 7907.5 92700.0 ;
      RECT  7962.5 92905.0 8097.5 92840.0 ;
      RECT  8092.5 92660.0 8157.5 92525.0 ;
      RECT  7455.0 91967.5 8465.0 91902.5 ;
      RECT  7455.0 93312.5 8465.0 93247.5 ;
      RECT  7522.5 93442.5 7587.5 93247.5 ;
      RECT  7522.5 94282.5 7587.5 94657.5 ;
      RECT  7902.5 94282.5 7967.5 94657.5 ;
      RECT  8262.5 94440.0 8327.5 94625.0 ;
      RECT  8262.5 93280.0 8327.5 93465.0 ;
      RECT  7522.5 94282.5 7587.5 94417.5 ;
      RECT  7712.5 94282.5 7777.5 94417.5 ;
      RECT  7712.5 94282.5 7777.5 94417.5 ;
      RECT  7522.5 94282.5 7587.5 94417.5 ;
      RECT  7712.5 94282.5 7777.5 94417.5 ;
      RECT  7902.5 94282.5 7967.5 94417.5 ;
      RECT  7902.5 94282.5 7967.5 94417.5 ;
      RECT  7712.5 94282.5 7777.5 94417.5 ;
      RECT  7902.5 94282.5 7967.5 94417.5 ;
      RECT  8092.5 94282.5 8157.5 94417.5 ;
      RECT  8092.5 94282.5 8157.5 94417.5 ;
      RECT  7902.5 94282.5 7967.5 94417.5 ;
      RECT  7522.5 93442.5 7587.5 93577.5 ;
      RECT  7712.5 93442.5 7777.5 93577.5 ;
      RECT  7712.5 93442.5 7777.5 93577.5 ;
      RECT  7522.5 93442.5 7587.5 93577.5 ;
      RECT  7712.5 93442.5 7777.5 93577.5 ;
      RECT  7902.5 93442.5 7967.5 93577.5 ;
      RECT  7902.5 93442.5 7967.5 93577.5 ;
      RECT  7712.5 93442.5 7777.5 93577.5 ;
      RECT  7902.5 93442.5 7967.5 93577.5 ;
      RECT  8092.5 93442.5 8157.5 93577.5 ;
      RECT  8092.5 93442.5 8157.5 93577.5 ;
      RECT  7902.5 93442.5 7967.5 93577.5 ;
      RECT  8262.5 94372.5 8327.5 94507.5 ;
      RECT  8262.5 93397.5 8327.5 93532.5 ;
      RECT  8097.5 93655.0 7962.5 93720.0 ;
      RECT  7907.5 93795.0 7772.5 93860.0 ;
      RECT  7717.5 93935.0 7582.5 94000.0 ;
      RECT  7712.5 94282.5 7777.5 94417.5 ;
      RECT  8092.5 94282.5 8157.5 94417.5 ;
      RECT  8092.5 93442.5 8157.5 93577.5 ;
      RECT  8092.5 93900.0 8157.5 94035.0 ;
      RECT  7582.5 93935.0 7717.5 94000.0 ;
      RECT  7772.5 93795.0 7907.5 93860.0 ;
      RECT  7962.5 93655.0 8097.5 93720.0 ;
      RECT  8092.5 93900.0 8157.5 94035.0 ;
      RECT  7455.0 94592.5 8465.0 94657.5 ;
      RECT  7455.0 93247.5 8465.0 93312.5 ;
      RECT  7522.5 95807.5 7587.5 96002.5 ;
      RECT  7522.5 94967.5 7587.5 94592.5 ;
      RECT  7902.5 94967.5 7967.5 94592.5 ;
      RECT  8262.5 94810.0 8327.5 94625.0 ;
      RECT  8262.5 95970.0 8327.5 95785.0 ;
      RECT  7522.5 94967.5 7587.5 94832.5 ;
      RECT  7712.5 94967.5 7777.5 94832.5 ;
      RECT  7712.5 94967.5 7777.5 94832.5 ;
      RECT  7522.5 94967.5 7587.5 94832.5 ;
      RECT  7712.5 94967.5 7777.5 94832.5 ;
      RECT  7902.5 94967.5 7967.5 94832.5 ;
      RECT  7902.5 94967.5 7967.5 94832.5 ;
      RECT  7712.5 94967.5 7777.5 94832.5 ;
      RECT  7902.5 94967.5 7967.5 94832.5 ;
      RECT  8092.5 94967.5 8157.5 94832.5 ;
      RECT  8092.5 94967.5 8157.5 94832.5 ;
      RECT  7902.5 94967.5 7967.5 94832.5 ;
      RECT  7522.5 95807.5 7587.5 95672.5 ;
      RECT  7712.5 95807.5 7777.5 95672.5 ;
      RECT  7712.5 95807.5 7777.5 95672.5 ;
      RECT  7522.5 95807.5 7587.5 95672.5 ;
      RECT  7712.5 95807.5 7777.5 95672.5 ;
      RECT  7902.5 95807.5 7967.5 95672.5 ;
      RECT  7902.5 95807.5 7967.5 95672.5 ;
      RECT  7712.5 95807.5 7777.5 95672.5 ;
      RECT  7902.5 95807.5 7967.5 95672.5 ;
      RECT  8092.5 95807.5 8157.5 95672.5 ;
      RECT  8092.5 95807.5 8157.5 95672.5 ;
      RECT  7902.5 95807.5 7967.5 95672.5 ;
      RECT  8262.5 94877.5 8327.5 94742.5 ;
      RECT  8262.5 95852.5 8327.5 95717.5 ;
      RECT  8097.5 95595.0 7962.5 95530.0 ;
      RECT  7907.5 95455.0 7772.5 95390.0 ;
      RECT  7717.5 95315.0 7582.5 95250.0 ;
      RECT  7712.5 94967.5 7777.5 94832.5 ;
      RECT  8092.5 94967.5 8157.5 94832.5 ;
      RECT  8092.5 95807.5 8157.5 95672.5 ;
      RECT  8092.5 95350.0 8157.5 95215.0 ;
      RECT  7582.5 95315.0 7717.5 95250.0 ;
      RECT  7772.5 95455.0 7907.5 95390.0 ;
      RECT  7962.5 95595.0 8097.5 95530.0 ;
      RECT  8092.5 95350.0 8157.5 95215.0 ;
      RECT  7455.0 94657.5 8465.0 94592.5 ;
      RECT  7455.0 96002.5 8465.0 95937.5 ;
      RECT  7522.5 96132.5 7587.5 95937.5 ;
      RECT  7522.5 96972.5 7587.5 97347.5 ;
      RECT  7902.5 96972.5 7967.5 97347.5 ;
      RECT  8262.5 97130.0 8327.5 97315.0 ;
      RECT  8262.5 95970.0 8327.5 96155.0 ;
      RECT  7522.5 96972.5 7587.5 97107.5 ;
      RECT  7712.5 96972.5 7777.5 97107.5 ;
      RECT  7712.5 96972.5 7777.5 97107.5 ;
      RECT  7522.5 96972.5 7587.5 97107.5 ;
      RECT  7712.5 96972.5 7777.5 97107.5 ;
      RECT  7902.5 96972.5 7967.5 97107.5 ;
      RECT  7902.5 96972.5 7967.5 97107.5 ;
      RECT  7712.5 96972.5 7777.5 97107.5 ;
      RECT  7902.5 96972.5 7967.5 97107.5 ;
      RECT  8092.5 96972.5 8157.5 97107.5 ;
      RECT  8092.5 96972.5 8157.5 97107.5 ;
      RECT  7902.5 96972.5 7967.5 97107.5 ;
      RECT  7522.5 96132.5 7587.5 96267.5 ;
      RECT  7712.5 96132.5 7777.5 96267.5 ;
      RECT  7712.5 96132.5 7777.5 96267.5 ;
      RECT  7522.5 96132.5 7587.5 96267.5 ;
      RECT  7712.5 96132.5 7777.5 96267.5 ;
      RECT  7902.5 96132.5 7967.5 96267.5 ;
      RECT  7902.5 96132.5 7967.5 96267.5 ;
      RECT  7712.5 96132.5 7777.5 96267.5 ;
      RECT  7902.5 96132.5 7967.5 96267.5 ;
      RECT  8092.5 96132.5 8157.5 96267.5 ;
      RECT  8092.5 96132.5 8157.5 96267.5 ;
      RECT  7902.5 96132.5 7967.5 96267.5 ;
      RECT  8262.5 97062.5 8327.5 97197.5 ;
      RECT  8262.5 96087.5 8327.5 96222.5 ;
      RECT  8097.5 96345.0 7962.5 96410.0 ;
      RECT  7907.5 96485.0 7772.5 96550.0 ;
      RECT  7717.5 96625.0 7582.5 96690.0 ;
      RECT  7712.5 96972.5 7777.5 97107.5 ;
      RECT  8092.5 96972.5 8157.5 97107.5 ;
      RECT  8092.5 96132.5 8157.5 96267.5 ;
      RECT  8092.5 96590.0 8157.5 96725.0 ;
      RECT  7582.5 96625.0 7717.5 96690.0 ;
      RECT  7772.5 96485.0 7907.5 96550.0 ;
      RECT  7962.5 96345.0 8097.5 96410.0 ;
      RECT  8092.5 96590.0 8157.5 96725.0 ;
      RECT  7455.0 97282.5 8465.0 97347.5 ;
      RECT  7455.0 95937.5 8465.0 96002.5 ;
      RECT  7522.5 98497.5 7587.5 98692.5 ;
      RECT  7522.5 97657.5 7587.5 97282.5 ;
      RECT  7902.5 97657.5 7967.5 97282.5 ;
      RECT  8262.5 97500.0 8327.5 97315.0 ;
      RECT  8262.5 98660.0 8327.5 98475.0 ;
      RECT  7522.5 97657.5 7587.5 97522.5 ;
      RECT  7712.5 97657.5 7777.5 97522.5 ;
      RECT  7712.5 97657.5 7777.5 97522.5 ;
      RECT  7522.5 97657.5 7587.5 97522.5 ;
      RECT  7712.5 97657.5 7777.5 97522.5 ;
      RECT  7902.5 97657.5 7967.5 97522.5 ;
      RECT  7902.5 97657.5 7967.5 97522.5 ;
      RECT  7712.5 97657.5 7777.5 97522.5 ;
      RECT  7902.5 97657.5 7967.5 97522.5 ;
      RECT  8092.5 97657.5 8157.5 97522.5 ;
      RECT  8092.5 97657.5 8157.5 97522.5 ;
      RECT  7902.5 97657.5 7967.5 97522.5 ;
      RECT  7522.5 98497.5 7587.5 98362.5 ;
      RECT  7712.5 98497.5 7777.5 98362.5 ;
      RECT  7712.5 98497.5 7777.5 98362.5 ;
      RECT  7522.5 98497.5 7587.5 98362.5 ;
      RECT  7712.5 98497.5 7777.5 98362.5 ;
      RECT  7902.5 98497.5 7967.5 98362.5 ;
      RECT  7902.5 98497.5 7967.5 98362.5 ;
      RECT  7712.5 98497.5 7777.5 98362.5 ;
      RECT  7902.5 98497.5 7967.5 98362.5 ;
      RECT  8092.5 98497.5 8157.5 98362.5 ;
      RECT  8092.5 98497.5 8157.5 98362.5 ;
      RECT  7902.5 98497.5 7967.5 98362.5 ;
      RECT  8262.5 97567.5 8327.5 97432.5 ;
      RECT  8262.5 98542.5 8327.5 98407.5 ;
      RECT  8097.5 98285.0 7962.5 98220.0 ;
      RECT  7907.5 98145.0 7772.5 98080.0 ;
      RECT  7717.5 98005.0 7582.5 97940.0 ;
      RECT  7712.5 97657.5 7777.5 97522.5 ;
      RECT  8092.5 97657.5 8157.5 97522.5 ;
      RECT  8092.5 98497.5 8157.5 98362.5 ;
      RECT  8092.5 98040.0 8157.5 97905.0 ;
      RECT  7582.5 98005.0 7717.5 97940.0 ;
      RECT  7772.5 98145.0 7907.5 98080.0 ;
      RECT  7962.5 98285.0 8097.5 98220.0 ;
      RECT  8092.5 98040.0 8157.5 97905.0 ;
      RECT  7455.0 97347.5 8465.0 97282.5 ;
      RECT  7455.0 98692.5 8465.0 98627.5 ;
      RECT  7522.5 98822.5 7587.5 98627.5 ;
      RECT  7522.5 99662.5 7587.5 100037.5 ;
      RECT  7902.5 99662.5 7967.5 100037.5 ;
      RECT  8262.5 99820.0 8327.5 100005.0 ;
      RECT  8262.5 98660.0 8327.5 98845.0 ;
      RECT  7522.5 99662.5 7587.5 99797.5 ;
      RECT  7712.5 99662.5 7777.5 99797.5 ;
      RECT  7712.5 99662.5 7777.5 99797.5 ;
      RECT  7522.5 99662.5 7587.5 99797.5 ;
      RECT  7712.5 99662.5 7777.5 99797.5 ;
      RECT  7902.5 99662.5 7967.5 99797.5 ;
      RECT  7902.5 99662.5 7967.5 99797.5 ;
      RECT  7712.5 99662.5 7777.5 99797.5 ;
      RECT  7902.5 99662.5 7967.5 99797.5 ;
      RECT  8092.5 99662.5 8157.5 99797.5 ;
      RECT  8092.5 99662.5 8157.5 99797.5 ;
      RECT  7902.5 99662.5 7967.5 99797.5 ;
      RECT  7522.5 98822.5 7587.5 98957.5 ;
      RECT  7712.5 98822.5 7777.5 98957.5 ;
      RECT  7712.5 98822.5 7777.5 98957.5 ;
      RECT  7522.5 98822.5 7587.5 98957.5 ;
      RECT  7712.5 98822.5 7777.5 98957.5 ;
      RECT  7902.5 98822.5 7967.5 98957.5 ;
      RECT  7902.5 98822.5 7967.5 98957.5 ;
      RECT  7712.5 98822.5 7777.5 98957.5 ;
      RECT  7902.5 98822.5 7967.5 98957.5 ;
      RECT  8092.5 98822.5 8157.5 98957.5 ;
      RECT  8092.5 98822.5 8157.5 98957.5 ;
      RECT  7902.5 98822.5 7967.5 98957.5 ;
      RECT  8262.5 99752.5 8327.5 99887.5 ;
      RECT  8262.5 98777.5 8327.5 98912.5 ;
      RECT  8097.5 99035.0 7962.5 99100.0 ;
      RECT  7907.5 99175.0 7772.5 99240.0 ;
      RECT  7717.5 99315.0 7582.5 99380.0 ;
      RECT  7712.5 99662.5 7777.5 99797.5 ;
      RECT  8092.5 99662.5 8157.5 99797.5 ;
      RECT  8092.5 98822.5 8157.5 98957.5 ;
      RECT  8092.5 99280.0 8157.5 99415.0 ;
      RECT  7582.5 99315.0 7717.5 99380.0 ;
      RECT  7772.5 99175.0 7907.5 99240.0 ;
      RECT  7962.5 99035.0 8097.5 99100.0 ;
      RECT  8092.5 99280.0 8157.5 99415.0 ;
      RECT  7455.0 99972.5 8465.0 100037.5 ;
      RECT  7455.0 98627.5 8465.0 98692.5 ;
      RECT  7522.5 101187.5 7587.5 101382.5 ;
      RECT  7522.5 100347.5 7587.5 99972.5 ;
      RECT  7902.5 100347.5 7967.5 99972.5 ;
      RECT  8262.5 100190.0 8327.5 100005.0 ;
      RECT  8262.5 101350.0 8327.5 101165.0 ;
      RECT  7522.5 100347.5 7587.5 100212.5 ;
      RECT  7712.5 100347.5 7777.5 100212.5 ;
      RECT  7712.5 100347.5 7777.5 100212.5 ;
      RECT  7522.5 100347.5 7587.5 100212.5 ;
      RECT  7712.5 100347.5 7777.5 100212.5 ;
      RECT  7902.5 100347.5 7967.5 100212.5 ;
      RECT  7902.5 100347.5 7967.5 100212.5 ;
      RECT  7712.5 100347.5 7777.5 100212.5 ;
      RECT  7902.5 100347.5 7967.5 100212.5 ;
      RECT  8092.5 100347.5 8157.5 100212.5 ;
      RECT  8092.5 100347.5 8157.5 100212.5 ;
      RECT  7902.5 100347.5 7967.5 100212.5 ;
      RECT  7522.5 101187.5 7587.5 101052.5 ;
      RECT  7712.5 101187.5 7777.5 101052.5 ;
      RECT  7712.5 101187.5 7777.5 101052.5 ;
      RECT  7522.5 101187.5 7587.5 101052.5 ;
      RECT  7712.5 101187.5 7777.5 101052.5 ;
      RECT  7902.5 101187.5 7967.5 101052.5 ;
      RECT  7902.5 101187.5 7967.5 101052.5 ;
      RECT  7712.5 101187.5 7777.5 101052.5 ;
      RECT  7902.5 101187.5 7967.5 101052.5 ;
      RECT  8092.5 101187.5 8157.5 101052.5 ;
      RECT  8092.5 101187.5 8157.5 101052.5 ;
      RECT  7902.5 101187.5 7967.5 101052.5 ;
      RECT  8262.5 100257.5 8327.5 100122.5 ;
      RECT  8262.5 101232.5 8327.5 101097.5 ;
      RECT  8097.5 100975.0 7962.5 100910.0 ;
      RECT  7907.5 100835.0 7772.5 100770.0 ;
      RECT  7717.5 100695.0 7582.5 100630.0 ;
      RECT  7712.5 100347.5 7777.5 100212.5 ;
      RECT  8092.5 100347.5 8157.5 100212.5 ;
      RECT  8092.5 101187.5 8157.5 101052.5 ;
      RECT  8092.5 100730.0 8157.5 100595.0 ;
      RECT  7582.5 100695.0 7717.5 100630.0 ;
      RECT  7772.5 100835.0 7907.5 100770.0 ;
      RECT  7962.5 100975.0 8097.5 100910.0 ;
      RECT  8092.5 100730.0 8157.5 100595.0 ;
      RECT  7455.0 100037.5 8465.0 99972.5 ;
      RECT  7455.0 101382.5 8465.0 101317.5 ;
      RECT  7522.5 101512.5 7587.5 101317.5 ;
      RECT  7522.5 102352.5 7587.5 102727.5 ;
      RECT  7902.5 102352.5 7967.5 102727.5 ;
      RECT  8262.5 102510.0 8327.5 102695.0 ;
      RECT  8262.5 101350.0 8327.5 101535.0 ;
      RECT  7522.5 102352.5 7587.5 102487.5 ;
      RECT  7712.5 102352.5 7777.5 102487.5 ;
      RECT  7712.5 102352.5 7777.5 102487.5 ;
      RECT  7522.5 102352.5 7587.5 102487.5 ;
      RECT  7712.5 102352.5 7777.5 102487.5 ;
      RECT  7902.5 102352.5 7967.5 102487.5 ;
      RECT  7902.5 102352.5 7967.5 102487.5 ;
      RECT  7712.5 102352.5 7777.5 102487.5 ;
      RECT  7902.5 102352.5 7967.5 102487.5 ;
      RECT  8092.5 102352.5 8157.5 102487.5 ;
      RECT  8092.5 102352.5 8157.5 102487.5 ;
      RECT  7902.5 102352.5 7967.5 102487.5 ;
      RECT  7522.5 101512.5 7587.5 101647.5 ;
      RECT  7712.5 101512.5 7777.5 101647.5 ;
      RECT  7712.5 101512.5 7777.5 101647.5 ;
      RECT  7522.5 101512.5 7587.5 101647.5 ;
      RECT  7712.5 101512.5 7777.5 101647.5 ;
      RECT  7902.5 101512.5 7967.5 101647.5 ;
      RECT  7902.5 101512.5 7967.5 101647.5 ;
      RECT  7712.5 101512.5 7777.5 101647.5 ;
      RECT  7902.5 101512.5 7967.5 101647.5 ;
      RECT  8092.5 101512.5 8157.5 101647.5 ;
      RECT  8092.5 101512.5 8157.5 101647.5 ;
      RECT  7902.5 101512.5 7967.5 101647.5 ;
      RECT  8262.5 102442.5 8327.5 102577.5 ;
      RECT  8262.5 101467.5 8327.5 101602.5 ;
      RECT  8097.5 101725.0 7962.5 101790.0 ;
      RECT  7907.5 101865.0 7772.5 101930.0 ;
      RECT  7717.5 102005.0 7582.5 102070.0 ;
      RECT  7712.5 102352.5 7777.5 102487.5 ;
      RECT  8092.5 102352.5 8157.5 102487.5 ;
      RECT  8092.5 101512.5 8157.5 101647.5 ;
      RECT  8092.5 101970.0 8157.5 102105.0 ;
      RECT  7582.5 102005.0 7717.5 102070.0 ;
      RECT  7772.5 101865.0 7907.5 101930.0 ;
      RECT  7962.5 101725.0 8097.5 101790.0 ;
      RECT  8092.5 101970.0 8157.5 102105.0 ;
      RECT  7455.0 102662.5 8465.0 102727.5 ;
      RECT  7455.0 101317.5 8465.0 101382.5 ;
      RECT  7522.5 103877.5 7587.5 104072.5 ;
      RECT  7522.5 103037.5 7587.5 102662.5 ;
      RECT  7902.5 103037.5 7967.5 102662.5 ;
      RECT  8262.5 102880.0 8327.5 102695.0 ;
      RECT  8262.5 104040.0 8327.5 103855.0 ;
      RECT  7522.5 103037.5 7587.5 102902.5 ;
      RECT  7712.5 103037.5 7777.5 102902.5 ;
      RECT  7712.5 103037.5 7777.5 102902.5 ;
      RECT  7522.5 103037.5 7587.5 102902.5 ;
      RECT  7712.5 103037.5 7777.5 102902.5 ;
      RECT  7902.5 103037.5 7967.5 102902.5 ;
      RECT  7902.5 103037.5 7967.5 102902.5 ;
      RECT  7712.5 103037.5 7777.5 102902.5 ;
      RECT  7902.5 103037.5 7967.5 102902.5 ;
      RECT  8092.5 103037.5 8157.5 102902.5 ;
      RECT  8092.5 103037.5 8157.5 102902.5 ;
      RECT  7902.5 103037.5 7967.5 102902.5 ;
      RECT  7522.5 103877.5 7587.5 103742.5 ;
      RECT  7712.5 103877.5 7777.5 103742.5 ;
      RECT  7712.5 103877.5 7777.5 103742.5 ;
      RECT  7522.5 103877.5 7587.5 103742.5 ;
      RECT  7712.5 103877.5 7777.5 103742.5 ;
      RECT  7902.5 103877.5 7967.5 103742.5 ;
      RECT  7902.5 103877.5 7967.5 103742.5 ;
      RECT  7712.5 103877.5 7777.5 103742.5 ;
      RECT  7902.5 103877.5 7967.5 103742.5 ;
      RECT  8092.5 103877.5 8157.5 103742.5 ;
      RECT  8092.5 103877.5 8157.5 103742.5 ;
      RECT  7902.5 103877.5 7967.5 103742.5 ;
      RECT  8262.5 102947.5 8327.5 102812.5 ;
      RECT  8262.5 103922.5 8327.5 103787.5 ;
      RECT  8097.5 103665.0 7962.5 103600.0 ;
      RECT  7907.5 103525.0 7772.5 103460.0 ;
      RECT  7717.5 103385.0 7582.5 103320.0 ;
      RECT  7712.5 103037.5 7777.5 102902.5 ;
      RECT  8092.5 103037.5 8157.5 102902.5 ;
      RECT  8092.5 103877.5 8157.5 103742.5 ;
      RECT  8092.5 103420.0 8157.5 103285.0 ;
      RECT  7582.5 103385.0 7717.5 103320.0 ;
      RECT  7772.5 103525.0 7907.5 103460.0 ;
      RECT  7962.5 103665.0 8097.5 103600.0 ;
      RECT  8092.5 103420.0 8157.5 103285.0 ;
      RECT  7455.0 102727.5 8465.0 102662.5 ;
      RECT  7455.0 104072.5 8465.0 104007.5 ;
      RECT  7522.5 104202.5 7587.5 104007.5 ;
      RECT  7522.5 105042.5 7587.5 105417.5 ;
      RECT  7902.5 105042.5 7967.5 105417.5 ;
      RECT  8262.5 105200.0 8327.5 105385.0 ;
      RECT  8262.5 104040.0 8327.5 104225.0 ;
      RECT  7522.5 105042.5 7587.5 105177.5 ;
      RECT  7712.5 105042.5 7777.5 105177.5 ;
      RECT  7712.5 105042.5 7777.5 105177.5 ;
      RECT  7522.5 105042.5 7587.5 105177.5 ;
      RECT  7712.5 105042.5 7777.5 105177.5 ;
      RECT  7902.5 105042.5 7967.5 105177.5 ;
      RECT  7902.5 105042.5 7967.5 105177.5 ;
      RECT  7712.5 105042.5 7777.5 105177.5 ;
      RECT  7902.5 105042.5 7967.5 105177.5 ;
      RECT  8092.5 105042.5 8157.5 105177.5 ;
      RECT  8092.5 105042.5 8157.5 105177.5 ;
      RECT  7902.5 105042.5 7967.5 105177.5 ;
      RECT  7522.5 104202.5 7587.5 104337.5 ;
      RECT  7712.5 104202.5 7777.5 104337.5 ;
      RECT  7712.5 104202.5 7777.5 104337.5 ;
      RECT  7522.5 104202.5 7587.5 104337.5 ;
      RECT  7712.5 104202.5 7777.5 104337.5 ;
      RECT  7902.5 104202.5 7967.5 104337.5 ;
      RECT  7902.5 104202.5 7967.5 104337.5 ;
      RECT  7712.5 104202.5 7777.5 104337.5 ;
      RECT  7902.5 104202.5 7967.5 104337.5 ;
      RECT  8092.5 104202.5 8157.5 104337.5 ;
      RECT  8092.5 104202.5 8157.5 104337.5 ;
      RECT  7902.5 104202.5 7967.5 104337.5 ;
      RECT  8262.5 105132.5 8327.5 105267.5 ;
      RECT  8262.5 104157.5 8327.5 104292.5 ;
      RECT  8097.5 104415.0 7962.5 104480.0 ;
      RECT  7907.5 104555.0 7772.5 104620.0 ;
      RECT  7717.5 104695.0 7582.5 104760.0 ;
      RECT  7712.5 105042.5 7777.5 105177.5 ;
      RECT  8092.5 105042.5 8157.5 105177.5 ;
      RECT  8092.5 104202.5 8157.5 104337.5 ;
      RECT  8092.5 104660.0 8157.5 104795.0 ;
      RECT  7582.5 104695.0 7717.5 104760.0 ;
      RECT  7772.5 104555.0 7907.5 104620.0 ;
      RECT  7962.5 104415.0 8097.5 104480.0 ;
      RECT  8092.5 104660.0 8157.5 104795.0 ;
      RECT  7455.0 105352.5 8465.0 105417.5 ;
      RECT  7455.0 104007.5 8465.0 104072.5 ;
      RECT  7522.5 106567.5 7587.5 106762.5 ;
      RECT  7522.5 105727.5 7587.5 105352.5 ;
      RECT  7902.5 105727.5 7967.5 105352.5 ;
      RECT  8262.5 105570.0 8327.5 105385.0 ;
      RECT  8262.5 106730.0 8327.5 106545.0 ;
      RECT  7522.5 105727.5 7587.5 105592.5 ;
      RECT  7712.5 105727.5 7777.5 105592.5 ;
      RECT  7712.5 105727.5 7777.5 105592.5 ;
      RECT  7522.5 105727.5 7587.5 105592.5 ;
      RECT  7712.5 105727.5 7777.5 105592.5 ;
      RECT  7902.5 105727.5 7967.5 105592.5 ;
      RECT  7902.5 105727.5 7967.5 105592.5 ;
      RECT  7712.5 105727.5 7777.5 105592.5 ;
      RECT  7902.5 105727.5 7967.5 105592.5 ;
      RECT  8092.5 105727.5 8157.5 105592.5 ;
      RECT  8092.5 105727.5 8157.5 105592.5 ;
      RECT  7902.5 105727.5 7967.5 105592.5 ;
      RECT  7522.5 106567.5 7587.5 106432.5 ;
      RECT  7712.5 106567.5 7777.5 106432.5 ;
      RECT  7712.5 106567.5 7777.5 106432.5 ;
      RECT  7522.5 106567.5 7587.5 106432.5 ;
      RECT  7712.5 106567.5 7777.5 106432.5 ;
      RECT  7902.5 106567.5 7967.5 106432.5 ;
      RECT  7902.5 106567.5 7967.5 106432.5 ;
      RECT  7712.5 106567.5 7777.5 106432.5 ;
      RECT  7902.5 106567.5 7967.5 106432.5 ;
      RECT  8092.5 106567.5 8157.5 106432.5 ;
      RECT  8092.5 106567.5 8157.5 106432.5 ;
      RECT  7902.5 106567.5 7967.5 106432.5 ;
      RECT  8262.5 105637.5 8327.5 105502.5 ;
      RECT  8262.5 106612.5 8327.5 106477.5 ;
      RECT  8097.5 106355.0 7962.5 106290.0 ;
      RECT  7907.5 106215.0 7772.5 106150.0 ;
      RECT  7717.5 106075.0 7582.5 106010.0 ;
      RECT  7712.5 105727.5 7777.5 105592.5 ;
      RECT  8092.5 105727.5 8157.5 105592.5 ;
      RECT  8092.5 106567.5 8157.5 106432.5 ;
      RECT  8092.5 106110.0 8157.5 105975.0 ;
      RECT  7582.5 106075.0 7717.5 106010.0 ;
      RECT  7772.5 106215.0 7907.5 106150.0 ;
      RECT  7962.5 106355.0 8097.5 106290.0 ;
      RECT  8092.5 106110.0 8157.5 105975.0 ;
      RECT  7455.0 105417.5 8465.0 105352.5 ;
      RECT  7455.0 106762.5 8465.0 106697.5 ;
      RECT  7522.5 106892.5 7587.5 106697.5 ;
      RECT  7522.5 107732.5 7587.5 108107.5 ;
      RECT  7902.5 107732.5 7967.5 108107.5 ;
      RECT  8262.5 107890.0 8327.5 108075.0 ;
      RECT  8262.5 106730.0 8327.5 106915.0 ;
      RECT  7522.5 107732.5 7587.5 107867.5 ;
      RECT  7712.5 107732.5 7777.5 107867.5 ;
      RECT  7712.5 107732.5 7777.5 107867.5 ;
      RECT  7522.5 107732.5 7587.5 107867.5 ;
      RECT  7712.5 107732.5 7777.5 107867.5 ;
      RECT  7902.5 107732.5 7967.5 107867.5 ;
      RECT  7902.5 107732.5 7967.5 107867.5 ;
      RECT  7712.5 107732.5 7777.5 107867.5 ;
      RECT  7902.5 107732.5 7967.5 107867.5 ;
      RECT  8092.5 107732.5 8157.5 107867.5 ;
      RECT  8092.5 107732.5 8157.5 107867.5 ;
      RECT  7902.5 107732.5 7967.5 107867.5 ;
      RECT  7522.5 106892.5 7587.5 107027.5 ;
      RECT  7712.5 106892.5 7777.5 107027.5 ;
      RECT  7712.5 106892.5 7777.5 107027.5 ;
      RECT  7522.5 106892.5 7587.5 107027.5 ;
      RECT  7712.5 106892.5 7777.5 107027.5 ;
      RECT  7902.5 106892.5 7967.5 107027.5 ;
      RECT  7902.5 106892.5 7967.5 107027.5 ;
      RECT  7712.5 106892.5 7777.5 107027.5 ;
      RECT  7902.5 106892.5 7967.5 107027.5 ;
      RECT  8092.5 106892.5 8157.5 107027.5 ;
      RECT  8092.5 106892.5 8157.5 107027.5 ;
      RECT  7902.5 106892.5 7967.5 107027.5 ;
      RECT  8262.5 107822.5 8327.5 107957.5 ;
      RECT  8262.5 106847.5 8327.5 106982.5 ;
      RECT  8097.5 107105.0 7962.5 107170.0 ;
      RECT  7907.5 107245.0 7772.5 107310.0 ;
      RECT  7717.5 107385.0 7582.5 107450.0 ;
      RECT  7712.5 107732.5 7777.5 107867.5 ;
      RECT  8092.5 107732.5 8157.5 107867.5 ;
      RECT  8092.5 106892.5 8157.5 107027.5 ;
      RECT  8092.5 107350.0 8157.5 107485.0 ;
      RECT  7582.5 107385.0 7717.5 107450.0 ;
      RECT  7772.5 107245.0 7907.5 107310.0 ;
      RECT  7962.5 107105.0 8097.5 107170.0 ;
      RECT  8092.5 107350.0 8157.5 107485.0 ;
      RECT  7455.0 108042.5 8465.0 108107.5 ;
      RECT  7455.0 106697.5 8465.0 106762.5 ;
      RECT  7522.5 109257.5 7587.5 109452.5 ;
      RECT  7522.5 108417.5 7587.5 108042.5 ;
      RECT  7902.5 108417.5 7967.5 108042.5 ;
      RECT  8262.5 108260.0 8327.5 108075.0 ;
      RECT  8262.5 109420.0 8327.5 109235.0 ;
      RECT  7522.5 108417.5 7587.5 108282.5 ;
      RECT  7712.5 108417.5 7777.5 108282.5 ;
      RECT  7712.5 108417.5 7777.5 108282.5 ;
      RECT  7522.5 108417.5 7587.5 108282.5 ;
      RECT  7712.5 108417.5 7777.5 108282.5 ;
      RECT  7902.5 108417.5 7967.5 108282.5 ;
      RECT  7902.5 108417.5 7967.5 108282.5 ;
      RECT  7712.5 108417.5 7777.5 108282.5 ;
      RECT  7902.5 108417.5 7967.5 108282.5 ;
      RECT  8092.5 108417.5 8157.5 108282.5 ;
      RECT  8092.5 108417.5 8157.5 108282.5 ;
      RECT  7902.5 108417.5 7967.5 108282.5 ;
      RECT  7522.5 109257.5 7587.5 109122.5 ;
      RECT  7712.5 109257.5 7777.5 109122.5 ;
      RECT  7712.5 109257.5 7777.5 109122.5 ;
      RECT  7522.5 109257.5 7587.5 109122.5 ;
      RECT  7712.5 109257.5 7777.5 109122.5 ;
      RECT  7902.5 109257.5 7967.5 109122.5 ;
      RECT  7902.5 109257.5 7967.5 109122.5 ;
      RECT  7712.5 109257.5 7777.5 109122.5 ;
      RECT  7902.5 109257.5 7967.5 109122.5 ;
      RECT  8092.5 109257.5 8157.5 109122.5 ;
      RECT  8092.5 109257.5 8157.5 109122.5 ;
      RECT  7902.5 109257.5 7967.5 109122.5 ;
      RECT  8262.5 108327.5 8327.5 108192.5 ;
      RECT  8262.5 109302.5 8327.5 109167.5 ;
      RECT  8097.5 109045.0 7962.5 108980.0 ;
      RECT  7907.5 108905.0 7772.5 108840.0 ;
      RECT  7717.5 108765.0 7582.5 108700.0 ;
      RECT  7712.5 108417.5 7777.5 108282.5 ;
      RECT  8092.5 108417.5 8157.5 108282.5 ;
      RECT  8092.5 109257.5 8157.5 109122.5 ;
      RECT  8092.5 108800.0 8157.5 108665.0 ;
      RECT  7582.5 108765.0 7717.5 108700.0 ;
      RECT  7772.5 108905.0 7907.5 108840.0 ;
      RECT  7962.5 109045.0 8097.5 108980.0 ;
      RECT  8092.5 108800.0 8157.5 108665.0 ;
      RECT  7455.0 108107.5 8465.0 108042.5 ;
      RECT  7455.0 109452.5 8465.0 109387.5 ;
      RECT  7522.5 109582.5 7587.5 109387.5 ;
      RECT  7522.5 110422.5 7587.5 110797.5 ;
      RECT  7902.5 110422.5 7967.5 110797.5 ;
      RECT  8262.5 110580.0 8327.5 110765.0 ;
      RECT  8262.5 109420.0 8327.5 109605.0 ;
      RECT  7522.5 110422.5 7587.5 110557.5 ;
      RECT  7712.5 110422.5 7777.5 110557.5 ;
      RECT  7712.5 110422.5 7777.5 110557.5 ;
      RECT  7522.5 110422.5 7587.5 110557.5 ;
      RECT  7712.5 110422.5 7777.5 110557.5 ;
      RECT  7902.5 110422.5 7967.5 110557.5 ;
      RECT  7902.5 110422.5 7967.5 110557.5 ;
      RECT  7712.5 110422.5 7777.5 110557.5 ;
      RECT  7902.5 110422.5 7967.5 110557.5 ;
      RECT  8092.5 110422.5 8157.5 110557.5 ;
      RECT  8092.5 110422.5 8157.5 110557.5 ;
      RECT  7902.5 110422.5 7967.5 110557.5 ;
      RECT  7522.5 109582.5 7587.5 109717.5 ;
      RECT  7712.5 109582.5 7777.5 109717.5 ;
      RECT  7712.5 109582.5 7777.5 109717.5 ;
      RECT  7522.5 109582.5 7587.5 109717.5 ;
      RECT  7712.5 109582.5 7777.5 109717.5 ;
      RECT  7902.5 109582.5 7967.5 109717.5 ;
      RECT  7902.5 109582.5 7967.5 109717.5 ;
      RECT  7712.5 109582.5 7777.5 109717.5 ;
      RECT  7902.5 109582.5 7967.5 109717.5 ;
      RECT  8092.5 109582.5 8157.5 109717.5 ;
      RECT  8092.5 109582.5 8157.5 109717.5 ;
      RECT  7902.5 109582.5 7967.5 109717.5 ;
      RECT  8262.5 110512.5 8327.5 110647.5 ;
      RECT  8262.5 109537.5 8327.5 109672.5 ;
      RECT  8097.5 109795.0 7962.5 109860.0 ;
      RECT  7907.5 109935.0 7772.5 110000.0 ;
      RECT  7717.5 110075.0 7582.5 110140.0 ;
      RECT  7712.5 110422.5 7777.5 110557.5 ;
      RECT  8092.5 110422.5 8157.5 110557.5 ;
      RECT  8092.5 109582.5 8157.5 109717.5 ;
      RECT  8092.5 110040.0 8157.5 110175.0 ;
      RECT  7582.5 110075.0 7717.5 110140.0 ;
      RECT  7772.5 109935.0 7907.5 110000.0 ;
      RECT  7962.5 109795.0 8097.5 109860.0 ;
      RECT  8092.5 110040.0 8157.5 110175.0 ;
      RECT  7455.0 110732.5 8465.0 110797.5 ;
      RECT  7455.0 109387.5 8465.0 109452.5 ;
      RECT  7522.5 111947.5 7587.5 112142.5 ;
      RECT  7522.5 111107.5 7587.5 110732.5 ;
      RECT  7902.5 111107.5 7967.5 110732.5 ;
      RECT  8262.5 110950.0 8327.5 110765.0 ;
      RECT  8262.5 112110.0 8327.5 111925.0 ;
      RECT  7522.5 111107.5 7587.5 110972.5 ;
      RECT  7712.5 111107.5 7777.5 110972.5 ;
      RECT  7712.5 111107.5 7777.5 110972.5 ;
      RECT  7522.5 111107.5 7587.5 110972.5 ;
      RECT  7712.5 111107.5 7777.5 110972.5 ;
      RECT  7902.5 111107.5 7967.5 110972.5 ;
      RECT  7902.5 111107.5 7967.5 110972.5 ;
      RECT  7712.5 111107.5 7777.5 110972.5 ;
      RECT  7902.5 111107.5 7967.5 110972.5 ;
      RECT  8092.5 111107.5 8157.5 110972.5 ;
      RECT  8092.5 111107.5 8157.5 110972.5 ;
      RECT  7902.5 111107.5 7967.5 110972.5 ;
      RECT  7522.5 111947.5 7587.5 111812.5 ;
      RECT  7712.5 111947.5 7777.5 111812.5 ;
      RECT  7712.5 111947.5 7777.5 111812.5 ;
      RECT  7522.5 111947.5 7587.5 111812.5 ;
      RECT  7712.5 111947.5 7777.5 111812.5 ;
      RECT  7902.5 111947.5 7967.5 111812.5 ;
      RECT  7902.5 111947.5 7967.5 111812.5 ;
      RECT  7712.5 111947.5 7777.5 111812.5 ;
      RECT  7902.5 111947.5 7967.5 111812.5 ;
      RECT  8092.5 111947.5 8157.5 111812.5 ;
      RECT  8092.5 111947.5 8157.5 111812.5 ;
      RECT  7902.5 111947.5 7967.5 111812.5 ;
      RECT  8262.5 111017.5 8327.5 110882.5 ;
      RECT  8262.5 111992.5 8327.5 111857.5 ;
      RECT  8097.5 111735.0 7962.5 111670.0 ;
      RECT  7907.5 111595.0 7772.5 111530.0 ;
      RECT  7717.5 111455.0 7582.5 111390.0 ;
      RECT  7712.5 111107.5 7777.5 110972.5 ;
      RECT  8092.5 111107.5 8157.5 110972.5 ;
      RECT  8092.5 111947.5 8157.5 111812.5 ;
      RECT  8092.5 111490.0 8157.5 111355.0 ;
      RECT  7582.5 111455.0 7717.5 111390.0 ;
      RECT  7772.5 111595.0 7907.5 111530.0 ;
      RECT  7962.5 111735.0 8097.5 111670.0 ;
      RECT  8092.5 111490.0 8157.5 111355.0 ;
      RECT  7455.0 110797.5 8465.0 110732.5 ;
      RECT  7455.0 112142.5 8465.0 112077.5 ;
      RECT  7522.5 112272.5 7587.5 112077.5 ;
      RECT  7522.5 113112.5 7587.5 113487.5 ;
      RECT  7902.5 113112.5 7967.5 113487.5 ;
      RECT  8262.5 113270.0 8327.5 113455.0 ;
      RECT  8262.5 112110.0 8327.5 112295.0 ;
      RECT  7522.5 113112.5 7587.5 113247.5 ;
      RECT  7712.5 113112.5 7777.5 113247.5 ;
      RECT  7712.5 113112.5 7777.5 113247.5 ;
      RECT  7522.5 113112.5 7587.5 113247.5 ;
      RECT  7712.5 113112.5 7777.5 113247.5 ;
      RECT  7902.5 113112.5 7967.5 113247.5 ;
      RECT  7902.5 113112.5 7967.5 113247.5 ;
      RECT  7712.5 113112.5 7777.5 113247.5 ;
      RECT  7902.5 113112.5 7967.5 113247.5 ;
      RECT  8092.5 113112.5 8157.5 113247.5 ;
      RECT  8092.5 113112.5 8157.5 113247.5 ;
      RECT  7902.5 113112.5 7967.5 113247.5 ;
      RECT  7522.5 112272.5 7587.5 112407.5 ;
      RECT  7712.5 112272.5 7777.5 112407.5 ;
      RECT  7712.5 112272.5 7777.5 112407.5 ;
      RECT  7522.5 112272.5 7587.5 112407.5 ;
      RECT  7712.5 112272.5 7777.5 112407.5 ;
      RECT  7902.5 112272.5 7967.5 112407.5 ;
      RECT  7902.5 112272.5 7967.5 112407.5 ;
      RECT  7712.5 112272.5 7777.5 112407.5 ;
      RECT  7902.5 112272.5 7967.5 112407.5 ;
      RECT  8092.5 112272.5 8157.5 112407.5 ;
      RECT  8092.5 112272.5 8157.5 112407.5 ;
      RECT  7902.5 112272.5 7967.5 112407.5 ;
      RECT  8262.5 113202.5 8327.5 113337.5 ;
      RECT  8262.5 112227.5 8327.5 112362.5 ;
      RECT  8097.5 112485.0 7962.5 112550.0 ;
      RECT  7907.5 112625.0 7772.5 112690.0 ;
      RECT  7717.5 112765.0 7582.5 112830.0 ;
      RECT  7712.5 113112.5 7777.5 113247.5 ;
      RECT  8092.5 113112.5 8157.5 113247.5 ;
      RECT  8092.5 112272.5 8157.5 112407.5 ;
      RECT  8092.5 112730.0 8157.5 112865.0 ;
      RECT  7582.5 112765.0 7717.5 112830.0 ;
      RECT  7772.5 112625.0 7907.5 112690.0 ;
      RECT  7962.5 112485.0 8097.5 112550.0 ;
      RECT  8092.5 112730.0 8157.5 112865.0 ;
      RECT  7455.0 113422.5 8465.0 113487.5 ;
      RECT  7455.0 112077.5 8465.0 112142.5 ;
      RECT  7522.5 114637.5 7587.5 114832.5 ;
      RECT  7522.5 113797.5 7587.5 113422.5 ;
      RECT  7902.5 113797.5 7967.5 113422.5 ;
      RECT  8262.5 113640.0 8327.5 113455.0 ;
      RECT  8262.5 114800.0 8327.5 114615.0 ;
      RECT  7522.5 113797.5 7587.5 113662.5 ;
      RECT  7712.5 113797.5 7777.5 113662.5 ;
      RECT  7712.5 113797.5 7777.5 113662.5 ;
      RECT  7522.5 113797.5 7587.5 113662.5 ;
      RECT  7712.5 113797.5 7777.5 113662.5 ;
      RECT  7902.5 113797.5 7967.5 113662.5 ;
      RECT  7902.5 113797.5 7967.5 113662.5 ;
      RECT  7712.5 113797.5 7777.5 113662.5 ;
      RECT  7902.5 113797.5 7967.5 113662.5 ;
      RECT  8092.5 113797.5 8157.5 113662.5 ;
      RECT  8092.5 113797.5 8157.5 113662.5 ;
      RECT  7902.5 113797.5 7967.5 113662.5 ;
      RECT  7522.5 114637.5 7587.5 114502.5 ;
      RECT  7712.5 114637.5 7777.5 114502.5 ;
      RECT  7712.5 114637.5 7777.5 114502.5 ;
      RECT  7522.5 114637.5 7587.5 114502.5 ;
      RECT  7712.5 114637.5 7777.5 114502.5 ;
      RECT  7902.5 114637.5 7967.5 114502.5 ;
      RECT  7902.5 114637.5 7967.5 114502.5 ;
      RECT  7712.5 114637.5 7777.5 114502.5 ;
      RECT  7902.5 114637.5 7967.5 114502.5 ;
      RECT  8092.5 114637.5 8157.5 114502.5 ;
      RECT  8092.5 114637.5 8157.5 114502.5 ;
      RECT  7902.5 114637.5 7967.5 114502.5 ;
      RECT  8262.5 113707.5 8327.5 113572.5 ;
      RECT  8262.5 114682.5 8327.5 114547.5 ;
      RECT  8097.5 114425.0 7962.5 114360.0 ;
      RECT  7907.5 114285.0 7772.5 114220.0 ;
      RECT  7717.5 114145.0 7582.5 114080.0 ;
      RECT  7712.5 113797.5 7777.5 113662.5 ;
      RECT  8092.5 113797.5 8157.5 113662.5 ;
      RECT  8092.5 114637.5 8157.5 114502.5 ;
      RECT  8092.5 114180.0 8157.5 114045.0 ;
      RECT  7582.5 114145.0 7717.5 114080.0 ;
      RECT  7772.5 114285.0 7907.5 114220.0 ;
      RECT  7962.5 114425.0 8097.5 114360.0 ;
      RECT  8092.5 114180.0 8157.5 114045.0 ;
      RECT  7455.0 113487.5 8465.0 113422.5 ;
      RECT  7455.0 114832.5 8465.0 114767.5 ;
      RECT  7522.5 114962.5 7587.5 114767.5 ;
      RECT  7522.5 115802.5 7587.5 116177.5 ;
      RECT  7902.5 115802.5 7967.5 116177.5 ;
      RECT  8262.5 115960.0 8327.5 116145.0 ;
      RECT  8262.5 114800.0 8327.5 114985.0 ;
      RECT  7522.5 115802.5 7587.5 115937.5 ;
      RECT  7712.5 115802.5 7777.5 115937.5 ;
      RECT  7712.5 115802.5 7777.5 115937.5 ;
      RECT  7522.5 115802.5 7587.5 115937.5 ;
      RECT  7712.5 115802.5 7777.5 115937.5 ;
      RECT  7902.5 115802.5 7967.5 115937.5 ;
      RECT  7902.5 115802.5 7967.5 115937.5 ;
      RECT  7712.5 115802.5 7777.5 115937.5 ;
      RECT  7902.5 115802.5 7967.5 115937.5 ;
      RECT  8092.5 115802.5 8157.5 115937.5 ;
      RECT  8092.5 115802.5 8157.5 115937.5 ;
      RECT  7902.5 115802.5 7967.5 115937.5 ;
      RECT  7522.5 114962.5 7587.5 115097.5 ;
      RECT  7712.5 114962.5 7777.5 115097.5 ;
      RECT  7712.5 114962.5 7777.5 115097.5 ;
      RECT  7522.5 114962.5 7587.5 115097.5 ;
      RECT  7712.5 114962.5 7777.5 115097.5 ;
      RECT  7902.5 114962.5 7967.5 115097.5 ;
      RECT  7902.5 114962.5 7967.5 115097.5 ;
      RECT  7712.5 114962.5 7777.5 115097.5 ;
      RECT  7902.5 114962.5 7967.5 115097.5 ;
      RECT  8092.5 114962.5 8157.5 115097.5 ;
      RECT  8092.5 114962.5 8157.5 115097.5 ;
      RECT  7902.5 114962.5 7967.5 115097.5 ;
      RECT  8262.5 115892.5 8327.5 116027.5 ;
      RECT  8262.5 114917.5 8327.5 115052.5 ;
      RECT  8097.5 115175.0 7962.5 115240.0 ;
      RECT  7907.5 115315.0 7772.5 115380.0 ;
      RECT  7717.5 115455.0 7582.5 115520.0 ;
      RECT  7712.5 115802.5 7777.5 115937.5 ;
      RECT  8092.5 115802.5 8157.5 115937.5 ;
      RECT  8092.5 114962.5 8157.5 115097.5 ;
      RECT  8092.5 115420.0 8157.5 115555.0 ;
      RECT  7582.5 115455.0 7717.5 115520.0 ;
      RECT  7772.5 115315.0 7907.5 115380.0 ;
      RECT  7962.5 115175.0 8097.5 115240.0 ;
      RECT  8092.5 115420.0 8157.5 115555.0 ;
      RECT  7455.0 116112.5 8465.0 116177.5 ;
      RECT  7455.0 114767.5 8465.0 114832.5 ;
      RECT  7522.5 117327.5 7587.5 117522.5 ;
      RECT  7522.5 116487.5 7587.5 116112.5 ;
      RECT  7902.5 116487.5 7967.5 116112.5 ;
      RECT  8262.5 116330.0 8327.5 116145.0 ;
      RECT  8262.5 117490.0 8327.5 117305.0 ;
      RECT  7522.5 116487.5 7587.5 116352.5 ;
      RECT  7712.5 116487.5 7777.5 116352.5 ;
      RECT  7712.5 116487.5 7777.5 116352.5 ;
      RECT  7522.5 116487.5 7587.5 116352.5 ;
      RECT  7712.5 116487.5 7777.5 116352.5 ;
      RECT  7902.5 116487.5 7967.5 116352.5 ;
      RECT  7902.5 116487.5 7967.5 116352.5 ;
      RECT  7712.5 116487.5 7777.5 116352.5 ;
      RECT  7902.5 116487.5 7967.5 116352.5 ;
      RECT  8092.5 116487.5 8157.5 116352.5 ;
      RECT  8092.5 116487.5 8157.5 116352.5 ;
      RECT  7902.5 116487.5 7967.5 116352.5 ;
      RECT  7522.5 117327.5 7587.5 117192.5 ;
      RECT  7712.5 117327.5 7777.5 117192.5 ;
      RECT  7712.5 117327.5 7777.5 117192.5 ;
      RECT  7522.5 117327.5 7587.5 117192.5 ;
      RECT  7712.5 117327.5 7777.5 117192.5 ;
      RECT  7902.5 117327.5 7967.5 117192.5 ;
      RECT  7902.5 117327.5 7967.5 117192.5 ;
      RECT  7712.5 117327.5 7777.5 117192.5 ;
      RECT  7902.5 117327.5 7967.5 117192.5 ;
      RECT  8092.5 117327.5 8157.5 117192.5 ;
      RECT  8092.5 117327.5 8157.5 117192.5 ;
      RECT  7902.5 117327.5 7967.5 117192.5 ;
      RECT  8262.5 116397.5 8327.5 116262.5 ;
      RECT  8262.5 117372.5 8327.5 117237.5 ;
      RECT  8097.5 117115.0 7962.5 117050.0 ;
      RECT  7907.5 116975.0 7772.5 116910.0 ;
      RECT  7717.5 116835.0 7582.5 116770.0 ;
      RECT  7712.5 116487.5 7777.5 116352.5 ;
      RECT  8092.5 116487.5 8157.5 116352.5 ;
      RECT  8092.5 117327.5 8157.5 117192.5 ;
      RECT  8092.5 116870.0 8157.5 116735.0 ;
      RECT  7582.5 116835.0 7717.5 116770.0 ;
      RECT  7772.5 116975.0 7907.5 116910.0 ;
      RECT  7962.5 117115.0 8097.5 117050.0 ;
      RECT  8092.5 116870.0 8157.5 116735.0 ;
      RECT  7455.0 116177.5 8465.0 116112.5 ;
      RECT  7455.0 117522.5 8465.0 117457.5 ;
      RECT  7522.5 117652.5 7587.5 117457.5 ;
      RECT  7522.5 118492.5 7587.5 118867.5 ;
      RECT  7902.5 118492.5 7967.5 118867.5 ;
      RECT  8262.5 118650.0 8327.5 118835.0 ;
      RECT  8262.5 117490.0 8327.5 117675.0 ;
      RECT  7522.5 118492.5 7587.5 118627.5 ;
      RECT  7712.5 118492.5 7777.5 118627.5 ;
      RECT  7712.5 118492.5 7777.5 118627.5 ;
      RECT  7522.5 118492.5 7587.5 118627.5 ;
      RECT  7712.5 118492.5 7777.5 118627.5 ;
      RECT  7902.5 118492.5 7967.5 118627.5 ;
      RECT  7902.5 118492.5 7967.5 118627.5 ;
      RECT  7712.5 118492.5 7777.5 118627.5 ;
      RECT  7902.5 118492.5 7967.5 118627.5 ;
      RECT  8092.5 118492.5 8157.5 118627.5 ;
      RECT  8092.5 118492.5 8157.5 118627.5 ;
      RECT  7902.5 118492.5 7967.5 118627.5 ;
      RECT  7522.5 117652.5 7587.5 117787.5 ;
      RECT  7712.5 117652.5 7777.5 117787.5 ;
      RECT  7712.5 117652.5 7777.5 117787.5 ;
      RECT  7522.5 117652.5 7587.5 117787.5 ;
      RECT  7712.5 117652.5 7777.5 117787.5 ;
      RECT  7902.5 117652.5 7967.5 117787.5 ;
      RECT  7902.5 117652.5 7967.5 117787.5 ;
      RECT  7712.5 117652.5 7777.5 117787.5 ;
      RECT  7902.5 117652.5 7967.5 117787.5 ;
      RECT  8092.5 117652.5 8157.5 117787.5 ;
      RECT  8092.5 117652.5 8157.5 117787.5 ;
      RECT  7902.5 117652.5 7967.5 117787.5 ;
      RECT  8262.5 118582.5 8327.5 118717.5 ;
      RECT  8262.5 117607.5 8327.5 117742.5 ;
      RECT  8097.5 117865.0 7962.5 117930.0 ;
      RECT  7907.5 118005.0 7772.5 118070.0 ;
      RECT  7717.5 118145.0 7582.5 118210.0 ;
      RECT  7712.5 118492.5 7777.5 118627.5 ;
      RECT  8092.5 118492.5 8157.5 118627.5 ;
      RECT  8092.5 117652.5 8157.5 117787.5 ;
      RECT  8092.5 118110.0 8157.5 118245.0 ;
      RECT  7582.5 118145.0 7717.5 118210.0 ;
      RECT  7772.5 118005.0 7907.5 118070.0 ;
      RECT  7962.5 117865.0 8097.5 117930.0 ;
      RECT  8092.5 118110.0 8157.5 118245.0 ;
      RECT  7455.0 118802.5 8465.0 118867.5 ;
      RECT  7455.0 117457.5 8465.0 117522.5 ;
      RECT  7522.5 120017.5 7587.5 120212.5 ;
      RECT  7522.5 119177.5 7587.5 118802.5 ;
      RECT  7902.5 119177.5 7967.5 118802.5 ;
      RECT  8262.5 119020.0 8327.5 118835.0 ;
      RECT  8262.5 120180.0 8327.5 119995.0 ;
      RECT  7522.5 119177.5 7587.5 119042.5 ;
      RECT  7712.5 119177.5 7777.5 119042.5 ;
      RECT  7712.5 119177.5 7777.5 119042.5 ;
      RECT  7522.5 119177.5 7587.5 119042.5 ;
      RECT  7712.5 119177.5 7777.5 119042.5 ;
      RECT  7902.5 119177.5 7967.5 119042.5 ;
      RECT  7902.5 119177.5 7967.5 119042.5 ;
      RECT  7712.5 119177.5 7777.5 119042.5 ;
      RECT  7902.5 119177.5 7967.5 119042.5 ;
      RECT  8092.5 119177.5 8157.5 119042.5 ;
      RECT  8092.5 119177.5 8157.5 119042.5 ;
      RECT  7902.5 119177.5 7967.5 119042.5 ;
      RECT  7522.5 120017.5 7587.5 119882.5 ;
      RECT  7712.5 120017.5 7777.5 119882.5 ;
      RECT  7712.5 120017.5 7777.5 119882.5 ;
      RECT  7522.5 120017.5 7587.5 119882.5 ;
      RECT  7712.5 120017.5 7777.5 119882.5 ;
      RECT  7902.5 120017.5 7967.5 119882.5 ;
      RECT  7902.5 120017.5 7967.5 119882.5 ;
      RECT  7712.5 120017.5 7777.5 119882.5 ;
      RECT  7902.5 120017.5 7967.5 119882.5 ;
      RECT  8092.5 120017.5 8157.5 119882.5 ;
      RECT  8092.5 120017.5 8157.5 119882.5 ;
      RECT  7902.5 120017.5 7967.5 119882.5 ;
      RECT  8262.5 119087.5 8327.5 118952.5 ;
      RECT  8262.5 120062.5 8327.5 119927.5 ;
      RECT  8097.5 119805.0 7962.5 119740.0 ;
      RECT  7907.5 119665.0 7772.5 119600.0 ;
      RECT  7717.5 119525.0 7582.5 119460.0 ;
      RECT  7712.5 119177.5 7777.5 119042.5 ;
      RECT  8092.5 119177.5 8157.5 119042.5 ;
      RECT  8092.5 120017.5 8157.5 119882.5 ;
      RECT  8092.5 119560.0 8157.5 119425.0 ;
      RECT  7582.5 119525.0 7717.5 119460.0 ;
      RECT  7772.5 119665.0 7907.5 119600.0 ;
      RECT  7962.5 119805.0 8097.5 119740.0 ;
      RECT  8092.5 119560.0 8157.5 119425.0 ;
      RECT  7455.0 118867.5 8465.0 118802.5 ;
      RECT  7455.0 120212.5 8465.0 120147.5 ;
      RECT  7522.5 120342.5 7587.5 120147.5 ;
      RECT  7522.5 121182.5 7587.5 121557.5 ;
      RECT  7902.5 121182.5 7967.5 121557.5 ;
      RECT  8262.5 121340.0 8327.5 121525.0 ;
      RECT  8262.5 120180.0 8327.5 120365.0 ;
      RECT  7522.5 121182.5 7587.5 121317.5 ;
      RECT  7712.5 121182.5 7777.5 121317.5 ;
      RECT  7712.5 121182.5 7777.5 121317.5 ;
      RECT  7522.5 121182.5 7587.5 121317.5 ;
      RECT  7712.5 121182.5 7777.5 121317.5 ;
      RECT  7902.5 121182.5 7967.5 121317.5 ;
      RECT  7902.5 121182.5 7967.5 121317.5 ;
      RECT  7712.5 121182.5 7777.5 121317.5 ;
      RECT  7902.5 121182.5 7967.5 121317.5 ;
      RECT  8092.5 121182.5 8157.5 121317.5 ;
      RECT  8092.5 121182.5 8157.5 121317.5 ;
      RECT  7902.5 121182.5 7967.5 121317.5 ;
      RECT  7522.5 120342.5 7587.5 120477.5 ;
      RECT  7712.5 120342.5 7777.5 120477.5 ;
      RECT  7712.5 120342.5 7777.5 120477.5 ;
      RECT  7522.5 120342.5 7587.5 120477.5 ;
      RECT  7712.5 120342.5 7777.5 120477.5 ;
      RECT  7902.5 120342.5 7967.5 120477.5 ;
      RECT  7902.5 120342.5 7967.5 120477.5 ;
      RECT  7712.5 120342.5 7777.5 120477.5 ;
      RECT  7902.5 120342.5 7967.5 120477.5 ;
      RECT  8092.5 120342.5 8157.5 120477.5 ;
      RECT  8092.5 120342.5 8157.5 120477.5 ;
      RECT  7902.5 120342.5 7967.5 120477.5 ;
      RECT  8262.5 121272.5 8327.5 121407.5 ;
      RECT  8262.5 120297.5 8327.5 120432.5 ;
      RECT  8097.5 120555.0 7962.5 120620.0 ;
      RECT  7907.5 120695.0 7772.5 120760.0 ;
      RECT  7717.5 120835.0 7582.5 120900.0 ;
      RECT  7712.5 121182.5 7777.5 121317.5 ;
      RECT  8092.5 121182.5 8157.5 121317.5 ;
      RECT  8092.5 120342.5 8157.5 120477.5 ;
      RECT  8092.5 120800.0 8157.5 120935.0 ;
      RECT  7582.5 120835.0 7717.5 120900.0 ;
      RECT  7772.5 120695.0 7907.5 120760.0 ;
      RECT  7962.5 120555.0 8097.5 120620.0 ;
      RECT  8092.5 120800.0 8157.5 120935.0 ;
      RECT  7455.0 121492.5 8465.0 121557.5 ;
      RECT  7455.0 120147.5 8465.0 120212.5 ;
      RECT  7522.5 122707.5 7587.5 122902.5 ;
      RECT  7522.5 121867.5 7587.5 121492.5 ;
      RECT  7902.5 121867.5 7967.5 121492.5 ;
      RECT  8262.5 121710.0 8327.5 121525.0 ;
      RECT  8262.5 122870.0 8327.5 122685.0 ;
      RECT  7522.5 121867.5 7587.5 121732.5 ;
      RECT  7712.5 121867.5 7777.5 121732.5 ;
      RECT  7712.5 121867.5 7777.5 121732.5 ;
      RECT  7522.5 121867.5 7587.5 121732.5 ;
      RECT  7712.5 121867.5 7777.5 121732.5 ;
      RECT  7902.5 121867.5 7967.5 121732.5 ;
      RECT  7902.5 121867.5 7967.5 121732.5 ;
      RECT  7712.5 121867.5 7777.5 121732.5 ;
      RECT  7902.5 121867.5 7967.5 121732.5 ;
      RECT  8092.5 121867.5 8157.5 121732.5 ;
      RECT  8092.5 121867.5 8157.5 121732.5 ;
      RECT  7902.5 121867.5 7967.5 121732.5 ;
      RECT  7522.5 122707.5 7587.5 122572.5 ;
      RECT  7712.5 122707.5 7777.5 122572.5 ;
      RECT  7712.5 122707.5 7777.5 122572.5 ;
      RECT  7522.5 122707.5 7587.5 122572.5 ;
      RECT  7712.5 122707.5 7777.5 122572.5 ;
      RECT  7902.5 122707.5 7967.5 122572.5 ;
      RECT  7902.5 122707.5 7967.5 122572.5 ;
      RECT  7712.5 122707.5 7777.5 122572.5 ;
      RECT  7902.5 122707.5 7967.5 122572.5 ;
      RECT  8092.5 122707.5 8157.5 122572.5 ;
      RECT  8092.5 122707.5 8157.5 122572.5 ;
      RECT  7902.5 122707.5 7967.5 122572.5 ;
      RECT  8262.5 121777.5 8327.5 121642.5 ;
      RECT  8262.5 122752.5 8327.5 122617.5 ;
      RECT  8097.5 122495.0 7962.5 122430.0 ;
      RECT  7907.5 122355.0 7772.5 122290.0 ;
      RECT  7717.5 122215.0 7582.5 122150.0 ;
      RECT  7712.5 121867.5 7777.5 121732.5 ;
      RECT  8092.5 121867.5 8157.5 121732.5 ;
      RECT  8092.5 122707.5 8157.5 122572.5 ;
      RECT  8092.5 122250.0 8157.5 122115.0 ;
      RECT  7582.5 122215.0 7717.5 122150.0 ;
      RECT  7772.5 122355.0 7907.5 122290.0 ;
      RECT  7962.5 122495.0 8097.5 122430.0 ;
      RECT  8092.5 122250.0 8157.5 122115.0 ;
      RECT  7455.0 121557.5 8465.0 121492.5 ;
      RECT  7455.0 122902.5 8465.0 122837.5 ;
      RECT  7522.5 123032.5 7587.5 122837.5 ;
      RECT  7522.5 123872.5 7587.5 124247.5 ;
      RECT  7902.5 123872.5 7967.5 124247.5 ;
      RECT  8262.5 124030.0 8327.5 124215.0 ;
      RECT  8262.5 122870.0 8327.5 123055.0 ;
      RECT  7522.5 123872.5 7587.5 124007.5 ;
      RECT  7712.5 123872.5 7777.5 124007.5 ;
      RECT  7712.5 123872.5 7777.5 124007.5 ;
      RECT  7522.5 123872.5 7587.5 124007.5 ;
      RECT  7712.5 123872.5 7777.5 124007.5 ;
      RECT  7902.5 123872.5 7967.5 124007.5 ;
      RECT  7902.5 123872.5 7967.5 124007.5 ;
      RECT  7712.5 123872.5 7777.5 124007.5 ;
      RECT  7902.5 123872.5 7967.5 124007.5 ;
      RECT  8092.5 123872.5 8157.5 124007.5 ;
      RECT  8092.5 123872.5 8157.5 124007.5 ;
      RECT  7902.5 123872.5 7967.5 124007.5 ;
      RECT  7522.5 123032.5 7587.5 123167.5 ;
      RECT  7712.5 123032.5 7777.5 123167.5 ;
      RECT  7712.5 123032.5 7777.5 123167.5 ;
      RECT  7522.5 123032.5 7587.5 123167.5 ;
      RECT  7712.5 123032.5 7777.5 123167.5 ;
      RECT  7902.5 123032.5 7967.5 123167.5 ;
      RECT  7902.5 123032.5 7967.5 123167.5 ;
      RECT  7712.5 123032.5 7777.5 123167.5 ;
      RECT  7902.5 123032.5 7967.5 123167.5 ;
      RECT  8092.5 123032.5 8157.5 123167.5 ;
      RECT  8092.5 123032.5 8157.5 123167.5 ;
      RECT  7902.5 123032.5 7967.5 123167.5 ;
      RECT  8262.5 123962.5 8327.5 124097.5 ;
      RECT  8262.5 122987.5 8327.5 123122.5 ;
      RECT  8097.5 123245.0 7962.5 123310.0 ;
      RECT  7907.5 123385.0 7772.5 123450.0 ;
      RECT  7717.5 123525.0 7582.5 123590.0 ;
      RECT  7712.5 123872.5 7777.5 124007.5 ;
      RECT  8092.5 123872.5 8157.5 124007.5 ;
      RECT  8092.5 123032.5 8157.5 123167.5 ;
      RECT  8092.5 123490.0 8157.5 123625.0 ;
      RECT  7582.5 123525.0 7717.5 123590.0 ;
      RECT  7772.5 123385.0 7907.5 123450.0 ;
      RECT  7962.5 123245.0 8097.5 123310.0 ;
      RECT  8092.5 123490.0 8157.5 123625.0 ;
      RECT  7455.0 124182.5 8465.0 124247.5 ;
      RECT  7455.0 122837.5 8465.0 122902.5 ;
      RECT  7522.5 125397.5 7587.5 125592.5 ;
      RECT  7522.5 124557.5 7587.5 124182.5 ;
      RECT  7902.5 124557.5 7967.5 124182.5 ;
      RECT  8262.5 124400.0 8327.5 124215.0 ;
      RECT  8262.5 125560.0 8327.5 125375.0 ;
      RECT  7522.5 124557.5 7587.5 124422.5 ;
      RECT  7712.5 124557.5 7777.5 124422.5 ;
      RECT  7712.5 124557.5 7777.5 124422.5 ;
      RECT  7522.5 124557.5 7587.5 124422.5 ;
      RECT  7712.5 124557.5 7777.5 124422.5 ;
      RECT  7902.5 124557.5 7967.5 124422.5 ;
      RECT  7902.5 124557.5 7967.5 124422.5 ;
      RECT  7712.5 124557.5 7777.5 124422.5 ;
      RECT  7902.5 124557.5 7967.5 124422.5 ;
      RECT  8092.5 124557.5 8157.5 124422.5 ;
      RECT  8092.5 124557.5 8157.5 124422.5 ;
      RECT  7902.5 124557.5 7967.5 124422.5 ;
      RECT  7522.5 125397.5 7587.5 125262.5 ;
      RECT  7712.5 125397.5 7777.5 125262.5 ;
      RECT  7712.5 125397.5 7777.5 125262.5 ;
      RECT  7522.5 125397.5 7587.5 125262.5 ;
      RECT  7712.5 125397.5 7777.5 125262.5 ;
      RECT  7902.5 125397.5 7967.5 125262.5 ;
      RECT  7902.5 125397.5 7967.5 125262.5 ;
      RECT  7712.5 125397.5 7777.5 125262.5 ;
      RECT  7902.5 125397.5 7967.5 125262.5 ;
      RECT  8092.5 125397.5 8157.5 125262.5 ;
      RECT  8092.5 125397.5 8157.5 125262.5 ;
      RECT  7902.5 125397.5 7967.5 125262.5 ;
      RECT  8262.5 124467.5 8327.5 124332.5 ;
      RECT  8262.5 125442.5 8327.5 125307.5 ;
      RECT  8097.5 125185.0 7962.5 125120.0 ;
      RECT  7907.5 125045.0 7772.5 124980.0 ;
      RECT  7717.5 124905.0 7582.5 124840.0 ;
      RECT  7712.5 124557.5 7777.5 124422.5 ;
      RECT  8092.5 124557.5 8157.5 124422.5 ;
      RECT  8092.5 125397.5 8157.5 125262.5 ;
      RECT  8092.5 124940.0 8157.5 124805.0 ;
      RECT  7582.5 124905.0 7717.5 124840.0 ;
      RECT  7772.5 125045.0 7907.5 124980.0 ;
      RECT  7962.5 125185.0 8097.5 125120.0 ;
      RECT  8092.5 124940.0 8157.5 124805.0 ;
      RECT  7455.0 124247.5 8465.0 124182.5 ;
      RECT  7455.0 125592.5 8465.0 125527.5 ;
      RECT  7522.5 125722.5 7587.5 125527.5 ;
      RECT  7522.5 126562.5 7587.5 126937.5 ;
      RECT  7902.5 126562.5 7967.5 126937.5 ;
      RECT  8262.5 126720.0 8327.5 126905.0 ;
      RECT  8262.5 125560.0 8327.5 125745.0 ;
      RECT  7522.5 126562.5 7587.5 126697.5 ;
      RECT  7712.5 126562.5 7777.5 126697.5 ;
      RECT  7712.5 126562.5 7777.5 126697.5 ;
      RECT  7522.5 126562.5 7587.5 126697.5 ;
      RECT  7712.5 126562.5 7777.5 126697.5 ;
      RECT  7902.5 126562.5 7967.5 126697.5 ;
      RECT  7902.5 126562.5 7967.5 126697.5 ;
      RECT  7712.5 126562.5 7777.5 126697.5 ;
      RECT  7902.5 126562.5 7967.5 126697.5 ;
      RECT  8092.5 126562.5 8157.5 126697.5 ;
      RECT  8092.5 126562.5 8157.5 126697.5 ;
      RECT  7902.5 126562.5 7967.5 126697.5 ;
      RECT  7522.5 125722.5 7587.5 125857.5 ;
      RECT  7712.5 125722.5 7777.5 125857.5 ;
      RECT  7712.5 125722.5 7777.5 125857.5 ;
      RECT  7522.5 125722.5 7587.5 125857.5 ;
      RECT  7712.5 125722.5 7777.5 125857.5 ;
      RECT  7902.5 125722.5 7967.5 125857.5 ;
      RECT  7902.5 125722.5 7967.5 125857.5 ;
      RECT  7712.5 125722.5 7777.5 125857.5 ;
      RECT  7902.5 125722.5 7967.5 125857.5 ;
      RECT  8092.5 125722.5 8157.5 125857.5 ;
      RECT  8092.5 125722.5 8157.5 125857.5 ;
      RECT  7902.5 125722.5 7967.5 125857.5 ;
      RECT  8262.5 126652.5 8327.5 126787.5 ;
      RECT  8262.5 125677.5 8327.5 125812.5 ;
      RECT  8097.5 125935.0 7962.5 126000.0 ;
      RECT  7907.5 126075.0 7772.5 126140.0 ;
      RECT  7717.5 126215.0 7582.5 126280.0 ;
      RECT  7712.5 126562.5 7777.5 126697.5 ;
      RECT  8092.5 126562.5 8157.5 126697.5 ;
      RECT  8092.5 125722.5 8157.5 125857.5 ;
      RECT  8092.5 126180.0 8157.5 126315.0 ;
      RECT  7582.5 126215.0 7717.5 126280.0 ;
      RECT  7772.5 126075.0 7907.5 126140.0 ;
      RECT  7962.5 125935.0 8097.5 126000.0 ;
      RECT  8092.5 126180.0 8157.5 126315.0 ;
      RECT  7455.0 126872.5 8465.0 126937.5 ;
      RECT  7455.0 125527.5 8465.0 125592.5 ;
      RECT  7522.5 128087.5 7587.5 128282.5 ;
      RECT  7522.5 127247.5 7587.5 126872.5 ;
      RECT  7902.5 127247.5 7967.5 126872.5 ;
      RECT  8262.5 127090.0 8327.5 126905.0 ;
      RECT  8262.5 128250.0 8327.5 128065.0 ;
      RECT  7522.5 127247.5 7587.5 127112.5 ;
      RECT  7712.5 127247.5 7777.5 127112.5 ;
      RECT  7712.5 127247.5 7777.5 127112.5 ;
      RECT  7522.5 127247.5 7587.5 127112.5 ;
      RECT  7712.5 127247.5 7777.5 127112.5 ;
      RECT  7902.5 127247.5 7967.5 127112.5 ;
      RECT  7902.5 127247.5 7967.5 127112.5 ;
      RECT  7712.5 127247.5 7777.5 127112.5 ;
      RECT  7902.5 127247.5 7967.5 127112.5 ;
      RECT  8092.5 127247.5 8157.5 127112.5 ;
      RECT  8092.5 127247.5 8157.5 127112.5 ;
      RECT  7902.5 127247.5 7967.5 127112.5 ;
      RECT  7522.5 128087.5 7587.5 127952.5 ;
      RECT  7712.5 128087.5 7777.5 127952.5 ;
      RECT  7712.5 128087.5 7777.5 127952.5 ;
      RECT  7522.5 128087.5 7587.5 127952.5 ;
      RECT  7712.5 128087.5 7777.5 127952.5 ;
      RECT  7902.5 128087.5 7967.5 127952.5 ;
      RECT  7902.5 128087.5 7967.5 127952.5 ;
      RECT  7712.5 128087.5 7777.5 127952.5 ;
      RECT  7902.5 128087.5 7967.5 127952.5 ;
      RECT  8092.5 128087.5 8157.5 127952.5 ;
      RECT  8092.5 128087.5 8157.5 127952.5 ;
      RECT  7902.5 128087.5 7967.5 127952.5 ;
      RECT  8262.5 127157.5 8327.5 127022.5 ;
      RECT  8262.5 128132.5 8327.5 127997.5 ;
      RECT  8097.5 127875.0 7962.5 127810.0 ;
      RECT  7907.5 127735.0 7772.5 127670.0 ;
      RECT  7717.5 127595.0 7582.5 127530.0 ;
      RECT  7712.5 127247.5 7777.5 127112.5 ;
      RECT  8092.5 127247.5 8157.5 127112.5 ;
      RECT  8092.5 128087.5 8157.5 127952.5 ;
      RECT  8092.5 127630.0 8157.5 127495.0 ;
      RECT  7582.5 127595.0 7717.5 127530.0 ;
      RECT  7772.5 127735.0 7907.5 127670.0 ;
      RECT  7962.5 127875.0 8097.5 127810.0 ;
      RECT  8092.5 127630.0 8157.5 127495.0 ;
      RECT  7455.0 126937.5 8465.0 126872.5 ;
      RECT  7455.0 128282.5 8465.0 128217.5 ;
      RECT  7522.5 128412.5 7587.5 128217.5 ;
      RECT  7522.5 129252.5 7587.5 129627.5 ;
      RECT  7902.5 129252.5 7967.5 129627.5 ;
      RECT  8262.5 129410.0 8327.5 129595.0 ;
      RECT  8262.5 128250.0 8327.5 128435.0 ;
      RECT  7522.5 129252.5 7587.5 129387.5 ;
      RECT  7712.5 129252.5 7777.5 129387.5 ;
      RECT  7712.5 129252.5 7777.5 129387.5 ;
      RECT  7522.5 129252.5 7587.5 129387.5 ;
      RECT  7712.5 129252.5 7777.5 129387.5 ;
      RECT  7902.5 129252.5 7967.5 129387.5 ;
      RECT  7902.5 129252.5 7967.5 129387.5 ;
      RECT  7712.5 129252.5 7777.5 129387.5 ;
      RECT  7902.5 129252.5 7967.5 129387.5 ;
      RECT  8092.5 129252.5 8157.5 129387.5 ;
      RECT  8092.5 129252.5 8157.5 129387.5 ;
      RECT  7902.5 129252.5 7967.5 129387.5 ;
      RECT  7522.5 128412.5 7587.5 128547.5 ;
      RECT  7712.5 128412.5 7777.5 128547.5 ;
      RECT  7712.5 128412.5 7777.5 128547.5 ;
      RECT  7522.5 128412.5 7587.5 128547.5 ;
      RECT  7712.5 128412.5 7777.5 128547.5 ;
      RECT  7902.5 128412.5 7967.5 128547.5 ;
      RECT  7902.5 128412.5 7967.5 128547.5 ;
      RECT  7712.5 128412.5 7777.5 128547.5 ;
      RECT  7902.5 128412.5 7967.5 128547.5 ;
      RECT  8092.5 128412.5 8157.5 128547.5 ;
      RECT  8092.5 128412.5 8157.5 128547.5 ;
      RECT  7902.5 128412.5 7967.5 128547.5 ;
      RECT  8262.5 129342.5 8327.5 129477.5 ;
      RECT  8262.5 128367.5 8327.5 128502.5 ;
      RECT  8097.5 128625.0 7962.5 128690.0 ;
      RECT  7907.5 128765.0 7772.5 128830.0 ;
      RECT  7717.5 128905.0 7582.5 128970.0 ;
      RECT  7712.5 129252.5 7777.5 129387.5 ;
      RECT  8092.5 129252.5 8157.5 129387.5 ;
      RECT  8092.5 128412.5 8157.5 128547.5 ;
      RECT  8092.5 128870.0 8157.5 129005.0 ;
      RECT  7582.5 128905.0 7717.5 128970.0 ;
      RECT  7772.5 128765.0 7907.5 128830.0 ;
      RECT  7962.5 128625.0 8097.5 128690.0 ;
      RECT  8092.5 128870.0 8157.5 129005.0 ;
      RECT  7455.0 129562.5 8465.0 129627.5 ;
      RECT  7455.0 128217.5 8465.0 128282.5 ;
      RECT  7522.5 130777.5 7587.5 130972.5 ;
      RECT  7522.5 129937.5 7587.5 129562.5 ;
      RECT  7902.5 129937.5 7967.5 129562.5 ;
      RECT  8262.5 129780.0 8327.5 129595.0 ;
      RECT  8262.5 130940.0 8327.5 130755.0 ;
      RECT  7522.5 129937.5 7587.5 129802.5 ;
      RECT  7712.5 129937.5 7777.5 129802.5 ;
      RECT  7712.5 129937.5 7777.5 129802.5 ;
      RECT  7522.5 129937.5 7587.5 129802.5 ;
      RECT  7712.5 129937.5 7777.5 129802.5 ;
      RECT  7902.5 129937.5 7967.5 129802.5 ;
      RECT  7902.5 129937.5 7967.5 129802.5 ;
      RECT  7712.5 129937.5 7777.5 129802.5 ;
      RECT  7902.5 129937.5 7967.5 129802.5 ;
      RECT  8092.5 129937.5 8157.5 129802.5 ;
      RECT  8092.5 129937.5 8157.5 129802.5 ;
      RECT  7902.5 129937.5 7967.5 129802.5 ;
      RECT  7522.5 130777.5 7587.5 130642.5 ;
      RECT  7712.5 130777.5 7777.5 130642.5 ;
      RECT  7712.5 130777.5 7777.5 130642.5 ;
      RECT  7522.5 130777.5 7587.5 130642.5 ;
      RECT  7712.5 130777.5 7777.5 130642.5 ;
      RECT  7902.5 130777.5 7967.5 130642.5 ;
      RECT  7902.5 130777.5 7967.5 130642.5 ;
      RECT  7712.5 130777.5 7777.5 130642.5 ;
      RECT  7902.5 130777.5 7967.5 130642.5 ;
      RECT  8092.5 130777.5 8157.5 130642.5 ;
      RECT  8092.5 130777.5 8157.5 130642.5 ;
      RECT  7902.5 130777.5 7967.5 130642.5 ;
      RECT  8262.5 129847.5 8327.5 129712.5 ;
      RECT  8262.5 130822.5 8327.5 130687.5 ;
      RECT  8097.5 130565.0 7962.5 130500.0 ;
      RECT  7907.5 130425.0 7772.5 130360.0 ;
      RECT  7717.5 130285.0 7582.5 130220.0 ;
      RECT  7712.5 129937.5 7777.5 129802.5 ;
      RECT  8092.5 129937.5 8157.5 129802.5 ;
      RECT  8092.5 130777.5 8157.5 130642.5 ;
      RECT  8092.5 130320.0 8157.5 130185.0 ;
      RECT  7582.5 130285.0 7717.5 130220.0 ;
      RECT  7772.5 130425.0 7907.5 130360.0 ;
      RECT  7962.5 130565.0 8097.5 130500.0 ;
      RECT  8092.5 130320.0 8157.5 130185.0 ;
      RECT  7455.0 129627.5 8465.0 129562.5 ;
      RECT  7455.0 130972.5 8465.0 130907.5 ;
      RECT  7522.5 131102.5 7587.5 130907.5 ;
      RECT  7522.5 131942.5 7587.5 132317.5 ;
      RECT  7902.5 131942.5 7967.5 132317.5 ;
      RECT  8262.5 132100.0 8327.5 132285.0 ;
      RECT  8262.5 130940.0 8327.5 131125.0 ;
      RECT  7522.5 131942.5 7587.5 132077.5 ;
      RECT  7712.5 131942.5 7777.5 132077.5 ;
      RECT  7712.5 131942.5 7777.5 132077.5 ;
      RECT  7522.5 131942.5 7587.5 132077.5 ;
      RECT  7712.5 131942.5 7777.5 132077.5 ;
      RECT  7902.5 131942.5 7967.5 132077.5 ;
      RECT  7902.5 131942.5 7967.5 132077.5 ;
      RECT  7712.5 131942.5 7777.5 132077.5 ;
      RECT  7902.5 131942.5 7967.5 132077.5 ;
      RECT  8092.5 131942.5 8157.5 132077.5 ;
      RECT  8092.5 131942.5 8157.5 132077.5 ;
      RECT  7902.5 131942.5 7967.5 132077.5 ;
      RECT  7522.5 131102.5 7587.5 131237.5 ;
      RECT  7712.5 131102.5 7777.5 131237.5 ;
      RECT  7712.5 131102.5 7777.5 131237.5 ;
      RECT  7522.5 131102.5 7587.5 131237.5 ;
      RECT  7712.5 131102.5 7777.5 131237.5 ;
      RECT  7902.5 131102.5 7967.5 131237.5 ;
      RECT  7902.5 131102.5 7967.5 131237.5 ;
      RECT  7712.5 131102.5 7777.5 131237.5 ;
      RECT  7902.5 131102.5 7967.5 131237.5 ;
      RECT  8092.5 131102.5 8157.5 131237.5 ;
      RECT  8092.5 131102.5 8157.5 131237.5 ;
      RECT  7902.5 131102.5 7967.5 131237.5 ;
      RECT  8262.5 132032.5 8327.5 132167.5 ;
      RECT  8262.5 131057.5 8327.5 131192.5 ;
      RECT  8097.5 131315.0 7962.5 131380.0 ;
      RECT  7907.5 131455.0 7772.5 131520.0 ;
      RECT  7717.5 131595.0 7582.5 131660.0 ;
      RECT  7712.5 131942.5 7777.5 132077.5 ;
      RECT  8092.5 131942.5 8157.5 132077.5 ;
      RECT  8092.5 131102.5 8157.5 131237.5 ;
      RECT  8092.5 131560.0 8157.5 131695.0 ;
      RECT  7582.5 131595.0 7717.5 131660.0 ;
      RECT  7772.5 131455.0 7907.5 131520.0 ;
      RECT  7962.5 131315.0 8097.5 131380.0 ;
      RECT  8092.5 131560.0 8157.5 131695.0 ;
      RECT  7455.0 132252.5 8465.0 132317.5 ;
      RECT  7455.0 130907.5 8465.0 130972.5 ;
      RECT  7522.5 133467.5 7587.5 133662.5 ;
      RECT  7522.5 132627.5 7587.5 132252.5 ;
      RECT  7902.5 132627.5 7967.5 132252.5 ;
      RECT  8262.5 132470.0 8327.5 132285.0 ;
      RECT  8262.5 133630.0 8327.5 133445.0 ;
      RECT  7522.5 132627.5 7587.5 132492.5 ;
      RECT  7712.5 132627.5 7777.5 132492.5 ;
      RECT  7712.5 132627.5 7777.5 132492.5 ;
      RECT  7522.5 132627.5 7587.5 132492.5 ;
      RECT  7712.5 132627.5 7777.5 132492.5 ;
      RECT  7902.5 132627.5 7967.5 132492.5 ;
      RECT  7902.5 132627.5 7967.5 132492.5 ;
      RECT  7712.5 132627.5 7777.5 132492.5 ;
      RECT  7902.5 132627.5 7967.5 132492.5 ;
      RECT  8092.5 132627.5 8157.5 132492.5 ;
      RECT  8092.5 132627.5 8157.5 132492.5 ;
      RECT  7902.5 132627.5 7967.5 132492.5 ;
      RECT  7522.5 133467.5 7587.5 133332.5 ;
      RECT  7712.5 133467.5 7777.5 133332.5 ;
      RECT  7712.5 133467.5 7777.5 133332.5 ;
      RECT  7522.5 133467.5 7587.5 133332.5 ;
      RECT  7712.5 133467.5 7777.5 133332.5 ;
      RECT  7902.5 133467.5 7967.5 133332.5 ;
      RECT  7902.5 133467.5 7967.5 133332.5 ;
      RECT  7712.5 133467.5 7777.5 133332.5 ;
      RECT  7902.5 133467.5 7967.5 133332.5 ;
      RECT  8092.5 133467.5 8157.5 133332.5 ;
      RECT  8092.5 133467.5 8157.5 133332.5 ;
      RECT  7902.5 133467.5 7967.5 133332.5 ;
      RECT  8262.5 132537.5 8327.5 132402.5 ;
      RECT  8262.5 133512.5 8327.5 133377.5 ;
      RECT  8097.5 133255.0 7962.5 133190.0 ;
      RECT  7907.5 133115.0 7772.5 133050.0 ;
      RECT  7717.5 132975.0 7582.5 132910.0 ;
      RECT  7712.5 132627.5 7777.5 132492.5 ;
      RECT  8092.5 132627.5 8157.5 132492.5 ;
      RECT  8092.5 133467.5 8157.5 133332.5 ;
      RECT  8092.5 133010.0 8157.5 132875.0 ;
      RECT  7582.5 132975.0 7717.5 132910.0 ;
      RECT  7772.5 133115.0 7907.5 133050.0 ;
      RECT  7962.5 133255.0 8097.5 133190.0 ;
      RECT  8092.5 133010.0 8157.5 132875.0 ;
      RECT  7455.0 132317.5 8465.0 132252.5 ;
      RECT  7455.0 133662.5 8465.0 133597.5 ;
      RECT  7522.5 133792.5 7587.5 133597.5 ;
      RECT  7522.5 134632.5 7587.5 135007.5 ;
      RECT  7902.5 134632.5 7967.5 135007.5 ;
      RECT  8262.5 134790.0 8327.5 134975.0 ;
      RECT  8262.5 133630.0 8327.5 133815.0 ;
      RECT  7522.5 134632.5 7587.5 134767.5 ;
      RECT  7712.5 134632.5 7777.5 134767.5 ;
      RECT  7712.5 134632.5 7777.5 134767.5 ;
      RECT  7522.5 134632.5 7587.5 134767.5 ;
      RECT  7712.5 134632.5 7777.5 134767.5 ;
      RECT  7902.5 134632.5 7967.5 134767.5 ;
      RECT  7902.5 134632.5 7967.5 134767.5 ;
      RECT  7712.5 134632.5 7777.5 134767.5 ;
      RECT  7902.5 134632.5 7967.5 134767.5 ;
      RECT  8092.5 134632.5 8157.5 134767.5 ;
      RECT  8092.5 134632.5 8157.5 134767.5 ;
      RECT  7902.5 134632.5 7967.5 134767.5 ;
      RECT  7522.5 133792.5 7587.5 133927.5 ;
      RECT  7712.5 133792.5 7777.5 133927.5 ;
      RECT  7712.5 133792.5 7777.5 133927.5 ;
      RECT  7522.5 133792.5 7587.5 133927.5 ;
      RECT  7712.5 133792.5 7777.5 133927.5 ;
      RECT  7902.5 133792.5 7967.5 133927.5 ;
      RECT  7902.5 133792.5 7967.5 133927.5 ;
      RECT  7712.5 133792.5 7777.5 133927.5 ;
      RECT  7902.5 133792.5 7967.5 133927.5 ;
      RECT  8092.5 133792.5 8157.5 133927.5 ;
      RECT  8092.5 133792.5 8157.5 133927.5 ;
      RECT  7902.5 133792.5 7967.5 133927.5 ;
      RECT  8262.5 134722.5 8327.5 134857.5 ;
      RECT  8262.5 133747.5 8327.5 133882.5 ;
      RECT  8097.5 134005.0 7962.5 134070.0 ;
      RECT  7907.5 134145.0 7772.5 134210.0 ;
      RECT  7717.5 134285.0 7582.5 134350.0 ;
      RECT  7712.5 134632.5 7777.5 134767.5 ;
      RECT  8092.5 134632.5 8157.5 134767.5 ;
      RECT  8092.5 133792.5 8157.5 133927.5 ;
      RECT  8092.5 134250.0 8157.5 134385.0 ;
      RECT  7582.5 134285.0 7717.5 134350.0 ;
      RECT  7772.5 134145.0 7907.5 134210.0 ;
      RECT  7962.5 134005.0 8097.5 134070.0 ;
      RECT  8092.5 134250.0 8157.5 134385.0 ;
      RECT  7455.0 134942.5 8465.0 135007.5 ;
      RECT  7455.0 133597.5 8465.0 133662.5 ;
      RECT  7522.5 136157.5 7587.5 136352.5 ;
      RECT  7522.5 135317.5 7587.5 134942.5 ;
      RECT  7902.5 135317.5 7967.5 134942.5 ;
      RECT  8262.5 135160.0 8327.5 134975.0 ;
      RECT  8262.5 136320.0 8327.5 136135.0 ;
      RECT  7522.5 135317.5 7587.5 135182.5 ;
      RECT  7712.5 135317.5 7777.5 135182.5 ;
      RECT  7712.5 135317.5 7777.5 135182.5 ;
      RECT  7522.5 135317.5 7587.5 135182.5 ;
      RECT  7712.5 135317.5 7777.5 135182.5 ;
      RECT  7902.5 135317.5 7967.5 135182.5 ;
      RECT  7902.5 135317.5 7967.5 135182.5 ;
      RECT  7712.5 135317.5 7777.5 135182.5 ;
      RECT  7902.5 135317.5 7967.5 135182.5 ;
      RECT  8092.5 135317.5 8157.5 135182.5 ;
      RECT  8092.5 135317.5 8157.5 135182.5 ;
      RECT  7902.5 135317.5 7967.5 135182.5 ;
      RECT  7522.5 136157.5 7587.5 136022.5 ;
      RECT  7712.5 136157.5 7777.5 136022.5 ;
      RECT  7712.5 136157.5 7777.5 136022.5 ;
      RECT  7522.5 136157.5 7587.5 136022.5 ;
      RECT  7712.5 136157.5 7777.5 136022.5 ;
      RECT  7902.5 136157.5 7967.5 136022.5 ;
      RECT  7902.5 136157.5 7967.5 136022.5 ;
      RECT  7712.5 136157.5 7777.5 136022.5 ;
      RECT  7902.5 136157.5 7967.5 136022.5 ;
      RECT  8092.5 136157.5 8157.5 136022.5 ;
      RECT  8092.5 136157.5 8157.5 136022.5 ;
      RECT  7902.5 136157.5 7967.5 136022.5 ;
      RECT  8262.5 135227.5 8327.5 135092.5 ;
      RECT  8262.5 136202.5 8327.5 136067.5 ;
      RECT  8097.5 135945.0 7962.5 135880.0 ;
      RECT  7907.5 135805.0 7772.5 135740.0 ;
      RECT  7717.5 135665.0 7582.5 135600.0 ;
      RECT  7712.5 135317.5 7777.5 135182.5 ;
      RECT  8092.5 135317.5 8157.5 135182.5 ;
      RECT  8092.5 136157.5 8157.5 136022.5 ;
      RECT  8092.5 135700.0 8157.5 135565.0 ;
      RECT  7582.5 135665.0 7717.5 135600.0 ;
      RECT  7772.5 135805.0 7907.5 135740.0 ;
      RECT  7962.5 135945.0 8097.5 135880.0 ;
      RECT  8092.5 135700.0 8157.5 135565.0 ;
      RECT  7455.0 135007.5 8465.0 134942.5 ;
      RECT  7455.0 136352.5 8465.0 136287.5 ;
      RECT  7522.5 136482.5 7587.5 136287.5 ;
      RECT  7522.5 137322.5 7587.5 137697.5 ;
      RECT  7902.5 137322.5 7967.5 137697.5 ;
      RECT  8262.5 137480.0 8327.5 137665.0 ;
      RECT  8262.5 136320.0 8327.5 136505.0 ;
      RECT  7522.5 137322.5 7587.5 137457.5 ;
      RECT  7712.5 137322.5 7777.5 137457.5 ;
      RECT  7712.5 137322.5 7777.5 137457.5 ;
      RECT  7522.5 137322.5 7587.5 137457.5 ;
      RECT  7712.5 137322.5 7777.5 137457.5 ;
      RECT  7902.5 137322.5 7967.5 137457.5 ;
      RECT  7902.5 137322.5 7967.5 137457.5 ;
      RECT  7712.5 137322.5 7777.5 137457.5 ;
      RECT  7902.5 137322.5 7967.5 137457.5 ;
      RECT  8092.5 137322.5 8157.5 137457.5 ;
      RECT  8092.5 137322.5 8157.5 137457.5 ;
      RECT  7902.5 137322.5 7967.5 137457.5 ;
      RECT  7522.5 136482.5 7587.5 136617.5 ;
      RECT  7712.5 136482.5 7777.5 136617.5 ;
      RECT  7712.5 136482.5 7777.5 136617.5 ;
      RECT  7522.5 136482.5 7587.5 136617.5 ;
      RECT  7712.5 136482.5 7777.5 136617.5 ;
      RECT  7902.5 136482.5 7967.5 136617.5 ;
      RECT  7902.5 136482.5 7967.5 136617.5 ;
      RECT  7712.5 136482.5 7777.5 136617.5 ;
      RECT  7902.5 136482.5 7967.5 136617.5 ;
      RECT  8092.5 136482.5 8157.5 136617.5 ;
      RECT  8092.5 136482.5 8157.5 136617.5 ;
      RECT  7902.5 136482.5 7967.5 136617.5 ;
      RECT  8262.5 137412.5 8327.5 137547.5 ;
      RECT  8262.5 136437.5 8327.5 136572.5 ;
      RECT  8097.5 136695.0 7962.5 136760.0 ;
      RECT  7907.5 136835.0 7772.5 136900.0 ;
      RECT  7717.5 136975.0 7582.5 137040.0 ;
      RECT  7712.5 137322.5 7777.5 137457.5 ;
      RECT  8092.5 137322.5 8157.5 137457.5 ;
      RECT  8092.5 136482.5 8157.5 136617.5 ;
      RECT  8092.5 136940.0 8157.5 137075.0 ;
      RECT  7582.5 136975.0 7717.5 137040.0 ;
      RECT  7772.5 136835.0 7907.5 136900.0 ;
      RECT  7962.5 136695.0 8097.5 136760.0 ;
      RECT  8092.5 136940.0 8157.5 137075.0 ;
      RECT  7455.0 137632.5 8465.0 137697.5 ;
      RECT  7455.0 136287.5 8465.0 136352.5 ;
      RECT  7522.5 138847.5 7587.5 139042.5 ;
      RECT  7522.5 138007.5 7587.5 137632.5 ;
      RECT  7902.5 138007.5 7967.5 137632.5 ;
      RECT  8262.5 137850.0 8327.5 137665.0 ;
      RECT  8262.5 139010.0 8327.5 138825.0 ;
      RECT  7522.5 138007.5 7587.5 137872.5 ;
      RECT  7712.5 138007.5 7777.5 137872.5 ;
      RECT  7712.5 138007.5 7777.5 137872.5 ;
      RECT  7522.5 138007.5 7587.5 137872.5 ;
      RECT  7712.5 138007.5 7777.5 137872.5 ;
      RECT  7902.5 138007.5 7967.5 137872.5 ;
      RECT  7902.5 138007.5 7967.5 137872.5 ;
      RECT  7712.5 138007.5 7777.5 137872.5 ;
      RECT  7902.5 138007.5 7967.5 137872.5 ;
      RECT  8092.5 138007.5 8157.5 137872.5 ;
      RECT  8092.5 138007.5 8157.5 137872.5 ;
      RECT  7902.5 138007.5 7967.5 137872.5 ;
      RECT  7522.5 138847.5 7587.5 138712.5 ;
      RECT  7712.5 138847.5 7777.5 138712.5 ;
      RECT  7712.5 138847.5 7777.5 138712.5 ;
      RECT  7522.5 138847.5 7587.5 138712.5 ;
      RECT  7712.5 138847.5 7777.5 138712.5 ;
      RECT  7902.5 138847.5 7967.5 138712.5 ;
      RECT  7902.5 138847.5 7967.5 138712.5 ;
      RECT  7712.5 138847.5 7777.5 138712.5 ;
      RECT  7902.5 138847.5 7967.5 138712.5 ;
      RECT  8092.5 138847.5 8157.5 138712.5 ;
      RECT  8092.5 138847.5 8157.5 138712.5 ;
      RECT  7902.5 138847.5 7967.5 138712.5 ;
      RECT  8262.5 137917.5 8327.5 137782.5 ;
      RECT  8262.5 138892.5 8327.5 138757.5 ;
      RECT  8097.5 138635.0 7962.5 138570.0 ;
      RECT  7907.5 138495.0 7772.5 138430.0 ;
      RECT  7717.5 138355.0 7582.5 138290.0 ;
      RECT  7712.5 138007.5 7777.5 137872.5 ;
      RECT  8092.5 138007.5 8157.5 137872.5 ;
      RECT  8092.5 138847.5 8157.5 138712.5 ;
      RECT  8092.5 138390.0 8157.5 138255.0 ;
      RECT  7582.5 138355.0 7717.5 138290.0 ;
      RECT  7772.5 138495.0 7907.5 138430.0 ;
      RECT  7962.5 138635.0 8097.5 138570.0 ;
      RECT  8092.5 138390.0 8157.5 138255.0 ;
      RECT  7455.0 137697.5 8465.0 137632.5 ;
      RECT  7455.0 139042.5 8465.0 138977.5 ;
      RECT  7522.5 139172.5 7587.5 138977.5 ;
      RECT  7522.5 140012.5 7587.5 140387.5 ;
      RECT  7902.5 140012.5 7967.5 140387.5 ;
      RECT  8262.5 140170.0 8327.5 140355.0 ;
      RECT  8262.5 139010.0 8327.5 139195.0 ;
      RECT  7522.5 140012.5 7587.5 140147.5 ;
      RECT  7712.5 140012.5 7777.5 140147.5 ;
      RECT  7712.5 140012.5 7777.5 140147.5 ;
      RECT  7522.5 140012.5 7587.5 140147.5 ;
      RECT  7712.5 140012.5 7777.5 140147.5 ;
      RECT  7902.5 140012.5 7967.5 140147.5 ;
      RECT  7902.5 140012.5 7967.5 140147.5 ;
      RECT  7712.5 140012.5 7777.5 140147.5 ;
      RECT  7902.5 140012.5 7967.5 140147.5 ;
      RECT  8092.5 140012.5 8157.5 140147.5 ;
      RECT  8092.5 140012.5 8157.5 140147.5 ;
      RECT  7902.5 140012.5 7967.5 140147.5 ;
      RECT  7522.5 139172.5 7587.5 139307.5 ;
      RECT  7712.5 139172.5 7777.5 139307.5 ;
      RECT  7712.5 139172.5 7777.5 139307.5 ;
      RECT  7522.5 139172.5 7587.5 139307.5 ;
      RECT  7712.5 139172.5 7777.5 139307.5 ;
      RECT  7902.5 139172.5 7967.5 139307.5 ;
      RECT  7902.5 139172.5 7967.5 139307.5 ;
      RECT  7712.5 139172.5 7777.5 139307.5 ;
      RECT  7902.5 139172.5 7967.5 139307.5 ;
      RECT  8092.5 139172.5 8157.5 139307.5 ;
      RECT  8092.5 139172.5 8157.5 139307.5 ;
      RECT  7902.5 139172.5 7967.5 139307.5 ;
      RECT  8262.5 140102.5 8327.5 140237.5 ;
      RECT  8262.5 139127.5 8327.5 139262.5 ;
      RECT  8097.5 139385.0 7962.5 139450.0 ;
      RECT  7907.5 139525.0 7772.5 139590.0 ;
      RECT  7717.5 139665.0 7582.5 139730.0 ;
      RECT  7712.5 140012.5 7777.5 140147.5 ;
      RECT  8092.5 140012.5 8157.5 140147.5 ;
      RECT  8092.5 139172.5 8157.5 139307.5 ;
      RECT  8092.5 139630.0 8157.5 139765.0 ;
      RECT  7582.5 139665.0 7717.5 139730.0 ;
      RECT  7772.5 139525.0 7907.5 139590.0 ;
      RECT  7962.5 139385.0 8097.5 139450.0 ;
      RECT  8092.5 139630.0 8157.5 139765.0 ;
      RECT  7455.0 140322.5 8465.0 140387.5 ;
      RECT  7455.0 138977.5 8465.0 139042.5 ;
      RECT  7522.5 141537.5 7587.5 141732.5 ;
      RECT  7522.5 140697.5 7587.5 140322.5 ;
      RECT  7902.5 140697.5 7967.5 140322.5 ;
      RECT  8262.5 140540.0 8327.5 140355.0 ;
      RECT  8262.5 141700.0 8327.5 141515.0 ;
      RECT  7522.5 140697.5 7587.5 140562.5 ;
      RECT  7712.5 140697.5 7777.5 140562.5 ;
      RECT  7712.5 140697.5 7777.5 140562.5 ;
      RECT  7522.5 140697.5 7587.5 140562.5 ;
      RECT  7712.5 140697.5 7777.5 140562.5 ;
      RECT  7902.5 140697.5 7967.5 140562.5 ;
      RECT  7902.5 140697.5 7967.5 140562.5 ;
      RECT  7712.5 140697.5 7777.5 140562.5 ;
      RECT  7902.5 140697.5 7967.5 140562.5 ;
      RECT  8092.5 140697.5 8157.5 140562.5 ;
      RECT  8092.5 140697.5 8157.5 140562.5 ;
      RECT  7902.5 140697.5 7967.5 140562.5 ;
      RECT  7522.5 141537.5 7587.5 141402.5 ;
      RECT  7712.5 141537.5 7777.5 141402.5 ;
      RECT  7712.5 141537.5 7777.5 141402.5 ;
      RECT  7522.5 141537.5 7587.5 141402.5 ;
      RECT  7712.5 141537.5 7777.5 141402.5 ;
      RECT  7902.5 141537.5 7967.5 141402.5 ;
      RECT  7902.5 141537.5 7967.5 141402.5 ;
      RECT  7712.5 141537.5 7777.5 141402.5 ;
      RECT  7902.5 141537.5 7967.5 141402.5 ;
      RECT  8092.5 141537.5 8157.5 141402.5 ;
      RECT  8092.5 141537.5 8157.5 141402.5 ;
      RECT  7902.5 141537.5 7967.5 141402.5 ;
      RECT  8262.5 140607.5 8327.5 140472.5 ;
      RECT  8262.5 141582.5 8327.5 141447.5 ;
      RECT  8097.5 141325.0 7962.5 141260.0 ;
      RECT  7907.5 141185.0 7772.5 141120.0 ;
      RECT  7717.5 141045.0 7582.5 140980.0 ;
      RECT  7712.5 140697.5 7777.5 140562.5 ;
      RECT  8092.5 140697.5 8157.5 140562.5 ;
      RECT  8092.5 141537.5 8157.5 141402.5 ;
      RECT  8092.5 141080.0 8157.5 140945.0 ;
      RECT  7582.5 141045.0 7717.5 140980.0 ;
      RECT  7772.5 141185.0 7907.5 141120.0 ;
      RECT  7962.5 141325.0 8097.5 141260.0 ;
      RECT  8092.5 141080.0 8157.5 140945.0 ;
      RECT  7455.0 140387.5 8465.0 140322.5 ;
      RECT  7455.0 141732.5 8465.0 141667.5 ;
      RECT  7522.5 141862.5 7587.5 141667.5 ;
      RECT  7522.5 142702.5 7587.5 143077.5 ;
      RECT  7902.5 142702.5 7967.5 143077.5 ;
      RECT  8262.5 142860.0 8327.5 143045.0 ;
      RECT  8262.5 141700.0 8327.5 141885.0 ;
      RECT  7522.5 142702.5 7587.5 142837.5 ;
      RECT  7712.5 142702.5 7777.5 142837.5 ;
      RECT  7712.5 142702.5 7777.5 142837.5 ;
      RECT  7522.5 142702.5 7587.5 142837.5 ;
      RECT  7712.5 142702.5 7777.5 142837.5 ;
      RECT  7902.5 142702.5 7967.5 142837.5 ;
      RECT  7902.5 142702.5 7967.5 142837.5 ;
      RECT  7712.5 142702.5 7777.5 142837.5 ;
      RECT  7902.5 142702.5 7967.5 142837.5 ;
      RECT  8092.5 142702.5 8157.5 142837.5 ;
      RECT  8092.5 142702.5 8157.5 142837.5 ;
      RECT  7902.5 142702.5 7967.5 142837.5 ;
      RECT  7522.5 141862.5 7587.5 141997.5 ;
      RECT  7712.5 141862.5 7777.5 141997.5 ;
      RECT  7712.5 141862.5 7777.5 141997.5 ;
      RECT  7522.5 141862.5 7587.5 141997.5 ;
      RECT  7712.5 141862.5 7777.5 141997.5 ;
      RECT  7902.5 141862.5 7967.5 141997.5 ;
      RECT  7902.5 141862.5 7967.5 141997.5 ;
      RECT  7712.5 141862.5 7777.5 141997.5 ;
      RECT  7902.5 141862.5 7967.5 141997.5 ;
      RECT  8092.5 141862.5 8157.5 141997.5 ;
      RECT  8092.5 141862.5 8157.5 141997.5 ;
      RECT  7902.5 141862.5 7967.5 141997.5 ;
      RECT  8262.5 142792.5 8327.5 142927.5 ;
      RECT  8262.5 141817.5 8327.5 141952.5 ;
      RECT  8097.5 142075.0 7962.5 142140.0 ;
      RECT  7907.5 142215.0 7772.5 142280.0 ;
      RECT  7717.5 142355.0 7582.5 142420.0 ;
      RECT  7712.5 142702.5 7777.5 142837.5 ;
      RECT  8092.5 142702.5 8157.5 142837.5 ;
      RECT  8092.5 141862.5 8157.5 141997.5 ;
      RECT  8092.5 142320.0 8157.5 142455.0 ;
      RECT  7582.5 142355.0 7717.5 142420.0 ;
      RECT  7772.5 142215.0 7907.5 142280.0 ;
      RECT  7962.5 142075.0 8097.5 142140.0 ;
      RECT  8092.5 142320.0 8157.5 142455.0 ;
      RECT  7455.0 143012.5 8465.0 143077.5 ;
      RECT  7455.0 141667.5 8465.0 141732.5 ;
      RECT  7522.5 144227.5 7587.5 144422.5 ;
      RECT  7522.5 143387.5 7587.5 143012.5 ;
      RECT  7902.5 143387.5 7967.5 143012.5 ;
      RECT  8262.5 143230.0 8327.5 143045.0 ;
      RECT  8262.5 144390.0 8327.5 144205.0 ;
      RECT  7522.5 143387.5 7587.5 143252.5 ;
      RECT  7712.5 143387.5 7777.5 143252.5 ;
      RECT  7712.5 143387.5 7777.5 143252.5 ;
      RECT  7522.5 143387.5 7587.5 143252.5 ;
      RECT  7712.5 143387.5 7777.5 143252.5 ;
      RECT  7902.5 143387.5 7967.5 143252.5 ;
      RECT  7902.5 143387.5 7967.5 143252.5 ;
      RECT  7712.5 143387.5 7777.5 143252.5 ;
      RECT  7902.5 143387.5 7967.5 143252.5 ;
      RECT  8092.5 143387.5 8157.5 143252.5 ;
      RECT  8092.5 143387.5 8157.5 143252.5 ;
      RECT  7902.5 143387.5 7967.5 143252.5 ;
      RECT  7522.5 144227.5 7587.5 144092.5 ;
      RECT  7712.5 144227.5 7777.5 144092.5 ;
      RECT  7712.5 144227.5 7777.5 144092.5 ;
      RECT  7522.5 144227.5 7587.5 144092.5 ;
      RECT  7712.5 144227.5 7777.5 144092.5 ;
      RECT  7902.5 144227.5 7967.5 144092.5 ;
      RECT  7902.5 144227.5 7967.5 144092.5 ;
      RECT  7712.5 144227.5 7777.5 144092.5 ;
      RECT  7902.5 144227.5 7967.5 144092.5 ;
      RECT  8092.5 144227.5 8157.5 144092.5 ;
      RECT  8092.5 144227.5 8157.5 144092.5 ;
      RECT  7902.5 144227.5 7967.5 144092.5 ;
      RECT  8262.5 143297.5 8327.5 143162.5 ;
      RECT  8262.5 144272.5 8327.5 144137.5 ;
      RECT  8097.5 144015.0 7962.5 143950.0 ;
      RECT  7907.5 143875.0 7772.5 143810.0 ;
      RECT  7717.5 143735.0 7582.5 143670.0 ;
      RECT  7712.5 143387.5 7777.5 143252.5 ;
      RECT  8092.5 143387.5 8157.5 143252.5 ;
      RECT  8092.5 144227.5 8157.5 144092.5 ;
      RECT  8092.5 143770.0 8157.5 143635.0 ;
      RECT  7582.5 143735.0 7717.5 143670.0 ;
      RECT  7772.5 143875.0 7907.5 143810.0 ;
      RECT  7962.5 144015.0 8097.5 143950.0 ;
      RECT  8092.5 143770.0 8157.5 143635.0 ;
      RECT  7455.0 143077.5 8465.0 143012.5 ;
      RECT  7455.0 144422.5 8465.0 144357.5 ;
      RECT  7522.5 144552.5 7587.5 144357.5 ;
      RECT  7522.5 145392.5 7587.5 145767.5 ;
      RECT  7902.5 145392.5 7967.5 145767.5 ;
      RECT  8262.5 145550.0 8327.5 145735.0 ;
      RECT  8262.5 144390.0 8327.5 144575.0 ;
      RECT  7522.5 145392.5 7587.5 145527.5 ;
      RECT  7712.5 145392.5 7777.5 145527.5 ;
      RECT  7712.5 145392.5 7777.5 145527.5 ;
      RECT  7522.5 145392.5 7587.5 145527.5 ;
      RECT  7712.5 145392.5 7777.5 145527.5 ;
      RECT  7902.5 145392.5 7967.5 145527.5 ;
      RECT  7902.5 145392.5 7967.5 145527.5 ;
      RECT  7712.5 145392.5 7777.5 145527.5 ;
      RECT  7902.5 145392.5 7967.5 145527.5 ;
      RECT  8092.5 145392.5 8157.5 145527.5 ;
      RECT  8092.5 145392.5 8157.5 145527.5 ;
      RECT  7902.5 145392.5 7967.5 145527.5 ;
      RECT  7522.5 144552.5 7587.5 144687.5 ;
      RECT  7712.5 144552.5 7777.5 144687.5 ;
      RECT  7712.5 144552.5 7777.5 144687.5 ;
      RECT  7522.5 144552.5 7587.5 144687.5 ;
      RECT  7712.5 144552.5 7777.5 144687.5 ;
      RECT  7902.5 144552.5 7967.5 144687.5 ;
      RECT  7902.5 144552.5 7967.5 144687.5 ;
      RECT  7712.5 144552.5 7777.5 144687.5 ;
      RECT  7902.5 144552.5 7967.5 144687.5 ;
      RECT  8092.5 144552.5 8157.5 144687.5 ;
      RECT  8092.5 144552.5 8157.5 144687.5 ;
      RECT  7902.5 144552.5 7967.5 144687.5 ;
      RECT  8262.5 145482.5 8327.5 145617.5 ;
      RECT  8262.5 144507.5 8327.5 144642.5 ;
      RECT  8097.5 144765.0 7962.5 144830.0 ;
      RECT  7907.5 144905.0 7772.5 144970.0 ;
      RECT  7717.5 145045.0 7582.5 145110.0 ;
      RECT  7712.5 145392.5 7777.5 145527.5 ;
      RECT  8092.5 145392.5 8157.5 145527.5 ;
      RECT  8092.5 144552.5 8157.5 144687.5 ;
      RECT  8092.5 145010.0 8157.5 145145.0 ;
      RECT  7582.5 145045.0 7717.5 145110.0 ;
      RECT  7772.5 144905.0 7907.5 144970.0 ;
      RECT  7962.5 144765.0 8097.5 144830.0 ;
      RECT  8092.5 145010.0 8157.5 145145.0 ;
      RECT  7455.0 145702.5 8465.0 145767.5 ;
      RECT  7455.0 144357.5 8465.0 144422.5 ;
      RECT  7522.5 146917.5 7587.5 147112.5 ;
      RECT  7522.5 146077.5 7587.5 145702.5 ;
      RECT  7902.5 146077.5 7967.5 145702.5 ;
      RECT  8262.5 145920.0 8327.5 145735.0 ;
      RECT  8262.5 147080.0 8327.5 146895.0 ;
      RECT  7522.5 146077.5 7587.5 145942.5 ;
      RECT  7712.5 146077.5 7777.5 145942.5 ;
      RECT  7712.5 146077.5 7777.5 145942.5 ;
      RECT  7522.5 146077.5 7587.5 145942.5 ;
      RECT  7712.5 146077.5 7777.5 145942.5 ;
      RECT  7902.5 146077.5 7967.5 145942.5 ;
      RECT  7902.5 146077.5 7967.5 145942.5 ;
      RECT  7712.5 146077.5 7777.5 145942.5 ;
      RECT  7902.5 146077.5 7967.5 145942.5 ;
      RECT  8092.5 146077.5 8157.5 145942.5 ;
      RECT  8092.5 146077.5 8157.5 145942.5 ;
      RECT  7902.5 146077.5 7967.5 145942.5 ;
      RECT  7522.5 146917.5 7587.5 146782.5 ;
      RECT  7712.5 146917.5 7777.5 146782.5 ;
      RECT  7712.5 146917.5 7777.5 146782.5 ;
      RECT  7522.5 146917.5 7587.5 146782.5 ;
      RECT  7712.5 146917.5 7777.5 146782.5 ;
      RECT  7902.5 146917.5 7967.5 146782.5 ;
      RECT  7902.5 146917.5 7967.5 146782.5 ;
      RECT  7712.5 146917.5 7777.5 146782.5 ;
      RECT  7902.5 146917.5 7967.5 146782.5 ;
      RECT  8092.5 146917.5 8157.5 146782.5 ;
      RECT  8092.5 146917.5 8157.5 146782.5 ;
      RECT  7902.5 146917.5 7967.5 146782.5 ;
      RECT  8262.5 145987.5 8327.5 145852.5 ;
      RECT  8262.5 146962.5 8327.5 146827.5 ;
      RECT  8097.5 146705.0 7962.5 146640.0 ;
      RECT  7907.5 146565.0 7772.5 146500.0 ;
      RECT  7717.5 146425.0 7582.5 146360.0 ;
      RECT  7712.5 146077.5 7777.5 145942.5 ;
      RECT  8092.5 146077.5 8157.5 145942.5 ;
      RECT  8092.5 146917.5 8157.5 146782.5 ;
      RECT  8092.5 146460.0 8157.5 146325.0 ;
      RECT  7582.5 146425.0 7717.5 146360.0 ;
      RECT  7772.5 146565.0 7907.5 146500.0 ;
      RECT  7962.5 146705.0 8097.5 146640.0 ;
      RECT  8092.5 146460.0 8157.5 146325.0 ;
      RECT  7455.0 145767.5 8465.0 145702.5 ;
      RECT  7455.0 147112.5 8465.0 147047.5 ;
      RECT  7522.5 147242.5 7587.5 147047.5 ;
      RECT  7522.5 148082.5 7587.5 148457.5 ;
      RECT  7902.5 148082.5 7967.5 148457.5 ;
      RECT  8262.5 148240.0 8327.5 148425.0 ;
      RECT  8262.5 147080.0 8327.5 147265.0 ;
      RECT  7522.5 148082.5 7587.5 148217.5 ;
      RECT  7712.5 148082.5 7777.5 148217.5 ;
      RECT  7712.5 148082.5 7777.5 148217.5 ;
      RECT  7522.5 148082.5 7587.5 148217.5 ;
      RECT  7712.5 148082.5 7777.5 148217.5 ;
      RECT  7902.5 148082.5 7967.5 148217.5 ;
      RECT  7902.5 148082.5 7967.5 148217.5 ;
      RECT  7712.5 148082.5 7777.5 148217.5 ;
      RECT  7902.5 148082.5 7967.5 148217.5 ;
      RECT  8092.5 148082.5 8157.5 148217.5 ;
      RECT  8092.5 148082.5 8157.5 148217.5 ;
      RECT  7902.5 148082.5 7967.5 148217.5 ;
      RECT  7522.5 147242.5 7587.5 147377.5 ;
      RECT  7712.5 147242.5 7777.5 147377.5 ;
      RECT  7712.5 147242.5 7777.5 147377.5 ;
      RECT  7522.5 147242.5 7587.5 147377.5 ;
      RECT  7712.5 147242.5 7777.5 147377.5 ;
      RECT  7902.5 147242.5 7967.5 147377.5 ;
      RECT  7902.5 147242.5 7967.5 147377.5 ;
      RECT  7712.5 147242.5 7777.5 147377.5 ;
      RECT  7902.5 147242.5 7967.5 147377.5 ;
      RECT  8092.5 147242.5 8157.5 147377.5 ;
      RECT  8092.5 147242.5 8157.5 147377.5 ;
      RECT  7902.5 147242.5 7967.5 147377.5 ;
      RECT  8262.5 148172.5 8327.5 148307.5 ;
      RECT  8262.5 147197.5 8327.5 147332.5 ;
      RECT  8097.5 147455.0 7962.5 147520.0 ;
      RECT  7907.5 147595.0 7772.5 147660.0 ;
      RECT  7717.5 147735.0 7582.5 147800.0 ;
      RECT  7712.5 148082.5 7777.5 148217.5 ;
      RECT  8092.5 148082.5 8157.5 148217.5 ;
      RECT  8092.5 147242.5 8157.5 147377.5 ;
      RECT  8092.5 147700.0 8157.5 147835.0 ;
      RECT  7582.5 147735.0 7717.5 147800.0 ;
      RECT  7772.5 147595.0 7907.5 147660.0 ;
      RECT  7962.5 147455.0 8097.5 147520.0 ;
      RECT  8092.5 147700.0 8157.5 147835.0 ;
      RECT  7455.0 148392.5 8465.0 148457.5 ;
      RECT  7455.0 147047.5 8465.0 147112.5 ;
      RECT  7522.5 149607.5 7587.5 149802.5 ;
      RECT  7522.5 148767.5 7587.5 148392.5 ;
      RECT  7902.5 148767.5 7967.5 148392.5 ;
      RECT  8262.5 148610.0 8327.5 148425.0 ;
      RECT  8262.5 149770.0 8327.5 149585.0 ;
      RECT  7522.5 148767.5 7587.5 148632.5 ;
      RECT  7712.5 148767.5 7777.5 148632.5 ;
      RECT  7712.5 148767.5 7777.5 148632.5 ;
      RECT  7522.5 148767.5 7587.5 148632.5 ;
      RECT  7712.5 148767.5 7777.5 148632.5 ;
      RECT  7902.5 148767.5 7967.5 148632.5 ;
      RECT  7902.5 148767.5 7967.5 148632.5 ;
      RECT  7712.5 148767.5 7777.5 148632.5 ;
      RECT  7902.5 148767.5 7967.5 148632.5 ;
      RECT  8092.5 148767.5 8157.5 148632.5 ;
      RECT  8092.5 148767.5 8157.5 148632.5 ;
      RECT  7902.5 148767.5 7967.5 148632.5 ;
      RECT  7522.5 149607.5 7587.5 149472.5 ;
      RECT  7712.5 149607.5 7777.5 149472.5 ;
      RECT  7712.5 149607.5 7777.5 149472.5 ;
      RECT  7522.5 149607.5 7587.5 149472.5 ;
      RECT  7712.5 149607.5 7777.5 149472.5 ;
      RECT  7902.5 149607.5 7967.5 149472.5 ;
      RECT  7902.5 149607.5 7967.5 149472.5 ;
      RECT  7712.5 149607.5 7777.5 149472.5 ;
      RECT  7902.5 149607.5 7967.5 149472.5 ;
      RECT  8092.5 149607.5 8157.5 149472.5 ;
      RECT  8092.5 149607.5 8157.5 149472.5 ;
      RECT  7902.5 149607.5 7967.5 149472.5 ;
      RECT  8262.5 148677.5 8327.5 148542.5 ;
      RECT  8262.5 149652.5 8327.5 149517.5 ;
      RECT  8097.5 149395.0 7962.5 149330.0 ;
      RECT  7907.5 149255.0 7772.5 149190.0 ;
      RECT  7717.5 149115.0 7582.5 149050.0 ;
      RECT  7712.5 148767.5 7777.5 148632.5 ;
      RECT  8092.5 148767.5 8157.5 148632.5 ;
      RECT  8092.5 149607.5 8157.5 149472.5 ;
      RECT  8092.5 149150.0 8157.5 149015.0 ;
      RECT  7582.5 149115.0 7717.5 149050.0 ;
      RECT  7772.5 149255.0 7907.5 149190.0 ;
      RECT  7962.5 149395.0 8097.5 149330.0 ;
      RECT  8092.5 149150.0 8157.5 149015.0 ;
      RECT  7455.0 148457.5 8465.0 148392.5 ;
      RECT  7455.0 149802.5 8465.0 149737.5 ;
      RECT  7522.5 149932.5 7587.5 149737.5 ;
      RECT  7522.5 150772.5 7587.5 151147.5 ;
      RECT  7902.5 150772.5 7967.5 151147.5 ;
      RECT  8262.5 150930.0 8327.5 151115.0 ;
      RECT  8262.5 149770.0 8327.5 149955.0 ;
      RECT  7522.5 150772.5 7587.5 150907.5 ;
      RECT  7712.5 150772.5 7777.5 150907.5 ;
      RECT  7712.5 150772.5 7777.5 150907.5 ;
      RECT  7522.5 150772.5 7587.5 150907.5 ;
      RECT  7712.5 150772.5 7777.5 150907.5 ;
      RECT  7902.5 150772.5 7967.5 150907.5 ;
      RECT  7902.5 150772.5 7967.5 150907.5 ;
      RECT  7712.5 150772.5 7777.5 150907.5 ;
      RECT  7902.5 150772.5 7967.5 150907.5 ;
      RECT  8092.5 150772.5 8157.5 150907.5 ;
      RECT  8092.5 150772.5 8157.5 150907.5 ;
      RECT  7902.5 150772.5 7967.5 150907.5 ;
      RECT  7522.5 149932.5 7587.5 150067.5 ;
      RECT  7712.5 149932.5 7777.5 150067.5 ;
      RECT  7712.5 149932.5 7777.5 150067.5 ;
      RECT  7522.5 149932.5 7587.5 150067.5 ;
      RECT  7712.5 149932.5 7777.5 150067.5 ;
      RECT  7902.5 149932.5 7967.5 150067.5 ;
      RECT  7902.5 149932.5 7967.5 150067.5 ;
      RECT  7712.5 149932.5 7777.5 150067.5 ;
      RECT  7902.5 149932.5 7967.5 150067.5 ;
      RECT  8092.5 149932.5 8157.5 150067.5 ;
      RECT  8092.5 149932.5 8157.5 150067.5 ;
      RECT  7902.5 149932.5 7967.5 150067.5 ;
      RECT  8262.5 150862.5 8327.5 150997.5 ;
      RECT  8262.5 149887.5 8327.5 150022.5 ;
      RECT  8097.5 150145.0 7962.5 150210.0 ;
      RECT  7907.5 150285.0 7772.5 150350.0 ;
      RECT  7717.5 150425.0 7582.5 150490.0 ;
      RECT  7712.5 150772.5 7777.5 150907.5 ;
      RECT  8092.5 150772.5 8157.5 150907.5 ;
      RECT  8092.5 149932.5 8157.5 150067.5 ;
      RECT  8092.5 150390.0 8157.5 150525.0 ;
      RECT  7582.5 150425.0 7717.5 150490.0 ;
      RECT  7772.5 150285.0 7907.5 150350.0 ;
      RECT  7962.5 150145.0 8097.5 150210.0 ;
      RECT  8092.5 150390.0 8157.5 150525.0 ;
      RECT  7455.0 151082.5 8465.0 151147.5 ;
      RECT  7455.0 149737.5 8465.0 149802.5 ;
      RECT  7522.5 152297.5 7587.5 152492.5 ;
      RECT  7522.5 151457.5 7587.5 151082.5 ;
      RECT  7902.5 151457.5 7967.5 151082.5 ;
      RECT  8262.5 151300.0 8327.5 151115.0 ;
      RECT  8262.5 152460.0 8327.5 152275.0 ;
      RECT  7522.5 151457.5 7587.5 151322.5 ;
      RECT  7712.5 151457.5 7777.5 151322.5 ;
      RECT  7712.5 151457.5 7777.5 151322.5 ;
      RECT  7522.5 151457.5 7587.5 151322.5 ;
      RECT  7712.5 151457.5 7777.5 151322.5 ;
      RECT  7902.5 151457.5 7967.5 151322.5 ;
      RECT  7902.5 151457.5 7967.5 151322.5 ;
      RECT  7712.5 151457.5 7777.5 151322.5 ;
      RECT  7902.5 151457.5 7967.5 151322.5 ;
      RECT  8092.5 151457.5 8157.5 151322.5 ;
      RECT  8092.5 151457.5 8157.5 151322.5 ;
      RECT  7902.5 151457.5 7967.5 151322.5 ;
      RECT  7522.5 152297.5 7587.5 152162.5 ;
      RECT  7712.5 152297.5 7777.5 152162.5 ;
      RECT  7712.5 152297.5 7777.5 152162.5 ;
      RECT  7522.5 152297.5 7587.5 152162.5 ;
      RECT  7712.5 152297.5 7777.5 152162.5 ;
      RECT  7902.5 152297.5 7967.5 152162.5 ;
      RECT  7902.5 152297.5 7967.5 152162.5 ;
      RECT  7712.5 152297.5 7777.5 152162.5 ;
      RECT  7902.5 152297.5 7967.5 152162.5 ;
      RECT  8092.5 152297.5 8157.5 152162.5 ;
      RECT  8092.5 152297.5 8157.5 152162.5 ;
      RECT  7902.5 152297.5 7967.5 152162.5 ;
      RECT  8262.5 151367.5 8327.5 151232.5 ;
      RECT  8262.5 152342.5 8327.5 152207.5 ;
      RECT  8097.5 152085.0 7962.5 152020.0 ;
      RECT  7907.5 151945.0 7772.5 151880.0 ;
      RECT  7717.5 151805.0 7582.5 151740.0 ;
      RECT  7712.5 151457.5 7777.5 151322.5 ;
      RECT  8092.5 151457.5 8157.5 151322.5 ;
      RECT  8092.5 152297.5 8157.5 152162.5 ;
      RECT  8092.5 151840.0 8157.5 151705.0 ;
      RECT  7582.5 151805.0 7717.5 151740.0 ;
      RECT  7772.5 151945.0 7907.5 151880.0 ;
      RECT  7962.5 152085.0 8097.5 152020.0 ;
      RECT  8092.5 151840.0 8157.5 151705.0 ;
      RECT  7455.0 151147.5 8465.0 151082.5 ;
      RECT  7455.0 152492.5 8465.0 152427.5 ;
      RECT  7522.5 152622.5 7587.5 152427.5 ;
      RECT  7522.5 153462.5 7587.5 153837.5 ;
      RECT  7902.5 153462.5 7967.5 153837.5 ;
      RECT  8262.5 153620.0 8327.5 153805.0 ;
      RECT  8262.5 152460.0 8327.5 152645.0 ;
      RECT  7522.5 153462.5 7587.5 153597.5 ;
      RECT  7712.5 153462.5 7777.5 153597.5 ;
      RECT  7712.5 153462.5 7777.5 153597.5 ;
      RECT  7522.5 153462.5 7587.5 153597.5 ;
      RECT  7712.5 153462.5 7777.5 153597.5 ;
      RECT  7902.5 153462.5 7967.5 153597.5 ;
      RECT  7902.5 153462.5 7967.5 153597.5 ;
      RECT  7712.5 153462.5 7777.5 153597.5 ;
      RECT  7902.5 153462.5 7967.5 153597.5 ;
      RECT  8092.5 153462.5 8157.5 153597.5 ;
      RECT  8092.5 153462.5 8157.5 153597.5 ;
      RECT  7902.5 153462.5 7967.5 153597.5 ;
      RECT  7522.5 152622.5 7587.5 152757.5 ;
      RECT  7712.5 152622.5 7777.5 152757.5 ;
      RECT  7712.5 152622.5 7777.5 152757.5 ;
      RECT  7522.5 152622.5 7587.5 152757.5 ;
      RECT  7712.5 152622.5 7777.5 152757.5 ;
      RECT  7902.5 152622.5 7967.5 152757.5 ;
      RECT  7902.5 152622.5 7967.5 152757.5 ;
      RECT  7712.5 152622.5 7777.5 152757.5 ;
      RECT  7902.5 152622.5 7967.5 152757.5 ;
      RECT  8092.5 152622.5 8157.5 152757.5 ;
      RECT  8092.5 152622.5 8157.5 152757.5 ;
      RECT  7902.5 152622.5 7967.5 152757.5 ;
      RECT  8262.5 153552.5 8327.5 153687.5 ;
      RECT  8262.5 152577.5 8327.5 152712.5 ;
      RECT  8097.5 152835.0 7962.5 152900.0 ;
      RECT  7907.5 152975.0 7772.5 153040.0 ;
      RECT  7717.5 153115.0 7582.5 153180.0 ;
      RECT  7712.5 153462.5 7777.5 153597.5 ;
      RECT  8092.5 153462.5 8157.5 153597.5 ;
      RECT  8092.5 152622.5 8157.5 152757.5 ;
      RECT  8092.5 153080.0 8157.5 153215.0 ;
      RECT  7582.5 153115.0 7717.5 153180.0 ;
      RECT  7772.5 152975.0 7907.5 153040.0 ;
      RECT  7962.5 152835.0 8097.5 152900.0 ;
      RECT  8092.5 153080.0 8157.5 153215.0 ;
      RECT  7455.0 153772.5 8465.0 153837.5 ;
      RECT  7455.0 152427.5 8465.0 152492.5 ;
      RECT  7522.5 154987.5 7587.5 155182.5 ;
      RECT  7522.5 154147.5 7587.5 153772.5 ;
      RECT  7902.5 154147.5 7967.5 153772.5 ;
      RECT  8262.5 153990.0 8327.5 153805.0 ;
      RECT  8262.5 155150.0 8327.5 154965.0 ;
      RECT  7522.5 154147.5 7587.5 154012.5 ;
      RECT  7712.5 154147.5 7777.5 154012.5 ;
      RECT  7712.5 154147.5 7777.5 154012.5 ;
      RECT  7522.5 154147.5 7587.5 154012.5 ;
      RECT  7712.5 154147.5 7777.5 154012.5 ;
      RECT  7902.5 154147.5 7967.5 154012.5 ;
      RECT  7902.5 154147.5 7967.5 154012.5 ;
      RECT  7712.5 154147.5 7777.5 154012.5 ;
      RECT  7902.5 154147.5 7967.5 154012.5 ;
      RECT  8092.5 154147.5 8157.5 154012.5 ;
      RECT  8092.5 154147.5 8157.5 154012.5 ;
      RECT  7902.5 154147.5 7967.5 154012.5 ;
      RECT  7522.5 154987.5 7587.5 154852.5 ;
      RECT  7712.5 154987.5 7777.5 154852.5 ;
      RECT  7712.5 154987.5 7777.5 154852.5 ;
      RECT  7522.5 154987.5 7587.5 154852.5 ;
      RECT  7712.5 154987.5 7777.5 154852.5 ;
      RECT  7902.5 154987.5 7967.5 154852.5 ;
      RECT  7902.5 154987.5 7967.5 154852.5 ;
      RECT  7712.5 154987.5 7777.5 154852.5 ;
      RECT  7902.5 154987.5 7967.5 154852.5 ;
      RECT  8092.5 154987.5 8157.5 154852.5 ;
      RECT  8092.5 154987.5 8157.5 154852.5 ;
      RECT  7902.5 154987.5 7967.5 154852.5 ;
      RECT  8262.5 154057.5 8327.5 153922.5 ;
      RECT  8262.5 155032.5 8327.5 154897.5 ;
      RECT  8097.5 154775.0 7962.5 154710.0 ;
      RECT  7907.5 154635.0 7772.5 154570.0 ;
      RECT  7717.5 154495.0 7582.5 154430.0 ;
      RECT  7712.5 154147.5 7777.5 154012.5 ;
      RECT  8092.5 154147.5 8157.5 154012.5 ;
      RECT  8092.5 154987.5 8157.5 154852.5 ;
      RECT  8092.5 154530.0 8157.5 154395.0 ;
      RECT  7582.5 154495.0 7717.5 154430.0 ;
      RECT  7772.5 154635.0 7907.5 154570.0 ;
      RECT  7962.5 154775.0 8097.5 154710.0 ;
      RECT  8092.5 154530.0 8157.5 154395.0 ;
      RECT  7455.0 153837.5 8465.0 153772.5 ;
      RECT  7455.0 155182.5 8465.0 155117.5 ;
      RECT  7522.5 155312.5 7587.5 155117.5 ;
      RECT  7522.5 156152.5 7587.5 156527.5 ;
      RECT  7902.5 156152.5 7967.5 156527.5 ;
      RECT  8262.5 156310.0 8327.5 156495.0 ;
      RECT  8262.5 155150.0 8327.5 155335.0 ;
      RECT  7522.5 156152.5 7587.5 156287.5 ;
      RECT  7712.5 156152.5 7777.5 156287.5 ;
      RECT  7712.5 156152.5 7777.5 156287.5 ;
      RECT  7522.5 156152.5 7587.5 156287.5 ;
      RECT  7712.5 156152.5 7777.5 156287.5 ;
      RECT  7902.5 156152.5 7967.5 156287.5 ;
      RECT  7902.5 156152.5 7967.5 156287.5 ;
      RECT  7712.5 156152.5 7777.5 156287.5 ;
      RECT  7902.5 156152.5 7967.5 156287.5 ;
      RECT  8092.5 156152.5 8157.5 156287.5 ;
      RECT  8092.5 156152.5 8157.5 156287.5 ;
      RECT  7902.5 156152.5 7967.5 156287.5 ;
      RECT  7522.5 155312.5 7587.5 155447.5 ;
      RECT  7712.5 155312.5 7777.5 155447.5 ;
      RECT  7712.5 155312.5 7777.5 155447.5 ;
      RECT  7522.5 155312.5 7587.5 155447.5 ;
      RECT  7712.5 155312.5 7777.5 155447.5 ;
      RECT  7902.5 155312.5 7967.5 155447.5 ;
      RECT  7902.5 155312.5 7967.5 155447.5 ;
      RECT  7712.5 155312.5 7777.5 155447.5 ;
      RECT  7902.5 155312.5 7967.5 155447.5 ;
      RECT  8092.5 155312.5 8157.5 155447.5 ;
      RECT  8092.5 155312.5 8157.5 155447.5 ;
      RECT  7902.5 155312.5 7967.5 155447.5 ;
      RECT  8262.5 156242.5 8327.5 156377.5 ;
      RECT  8262.5 155267.5 8327.5 155402.5 ;
      RECT  8097.5 155525.0 7962.5 155590.0 ;
      RECT  7907.5 155665.0 7772.5 155730.0 ;
      RECT  7717.5 155805.0 7582.5 155870.0 ;
      RECT  7712.5 156152.5 7777.5 156287.5 ;
      RECT  8092.5 156152.5 8157.5 156287.5 ;
      RECT  8092.5 155312.5 8157.5 155447.5 ;
      RECT  8092.5 155770.0 8157.5 155905.0 ;
      RECT  7582.5 155805.0 7717.5 155870.0 ;
      RECT  7772.5 155665.0 7907.5 155730.0 ;
      RECT  7962.5 155525.0 8097.5 155590.0 ;
      RECT  8092.5 155770.0 8157.5 155905.0 ;
      RECT  7455.0 156462.5 8465.0 156527.5 ;
      RECT  7455.0 155117.5 8465.0 155182.5 ;
      RECT  7522.5 157677.5 7587.5 157872.5 ;
      RECT  7522.5 156837.5 7587.5 156462.5 ;
      RECT  7902.5 156837.5 7967.5 156462.5 ;
      RECT  8262.5 156680.0 8327.5 156495.0 ;
      RECT  8262.5 157840.0 8327.5 157655.0 ;
      RECT  7522.5 156837.5 7587.5 156702.5 ;
      RECT  7712.5 156837.5 7777.5 156702.5 ;
      RECT  7712.5 156837.5 7777.5 156702.5 ;
      RECT  7522.5 156837.5 7587.5 156702.5 ;
      RECT  7712.5 156837.5 7777.5 156702.5 ;
      RECT  7902.5 156837.5 7967.5 156702.5 ;
      RECT  7902.5 156837.5 7967.5 156702.5 ;
      RECT  7712.5 156837.5 7777.5 156702.5 ;
      RECT  7902.5 156837.5 7967.5 156702.5 ;
      RECT  8092.5 156837.5 8157.5 156702.5 ;
      RECT  8092.5 156837.5 8157.5 156702.5 ;
      RECT  7902.5 156837.5 7967.5 156702.5 ;
      RECT  7522.5 157677.5 7587.5 157542.5 ;
      RECT  7712.5 157677.5 7777.5 157542.5 ;
      RECT  7712.5 157677.5 7777.5 157542.5 ;
      RECT  7522.5 157677.5 7587.5 157542.5 ;
      RECT  7712.5 157677.5 7777.5 157542.5 ;
      RECT  7902.5 157677.5 7967.5 157542.5 ;
      RECT  7902.5 157677.5 7967.5 157542.5 ;
      RECT  7712.5 157677.5 7777.5 157542.5 ;
      RECT  7902.5 157677.5 7967.5 157542.5 ;
      RECT  8092.5 157677.5 8157.5 157542.5 ;
      RECT  8092.5 157677.5 8157.5 157542.5 ;
      RECT  7902.5 157677.5 7967.5 157542.5 ;
      RECT  8262.5 156747.5 8327.5 156612.5 ;
      RECT  8262.5 157722.5 8327.5 157587.5 ;
      RECT  8097.5 157465.0 7962.5 157400.0 ;
      RECT  7907.5 157325.0 7772.5 157260.0 ;
      RECT  7717.5 157185.0 7582.5 157120.0 ;
      RECT  7712.5 156837.5 7777.5 156702.5 ;
      RECT  8092.5 156837.5 8157.5 156702.5 ;
      RECT  8092.5 157677.5 8157.5 157542.5 ;
      RECT  8092.5 157220.0 8157.5 157085.0 ;
      RECT  7582.5 157185.0 7717.5 157120.0 ;
      RECT  7772.5 157325.0 7907.5 157260.0 ;
      RECT  7962.5 157465.0 8097.5 157400.0 ;
      RECT  8092.5 157220.0 8157.5 157085.0 ;
      RECT  7455.0 156527.5 8465.0 156462.5 ;
      RECT  7455.0 157872.5 8465.0 157807.5 ;
      RECT  7522.5 158002.5 7587.5 157807.5 ;
      RECT  7522.5 158842.5 7587.5 159217.5 ;
      RECT  7902.5 158842.5 7967.5 159217.5 ;
      RECT  8262.5 159000.0 8327.5 159185.0 ;
      RECT  8262.5 157840.0 8327.5 158025.0 ;
      RECT  7522.5 158842.5 7587.5 158977.5 ;
      RECT  7712.5 158842.5 7777.5 158977.5 ;
      RECT  7712.5 158842.5 7777.5 158977.5 ;
      RECT  7522.5 158842.5 7587.5 158977.5 ;
      RECT  7712.5 158842.5 7777.5 158977.5 ;
      RECT  7902.5 158842.5 7967.5 158977.5 ;
      RECT  7902.5 158842.5 7967.5 158977.5 ;
      RECT  7712.5 158842.5 7777.5 158977.5 ;
      RECT  7902.5 158842.5 7967.5 158977.5 ;
      RECT  8092.5 158842.5 8157.5 158977.5 ;
      RECT  8092.5 158842.5 8157.5 158977.5 ;
      RECT  7902.5 158842.5 7967.5 158977.5 ;
      RECT  7522.5 158002.5 7587.5 158137.5 ;
      RECT  7712.5 158002.5 7777.5 158137.5 ;
      RECT  7712.5 158002.5 7777.5 158137.5 ;
      RECT  7522.5 158002.5 7587.5 158137.5 ;
      RECT  7712.5 158002.5 7777.5 158137.5 ;
      RECT  7902.5 158002.5 7967.5 158137.5 ;
      RECT  7902.5 158002.5 7967.5 158137.5 ;
      RECT  7712.5 158002.5 7777.5 158137.5 ;
      RECT  7902.5 158002.5 7967.5 158137.5 ;
      RECT  8092.5 158002.5 8157.5 158137.5 ;
      RECT  8092.5 158002.5 8157.5 158137.5 ;
      RECT  7902.5 158002.5 7967.5 158137.5 ;
      RECT  8262.5 158932.5 8327.5 159067.5 ;
      RECT  8262.5 157957.5 8327.5 158092.5 ;
      RECT  8097.5 158215.0 7962.5 158280.0 ;
      RECT  7907.5 158355.0 7772.5 158420.0 ;
      RECT  7717.5 158495.0 7582.5 158560.0 ;
      RECT  7712.5 158842.5 7777.5 158977.5 ;
      RECT  8092.5 158842.5 8157.5 158977.5 ;
      RECT  8092.5 158002.5 8157.5 158137.5 ;
      RECT  8092.5 158460.0 8157.5 158595.0 ;
      RECT  7582.5 158495.0 7717.5 158560.0 ;
      RECT  7772.5 158355.0 7907.5 158420.0 ;
      RECT  7962.5 158215.0 8097.5 158280.0 ;
      RECT  8092.5 158460.0 8157.5 158595.0 ;
      RECT  7455.0 159152.5 8465.0 159217.5 ;
      RECT  7455.0 157807.5 8465.0 157872.5 ;
      RECT  7522.5 160367.5 7587.5 160562.5 ;
      RECT  7522.5 159527.5 7587.5 159152.5 ;
      RECT  7902.5 159527.5 7967.5 159152.5 ;
      RECT  8262.5 159370.0 8327.5 159185.0 ;
      RECT  8262.5 160530.0 8327.5 160345.0 ;
      RECT  7522.5 159527.5 7587.5 159392.5 ;
      RECT  7712.5 159527.5 7777.5 159392.5 ;
      RECT  7712.5 159527.5 7777.5 159392.5 ;
      RECT  7522.5 159527.5 7587.5 159392.5 ;
      RECT  7712.5 159527.5 7777.5 159392.5 ;
      RECT  7902.5 159527.5 7967.5 159392.5 ;
      RECT  7902.5 159527.5 7967.5 159392.5 ;
      RECT  7712.5 159527.5 7777.5 159392.5 ;
      RECT  7902.5 159527.5 7967.5 159392.5 ;
      RECT  8092.5 159527.5 8157.5 159392.5 ;
      RECT  8092.5 159527.5 8157.5 159392.5 ;
      RECT  7902.5 159527.5 7967.5 159392.5 ;
      RECT  7522.5 160367.5 7587.5 160232.5 ;
      RECT  7712.5 160367.5 7777.5 160232.5 ;
      RECT  7712.5 160367.5 7777.5 160232.5 ;
      RECT  7522.5 160367.5 7587.5 160232.5 ;
      RECT  7712.5 160367.5 7777.5 160232.5 ;
      RECT  7902.5 160367.5 7967.5 160232.5 ;
      RECT  7902.5 160367.5 7967.5 160232.5 ;
      RECT  7712.5 160367.5 7777.5 160232.5 ;
      RECT  7902.5 160367.5 7967.5 160232.5 ;
      RECT  8092.5 160367.5 8157.5 160232.5 ;
      RECT  8092.5 160367.5 8157.5 160232.5 ;
      RECT  7902.5 160367.5 7967.5 160232.5 ;
      RECT  8262.5 159437.5 8327.5 159302.5 ;
      RECT  8262.5 160412.5 8327.5 160277.5 ;
      RECT  8097.5 160155.0 7962.5 160090.0 ;
      RECT  7907.5 160015.0 7772.5 159950.0 ;
      RECT  7717.5 159875.0 7582.5 159810.0 ;
      RECT  7712.5 159527.5 7777.5 159392.5 ;
      RECT  8092.5 159527.5 8157.5 159392.5 ;
      RECT  8092.5 160367.5 8157.5 160232.5 ;
      RECT  8092.5 159910.0 8157.5 159775.0 ;
      RECT  7582.5 159875.0 7717.5 159810.0 ;
      RECT  7772.5 160015.0 7907.5 159950.0 ;
      RECT  7962.5 160155.0 8097.5 160090.0 ;
      RECT  8092.5 159910.0 8157.5 159775.0 ;
      RECT  7455.0 159217.5 8465.0 159152.5 ;
      RECT  7455.0 160562.5 8465.0 160497.5 ;
      RECT  7522.5 160692.5 7587.5 160497.5 ;
      RECT  7522.5 161532.5 7587.5 161907.5 ;
      RECT  7902.5 161532.5 7967.5 161907.5 ;
      RECT  8262.5 161690.0 8327.5 161875.0 ;
      RECT  8262.5 160530.0 8327.5 160715.0 ;
      RECT  7522.5 161532.5 7587.5 161667.5 ;
      RECT  7712.5 161532.5 7777.5 161667.5 ;
      RECT  7712.5 161532.5 7777.5 161667.5 ;
      RECT  7522.5 161532.5 7587.5 161667.5 ;
      RECT  7712.5 161532.5 7777.5 161667.5 ;
      RECT  7902.5 161532.5 7967.5 161667.5 ;
      RECT  7902.5 161532.5 7967.5 161667.5 ;
      RECT  7712.5 161532.5 7777.5 161667.5 ;
      RECT  7902.5 161532.5 7967.5 161667.5 ;
      RECT  8092.5 161532.5 8157.5 161667.5 ;
      RECT  8092.5 161532.5 8157.5 161667.5 ;
      RECT  7902.5 161532.5 7967.5 161667.5 ;
      RECT  7522.5 160692.5 7587.5 160827.5 ;
      RECT  7712.5 160692.5 7777.5 160827.5 ;
      RECT  7712.5 160692.5 7777.5 160827.5 ;
      RECT  7522.5 160692.5 7587.5 160827.5 ;
      RECT  7712.5 160692.5 7777.5 160827.5 ;
      RECT  7902.5 160692.5 7967.5 160827.5 ;
      RECT  7902.5 160692.5 7967.5 160827.5 ;
      RECT  7712.5 160692.5 7777.5 160827.5 ;
      RECT  7902.5 160692.5 7967.5 160827.5 ;
      RECT  8092.5 160692.5 8157.5 160827.5 ;
      RECT  8092.5 160692.5 8157.5 160827.5 ;
      RECT  7902.5 160692.5 7967.5 160827.5 ;
      RECT  8262.5 161622.5 8327.5 161757.5 ;
      RECT  8262.5 160647.5 8327.5 160782.5 ;
      RECT  8097.5 160905.0 7962.5 160970.0 ;
      RECT  7907.5 161045.0 7772.5 161110.0 ;
      RECT  7717.5 161185.0 7582.5 161250.0 ;
      RECT  7712.5 161532.5 7777.5 161667.5 ;
      RECT  8092.5 161532.5 8157.5 161667.5 ;
      RECT  8092.5 160692.5 8157.5 160827.5 ;
      RECT  8092.5 161150.0 8157.5 161285.0 ;
      RECT  7582.5 161185.0 7717.5 161250.0 ;
      RECT  7772.5 161045.0 7907.5 161110.0 ;
      RECT  7962.5 160905.0 8097.5 160970.0 ;
      RECT  8092.5 161150.0 8157.5 161285.0 ;
      RECT  7455.0 161842.5 8465.0 161907.5 ;
      RECT  7455.0 160497.5 8465.0 160562.5 ;
      RECT  7522.5 163057.5 7587.5 163252.5 ;
      RECT  7522.5 162217.5 7587.5 161842.5 ;
      RECT  7902.5 162217.5 7967.5 161842.5 ;
      RECT  8262.5 162060.0 8327.5 161875.0 ;
      RECT  8262.5 163220.0 8327.5 163035.0 ;
      RECT  7522.5 162217.5 7587.5 162082.5 ;
      RECT  7712.5 162217.5 7777.5 162082.5 ;
      RECT  7712.5 162217.5 7777.5 162082.5 ;
      RECT  7522.5 162217.5 7587.5 162082.5 ;
      RECT  7712.5 162217.5 7777.5 162082.5 ;
      RECT  7902.5 162217.5 7967.5 162082.5 ;
      RECT  7902.5 162217.5 7967.5 162082.5 ;
      RECT  7712.5 162217.5 7777.5 162082.5 ;
      RECT  7902.5 162217.5 7967.5 162082.5 ;
      RECT  8092.5 162217.5 8157.5 162082.5 ;
      RECT  8092.5 162217.5 8157.5 162082.5 ;
      RECT  7902.5 162217.5 7967.5 162082.5 ;
      RECT  7522.5 163057.5 7587.5 162922.5 ;
      RECT  7712.5 163057.5 7777.5 162922.5 ;
      RECT  7712.5 163057.5 7777.5 162922.5 ;
      RECT  7522.5 163057.5 7587.5 162922.5 ;
      RECT  7712.5 163057.5 7777.5 162922.5 ;
      RECT  7902.5 163057.5 7967.5 162922.5 ;
      RECT  7902.5 163057.5 7967.5 162922.5 ;
      RECT  7712.5 163057.5 7777.5 162922.5 ;
      RECT  7902.5 163057.5 7967.5 162922.5 ;
      RECT  8092.5 163057.5 8157.5 162922.5 ;
      RECT  8092.5 163057.5 8157.5 162922.5 ;
      RECT  7902.5 163057.5 7967.5 162922.5 ;
      RECT  8262.5 162127.5 8327.5 161992.5 ;
      RECT  8262.5 163102.5 8327.5 162967.5 ;
      RECT  8097.5 162845.0 7962.5 162780.0 ;
      RECT  7907.5 162705.0 7772.5 162640.0 ;
      RECT  7717.5 162565.0 7582.5 162500.0 ;
      RECT  7712.5 162217.5 7777.5 162082.5 ;
      RECT  8092.5 162217.5 8157.5 162082.5 ;
      RECT  8092.5 163057.5 8157.5 162922.5 ;
      RECT  8092.5 162600.0 8157.5 162465.0 ;
      RECT  7582.5 162565.0 7717.5 162500.0 ;
      RECT  7772.5 162705.0 7907.5 162640.0 ;
      RECT  7962.5 162845.0 8097.5 162780.0 ;
      RECT  8092.5 162600.0 8157.5 162465.0 ;
      RECT  7455.0 161907.5 8465.0 161842.5 ;
      RECT  7455.0 163252.5 8465.0 163187.5 ;
      RECT  7522.5 163382.5 7587.5 163187.5 ;
      RECT  7522.5 164222.5 7587.5 164597.5 ;
      RECT  7902.5 164222.5 7967.5 164597.5 ;
      RECT  8262.5 164380.0 8327.5 164565.0 ;
      RECT  8262.5 163220.0 8327.5 163405.0 ;
      RECT  7522.5 164222.5 7587.5 164357.5 ;
      RECT  7712.5 164222.5 7777.5 164357.5 ;
      RECT  7712.5 164222.5 7777.5 164357.5 ;
      RECT  7522.5 164222.5 7587.5 164357.5 ;
      RECT  7712.5 164222.5 7777.5 164357.5 ;
      RECT  7902.5 164222.5 7967.5 164357.5 ;
      RECT  7902.5 164222.5 7967.5 164357.5 ;
      RECT  7712.5 164222.5 7777.5 164357.5 ;
      RECT  7902.5 164222.5 7967.5 164357.5 ;
      RECT  8092.5 164222.5 8157.5 164357.5 ;
      RECT  8092.5 164222.5 8157.5 164357.5 ;
      RECT  7902.5 164222.5 7967.5 164357.5 ;
      RECT  7522.5 163382.5 7587.5 163517.5 ;
      RECT  7712.5 163382.5 7777.5 163517.5 ;
      RECT  7712.5 163382.5 7777.5 163517.5 ;
      RECT  7522.5 163382.5 7587.5 163517.5 ;
      RECT  7712.5 163382.5 7777.5 163517.5 ;
      RECT  7902.5 163382.5 7967.5 163517.5 ;
      RECT  7902.5 163382.5 7967.5 163517.5 ;
      RECT  7712.5 163382.5 7777.5 163517.5 ;
      RECT  7902.5 163382.5 7967.5 163517.5 ;
      RECT  8092.5 163382.5 8157.5 163517.5 ;
      RECT  8092.5 163382.5 8157.5 163517.5 ;
      RECT  7902.5 163382.5 7967.5 163517.5 ;
      RECT  8262.5 164312.5 8327.5 164447.5 ;
      RECT  8262.5 163337.5 8327.5 163472.5 ;
      RECT  8097.5 163595.0 7962.5 163660.0 ;
      RECT  7907.5 163735.0 7772.5 163800.0 ;
      RECT  7717.5 163875.0 7582.5 163940.0 ;
      RECT  7712.5 164222.5 7777.5 164357.5 ;
      RECT  8092.5 164222.5 8157.5 164357.5 ;
      RECT  8092.5 163382.5 8157.5 163517.5 ;
      RECT  8092.5 163840.0 8157.5 163975.0 ;
      RECT  7582.5 163875.0 7717.5 163940.0 ;
      RECT  7772.5 163735.0 7907.5 163800.0 ;
      RECT  7962.5 163595.0 8097.5 163660.0 ;
      RECT  8092.5 163840.0 8157.5 163975.0 ;
      RECT  7455.0 164532.5 8465.0 164597.5 ;
      RECT  7455.0 163187.5 8465.0 163252.5 ;
      RECT  7522.5 165747.5 7587.5 165942.5 ;
      RECT  7522.5 164907.5 7587.5 164532.5 ;
      RECT  7902.5 164907.5 7967.5 164532.5 ;
      RECT  8262.5 164750.0 8327.5 164565.0 ;
      RECT  8262.5 165910.0 8327.5 165725.0 ;
      RECT  7522.5 164907.5 7587.5 164772.5 ;
      RECT  7712.5 164907.5 7777.5 164772.5 ;
      RECT  7712.5 164907.5 7777.5 164772.5 ;
      RECT  7522.5 164907.5 7587.5 164772.5 ;
      RECT  7712.5 164907.5 7777.5 164772.5 ;
      RECT  7902.5 164907.5 7967.5 164772.5 ;
      RECT  7902.5 164907.5 7967.5 164772.5 ;
      RECT  7712.5 164907.5 7777.5 164772.5 ;
      RECT  7902.5 164907.5 7967.5 164772.5 ;
      RECT  8092.5 164907.5 8157.5 164772.5 ;
      RECT  8092.5 164907.5 8157.5 164772.5 ;
      RECT  7902.5 164907.5 7967.5 164772.5 ;
      RECT  7522.5 165747.5 7587.5 165612.5 ;
      RECT  7712.5 165747.5 7777.5 165612.5 ;
      RECT  7712.5 165747.5 7777.5 165612.5 ;
      RECT  7522.5 165747.5 7587.5 165612.5 ;
      RECT  7712.5 165747.5 7777.5 165612.5 ;
      RECT  7902.5 165747.5 7967.5 165612.5 ;
      RECT  7902.5 165747.5 7967.5 165612.5 ;
      RECT  7712.5 165747.5 7777.5 165612.5 ;
      RECT  7902.5 165747.5 7967.5 165612.5 ;
      RECT  8092.5 165747.5 8157.5 165612.5 ;
      RECT  8092.5 165747.5 8157.5 165612.5 ;
      RECT  7902.5 165747.5 7967.5 165612.5 ;
      RECT  8262.5 164817.5 8327.5 164682.5 ;
      RECT  8262.5 165792.5 8327.5 165657.5 ;
      RECT  8097.5 165535.0 7962.5 165470.0 ;
      RECT  7907.5 165395.0 7772.5 165330.0 ;
      RECT  7717.5 165255.0 7582.5 165190.0 ;
      RECT  7712.5 164907.5 7777.5 164772.5 ;
      RECT  8092.5 164907.5 8157.5 164772.5 ;
      RECT  8092.5 165747.5 8157.5 165612.5 ;
      RECT  8092.5 165290.0 8157.5 165155.0 ;
      RECT  7582.5 165255.0 7717.5 165190.0 ;
      RECT  7772.5 165395.0 7907.5 165330.0 ;
      RECT  7962.5 165535.0 8097.5 165470.0 ;
      RECT  8092.5 165290.0 8157.5 165155.0 ;
      RECT  7455.0 164597.5 8465.0 164532.5 ;
      RECT  7455.0 165942.5 8465.0 165877.5 ;
      RECT  7522.5 166072.5 7587.5 165877.5 ;
      RECT  7522.5 166912.5 7587.5 167287.5 ;
      RECT  7902.5 166912.5 7967.5 167287.5 ;
      RECT  8262.5 167070.0 8327.5 167255.0 ;
      RECT  8262.5 165910.0 8327.5 166095.0 ;
      RECT  7522.5 166912.5 7587.5 167047.5 ;
      RECT  7712.5 166912.5 7777.5 167047.5 ;
      RECT  7712.5 166912.5 7777.5 167047.5 ;
      RECT  7522.5 166912.5 7587.5 167047.5 ;
      RECT  7712.5 166912.5 7777.5 167047.5 ;
      RECT  7902.5 166912.5 7967.5 167047.5 ;
      RECT  7902.5 166912.5 7967.5 167047.5 ;
      RECT  7712.5 166912.5 7777.5 167047.5 ;
      RECT  7902.5 166912.5 7967.5 167047.5 ;
      RECT  8092.5 166912.5 8157.5 167047.5 ;
      RECT  8092.5 166912.5 8157.5 167047.5 ;
      RECT  7902.5 166912.5 7967.5 167047.5 ;
      RECT  7522.5 166072.5 7587.5 166207.5 ;
      RECT  7712.5 166072.5 7777.5 166207.5 ;
      RECT  7712.5 166072.5 7777.5 166207.5 ;
      RECT  7522.5 166072.5 7587.5 166207.5 ;
      RECT  7712.5 166072.5 7777.5 166207.5 ;
      RECT  7902.5 166072.5 7967.5 166207.5 ;
      RECT  7902.5 166072.5 7967.5 166207.5 ;
      RECT  7712.5 166072.5 7777.5 166207.5 ;
      RECT  7902.5 166072.5 7967.5 166207.5 ;
      RECT  8092.5 166072.5 8157.5 166207.5 ;
      RECT  8092.5 166072.5 8157.5 166207.5 ;
      RECT  7902.5 166072.5 7967.5 166207.5 ;
      RECT  8262.5 167002.5 8327.5 167137.5 ;
      RECT  8262.5 166027.5 8327.5 166162.5 ;
      RECT  8097.5 166285.0 7962.5 166350.0 ;
      RECT  7907.5 166425.0 7772.5 166490.0 ;
      RECT  7717.5 166565.0 7582.5 166630.0 ;
      RECT  7712.5 166912.5 7777.5 167047.5 ;
      RECT  8092.5 166912.5 8157.5 167047.5 ;
      RECT  8092.5 166072.5 8157.5 166207.5 ;
      RECT  8092.5 166530.0 8157.5 166665.0 ;
      RECT  7582.5 166565.0 7717.5 166630.0 ;
      RECT  7772.5 166425.0 7907.5 166490.0 ;
      RECT  7962.5 166285.0 8097.5 166350.0 ;
      RECT  8092.5 166530.0 8157.5 166665.0 ;
      RECT  7455.0 167222.5 8465.0 167287.5 ;
      RECT  7455.0 165877.5 8465.0 165942.5 ;
      RECT  7522.5 168437.5 7587.5 168632.5 ;
      RECT  7522.5 167597.5 7587.5 167222.5 ;
      RECT  7902.5 167597.5 7967.5 167222.5 ;
      RECT  8262.5 167440.0 8327.5 167255.0 ;
      RECT  8262.5 168600.0 8327.5 168415.0 ;
      RECT  7522.5 167597.5 7587.5 167462.5 ;
      RECT  7712.5 167597.5 7777.5 167462.5 ;
      RECT  7712.5 167597.5 7777.5 167462.5 ;
      RECT  7522.5 167597.5 7587.5 167462.5 ;
      RECT  7712.5 167597.5 7777.5 167462.5 ;
      RECT  7902.5 167597.5 7967.5 167462.5 ;
      RECT  7902.5 167597.5 7967.5 167462.5 ;
      RECT  7712.5 167597.5 7777.5 167462.5 ;
      RECT  7902.5 167597.5 7967.5 167462.5 ;
      RECT  8092.5 167597.5 8157.5 167462.5 ;
      RECT  8092.5 167597.5 8157.5 167462.5 ;
      RECT  7902.5 167597.5 7967.5 167462.5 ;
      RECT  7522.5 168437.5 7587.5 168302.5 ;
      RECT  7712.5 168437.5 7777.5 168302.5 ;
      RECT  7712.5 168437.5 7777.5 168302.5 ;
      RECT  7522.5 168437.5 7587.5 168302.5 ;
      RECT  7712.5 168437.5 7777.5 168302.5 ;
      RECT  7902.5 168437.5 7967.5 168302.5 ;
      RECT  7902.5 168437.5 7967.5 168302.5 ;
      RECT  7712.5 168437.5 7777.5 168302.5 ;
      RECT  7902.5 168437.5 7967.5 168302.5 ;
      RECT  8092.5 168437.5 8157.5 168302.5 ;
      RECT  8092.5 168437.5 8157.5 168302.5 ;
      RECT  7902.5 168437.5 7967.5 168302.5 ;
      RECT  8262.5 167507.5 8327.5 167372.5 ;
      RECT  8262.5 168482.5 8327.5 168347.5 ;
      RECT  8097.5 168225.0 7962.5 168160.0 ;
      RECT  7907.5 168085.0 7772.5 168020.0 ;
      RECT  7717.5 167945.0 7582.5 167880.0 ;
      RECT  7712.5 167597.5 7777.5 167462.5 ;
      RECT  8092.5 167597.5 8157.5 167462.5 ;
      RECT  8092.5 168437.5 8157.5 168302.5 ;
      RECT  8092.5 167980.0 8157.5 167845.0 ;
      RECT  7582.5 167945.0 7717.5 167880.0 ;
      RECT  7772.5 168085.0 7907.5 168020.0 ;
      RECT  7962.5 168225.0 8097.5 168160.0 ;
      RECT  8092.5 167980.0 8157.5 167845.0 ;
      RECT  7455.0 167287.5 8465.0 167222.5 ;
      RECT  7455.0 168632.5 8465.0 168567.5 ;
      RECT  7522.5 168762.5 7587.5 168567.5 ;
      RECT  7522.5 169602.5 7587.5 169977.5 ;
      RECT  7902.5 169602.5 7967.5 169977.5 ;
      RECT  8262.5 169760.0 8327.5 169945.0 ;
      RECT  8262.5 168600.0 8327.5 168785.0 ;
      RECT  7522.5 169602.5 7587.5 169737.5 ;
      RECT  7712.5 169602.5 7777.5 169737.5 ;
      RECT  7712.5 169602.5 7777.5 169737.5 ;
      RECT  7522.5 169602.5 7587.5 169737.5 ;
      RECT  7712.5 169602.5 7777.5 169737.5 ;
      RECT  7902.5 169602.5 7967.5 169737.5 ;
      RECT  7902.5 169602.5 7967.5 169737.5 ;
      RECT  7712.5 169602.5 7777.5 169737.5 ;
      RECT  7902.5 169602.5 7967.5 169737.5 ;
      RECT  8092.5 169602.5 8157.5 169737.5 ;
      RECT  8092.5 169602.5 8157.5 169737.5 ;
      RECT  7902.5 169602.5 7967.5 169737.5 ;
      RECT  7522.5 168762.5 7587.5 168897.5 ;
      RECT  7712.5 168762.5 7777.5 168897.5 ;
      RECT  7712.5 168762.5 7777.5 168897.5 ;
      RECT  7522.5 168762.5 7587.5 168897.5 ;
      RECT  7712.5 168762.5 7777.5 168897.5 ;
      RECT  7902.5 168762.5 7967.5 168897.5 ;
      RECT  7902.5 168762.5 7967.5 168897.5 ;
      RECT  7712.5 168762.5 7777.5 168897.5 ;
      RECT  7902.5 168762.5 7967.5 168897.5 ;
      RECT  8092.5 168762.5 8157.5 168897.5 ;
      RECT  8092.5 168762.5 8157.5 168897.5 ;
      RECT  7902.5 168762.5 7967.5 168897.5 ;
      RECT  8262.5 169692.5 8327.5 169827.5 ;
      RECT  8262.5 168717.5 8327.5 168852.5 ;
      RECT  8097.5 168975.0 7962.5 169040.0 ;
      RECT  7907.5 169115.0 7772.5 169180.0 ;
      RECT  7717.5 169255.0 7582.5 169320.0 ;
      RECT  7712.5 169602.5 7777.5 169737.5 ;
      RECT  8092.5 169602.5 8157.5 169737.5 ;
      RECT  8092.5 168762.5 8157.5 168897.5 ;
      RECT  8092.5 169220.0 8157.5 169355.0 ;
      RECT  7582.5 169255.0 7717.5 169320.0 ;
      RECT  7772.5 169115.0 7907.5 169180.0 ;
      RECT  7962.5 168975.0 8097.5 169040.0 ;
      RECT  8092.5 169220.0 8157.5 169355.0 ;
      RECT  7455.0 169912.5 8465.0 169977.5 ;
      RECT  7455.0 168567.5 8465.0 168632.5 ;
      RECT  7522.5 171127.5 7587.5 171322.5 ;
      RECT  7522.5 170287.5 7587.5 169912.5 ;
      RECT  7902.5 170287.5 7967.5 169912.5 ;
      RECT  8262.5 170130.0 8327.5 169945.0 ;
      RECT  8262.5 171290.0 8327.5 171105.0 ;
      RECT  7522.5 170287.5 7587.5 170152.5 ;
      RECT  7712.5 170287.5 7777.5 170152.5 ;
      RECT  7712.5 170287.5 7777.5 170152.5 ;
      RECT  7522.5 170287.5 7587.5 170152.5 ;
      RECT  7712.5 170287.5 7777.5 170152.5 ;
      RECT  7902.5 170287.5 7967.5 170152.5 ;
      RECT  7902.5 170287.5 7967.5 170152.5 ;
      RECT  7712.5 170287.5 7777.5 170152.5 ;
      RECT  7902.5 170287.5 7967.5 170152.5 ;
      RECT  8092.5 170287.5 8157.5 170152.5 ;
      RECT  8092.5 170287.5 8157.5 170152.5 ;
      RECT  7902.5 170287.5 7967.5 170152.5 ;
      RECT  7522.5 171127.5 7587.5 170992.5 ;
      RECT  7712.5 171127.5 7777.5 170992.5 ;
      RECT  7712.5 171127.5 7777.5 170992.5 ;
      RECT  7522.5 171127.5 7587.5 170992.5 ;
      RECT  7712.5 171127.5 7777.5 170992.5 ;
      RECT  7902.5 171127.5 7967.5 170992.5 ;
      RECT  7902.5 171127.5 7967.5 170992.5 ;
      RECT  7712.5 171127.5 7777.5 170992.5 ;
      RECT  7902.5 171127.5 7967.5 170992.5 ;
      RECT  8092.5 171127.5 8157.5 170992.5 ;
      RECT  8092.5 171127.5 8157.5 170992.5 ;
      RECT  7902.5 171127.5 7967.5 170992.5 ;
      RECT  8262.5 170197.5 8327.5 170062.5 ;
      RECT  8262.5 171172.5 8327.5 171037.5 ;
      RECT  8097.5 170915.0 7962.5 170850.0 ;
      RECT  7907.5 170775.0 7772.5 170710.0 ;
      RECT  7717.5 170635.0 7582.5 170570.0 ;
      RECT  7712.5 170287.5 7777.5 170152.5 ;
      RECT  8092.5 170287.5 8157.5 170152.5 ;
      RECT  8092.5 171127.5 8157.5 170992.5 ;
      RECT  8092.5 170670.0 8157.5 170535.0 ;
      RECT  7582.5 170635.0 7717.5 170570.0 ;
      RECT  7772.5 170775.0 7907.5 170710.0 ;
      RECT  7962.5 170915.0 8097.5 170850.0 ;
      RECT  8092.5 170670.0 8157.5 170535.0 ;
      RECT  7455.0 169977.5 8465.0 169912.5 ;
      RECT  7455.0 171322.5 8465.0 171257.5 ;
      RECT  7522.5 171452.5 7587.5 171257.5 ;
      RECT  7522.5 172292.5 7587.5 172667.5 ;
      RECT  7902.5 172292.5 7967.5 172667.5 ;
      RECT  8262.5 172450.0 8327.5 172635.0 ;
      RECT  8262.5 171290.0 8327.5 171475.0 ;
      RECT  7522.5 172292.5 7587.5 172427.5 ;
      RECT  7712.5 172292.5 7777.5 172427.5 ;
      RECT  7712.5 172292.5 7777.5 172427.5 ;
      RECT  7522.5 172292.5 7587.5 172427.5 ;
      RECT  7712.5 172292.5 7777.5 172427.5 ;
      RECT  7902.5 172292.5 7967.5 172427.5 ;
      RECT  7902.5 172292.5 7967.5 172427.5 ;
      RECT  7712.5 172292.5 7777.5 172427.5 ;
      RECT  7902.5 172292.5 7967.5 172427.5 ;
      RECT  8092.5 172292.5 8157.5 172427.5 ;
      RECT  8092.5 172292.5 8157.5 172427.5 ;
      RECT  7902.5 172292.5 7967.5 172427.5 ;
      RECT  7522.5 171452.5 7587.5 171587.5 ;
      RECT  7712.5 171452.5 7777.5 171587.5 ;
      RECT  7712.5 171452.5 7777.5 171587.5 ;
      RECT  7522.5 171452.5 7587.5 171587.5 ;
      RECT  7712.5 171452.5 7777.5 171587.5 ;
      RECT  7902.5 171452.5 7967.5 171587.5 ;
      RECT  7902.5 171452.5 7967.5 171587.5 ;
      RECT  7712.5 171452.5 7777.5 171587.5 ;
      RECT  7902.5 171452.5 7967.5 171587.5 ;
      RECT  8092.5 171452.5 8157.5 171587.5 ;
      RECT  8092.5 171452.5 8157.5 171587.5 ;
      RECT  7902.5 171452.5 7967.5 171587.5 ;
      RECT  8262.5 172382.5 8327.5 172517.5 ;
      RECT  8262.5 171407.5 8327.5 171542.5 ;
      RECT  8097.5 171665.0 7962.5 171730.0 ;
      RECT  7907.5 171805.0 7772.5 171870.0 ;
      RECT  7717.5 171945.0 7582.5 172010.0 ;
      RECT  7712.5 172292.5 7777.5 172427.5 ;
      RECT  8092.5 172292.5 8157.5 172427.5 ;
      RECT  8092.5 171452.5 8157.5 171587.5 ;
      RECT  8092.5 171910.0 8157.5 172045.0 ;
      RECT  7582.5 171945.0 7717.5 172010.0 ;
      RECT  7772.5 171805.0 7907.5 171870.0 ;
      RECT  7962.5 171665.0 8097.5 171730.0 ;
      RECT  8092.5 171910.0 8157.5 172045.0 ;
      RECT  7455.0 172602.5 8465.0 172667.5 ;
      RECT  7455.0 171257.5 8465.0 171322.5 ;
      RECT  7522.5 173817.5 7587.5 174012.5 ;
      RECT  7522.5 172977.5 7587.5 172602.5 ;
      RECT  7902.5 172977.5 7967.5 172602.5 ;
      RECT  8262.5 172820.0 8327.5 172635.0 ;
      RECT  8262.5 173980.0 8327.5 173795.0 ;
      RECT  7522.5 172977.5 7587.5 172842.5 ;
      RECT  7712.5 172977.5 7777.5 172842.5 ;
      RECT  7712.5 172977.5 7777.5 172842.5 ;
      RECT  7522.5 172977.5 7587.5 172842.5 ;
      RECT  7712.5 172977.5 7777.5 172842.5 ;
      RECT  7902.5 172977.5 7967.5 172842.5 ;
      RECT  7902.5 172977.5 7967.5 172842.5 ;
      RECT  7712.5 172977.5 7777.5 172842.5 ;
      RECT  7902.5 172977.5 7967.5 172842.5 ;
      RECT  8092.5 172977.5 8157.5 172842.5 ;
      RECT  8092.5 172977.5 8157.5 172842.5 ;
      RECT  7902.5 172977.5 7967.5 172842.5 ;
      RECT  7522.5 173817.5 7587.5 173682.5 ;
      RECT  7712.5 173817.5 7777.5 173682.5 ;
      RECT  7712.5 173817.5 7777.5 173682.5 ;
      RECT  7522.5 173817.5 7587.5 173682.5 ;
      RECT  7712.5 173817.5 7777.5 173682.5 ;
      RECT  7902.5 173817.5 7967.5 173682.5 ;
      RECT  7902.5 173817.5 7967.5 173682.5 ;
      RECT  7712.5 173817.5 7777.5 173682.5 ;
      RECT  7902.5 173817.5 7967.5 173682.5 ;
      RECT  8092.5 173817.5 8157.5 173682.5 ;
      RECT  8092.5 173817.5 8157.5 173682.5 ;
      RECT  7902.5 173817.5 7967.5 173682.5 ;
      RECT  8262.5 172887.5 8327.5 172752.5 ;
      RECT  8262.5 173862.5 8327.5 173727.5 ;
      RECT  8097.5 173605.0 7962.5 173540.0 ;
      RECT  7907.5 173465.0 7772.5 173400.0 ;
      RECT  7717.5 173325.0 7582.5 173260.0 ;
      RECT  7712.5 172977.5 7777.5 172842.5 ;
      RECT  8092.5 172977.5 8157.5 172842.5 ;
      RECT  8092.5 173817.5 8157.5 173682.5 ;
      RECT  8092.5 173360.0 8157.5 173225.0 ;
      RECT  7582.5 173325.0 7717.5 173260.0 ;
      RECT  7772.5 173465.0 7907.5 173400.0 ;
      RECT  7962.5 173605.0 8097.5 173540.0 ;
      RECT  8092.5 173360.0 8157.5 173225.0 ;
      RECT  7455.0 172667.5 8465.0 172602.5 ;
      RECT  7455.0 174012.5 8465.0 173947.5 ;
      RECT  7522.5 174142.5 7587.5 173947.5 ;
      RECT  7522.5 174982.5 7587.5 175357.5 ;
      RECT  7902.5 174982.5 7967.5 175357.5 ;
      RECT  8262.5 175140.0 8327.5 175325.0 ;
      RECT  8262.5 173980.0 8327.5 174165.0 ;
      RECT  7522.5 174982.5 7587.5 175117.5 ;
      RECT  7712.5 174982.5 7777.5 175117.5 ;
      RECT  7712.5 174982.5 7777.5 175117.5 ;
      RECT  7522.5 174982.5 7587.5 175117.5 ;
      RECT  7712.5 174982.5 7777.5 175117.5 ;
      RECT  7902.5 174982.5 7967.5 175117.5 ;
      RECT  7902.5 174982.5 7967.5 175117.5 ;
      RECT  7712.5 174982.5 7777.5 175117.5 ;
      RECT  7902.5 174982.5 7967.5 175117.5 ;
      RECT  8092.5 174982.5 8157.5 175117.5 ;
      RECT  8092.5 174982.5 8157.5 175117.5 ;
      RECT  7902.5 174982.5 7967.5 175117.5 ;
      RECT  7522.5 174142.5 7587.5 174277.5 ;
      RECT  7712.5 174142.5 7777.5 174277.5 ;
      RECT  7712.5 174142.5 7777.5 174277.5 ;
      RECT  7522.5 174142.5 7587.5 174277.5 ;
      RECT  7712.5 174142.5 7777.5 174277.5 ;
      RECT  7902.5 174142.5 7967.5 174277.5 ;
      RECT  7902.5 174142.5 7967.5 174277.5 ;
      RECT  7712.5 174142.5 7777.5 174277.5 ;
      RECT  7902.5 174142.5 7967.5 174277.5 ;
      RECT  8092.5 174142.5 8157.5 174277.5 ;
      RECT  8092.5 174142.5 8157.5 174277.5 ;
      RECT  7902.5 174142.5 7967.5 174277.5 ;
      RECT  8262.5 175072.5 8327.5 175207.5 ;
      RECT  8262.5 174097.5 8327.5 174232.5 ;
      RECT  8097.5 174355.0 7962.5 174420.0 ;
      RECT  7907.5 174495.0 7772.5 174560.0 ;
      RECT  7717.5 174635.0 7582.5 174700.0 ;
      RECT  7712.5 174982.5 7777.5 175117.5 ;
      RECT  8092.5 174982.5 8157.5 175117.5 ;
      RECT  8092.5 174142.5 8157.5 174277.5 ;
      RECT  8092.5 174600.0 8157.5 174735.0 ;
      RECT  7582.5 174635.0 7717.5 174700.0 ;
      RECT  7772.5 174495.0 7907.5 174560.0 ;
      RECT  7962.5 174355.0 8097.5 174420.0 ;
      RECT  8092.5 174600.0 8157.5 174735.0 ;
      RECT  7455.0 175292.5 8465.0 175357.5 ;
      RECT  7455.0 173947.5 8465.0 174012.5 ;
      RECT  7522.5 176507.5 7587.5 176702.5 ;
      RECT  7522.5 175667.5 7587.5 175292.5 ;
      RECT  7902.5 175667.5 7967.5 175292.5 ;
      RECT  8262.5 175510.0 8327.5 175325.0 ;
      RECT  8262.5 176670.0 8327.5 176485.0 ;
      RECT  7522.5 175667.5 7587.5 175532.5 ;
      RECT  7712.5 175667.5 7777.5 175532.5 ;
      RECT  7712.5 175667.5 7777.5 175532.5 ;
      RECT  7522.5 175667.5 7587.5 175532.5 ;
      RECT  7712.5 175667.5 7777.5 175532.5 ;
      RECT  7902.5 175667.5 7967.5 175532.5 ;
      RECT  7902.5 175667.5 7967.5 175532.5 ;
      RECT  7712.5 175667.5 7777.5 175532.5 ;
      RECT  7902.5 175667.5 7967.5 175532.5 ;
      RECT  8092.5 175667.5 8157.5 175532.5 ;
      RECT  8092.5 175667.5 8157.5 175532.5 ;
      RECT  7902.5 175667.5 7967.5 175532.5 ;
      RECT  7522.5 176507.5 7587.5 176372.5 ;
      RECT  7712.5 176507.5 7777.5 176372.5 ;
      RECT  7712.5 176507.5 7777.5 176372.5 ;
      RECT  7522.5 176507.5 7587.5 176372.5 ;
      RECT  7712.5 176507.5 7777.5 176372.5 ;
      RECT  7902.5 176507.5 7967.5 176372.5 ;
      RECT  7902.5 176507.5 7967.5 176372.5 ;
      RECT  7712.5 176507.5 7777.5 176372.5 ;
      RECT  7902.5 176507.5 7967.5 176372.5 ;
      RECT  8092.5 176507.5 8157.5 176372.5 ;
      RECT  8092.5 176507.5 8157.5 176372.5 ;
      RECT  7902.5 176507.5 7967.5 176372.5 ;
      RECT  8262.5 175577.5 8327.5 175442.5 ;
      RECT  8262.5 176552.5 8327.5 176417.5 ;
      RECT  8097.5 176295.0 7962.5 176230.0 ;
      RECT  7907.5 176155.0 7772.5 176090.0 ;
      RECT  7717.5 176015.0 7582.5 175950.0 ;
      RECT  7712.5 175667.5 7777.5 175532.5 ;
      RECT  8092.5 175667.5 8157.5 175532.5 ;
      RECT  8092.5 176507.5 8157.5 176372.5 ;
      RECT  8092.5 176050.0 8157.5 175915.0 ;
      RECT  7582.5 176015.0 7717.5 175950.0 ;
      RECT  7772.5 176155.0 7907.5 176090.0 ;
      RECT  7962.5 176295.0 8097.5 176230.0 ;
      RECT  8092.5 176050.0 8157.5 175915.0 ;
      RECT  7455.0 175357.5 8465.0 175292.5 ;
      RECT  7455.0 176702.5 8465.0 176637.5 ;
      RECT  7522.5 176832.5 7587.5 176637.5 ;
      RECT  7522.5 177672.5 7587.5 178047.5 ;
      RECT  7902.5 177672.5 7967.5 178047.5 ;
      RECT  8262.5 177830.0 8327.5 178015.0 ;
      RECT  8262.5 176670.0 8327.5 176855.0 ;
      RECT  7522.5 177672.5 7587.5 177807.5 ;
      RECT  7712.5 177672.5 7777.5 177807.5 ;
      RECT  7712.5 177672.5 7777.5 177807.5 ;
      RECT  7522.5 177672.5 7587.5 177807.5 ;
      RECT  7712.5 177672.5 7777.5 177807.5 ;
      RECT  7902.5 177672.5 7967.5 177807.5 ;
      RECT  7902.5 177672.5 7967.5 177807.5 ;
      RECT  7712.5 177672.5 7777.5 177807.5 ;
      RECT  7902.5 177672.5 7967.5 177807.5 ;
      RECT  8092.5 177672.5 8157.5 177807.5 ;
      RECT  8092.5 177672.5 8157.5 177807.5 ;
      RECT  7902.5 177672.5 7967.5 177807.5 ;
      RECT  7522.5 176832.5 7587.5 176967.5 ;
      RECT  7712.5 176832.5 7777.5 176967.5 ;
      RECT  7712.5 176832.5 7777.5 176967.5 ;
      RECT  7522.5 176832.5 7587.5 176967.5 ;
      RECT  7712.5 176832.5 7777.5 176967.5 ;
      RECT  7902.5 176832.5 7967.5 176967.5 ;
      RECT  7902.5 176832.5 7967.5 176967.5 ;
      RECT  7712.5 176832.5 7777.5 176967.5 ;
      RECT  7902.5 176832.5 7967.5 176967.5 ;
      RECT  8092.5 176832.5 8157.5 176967.5 ;
      RECT  8092.5 176832.5 8157.5 176967.5 ;
      RECT  7902.5 176832.5 7967.5 176967.5 ;
      RECT  8262.5 177762.5 8327.5 177897.5 ;
      RECT  8262.5 176787.5 8327.5 176922.5 ;
      RECT  8097.5 177045.0 7962.5 177110.0 ;
      RECT  7907.5 177185.0 7772.5 177250.0 ;
      RECT  7717.5 177325.0 7582.5 177390.0 ;
      RECT  7712.5 177672.5 7777.5 177807.5 ;
      RECT  8092.5 177672.5 8157.5 177807.5 ;
      RECT  8092.5 176832.5 8157.5 176967.5 ;
      RECT  8092.5 177290.0 8157.5 177425.0 ;
      RECT  7582.5 177325.0 7717.5 177390.0 ;
      RECT  7772.5 177185.0 7907.5 177250.0 ;
      RECT  7962.5 177045.0 8097.5 177110.0 ;
      RECT  8092.5 177290.0 8157.5 177425.0 ;
      RECT  7455.0 177982.5 8465.0 178047.5 ;
      RECT  7455.0 176637.5 8465.0 176702.5 ;
      RECT  7522.5 179197.5 7587.5 179392.5 ;
      RECT  7522.5 178357.5 7587.5 177982.5 ;
      RECT  7902.5 178357.5 7967.5 177982.5 ;
      RECT  8262.5 178200.0 8327.5 178015.0 ;
      RECT  8262.5 179360.0 8327.5 179175.0 ;
      RECT  7522.5 178357.5 7587.5 178222.5 ;
      RECT  7712.5 178357.5 7777.5 178222.5 ;
      RECT  7712.5 178357.5 7777.5 178222.5 ;
      RECT  7522.5 178357.5 7587.5 178222.5 ;
      RECT  7712.5 178357.5 7777.5 178222.5 ;
      RECT  7902.5 178357.5 7967.5 178222.5 ;
      RECT  7902.5 178357.5 7967.5 178222.5 ;
      RECT  7712.5 178357.5 7777.5 178222.5 ;
      RECT  7902.5 178357.5 7967.5 178222.5 ;
      RECT  8092.5 178357.5 8157.5 178222.5 ;
      RECT  8092.5 178357.5 8157.5 178222.5 ;
      RECT  7902.5 178357.5 7967.5 178222.5 ;
      RECT  7522.5 179197.5 7587.5 179062.5 ;
      RECT  7712.5 179197.5 7777.5 179062.5 ;
      RECT  7712.5 179197.5 7777.5 179062.5 ;
      RECT  7522.5 179197.5 7587.5 179062.5 ;
      RECT  7712.5 179197.5 7777.5 179062.5 ;
      RECT  7902.5 179197.5 7967.5 179062.5 ;
      RECT  7902.5 179197.5 7967.5 179062.5 ;
      RECT  7712.5 179197.5 7777.5 179062.5 ;
      RECT  7902.5 179197.5 7967.5 179062.5 ;
      RECT  8092.5 179197.5 8157.5 179062.5 ;
      RECT  8092.5 179197.5 8157.5 179062.5 ;
      RECT  7902.5 179197.5 7967.5 179062.5 ;
      RECT  8262.5 178267.5 8327.5 178132.5 ;
      RECT  8262.5 179242.5 8327.5 179107.5 ;
      RECT  8097.5 178985.0 7962.5 178920.0 ;
      RECT  7907.5 178845.0 7772.5 178780.0 ;
      RECT  7717.5 178705.0 7582.5 178640.0 ;
      RECT  7712.5 178357.5 7777.5 178222.5 ;
      RECT  8092.5 178357.5 8157.5 178222.5 ;
      RECT  8092.5 179197.5 8157.5 179062.5 ;
      RECT  8092.5 178740.0 8157.5 178605.0 ;
      RECT  7582.5 178705.0 7717.5 178640.0 ;
      RECT  7772.5 178845.0 7907.5 178780.0 ;
      RECT  7962.5 178985.0 8097.5 178920.0 ;
      RECT  8092.5 178740.0 8157.5 178605.0 ;
      RECT  7455.0 178047.5 8465.0 177982.5 ;
      RECT  7455.0 179392.5 8465.0 179327.5 ;
      RECT  7522.5 179522.5 7587.5 179327.5 ;
      RECT  7522.5 180362.5 7587.5 180737.5 ;
      RECT  7902.5 180362.5 7967.5 180737.5 ;
      RECT  8262.5 180520.0 8327.5 180705.0 ;
      RECT  8262.5 179360.0 8327.5 179545.0 ;
      RECT  7522.5 180362.5 7587.5 180497.5 ;
      RECT  7712.5 180362.5 7777.5 180497.5 ;
      RECT  7712.5 180362.5 7777.5 180497.5 ;
      RECT  7522.5 180362.5 7587.5 180497.5 ;
      RECT  7712.5 180362.5 7777.5 180497.5 ;
      RECT  7902.5 180362.5 7967.5 180497.5 ;
      RECT  7902.5 180362.5 7967.5 180497.5 ;
      RECT  7712.5 180362.5 7777.5 180497.5 ;
      RECT  7902.5 180362.5 7967.5 180497.5 ;
      RECT  8092.5 180362.5 8157.5 180497.5 ;
      RECT  8092.5 180362.5 8157.5 180497.5 ;
      RECT  7902.5 180362.5 7967.5 180497.5 ;
      RECT  7522.5 179522.5 7587.5 179657.5 ;
      RECT  7712.5 179522.5 7777.5 179657.5 ;
      RECT  7712.5 179522.5 7777.5 179657.5 ;
      RECT  7522.5 179522.5 7587.5 179657.5 ;
      RECT  7712.5 179522.5 7777.5 179657.5 ;
      RECT  7902.5 179522.5 7967.5 179657.5 ;
      RECT  7902.5 179522.5 7967.5 179657.5 ;
      RECT  7712.5 179522.5 7777.5 179657.5 ;
      RECT  7902.5 179522.5 7967.5 179657.5 ;
      RECT  8092.5 179522.5 8157.5 179657.5 ;
      RECT  8092.5 179522.5 8157.5 179657.5 ;
      RECT  7902.5 179522.5 7967.5 179657.5 ;
      RECT  8262.5 180452.5 8327.5 180587.5 ;
      RECT  8262.5 179477.5 8327.5 179612.5 ;
      RECT  8097.5 179735.0 7962.5 179800.0 ;
      RECT  7907.5 179875.0 7772.5 179940.0 ;
      RECT  7717.5 180015.0 7582.5 180080.0 ;
      RECT  7712.5 180362.5 7777.5 180497.5 ;
      RECT  8092.5 180362.5 8157.5 180497.5 ;
      RECT  8092.5 179522.5 8157.5 179657.5 ;
      RECT  8092.5 179980.0 8157.5 180115.0 ;
      RECT  7582.5 180015.0 7717.5 180080.0 ;
      RECT  7772.5 179875.0 7907.5 179940.0 ;
      RECT  7962.5 179735.0 8097.5 179800.0 ;
      RECT  8092.5 179980.0 8157.5 180115.0 ;
      RECT  7455.0 180672.5 8465.0 180737.5 ;
      RECT  7455.0 179327.5 8465.0 179392.5 ;
      RECT  7522.5 181887.5 7587.5 182082.5 ;
      RECT  7522.5 181047.5 7587.5 180672.5 ;
      RECT  7902.5 181047.5 7967.5 180672.5 ;
      RECT  8262.5 180890.0 8327.5 180705.0 ;
      RECT  8262.5 182050.0 8327.5 181865.0 ;
      RECT  7522.5 181047.5 7587.5 180912.5 ;
      RECT  7712.5 181047.5 7777.5 180912.5 ;
      RECT  7712.5 181047.5 7777.5 180912.5 ;
      RECT  7522.5 181047.5 7587.5 180912.5 ;
      RECT  7712.5 181047.5 7777.5 180912.5 ;
      RECT  7902.5 181047.5 7967.5 180912.5 ;
      RECT  7902.5 181047.5 7967.5 180912.5 ;
      RECT  7712.5 181047.5 7777.5 180912.5 ;
      RECT  7902.5 181047.5 7967.5 180912.5 ;
      RECT  8092.5 181047.5 8157.5 180912.5 ;
      RECT  8092.5 181047.5 8157.5 180912.5 ;
      RECT  7902.5 181047.5 7967.5 180912.5 ;
      RECT  7522.5 181887.5 7587.5 181752.5 ;
      RECT  7712.5 181887.5 7777.5 181752.5 ;
      RECT  7712.5 181887.5 7777.5 181752.5 ;
      RECT  7522.5 181887.5 7587.5 181752.5 ;
      RECT  7712.5 181887.5 7777.5 181752.5 ;
      RECT  7902.5 181887.5 7967.5 181752.5 ;
      RECT  7902.5 181887.5 7967.5 181752.5 ;
      RECT  7712.5 181887.5 7777.5 181752.5 ;
      RECT  7902.5 181887.5 7967.5 181752.5 ;
      RECT  8092.5 181887.5 8157.5 181752.5 ;
      RECT  8092.5 181887.5 8157.5 181752.5 ;
      RECT  7902.5 181887.5 7967.5 181752.5 ;
      RECT  8262.5 180957.5 8327.5 180822.5 ;
      RECT  8262.5 181932.5 8327.5 181797.5 ;
      RECT  8097.5 181675.0 7962.5 181610.0 ;
      RECT  7907.5 181535.0 7772.5 181470.0 ;
      RECT  7717.5 181395.0 7582.5 181330.0 ;
      RECT  7712.5 181047.5 7777.5 180912.5 ;
      RECT  8092.5 181047.5 8157.5 180912.5 ;
      RECT  8092.5 181887.5 8157.5 181752.5 ;
      RECT  8092.5 181430.0 8157.5 181295.0 ;
      RECT  7582.5 181395.0 7717.5 181330.0 ;
      RECT  7772.5 181535.0 7907.5 181470.0 ;
      RECT  7962.5 181675.0 8097.5 181610.0 ;
      RECT  8092.5 181430.0 8157.5 181295.0 ;
      RECT  7455.0 180737.5 8465.0 180672.5 ;
      RECT  7455.0 182082.5 8465.0 182017.5 ;
      RECT  7522.5 182212.5 7587.5 182017.5 ;
      RECT  7522.5 183052.5 7587.5 183427.5 ;
      RECT  7902.5 183052.5 7967.5 183427.5 ;
      RECT  8262.5 183210.0 8327.5 183395.0 ;
      RECT  8262.5 182050.0 8327.5 182235.0 ;
      RECT  7522.5 183052.5 7587.5 183187.5 ;
      RECT  7712.5 183052.5 7777.5 183187.5 ;
      RECT  7712.5 183052.5 7777.5 183187.5 ;
      RECT  7522.5 183052.5 7587.5 183187.5 ;
      RECT  7712.5 183052.5 7777.5 183187.5 ;
      RECT  7902.5 183052.5 7967.5 183187.5 ;
      RECT  7902.5 183052.5 7967.5 183187.5 ;
      RECT  7712.5 183052.5 7777.5 183187.5 ;
      RECT  7902.5 183052.5 7967.5 183187.5 ;
      RECT  8092.5 183052.5 8157.5 183187.5 ;
      RECT  8092.5 183052.5 8157.5 183187.5 ;
      RECT  7902.5 183052.5 7967.5 183187.5 ;
      RECT  7522.5 182212.5 7587.5 182347.5 ;
      RECT  7712.5 182212.5 7777.5 182347.5 ;
      RECT  7712.5 182212.5 7777.5 182347.5 ;
      RECT  7522.5 182212.5 7587.5 182347.5 ;
      RECT  7712.5 182212.5 7777.5 182347.5 ;
      RECT  7902.5 182212.5 7967.5 182347.5 ;
      RECT  7902.5 182212.5 7967.5 182347.5 ;
      RECT  7712.5 182212.5 7777.5 182347.5 ;
      RECT  7902.5 182212.5 7967.5 182347.5 ;
      RECT  8092.5 182212.5 8157.5 182347.5 ;
      RECT  8092.5 182212.5 8157.5 182347.5 ;
      RECT  7902.5 182212.5 7967.5 182347.5 ;
      RECT  8262.5 183142.5 8327.5 183277.5 ;
      RECT  8262.5 182167.5 8327.5 182302.5 ;
      RECT  8097.5 182425.0 7962.5 182490.0 ;
      RECT  7907.5 182565.0 7772.5 182630.0 ;
      RECT  7717.5 182705.0 7582.5 182770.0 ;
      RECT  7712.5 183052.5 7777.5 183187.5 ;
      RECT  8092.5 183052.5 8157.5 183187.5 ;
      RECT  8092.5 182212.5 8157.5 182347.5 ;
      RECT  8092.5 182670.0 8157.5 182805.0 ;
      RECT  7582.5 182705.0 7717.5 182770.0 ;
      RECT  7772.5 182565.0 7907.5 182630.0 ;
      RECT  7962.5 182425.0 8097.5 182490.0 ;
      RECT  8092.5 182670.0 8157.5 182805.0 ;
      RECT  7455.0 183362.5 8465.0 183427.5 ;
      RECT  7455.0 182017.5 8465.0 182082.5 ;
      RECT  7522.5 184577.5 7587.5 184772.5 ;
      RECT  7522.5 183737.5 7587.5 183362.5 ;
      RECT  7902.5 183737.5 7967.5 183362.5 ;
      RECT  8262.5 183580.0 8327.5 183395.0 ;
      RECT  8262.5 184740.0 8327.5 184555.0 ;
      RECT  7522.5 183737.5 7587.5 183602.5 ;
      RECT  7712.5 183737.5 7777.5 183602.5 ;
      RECT  7712.5 183737.5 7777.5 183602.5 ;
      RECT  7522.5 183737.5 7587.5 183602.5 ;
      RECT  7712.5 183737.5 7777.5 183602.5 ;
      RECT  7902.5 183737.5 7967.5 183602.5 ;
      RECT  7902.5 183737.5 7967.5 183602.5 ;
      RECT  7712.5 183737.5 7777.5 183602.5 ;
      RECT  7902.5 183737.5 7967.5 183602.5 ;
      RECT  8092.5 183737.5 8157.5 183602.5 ;
      RECT  8092.5 183737.5 8157.5 183602.5 ;
      RECT  7902.5 183737.5 7967.5 183602.5 ;
      RECT  7522.5 184577.5 7587.5 184442.5 ;
      RECT  7712.5 184577.5 7777.5 184442.5 ;
      RECT  7712.5 184577.5 7777.5 184442.5 ;
      RECT  7522.5 184577.5 7587.5 184442.5 ;
      RECT  7712.5 184577.5 7777.5 184442.5 ;
      RECT  7902.5 184577.5 7967.5 184442.5 ;
      RECT  7902.5 184577.5 7967.5 184442.5 ;
      RECT  7712.5 184577.5 7777.5 184442.5 ;
      RECT  7902.5 184577.5 7967.5 184442.5 ;
      RECT  8092.5 184577.5 8157.5 184442.5 ;
      RECT  8092.5 184577.5 8157.5 184442.5 ;
      RECT  7902.5 184577.5 7967.5 184442.5 ;
      RECT  8262.5 183647.5 8327.5 183512.5 ;
      RECT  8262.5 184622.5 8327.5 184487.5 ;
      RECT  8097.5 184365.0 7962.5 184300.0 ;
      RECT  7907.5 184225.0 7772.5 184160.0 ;
      RECT  7717.5 184085.0 7582.5 184020.0 ;
      RECT  7712.5 183737.5 7777.5 183602.5 ;
      RECT  8092.5 183737.5 8157.5 183602.5 ;
      RECT  8092.5 184577.5 8157.5 184442.5 ;
      RECT  8092.5 184120.0 8157.5 183985.0 ;
      RECT  7582.5 184085.0 7717.5 184020.0 ;
      RECT  7772.5 184225.0 7907.5 184160.0 ;
      RECT  7962.5 184365.0 8097.5 184300.0 ;
      RECT  8092.5 184120.0 8157.5 183985.0 ;
      RECT  7455.0 183427.5 8465.0 183362.5 ;
      RECT  7455.0 184772.5 8465.0 184707.5 ;
      RECT  7522.5 184902.5 7587.5 184707.5 ;
      RECT  7522.5 185742.5 7587.5 186117.5 ;
      RECT  7902.5 185742.5 7967.5 186117.5 ;
      RECT  8262.5 185900.0 8327.5 186085.0 ;
      RECT  8262.5 184740.0 8327.5 184925.0 ;
      RECT  7522.5 185742.5 7587.5 185877.5 ;
      RECT  7712.5 185742.5 7777.5 185877.5 ;
      RECT  7712.5 185742.5 7777.5 185877.5 ;
      RECT  7522.5 185742.5 7587.5 185877.5 ;
      RECT  7712.5 185742.5 7777.5 185877.5 ;
      RECT  7902.5 185742.5 7967.5 185877.5 ;
      RECT  7902.5 185742.5 7967.5 185877.5 ;
      RECT  7712.5 185742.5 7777.5 185877.5 ;
      RECT  7902.5 185742.5 7967.5 185877.5 ;
      RECT  8092.5 185742.5 8157.5 185877.5 ;
      RECT  8092.5 185742.5 8157.5 185877.5 ;
      RECT  7902.5 185742.5 7967.5 185877.5 ;
      RECT  7522.5 184902.5 7587.5 185037.5 ;
      RECT  7712.5 184902.5 7777.5 185037.5 ;
      RECT  7712.5 184902.5 7777.5 185037.5 ;
      RECT  7522.5 184902.5 7587.5 185037.5 ;
      RECT  7712.5 184902.5 7777.5 185037.5 ;
      RECT  7902.5 184902.5 7967.5 185037.5 ;
      RECT  7902.5 184902.5 7967.5 185037.5 ;
      RECT  7712.5 184902.5 7777.5 185037.5 ;
      RECT  7902.5 184902.5 7967.5 185037.5 ;
      RECT  8092.5 184902.5 8157.5 185037.5 ;
      RECT  8092.5 184902.5 8157.5 185037.5 ;
      RECT  7902.5 184902.5 7967.5 185037.5 ;
      RECT  8262.5 185832.5 8327.5 185967.5 ;
      RECT  8262.5 184857.5 8327.5 184992.5 ;
      RECT  8097.5 185115.0 7962.5 185180.0 ;
      RECT  7907.5 185255.0 7772.5 185320.0 ;
      RECT  7717.5 185395.0 7582.5 185460.0 ;
      RECT  7712.5 185742.5 7777.5 185877.5 ;
      RECT  8092.5 185742.5 8157.5 185877.5 ;
      RECT  8092.5 184902.5 8157.5 185037.5 ;
      RECT  8092.5 185360.0 8157.5 185495.0 ;
      RECT  7582.5 185395.0 7717.5 185460.0 ;
      RECT  7772.5 185255.0 7907.5 185320.0 ;
      RECT  7962.5 185115.0 8097.5 185180.0 ;
      RECT  8092.5 185360.0 8157.5 185495.0 ;
      RECT  7455.0 186052.5 8465.0 186117.5 ;
      RECT  7455.0 184707.5 8465.0 184772.5 ;
      RECT  7522.5 187267.5 7587.5 187462.5 ;
      RECT  7522.5 186427.5 7587.5 186052.5 ;
      RECT  7902.5 186427.5 7967.5 186052.5 ;
      RECT  8262.5 186270.0 8327.5 186085.0 ;
      RECT  8262.5 187430.0 8327.5 187245.0 ;
      RECT  7522.5 186427.5 7587.5 186292.5 ;
      RECT  7712.5 186427.5 7777.5 186292.5 ;
      RECT  7712.5 186427.5 7777.5 186292.5 ;
      RECT  7522.5 186427.5 7587.5 186292.5 ;
      RECT  7712.5 186427.5 7777.5 186292.5 ;
      RECT  7902.5 186427.5 7967.5 186292.5 ;
      RECT  7902.5 186427.5 7967.5 186292.5 ;
      RECT  7712.5 186427.5 7777.5 186292.5 ;
      RECT  7902.5 186427.5 7967.5 186292.5 ;
      RECT  8092.5 186427.5 8157.5 186292.5 ;
      RECT  8092.5 186427.5 8157.5 186292.5 ;
      RECT  7902.5 186427.5 7967.5 186292.5 ;
      RECT  7522.5 187267.5 7587.5 187132.5 ;
      RECT  7712.5 187267.5 7777.5 187132.5 ;
      RECT  7712.5 187267.5 7777.5 187132.5 ;
      RECT  7522.5 187267.5 7587.5 187132.5 ;
      RECT  7712.5 187267.5 7777.5 187132.5 ;
      RECT  7902.5 187267.5 7967.5 187132.5 ;
      RECT  7902.5 187267.5 7967.5 187132.5 ;
      RECT  7712.5 187267.5 7777.5 187132.5 ;
      RECT  7902.5 187267.5 7967.5 187132.5 ;
      RECT  8092.5 187267.5 8157.5 187132.5 ;
      RECT  8092.5 187267.5 8157.5 187132.5 ;
      RECT  7902.5 187267.5 7967.5 187132.5 ;
      RECT  8262.5 186337.5 8327.5 186202.5 ;
      RECT  8262.5 187312.5 8327.5 187177.5 ;
      RECT  8097.5 187055.0 7962.5 186990.0 ;
      RECT  7907.5 186915.0 7772.5 186850.0 ;
      RECT  7717.5 186775.0 7582.5 186710.0 ;
      RECT  7712.5 186427.5 7777.5 186292.5 ;
      RECT  8092.5 186427.5 8157.5 186292.5 ;
      RECT  8092.5 187267.5 8157.5 187132.5 ;
      RECT  8092.5 186810.0 8157.5 186675.0 ;
      RECT  7582.5 186775.0 7717.5 186710.0 ;
      RECT  7772.5 186915.0 7907.5 186850.0 ;
      RECT  7962.5 187055.0 8097.5 186990.0 ;
      RECT  8092.5 186810.0 8157.5 186675.0 ;
      RECT  7455.0 186117.5 8465.0 186052.5 ;
      RECT  7455.0 187462.5 8465.0 187397.5 ;
      RECT  7522.5 187592.5 7587.5 187397.5 ;
      RECT  7522.5 188432.5 7587.5 188807.5 ;
      RECT  7902.5 188432.5 7967.5 188807.5 ;
      RECT  8262.5 188590.0 8327.5 188775.0 ;
      RECT  8262.5 187430.0 8327.5 187615.0 ;
      RECT  7522.5 188432.5 7587.5 188567.5 ;
      RECT  7712.5 188432.5 7777.5 188567.5 ;
      RECT  7712.5 188432.5 7777.5 188567.5 ;
      RECT  7522.5 188432.5 7587.5 188567.5 ;
      RECT  7712.5 188432.5 7777.5 188567.5 ;
      RECT  7902.5 188432.5 7967.5 188567.5 ;
      RECT  7902.5 188432.5 7967.5 188567.5 ;
      RECT  7712.5 188432.5 7777.5 188567.5 ;
      RECT  7902.5 188432.5 7967.5 188567.5 ;
      RECT  8092.5 188432.5 8157.5 188567.5 ;
      RECT  8092.5 188432.5 8157.5 188567.5 ;
      RECT  7902.5 188432.5 7967.5 188567.5 ;
      RECT  7522.5 187592.5 7587.5 187727.5 ;
      RECT  7712.5 187592.5 7777.5 187727.5 ;
      RECT  7712.5 187592.5 7777.5 187727.5 ;
      RECT  7522.5 187592.5 7587.5 187727.5 ;
      RECT  7712.5 187592.5 7777.5 187727.5 ;
      RECT  7902.5 187592.5 7967.5 187727.5 ;
      RECT  7902.5 187592.5 7967.5 187727.5 ;
      RECT  7712.5 187592.5 7777.5 187727.5 ;
      RECT  7902.5 187592.5 7967.5 187727.5 ;
      RECT  8092.5 187592.5 8157.5 187727.5 ;
      RECT  8092.5 187592.5 8157.5 187727.5 ;
      RECT  7902.5 187592.5 7967.5 187727.5 ;
      RECT  8262.5 188522.5 8327.5 188657.5 ;
      RECT  8262.5 187547.5 8327.5 187682.5 ;
      RECT  8097.5 187805.0 7962.5 187870.0 ;
      RECT  7907.5 187945.0 7772.5 188010.0 ;
      RECT  7717.5 188085.0 7582.5 188150.0 ;
      RECT  7712.5 188432.5 7777.5 188567.5 ;
      RECT  8092.5 188432.5 8157.5 188567.5 ;
      RECT  8092.5 187592.5 8157.5 187727.5 ;
      RECT  8092.5 188050.0 8157.5 188185.0 ;
      RECT  7582.5 188085.0 7717.5 188150.0 ;
      RECT  7772.5 187945.0 7907.5 188010.0 ;
      RECT  7962.5 187805.0 8097.5 187870.0 ;
      RECT  8092.5 188050.0 8157.5 188185.0 ;
      RECT  7455.0 188742.5 8465.0 188807.5 ;
      RECT  7455.0 187397.5 8465.0 187462.5 ;
      RECT  7522.5 189957.5 7587.5 190152.5 ;
      RECT  7522.5 189117.5 7587.5 188742.5 ;
      RECT  7902.5 189117.5 7967.5 188742.5 ;
      RECT  8262.5 188960.0 8327.5 188775.0 ;
      RECT  8262.5 190120.0 8327.5 189935.0 ;
      RECT  7522.5 189117.5 7587.5 188982.5 ;
      RECT  7712.5 189117.5 7777.5 188982.5 ;
      RECT  7712.5 189117.5 7777.5 188982.5 ;
      RECT  7522.5 189117.5 7587.5 188982.5 ;
      RECT  7712.5 189117.5 7777.5 188982.5 ;
      RECT  7902.5 189117.5 7967.5 188982.5 ;
      RECT  7902.5 189117.5 7967.5 188982.5 ;
      RECT  7712.5 189117.5 7777.5 188982.5 ;
      RECT  7902.5 189117.5 7967.5 188982.5 ;
      RECT  8092.5 189117.5 8157.5 188982.5 ;
      RECT  8092.5 189117.5 8157.5 188982.5 ;
      RECT  7902.5 189117.5 7967.5 188982.5 ;
      RECT  7522.5 189957.5 7587.5 189822.5 ;
      RECT  7712.5 189957.5 7777.5 189822.5 ;
      RECT  7712.5 189957.5 7777.5 189822.5 ;
      RECT  7522.5 189957.5 7587.5 189822.5 ;
      RECT  7712.5 189957.5 7777.5 189822.5 ;
      RECT  7902.5 189957.5 7967.5 189822.5 ;
      RECT  7902.5 189957.5 7967.5 189822.5 ;
      RECT  7712.5 189957.5 7777.5 189822.5 ;
      RECT  7902.5 189957.5 7967.5 189822.5 ;
      RECT  8092.5 189957.5 8157.5 189822.5 ;
      RECT  8092.5 189957.5 8157.5 189822.5 ;
      RECT  7902.5 189957.5 7967.5 189822.5 ;
      RECT  8262.5 189027.5 8327.5 188892.5 ;
      RECT  8262.5 190002.5 8327.5 189867.5 ;
      RECT  8097.5 189745.0 7962.5 189680.0 ;
      RECT  7907.5 189605.0 7772.5 189540.0 ;
      RECT  7717.5 189465.0 7582.5 189400.0 ;
      RECT  7712.5 189117.5 7777.5 188982.5 ;
      RECT  8092.5 189117.5 8157.5 188982.5 ;
      RECT  8092.5 189957.5 8157.5 189822.5 ;
      RECT  8092.5 189500.0 8157.5 189365.0 ;
      RECT  7582.5 189465.0 7717.5 189400.0 ;
      RECT  7772.5 189605.0 7907.5 189540.0 ;
      RECT  7962.5 189745.0 8097.5 189680.0 ;
      RECT  8092.5 189500.0 8157.5 189365.0 ;
      RECT  7455.0 188807.5 8465.0 188742.5 ;
      RECT  7455.0 190152.5 8465.0 190087.5 ;
      RECT  7522.5 190282.5 7587.5 190087.5 ;
      RECT  7522.5 191122.5 7587.5 191497.5 ;
      RECT  7902.5 191122.5 7967.5 191497.5 ;
      RECT  8262.5 191280.0 8327.5 191465.0 ;
      RECT  8262.5 190120.0 8327.5 190305.0 ;
      RECT  7522.5 191122.5 7587.5 191257.5 ;
      RECT  7712.5 191122.5 7777.5 191257.5 ;
      RECT  7712.5 191122.5 7777.5 191257.5 ;
      RECT  7522.5 191122.5 7587.5 191257.5 ;
      RECT  7712.5 191122.5 7777.5 191257.5 ;
      RECT  7902.5 191122.5 7967.5 191257.5 ;
      RECT  7902.5 191122.5 7967.5 191257.5 ;
      RECT  7712.5 191122.5 7777.5 191257.5 ;
      RECT  7902.5 191122.5 7967.5 191257.5 ;
      RECT  8092.5 191122.5 8157.5 191257.5 ;
      RECT  8092.5 191122.5 8157.5 191257.5 ;
      RECT  7902.5 191122.5 7967.5 191257.5 ;
      RECT  7522.5 190282.5 7587.5 190417.5 ;
      RECT  7712.5 190282.5 7777.5 190417.5 ;
      RECT  7712.5 190282.5 7777.5 190417.5 ;
      RECT  7522.5 190282.5 7587.5 190417.5 ;
      RECT  7712.5 190282.5 7777.5 190417.5 ;
      RECT  7902.5 190282.5 7967.5 190417.5 ;
      RECT  7902.5 190282.5 7967.5 190417.5 ;
      RECT  7712.5 190282.5 7777.5 190417.5 ;
      RECT  7902.5 190282.5 7967.5 190417.5 ;
      RECT  8092.5 190282.5 8157.5 190417.5 ;
      RECT  8092.5 190282.5 8157.5 190417.5 ;
      RECT  7902.5 190282.5 7967.5 190417.5 ;
      RECT  8262.5 191212.5 8327.5 191347.5 ;
      RECT  8262.5 190237.5 8327.5 190372.5 ;
      RECT  8097.5 190495.0 7962.5 190560.0 ;
      RECT  7907.5 190635.0 7772.5 190700.0 ;
      RECT  7717.5 190775.0 7582.5 190840.0 ;
      RECT  7712.5 191122.5 7777.5 191257.5 ;
      RECT  8092.5 191122.5 8157.5 191257.5 ;
      RECT  8092.5 190282.5 8157.5 190417.5 ;
      RECT  8092.5 190740.0 8157.5 190875.0 ;
      RECT  7582.5 190775.0 7717.5 190840.0 ;
      RECT  7772.5 190635.0 7907.5 190700.0 ;
      RECT  7962.5 190495.0 8097.5 190560.0 ;
      RECT  8092.5 190740.0 8157.5 190875.0 ;
      RECT  7455.0 191432.5 8465.0 191497.5 ;
      RECT  7455.0 190087.5 8465.0 190152.5 ;
      RECT  7522.5 192647.5 7587.5 192842.5 ;
      RECT  7522.5 191807.5 7587.5 191432.5 ;
      RECT  7902.5 191807.5 7967.5 191432.5 ;
      RECT  8262.5 191650.0 8327.5 191465.0 ;
      RECT  8262.5 192810.0 8327.5 192625.0 ;
      RECT  7522.5 191807.5 7587.5 191672.5 ;
      RECT  7712.5 191807.5 7777.5 191672.5 ;
      RECT  7712.5 191807.5 7777.5 191672.5 ;
      RECT  7522.5 191807.5 7587.5 191672.5 ;
      RECT  7712.5 191807.5 7777.5 191672.5 ;
      RECT  7902.5 191807.5 7967.5 191672.5 ;
      RECT  7902.5 191807.5 7967.5 191672.5 ;
      RECT  7712.5 191807.5 7777.5 191672.5 ;
      RECT  7902.5 191807.5 7967.5 191672.5 ;
      RECT  8092.5 191807.5 8157.5 191672.5 ;
      RECT  8092.5 191807.5 8157.5 191672.5 ;
      RECT  7902.5 191807.5 7967.5 191672.5 ;
      RECT  7522.5 192647.5 7587.5 192512.5 ;
      RECT  7712.5 192647.5 7777.5 192512.5 ;
      RECT  7712.5 192647.5 7777.5 192512.5 ;
      RECT  7522.5 192647.5 7587.5 192512.5 ;
      RECT  7712.5 192647.5 7777.5 192512.5 ;
      RECT  7902.5 192647.5 7967.5 192512.5 ;
      RECT  7902.5 192647.5 7967.5 192512.5 ;
      RECT  7712.5 192647.5 7777.5 192512.5 ;
      RECT  7902.5 192647.5 7967.5 192512.5 ;
      RECT  8092.5 192647.5 8157.5 192512.5 ;
      RECT  8092.5 192647.5 8157.5 192512.5 ;
      RECT  7902.5 192647.5 7967.5 192512.5 ;
      RECT  8262.5 191717.5 8327.5 191582.5 ;
      RECT  8262.5 192692.5 8327.5 192557.5 ;
      RECT  8097.5 192435.0 7962.5 192370.0 ;
      RECT  7907.5 192295.0 7772.5 192230.0 ;
      RECT  7717.5 192155.0 7582.5 192090.0 ;
      RECT  7712.5 191807.5 7777.5 191672.5 ;
      RECT  8092.5 191807.5 8157.5 191672.5 ;
      RECT  8092.5 192647.5 8157.5 192512.5 ;
      RECT  8092.5 192190.0 8157.5 192055.0 ;
      RECT  7582.5 192155.0 7717.5 192090.0 ;
      RECT  7772.5 192295.0 7907.5 192230.0 ;
      RECT  7962.5 192435.0 8097.5 192370.0 ;
      RECT  8092.5 192190.0 8157.5 192055.0 ;
      RECT  7455.0 191497.5 8465.0 191432.5 ;
      RECT  7455.0 192842.5 8465.0 192777.5 ;
      RECT  7522.5 192972.5 7587.5 192777.5 ;
      RECT  7522.5 193812.5 7587.5 194187.5 ;
      RECT  7902.5 193812.5 7967.5 194187.5 ;
      RECT  8262.5 193970.0 8327.5 194155.0 ;
      RECT  8262.5 192810.0 8327.5 192995.0 ;
      RECT  7522.5 193812.5 7587.5 193947.5 ;
      RECT  7712.5 193812.5 7777.5 193947.5 ;
      RECT  7712.5 193812.5 7777.5 193947.5 ;
      RECT  7522.5 193812.5 7587.5 193947.5 ;
      RECT  7712.5 193812.5 7777.5 193947.5 ;
      RECT  7902.5 193812.5 7967.5 193947.5 ;
      RECT  7902.5 193812.5 7967.5 193947.5 ;
      RECT  7712.5 193812.5 7777.5 193947.5 ;
      RECT  7902.5 193812.5 7967.5 193947.5 ;
      RECT  8092.5 193812.5 8157.5 193947.5 ;
      RECT  8092.5 193812.5 8157.5 193947.5 ;
      RECT  7902.5 193812.5 7967.5 193947.5 ;
      RECT  7522.5 192972.5 7587.5 193107.5 ;
      RECT  7712.5 192972.5 7777.5 193107.5 ;
      RECT  7712.5 192972.5 7777.5 193107.5 ;
      RECT  7522.5 192972.5 7587.5 193107.5 ;
      RECT  7712.5 192972.5 7777.5 193107.5 ;
      RECT  7902.5 192972.5 7967.5 193107.5 ;
      RECT  7902.5 192972.5 7967.5 193107.5 ;
      RECT  7712.5 192972.5 7777.5 193107.5 ;
      RECT  7902.5 192972.5 7967.5 193107.5 ;
      RECT  8092.5 192972.5 8157.5 193107.5 ;
      RECT  8092.5 192972.5 8157.5 193107.5 ;
      RECT  7902.5 192972.5 7967.5 193107.5 ;
      RECT  8262.5 193902.5 8327.5 194037.5 ;
      RECT  8262.5 192927.5 8327.5 193062.5 ;
      RECT  8097.5 193185.0 7962.5 193250.0 ;
      RECT  7907.5 193325.0 7772.5 193390.0 ;
      RECT  7717.5 193465.0 7582.5 193530.0 ;
      RECT  7712.5 193812.5 7777.5 193947.5 ;
      RECT  8092.5 193812.5 8157.5 193947.5 ;
      RECT  8092.5 192972.5 8157.5 193107.5 ;
      RECT  8092.5 193430.0 8157.5 193565.0 ;
      RECT  7582.5 193465.0 7717.5 193530.0 ;
      RECT  7772.5 193325.0 7907.5 193390.0 ;
      RECT  7962.5 193185.0 8097.5 193250.0 ;
      RECT  8092.5 193430.0 8157.5 193565.0 ;
      RECT  7455.0 194122.5 8465.0 194187.5 ;
      RECT  7455.0 192777.5 8465.0 192842.5 ;
      RECT  7522.5 195337.5 7587.5 195532.5 ;
      RECT  7522.5 194497.5 7587.5 194122.5 ;
      RECT  7902.5 194497.5 7967.5 194122.5 ;
      RECT  8262.5 194340.0 8327.5 194155.0 ;
      RECT  8262.5 195500.0 8327.5 195315.0 ;
      RECT  7522.5 194497.5 7587.5 194362.5 ;
      RECT  7712.5 194497.5 7777.5 194362.5 ;
      RECT  7712.5 194497.5 7777.5 194362.5 ;
      RECT  7522.5 194497.5 7587.5 194362.5 ;
      RECT  7712.5 194497.5 7777.5 194362.5 ;
      RECT  7902.5 194497.5 7967.5 194362.5 ;
      RECT  7902.5 194497.5 7967.5 194362.5 ;
      RECT  7712.5 194497.5 7777.5 194362.5 ;
      RECT  7902.5 194497.5 7967.5 194362.5 ;
      RECT  8092.5 194497.5 8157.5 194362.5 ;
      RECT  8092.5 194497.5 8157.5 194362.5 ;
      RECT  7902.5 194497.5 7967.5 194362.5 ;
      RECT  7522.5 195337.5 7587.5 195202.5 ;
      RECT  7712.5 195337.5 7777.5 195202.5 ;
      RECT  7712.5 195337.5 7777.5 195202.5 ;
      RECT  7522.5 195337.5 7587.5 195202.5 ;
      RECT  7712.5 195337.5 7777.5 195202.5 ;
      RECT  7902.5 195337.5 7967.5 195202.5 ;
      RECT  7902.5 195337.5 7967.5 195202.5 ;
      RECT  7712.5 195337.5 7777.5 195202.5 ;
      RECT  7902.5 195337.5 7967.5 195202.5 ;
      RECT  8092.5 195337.5 8157.5 195202.5 ;
      RECT  8092.5 195337.5 8157.5 195202.5 ;
      RECT  7902.5 195337.5 7967.5 195202.5 ;
      RECT  8262.5 194407.5 8327.5 194272.5 ;
      RECT  8262.5 195382.5 8327.5 195247.5 ;
      RECT  8097.5 195125.0 7962.5 195060.0 ;
      RECT  7907.5 194985.0 7772.5 194920.0 ;
      RECT  7717.5 194845.0 7582.5 194780.0 ;
      RECT  7712.5 194497.5 7777.5 194362.5 ;
      RECT  8092.5 194497.5 8157.5 194362.5 ;
      RECT  8092.5 195337.5 8157.5 195202.5 ;
      RECT  8092.5 194880.0 8157.5 194745.0 ;
      RECT  7582.5 194845.0 7717.5 194780.0 ;
      RECT  7772.5 194985.0 7907.5 194920.0 ;
      RECT  7962.5 195125.0 8097.5 195060.0 ;
      RECT  8092.5 194880.0 8157.5 194745.0 ;
      RECT  7455.0 194187.5 8465.0 194122.5 ;
      RECT  7455.0 195532.5 8465.0 195467.5 ;
      RECT  7522.5 195662.5 7587.5 195467.5 ;
      RECT  7522.5 196502.5 7587.5 196877.5 ;
      RECT  7902.5 196502.5 7967.5 196877.5 ;
      RECT  8262.5 196660.0 8327.5 196845.0 ;
      RECT  8262.5 195500.0 8327.5 195685.0 ;
      RECT  7522.5 196502.5 7587.5 196637.5 ;
      RECT  7712.5 196502.5 7777.5 196637.5 ;
      RECT  7712.5 196502.5 7777.5 196637.5 ;
      RECT  7522.5 196502.5 7587.5 196637.5 ;
      RECT  7712.5 196502.5 7777.5 196637.5 ;
      RECT  7902.5 196502.5 7967.5 196637.5 ;
      RECT  7902.5 196502.5 7967.5 196637.5 ;
      RECT  7712.5 196502.5 7777.5 196637.5 ;
      RECT  7902.5 196502.5 7967.5 196637.5 ;
      RECT  8092.5 196502.5 8157.5 196637.5 ;
      RECT  8092.5 196502.5 8157.5 196637.5 ;
      RECT  7902.5 196502.5 7967.5 196637.5 ;
      RECT  7522.5 195662.5 7587.5 195797.5 ;
      RECT  7712.5 195662.5 7777.5 195797.5 ;
      RECT  7712.5 195662.5 7777.5 195797.5 ;
      RECT  7522.5 195662.5 7587.5 195797.5 ;
      RECT  7712.5 195662.5 7777.5 195797.5 ;
      RECT  7902.5 195662.5 7967.5 195797.5 ;
      RECT  7902.5 195662.5 7967.5 195797.5 ;
      RECT  7712.5 195662.5 7777.5 195797.5 ;
      RECT  7902.5 195662.5 7967.5 195797.5 ;
      RECT  8092.5 195662.5 8157.5 195797.5 ;
      RECT  8092.5 195662.5 8157.5 195797.5 ;
      RECT  7902.5 195662.5 7967.5 195797.5 ;
      RECT  8262.5 196592.5 8327.5 196727.5 ;
      RECT  8262.5 195617.5 8327.5 195752.5 ;
      RECT  8097.5 195875.0 7962.5 195940.0 ;
      RECT  7907.5 196015.0 7772.5 196080.0 ;
      RECT  7717.5 196155.0 7582.5 196220.0 ;
      RECT  7712.5 196502.5 7777.5 196637.5 ;
      RECT  8092.5 196502.5 8157.5 196637.5 ;
      RECT  8092.5 195662.5 8157.5 195797.5 ;
      RECT  8092.5 196120.0 8157.5 196255.0 ;
      RECT  7582.5 196155.0 7717.5 196220.0 ;
      RECT  7772.5 196015.0 7907.5 196080.0 ;
      RECT  7962.5 195875.0 8097.5 195940.0 ;
      RECT  8092.5 196120.0 8157.5 196255.0 ;
      RECT  7455.0 196812.5 8465.0 196877.5 ;
      RECT  7455.0 195467.5 8465.0 195532.5 ;
      RECT  7522.5 198027.5 7587.5 198222.5 ;
      RECT  7522.5 197187.5 7587.5 196812.5 ;
      RECT  7902.5 197187.5 7967.5 196812.5 ;
      RECT  8262.5 197030.0 8327.5 196845.0 ;
      RECT  8262.5 198190.0 8327.5 198005.0 ;
      RECT  7522.5 197187.5 7587.5 197052.5 ;
      RECT  7712.5 197187.5 7777.5 197052.5 ;
      RECT  7712.5 197187.5 7777.5 197052.5 ;
      RECT  7522.5 197187.5 7587.5 197052.5 ;
      RECT  7712.5 197187.5 7777.5 197052.5 ;
      RECT  7902.5 197187.5 7967.5 197052.5 ;
      RECT  7902.5 197187.5 7967.5 197052.5 ;
      RECT  7712.5 197187.5 7777.5 197052.5 ;
      RECT  7902.5 197187.5 7967.5 197052.5 ;
      RECT  8092.5 197187.5 8157.5 197052.5 ;
      RECT  8092.5 197187.5 8157.5 197052.5 ;
      RECT  7902.5 197187.5 7967.5 197052.5 ;
      RECT  7522.5 198027.5 7587.5 197892.5 ;
      RECT  7712.5 198027.5 7777.5 197892.5 ;
      RECT  7712.5 198027.5 7777.5 197892.5 ;
      RECT  7522.5 198027.5 7587.5 197892.5 ;
      RECT  7712.5 198027.5 7777.5 197892.5 ;
      RECT  7902.5 198027.5 7967.5 197892.5 ;
      RECT  7902.5 198027.5 7967.5 197892.5 ;
      RECT  7712.5 198027.5 7777.5 197892.5 ;
      RECT  7902.5 198027.5 7967.5 197892.5 ;
      RECT  8092.5 198027.5 8157.5 197892.5 ;
      RECT  8092.5 198027.5 8157.5 197892.5 ;
      RECT  7902.5 198027.5 7967.5 197892.5 ;
      RECT  8262.5 197097.5 8327.5 196962.5 ;
      RECT  8262.5 198072.5 8327.5 197937.5 ;
      RECT  8097.5 197815.0 7962.5 197750.0 ;
      RECT  7907.5 197675.0 7772.5 197610.0 ;
      RECT  7717.5 197535.0 7582.5 197470.0 ;
      RECT  7712.5 197187.5 7777.5 197052.5 ;
      RECT  8092.5 197187.5 8157.5 197052.5 ;
      RECT  8092.5 198027.5 8157.5 197892.5 ;
      RECT  8092.5 197570.0 8157.5 197435.0 ;
      RECT  7582.5 197535.0 7717.5 197470.0 ;
      RECT  7772.5 197675.0 7907.5 197610.0 ;
      RECT  7962.5 197815.0 8097.5 197750.0 ;
      RECT  8092.5 197570.0 8157.5 197435.0 ;
      RECT  7455.0 196877.5 8465.0 196812.5 ;
      RECT  7455.0 198222.5 8465.0 198157.5 ;
      RECT  7522.5 198352.5 7587.5 198157.5 ;
      RECT  7522.5 199192.5 7587.5 199567.5 ;
      RECT  7902.5 199192.5 7967.5 199567.5 ;
      RECT  8262.5 199350.0 8327.5 199535.0 ;
      RECT  8262.5 198190.0 8327.5 198375.0 ;
      RECT  7522.5 199192.5 7587.5 199327.5 ;
      RECT  7712.5 199192.5 7777.5 199327.5 ;
      RECT  7712.5 199192.5 7777.5 199327.5 ;
      RECT  7522.5 199192.5 7587.5 199327.5 ;
      RECT  7712.5 199192.5 7777.5 199327.5 ;
      RECT  7902.5 199192.5 7967.5 199327.5 ;
      RECT  7902.5 199192.5 7967.5 199327.5 ;
      RECT  7712.5 199192.5 7777.5 199327.5 ;
      RECT  7902.5 199192.5 7967.5 199327.5 ;
      RECT  8092.5 199192.5 8157.5 199327.5 ;
      RECT  8092.5 199192.5 8157.5 199327.5 ;
      RECT  7902.5 199192.5 7967.5 199327.5 ;
      RECT  7522.5 198352.5 7587.5 198487.5 ;
      RECT  7712.5 198352.5 7777.5 198487.5 ;
      RECT  7712.5 198352.5 7777.5 198487.5 ;
      RECT  7522.5 198352.5 7587.5 198487.5 ;
      RECT  7712.5 198352.5 7777.5 198487.5 ;
      RECT  7902.5 198352.5 7967.5 198487.5 ;
      RECT  7902.5 198352.5 7967.5 198487.5 ;
      RECT  7712.5 198352.5 7777.5 198487.5 ;
      RECT  7902.5 198352.5 7967.5 198487.5 ;
      RECT  8092.5 198352.5 8157.5 198487.5 ;
      RECT  8092.5 198352.5 8157.5 198487.5 ;
      RECT  7902.5 198352.5 7967.5 198487.5 ;
      RECT  8262.5 199282.5 8327.5 199417.5 ;
      RECT  8262.5 198307.5 8327.5 198442.5 ;
      RECT  8097.5 198565.0 7962.5 198630.0 ;
      RECT  7907.5 198705.0 7772.5 198770.0 ;
      RECT  7717.5 198845.0 7582.5 198910.0 ;
      RECT  7712.5 199192.5 7777.5 199327.5 ;
      RECT  8092.5 199192.5 8157.5 199327.5 ;
      RECT  8092.5 198352.5 8157.5 198487.5 ;
      RECT  8092.5 198810.0 8157.5 198945.0 ;
      RECT  7582.5 198845.0 7717.5 198910.0 ;
      RECT  7772.5 198705.0 7907.5 198770.0 ;
      RECT  7962.5 198565.0 8097.5 198630.0 ;
      RECT  8092.5 198810.0 8157.5 198945.0 ;
      RECT  7455.0 199502.5 8465.0 199567.5 ;
      RECT  7455.0 198157.5 8465.0 198222.5 ;
      RECT  7522.5 200717.5 7587.5 200912.5 ;
      RECT  7522.5 199877.5 7587.5 199502.5 ;
      RECT  7902.5 199877.5 7967.5 199502.5 ;
      RECT  8262.5 199720.0 8327.5 199535.0 ;
      RECT  8262.5 200880.0 8327.5 200695.0 ;
      RECT  7522.5 199877.5 7587.5 199742.5 ;
      RECT  7712.5 199877.5 7777.5 199742.5 ;
      RECT  7712.5 199877.5 7777.5 199742.5 ;
      RECT  7522.5 199877.5 7587.5 199742.5 ;
      RECT  7712.5 199877.5 7777.5 199742.5 ;
      RECT  7902.5 199877.5 7967.5 199742.5 ;
      RECT  7902.5 199877.5 7967.5 199742.5 ;
      RECT  7712.5 199877.5 7777.5 199742.5 ;
      RECT  7902.5 199877.5 7967.5 199742.5 ;
      RECT  8092.5 199877.5 8157.5 199742.5 ;
      RECT  8092.5 199877.5 8157.5 199742.5 ;
      RECT  7902.5 199877.5 7967.5 199742.5 ;
      RECT  7522.5 200717.5 7587.5 200582.5 ;
      RECT  7712.5 200717.5 7777.5 200582.5 ;
      RECT  7712.5 200717.5 7777.5 200582.5 ;
      RECT  7522.5 200717.5 7587.5 200582.5 ;
      RECT  7712.5 200717.5 7777.5 200582.5 ;
      RECT  7902.5 200717.5 7967.5 200582.5 ;
      RECT  7902.5 200717.5 7967.5 200582.5 ;
      RECT  7712.5 200717.5 7777.5 200582.5 ;
      RECT  7902.5 200717.5 7967.5 200582.5 ;
      RECT  8092.5 200717.5 8157.5 200582.5 ;
      RECT  8092.5 200717.5 8157.5 200582.5 ;
      RECT  7902.5 200717.5 7967.5 200582.5 ;
      RECT  8262.5 199787.5 8327.5 199652.5 ;
      RECT  8262.5 200762.5 8327.5 200627.5 ;
      RECT  8097.5 200505.0 7962.5 200440.0 ;
      RECT  7907.5 200365.0 7772.5 200300.0 ;
      RECT  7717.5 200225.0 7582.5 200160.0 ;
      RECT  7712.5 199877.5 7777.5 199742.5 ;
      RECT  8092.5 199877.5 8157.5 199742.5 ;
      RECT  8092.5 200717.5 8157.5 200582.5 ;
      RECT  8092.5 200260.0 8157.5 200125.0 ;
      RECT  7582.5 200225.0 7717.5 200160.0 ;
      RECT  7772.5 200365.0 7907.5 200300.0 ;
      RECT  7962.5 200505.0 8097.5 200440.0 ;
      RECT  8092.5 200260.0 8157.5 200125.0 ;
      RECT  7455.0 199567.5 8465.0 199502.5 ;
      RECT  7455.0 200912.5 8465.0 200847.5 ;
      RECT  7522.5 201042.5 7587.5 200847.5 ;
      RECT  7522.5 201882.5 7587.5 202257.5 ;
      RECT  7902.5 201882.5 7967.5 202257.5 ;
      RECT  8262.5 202040.0 8327.5 202225.0 ;
      RECT  8262.5 200880.0 8327.5 201065.0 ;
      RECT  7522.5 201882.5 7587.5 202017.5 ;
      RECT  7712.5 201882.5 7777.5 202017.5 ;
      RECT  7712.5 201882.5 7777.5 202017.5 ;
      RECT  7522.5 201882.5 7587.5 202017.5 ;
      RECT  7712.5 201882.5 7777.5 202017.5 ;
      RECT  7902.5 201882.5 7967.5 202017.5 ;
      RECT  7902.5 201882.5 7967.5 202017.5 ;
      RECT  7712.5 201882.5 7777.5 202017.5 ;
      RECT  7902.5 201882.5 7967.5 202017.5 ;
      RECT  8092.5 201882.5 8157.5 202017.5 ;
      RECT  8092.5 201882.5 8157.5 202017.5 ;
      RECT  7902.5 201882.5 7967.5 202017.5 ;
      RECT  7522.5 201042.5 7587.5 201177.5 ;
      RECT  7712.5 201042.5 7777.5 201177.5 ;
      RECT  7712.5 201042.5 7777.5 201177.5 ;
      RECT  7522.5 201042.5 7587.5 201177.5 ;
      RECT  7712.5 201042.5 7777.5 201177.5 ;
      RECT  7902.5 201042.5 7967.5 201177.5 ;
      RECT  7902.5 201042.5 7967.5 201177.5 ;
      RECT  7712.5 201042.5 7777.5 201177.5 ;
      RECT  7902.5 201042.5 7967.5 201177.5 ;
      RECT  8092.5 201042.5 8157.5 201177.5 ;
      RECT  8092.5 201042.5 8157.5 201177.5 ;
      RECT  7902.5 201042.5 7967.5 201177.5 ;
      RECT  8262.5 201972.5 8327.5 202107.5 ;
      RECT  8262.5 200997.5 8327.5 201132.5 ;
      RECT  8097.5 201255.0 7962.5 201320.0 ;
      RECT  7907.5 201395.0 7772.5 201460.0 ;
      RECT  7717.5 201535.0 7582.5 201600.0 ;
      RECT  7712.5 201882.5 7777.5 202017.5 ;
      RECT  8092.5 201882.5 8157.5 202017.5 ;
      RECT  8092.5 201042.5 8157.5 201177.5 ;
      RECT  8092.5 201500.0 8157.5 201635.0 ;
      RECT  7582.5 201535.0 7717.5 201600.0 ;
      RECT  7772.5 201395.0 7907.5 201460.0 ;
      RECT  7962.5 201255.0 8097.5 201320.0 ;
      RECT  8092.5 201500.0 8157.5 201635.0 ;
      RECT  7455.0 202192.5 8465.0 202257.5 ;
      RECT  7455.0 200847.5 8465.0 200912.5 ;
      RECT  7522.5 203407.5 7587.5 203602.5 ;
      RECT  7522.5 202567.5 7587.5 202192.5 ;
      RECT  7902.5 202567.5 7967.5 202192.5 ;
      RECT  8262.5 202410.0 8327.5 202225.0 ;
      RECT  8262.5 203570.0 8327.5 203385.0 ;
      RECT  7522.5 202567.5 7587.5 202432.5 ;
      RECT  7712.5 202567.5 7777.5 202432.5 ;
      RECT  7712.5 202567.5 7777.5 202432.5 ;
      RECT  7522.5 202567.5 7587.5 202432.5 ;
      RECT  7712.5 202567.5 7777.5 202432.5 ;
      RECT  7902.5 202567.5 7967.5 202432.5 ;
      RECT  7902.5 202567.5 7967.5 202432.5 ;
      RECT  7712.5 202567.5 7777.5 202432.5 ;
      RECT  7902.5 202567.5 7967.5 202432.5 ;
      RECT  8092.5 202567.5 8157.5 202432.5 ;
      RECT  8092.5 202567.5 8157.5 202432.5 ;
      RECT  7902.5 202567.5 7967.5 202432.5 ;
      RECT  7522.5 203407.5 7587.5 203272.5 ;
      RECT  7712.5 203407.5 7777.5 203272.5 ;
      RECT  7712.5 203407.5 7777.5 203272.5 ;
      RECT  7522.5 203407.5 7587.5 203272.5 ;
      RECT  7712.5 203407.5 7777.5 203272.5 ;
      RECT  7902.5 203407.5 7967.5 203272.5 ;
      RECT  7902.5 203407.5 7967.5 203272.5 ;
      RECT  7712.5 203407.5 7777.5 203272.5 ;
      RECT  7902.5 203407.5 7967.5 203272.5 ;
      RECT  8092.5 203407.5 8157.5 203272.5 ;
      RECT  8092.5 203407.5 8157.5 203272.5 ;
      RECT  7902.5 203407.5 7967.5 203272.5 ;
      RECT  8262.5 202477.5 8327.5 202342.5 ;
      RECT  8262.5 203452.5 8327.5 203317.5 ;
      RECT  8097.5 203195.0 7962.5 203130.0 ;
      RECT  7907.5 203055.0 7772.5 202990.0 ;
      RECT  7717.5 202915.0 7582.5 202850.0 ;
      RECT  7712.5 202567.5 7777.5 202432.5 ;
      RECT  8092.5 202567.5 8157.5 202432.5 ;
      RECT  8092.5 203407.5 8157.5 203272.5 ;
      RECT  8092.5 202950.0 8157.5 202815.0 ;
      RECT  7582.5 202915.0 7717.5 202850.0 ;
      RECT  7772.5 203055.0 7907.5 202990.0 ;
      RECT  7962.5 203195.0 8097.5 203130.0 ;
      RECT  8092.5 202950.0 8157.5 202815.0 ;
      RECT  7455.0 202257.5 8465.0 202192.5 ;
      RECT  7455.0 203602.5 8465.0 203537.5 ;
      RECT  7522.5 203732.5 7587.5 203537.5 ;
      RECT  7522.5 204572.5 7587.5 204947.5 ;
      RECT  7902.5 204572.5 7967.5 204947.5 ;
      RECT  8262.5 204730.0 8327.5 204915.0 ;
      RECT  8262.5 203570.0 8327.5 203755.0 ;
      RECT  7522.5 204572.5 7587.5 204707.5 ;
      RECT  7712.5 204572.5 7777.5 204707.5 ;
      RECT  7712.5 204572.5 7777.5 204707.5 ;
      RECT  7522.5 204572.5 7587.5 204707.5 ;
      RECT  7712.5 204572.5 7777.5 204707.5 ;
      RECT  7902.5 204572.5 7967.5 204707.5 ;
      RECT  7902.5 204572.5 7967.5 204707.5 ;
      RECT  7712.5 204572.5 7777.5 204707.5 ;
      RECT  7902.5 204572.5 7967.5 204707.5 ;
      RECT  8092.5 204572.5 8157.5 204707.5 ;
      RECT  8092.5 204572.5 8157.5 204707.5 ;
      RECT  7902.5 204572.5 7967.5 204707.5 ;
      RECT  7522.5 203732.5 7587.5 203867.5 ;
      RECT  7712.5 203732.5 7777.5 203867.5 ;
      RECT  7712.5 203732.5 7777.5 203867.5 ;
      RECT  7522.5 203732.5 7587.5 203867.5 ;
      RECT  7712.5 203732.5 7777.5 203867.5 ;
      RECT  7902.5 203732.5 7967.5 203867.5 ;
      RECT  7902.5 203732.5 7967.5 203867.5 ;
      RECT  7712.5 203732.5 7777.5 203867.5 ;
      RECT  7902.5 203732.5 7967.5 203867.5 ;
      RECT  8092.5 203732.5 8157.5 203867.5 ;
      RECT  8092.5 203732.5 8157.5 203867.5 ;
      RECT  7902.5 203732.5 7967.5 203867.5 ;
      RECT  8262.5 204662.5 8327.5 204797.5 ;
      RECT  8262.5 203687.5 8327.5 203822.5 ;
      RECT  8097.5 203945.0 7962.5 204010.0 ;
      RECT  7907.5 204085.0 7772.5 204150.0 ;
      RECT  7717.5 204225.0 7582.5 204290.0 ;
      RECT  7712.5 204572.5 7777.5 204707.5 ;
      RECT  8092.5 204572.5 8157.5 204707.5 ;
      RECT  8092.5 203732.5 8157.5 203867.5 ;
      RECT  8092.5 204190.0 8157.5 204325.0 ;
      RECT  7582.5 204225.0 7717.5 204290.0 ;
      RECT  7772.5 204085.0 7907.5 204150.0 ;
      RECT  7962.5 203945.0 8097.5 204010.0 ;
      RECT  8092.5 204190.0 8157.5 204325.0 ;
      RECT  7455.0 204882.5 8465.0 204947.5 ;
      RECT  7455.0 203537.5 8465.0 203602.5 ;
      RECT  7522.5 206097.5 7587.5 206292.5 ;
      RECT  7522.5 205257.5 7587.5 204882.5 ;
      RECT  7902.5 205257.5 7967.5 204882.5 ;
      RECT  8262.5 205100.0 8327.5 204915.0 ;
      RECT  8262.5 206260.0 8327.5 206075.0 ;
      RECT  7522.5 205257.5 7587.5 205122.5 ;
      RECT  7712.5 205257.5 7777.5 205122.5 ;
      RECT  7712.5 205257.5 7777.5 205122.5 ;
      RECT  7522.5 205257.5 7587.5 205122.5 ;
      RECT  7712.5 205257.5 7777.5 205122.5 ;
      RECT  7902.5 205257.5 7967.5 205122.5 ;
      RECT  7902.5 205257.5 7967.5 205122.5 ;
      RECT  7712.5 205257.5 7777.5 205122.5 ;
      RECT  7902.5 205257.5 7967.5 205122.5 ;
      RECT  8092.5 205257.5 8157.5 205122.5 ;
      RECT  8092.5 205257.5 8157.5 205122.5 ;
      RECT  7902.5 205257.5 7967.5 205122.5 ;
      RECT  7522.5 206097.5 7587.5 205962.5 ;
      RECT  7712.5 206097.5 7777.5 205962.5 ;
      RECT  7712.5 206097.5 7777.5 205962.5 ;
      RECT  7522.5 206097.5 7587.5 205962.5 ;
      RECT  7712.5 206097.5 7777.5 205962.5 ;
      RECT  7902.5 206097.5 7967.5 205962.5 ;
      RECT  7902.5 206097.5 7967.5 205962.5 ;
      RECT  7712.5 206097.5 7777.5 205962.5 ;
      RECT  7902.5 206097.5 7967.5 205962.5 ;
      RECT  8092.5 206097.5 8157.5 205962.5 ;
      RECT  8092.5 206097.5 8157.5 205962.5 ;
      RECT  7902.5 206097.5 7967.5 205962.5 ;
      RECT  8262.5 205167.5 8327.5 205032.5 ;
      RECT  8262.5 206142.5 8327.5 206007.5 ;
      RECT  8097.5 205885.0 7962.5 205820.0 ;
      RECT  7907.5 205745.0 7772.5 205680.0 ;
      RECT  7717.5 205605.0 7582.5 205540.0 ;
      RECT  7712.5 205257.5 7777.5 205122.5 ;
      RECT  8092.5 205257.5 8157.5 205122.5 ;
      RECT  8092.5 206097.5 8157.5 205962.5 ;
      RECT  8092.5 205640.0 8157.5 205505.0 ;
      RECT  7582.5 205605.0 7717.5 205540.0 ;
      RECT  7772.5 205745.0 7907.5 205680.0 ;
      RECT  7962.5 205885.0 8097.5 205820.0 ;
      RECT  8092.5 205640.0 8157.5 205505.0 ;
      RECT  7455.0 204947.5 8465.0 204882.5 ;
      RECT  7455.0 206292.5 8465.0 206227.5 ;
      RECT  8892.5 35260.0 8957.5 35445.0 ;
      RECT  8892.5 34100.0 8957.5 34285.0 ;
      RECT  8532.5 34217.5 8597.5 34067.5 ;
      RECT  8532.5 35102.5 8597.5 35477.5 ;
      RECT  8722.5 34217.5 8787.5 35102.5 ;
      RECT  8532.5 35102.5 8597.5 35237.5 ;
      RECT  8722.5 35102.5 8787.5 35237.5 ;
      RECT  8722.5 35102.5 8787.5 35237.5 ;
      RECT  8532.5 35102.5 8597.5 35237.5 ;
      RECT  8532.5 34217.5 8597.5 34352.5 ;
      RECT  8722.5 34217.5 8787.5 34352.5 ;
      RECT  8722.5 34217.5 8787.5 34352.5 ;
      RECT  8532.5 34217.5 8597.5 34352.5 ;
      RECT  8892.5 35192.5 8957.5 35327.5 ;
      RECT  8892.5 34217.5 8957.5 34352.5 ;
      RECT  8590.0 34660.0 8655.0 34795.0 ;
      RECT  8590.0 34660.0 8655.0 34795.0 ;
      RECT  8755.0 34695.0 8820.0 34760.0 ;
      RECT  8465.0 35412.5 9025.0 35477.5 ;
      RECT  8465.0 34067.5 9025.0 34132.5 ;
      RECT  8892.5 35630.0 8957.5 35445.0 ;
      RECT  8892.5 36790.0 8957.5 36605.0 ;
      RECT  8532.5 36672.5 8597.5 36822.5 ;
      RECT  8532.5 35787.5 8597.5 35412.5 ;
      RECT  8722.5 36672.5 8787.5 35787.5 ;
      RECT  8532.5 35787.5 8597.5 35652.5 ;
      RECT  8722.5 35787.5 8787.5 35652.5 ;
      RECT  8722.5 35787.5 8787.5 35652.5 ;
      RECT  8532.5 35787.5 8597.5 35652.5 ;
      RECT  8532.5 36672.5 8597.5 36537.5 ;
      RECT  8722.5 36672.5 8787.5 36537.5 ;
      RECT  8722.5 36672.5 8787.5 36537.5 ;
      RECT  8532.5 36672.5 8597.5 36537.5 ;
      RECT  8892.5 35697.5 8957.5 35562.5 ;
      RECT  8892.5 36672.5 8957.5 36537.5 ;
      RECT  8590.0 36230.0 8655.0 36095.0 ;
      RECT  8590.0 36230.0 8655.0 36095.0 ;
      RECT  8755.0 36195.0 8820.0 36130.0 ;
      RECT  8465.0 35477.5 9025.0 35412.5 ;
      RECT  8465.0 36822.5 9025.0 36757.5 ;
      RECT  8892.5 37950.0 8957.5 38135.0 ;
      RECT  8892.5 36790.0 8957.5 36975.0 ;
      RECT  8532.5 36907.5 8597.5 36757.5 ;
      RECT  8532.5 37792.5 8597.5 38167.5 ;
      RECT  8722.5 36907.5 8787.5 37792.5 ;
      RECT  8532.5 37792.5 8597.5 37927.5 ;
      RECT  8722.5 37792.5 8787.5 37927.5 ;
      RECT  8722.5 37792.5 8787.5 37927.5 ;
      RECT  8532.5 37792.5 8597.5 37927.5 ;
      RECT  8532.5 36907.5 8597.5 37042.5 ;
      RECT  8722.5 36907.5 8787.5 37042.5 ;
      RECT  8722.5 36907.5 8787.5 37042.5 ;
      RECT  8532.5 36907.5 8597.5 37042.5 ;
      RECT  8892.5 37882.5 8957.5 38017.5 ;
      RECT  8892.5 36907.5 8957.5 37042.5 ;
      RECT  8590.0 37350.0 8655.0 37485.0 ;
      RECT  8590.0 37350.0 8655.0 37485.0 ;
      RECT  8755.0 37385.0 8820.0 37450.0 ;
      RECT  8465.0 38102.5 9025.0 38167.5 ;
      RECT  8465.0 36757.5 9025.0 36822.5 ;
      RECT  8892.5 38320.0 8957.5 38135.0 ;
      RECT  8892.5 39480.0 8957.5 39295.0 ;
      RECT  8532.5 39362.5 8597.5 39512.5 ;
      RECT  8532.5 38477.5 8597.5 38102.5 ;
      RECT  8722.5 39362.5 8787.5 38477.5 ;
      RECT  8532.5 38477.5 8597.5 38342.5 ;
      RECT  8722.5 38477.5 8787.5 38342.5 ;
      RECT  8722.5 38477.5 8787.5 38342.5 ;
      RECT  8532.5 38477.5 8597.5 38342.5 ;
      RECT  8532.5 39362.5 8597.5 39227.5 ;
      RECT  8722.5 39362.5 8787.5 39227.5 ;
      RECT  8722.5 39362.5 8787.5 39227.5 ;
      RECT  8532.5 39362.5 8597.5 39227.5 ;
      RECT  8892.5 38387.5 8957.5 38252.5 ;
      RECT  8892.5 39362.5 8957.5 39227.5 ;
      RECT  8590.0 38920.0 8655.0 38785.0 ;
      RECT  8590.0 38920.0 8655.0 38785.0 ;
      RECT  8755.0 38885.0 8820.0 38820.0 ;
      RECT  8465.0 38167.5 9025.0 38102.5 ;
      RECT  8465.0 39512.5 9025.0 39447.5 ;
      RECT  8892.5 40640.0 8957.5 40825.0 ;
      RECT  8892.5 39480.0 8957.5 39665.0 ;
      RECT  8532.5 39597.5 8597.5 39447.5 ;
      RECT  8532.5 40482.5 8597.5 40857.5 ;
      RECT  8722.5 39597.5 8787.5 40482.5 ;
      RECT  8532.5 40482.5 8597.5 40617.5 ;
      RECT  8722.5 40482.5 8787.5 40617.5 ;
      RECT  8722.5 40482.5 8787.5 40617.5 ;
      RECT  8532.5 40482.5 8597.5 40617.5 ;
      RECT  8532.5 39597.5 8597.5 39732.5 ;
      RECT  8722.5 39597.5 8787.5 39732.5 ;
      RECT  8722.5 39597.5 8787.5 39732.5 ;
      RECT  8532.5 39597.5 8597.5 39732.5 ;
      RECT  8892.5 40572.5 8957.5 40707.5 ;
      RECT  8892.5 39597.5 8957.5 39732.5 ;
      RECT  8590.0 40040.0 8655.0 40175.0 ;
      RECT  8590.0 40040.0 8655.0 40175.0 ;
      RECT  8755.0 40075.0 8820.0 40140.0 ;
      RECT  8465.0 40792.5 9025.0 40857.5 ;
      RECT  8465.0 39447.5 9025.0 39512.5 ;
      RECT  8892.5 41010.0 8957.5 40825.0 ;
      RECT  8892.5 42170.0 8957.5 41985.0 ;
      RECT  8532.5 42052.5 8597.5 42202.5 ;
      RECT  8532.5 41167.5 8597.5 40792.5 ;
      RECT  8722.5 42052.5 8787.5 41167.5 ;
      RECT  8532.5 41167.5 8597.5 41032.5 ;
      RECT  8722.5 41167.5 8787.5 41032.5 ;
      RECT  8722.5 41167.5 8787.5 41032.5 ;
      RECT  8532.5 41167.5 8597.5 41032.5 ;
      RECT  8532.5 42052.5 8597.5 41917.5 ;
      RECT  8722.5 42052.5 8787.5 41917.5 ;
      RECT  8722.5 42052.5 8787.5 41917.5 ;
      RECT  8532.5 42052.5 8597.5 41917.5 ;
      RECT  8892.5 41077.5 8957.5 40942.5 ;
      RECT  8892.5 42052.5 8957.5 41917.5 ;
      RECT  8590.0 41610.0 8655.0 41475.0 ;
      RECT  8590.0 41610.0 8655.0 41475.0 ;
      RECT  8755.0 41575.0 8820.0 41510.0 ;
      RECT  8465.0 40857.5 9025.0 40792.5 ;
      RECT  8465.0 42202.5 9025.0 42137.5 ;
      RECT  8892.5 43330.0 8957.5 43515.0 ;
      RECT  8892.5 42170.0 8957.5 42355.0 ;
      RECT  8532.5 42287.5 8597.5 42137.5 ;
      RECT  8532.5 43172.5 8597.5 43547.5 ;
      RECT  8722.5 42287.5 8787.5 43172.5 ;
      RECT  8532.5 43172.5 8597.5 43307.5 ;
      RECT  8722.5 43172.5 8787.5 43307.5 ;
      RECT  8722.5 43172.5 8787.5 43307.5 ;
      RECT  8532.5 43172.5 8597.5 43307.5 ;
      RECT  8532.5 42287.5 8597.5 42422.5 ;
      RECT  8722.5 42287.5 8787.5 42422.5 ;
      RECT  8722.5 42287.5 8787.5 42422.5 ;
      RECT  8532.5 42287.5 8597.5 42422.5 ;
      RECT  8892.5 43262.5 8957.5 43397.5 ;
      RECT  8892.5 42287.5 8957.5 42422.5 ;
      RECT  8590.0 42730.0 8655.0 42865.0 ;
      RECT  8590.0 42730.0 8655.0 42865.0 ;
      RECT  8755.0 42765.0 8820.0 42830.0 ;
      RECT  8465.0 43482.5 9025.0 43547.5 ;
      RECT  8465.0 42137.5 9025.0 42202.5 ;
      RECT  8892.5 43700.0 8957.5 43515.0 ;
      RECT  8892.5 44860.0 8957.5 44675.0 ;
      RECT  8532.5 44742.5 8597.5 44892.5 ;
      RECT  8532.5 43857.5 8597.5 43482.5 ;
      RECT  8722.5 44742.5 8787.5 43857.5 ;
      RECT  8532.5 43857.5 8597.5 43722.5 ;
      RECT  8722.5 43857.5 8787.5 43722.5 ;
      RECT  8722.5 43857.5 8787.5 43722.5 ;
      RECT  8532.5 43857.5 8597.5 43722.5 ;
      RECT  8532.5 44742.5 8597.5 44607.5 ;
      RECT  8722.5 44742.5 8787.5 44607.5 ;
      RECT  8722.5 44742.5 8787.5 44607.5 ;
      RECT  8532.5 44742.5 8597.5 44607.5 ;
      RECT  8892.5 43767.5 8957.5 43632.5 ;
      RECT  8892.5 44742.5 8957.5 44607.5 ;
      RECT  8590.0 44300.0 8655.0 44165.0 ;
      RECT  8590.0 44300.0 8655.0 44165.0 ;
      RECT  8755.0 44265.0 8820.0 44200.0 ;
      RECT  8465.0 43547.5 9025.0 43482.5 ;
      RECT  8465.0 44892.5 9025.0 44827.5 ;
      RECT  8892.5 46020.0 8957.5 46205.0 ;
      RECT  8892.5 44860.0 8957.5 45045.0 ;
      RECT  8532.5 44977.5 8597.5 44827.5 ;
      RECT  8532.5 45862.5 8597.5 46237.5 ;
      RECT  8722.5 44977.5 8787.5 45862.5 ;
      RECT  8532.5 45862.5 8597.5 45997.5 ;
      RECT  8722.5 45862.5 8787.5 45997.5 ;
      RECT  8722.5 45862.5 8787.5 45997.5 ;
      RECT  8532.5 45862.5 8597.5 45997.5 ;
      RECT  8532.5 44977.5 8597.5 45112.5 ;
      RECT  8722.5 44977.5 8787.5 45112.5 ;
      RECT  8722.5 44977.5 8787.5 45112.5 ;
      RECT  8532.5 44977.5 8597.5 45112.5 ;
      RECT  8892.5 45952.5 8957.5 46087.5 ;
      RECT  8892.5 44977.5 8957.5 45112.5 ;
      RECT  8590.0 45420.0 8655.0 45555.0 ;
      RECT  8590.0 45420.0 8655.0 45555.0 ;
      RECT  8755.0 45455.0 8820.0 45520.0 ;
      RECT  8465.0 46172.5 9025.0 46237.5 ;
      RECT  8465.0 44827.5 9025.0 44892.5 ;
      RECT  8892.5 46390.0 8957.5 46205.0 ;
      RECT  8892.5 47550.0 8957.5 47365.0 ;
      RECT  8532.5 47432.5 8597.5 47582.5 ;
      RECT  8532.5 46547.5 8597.5 46172.5 ;
      RECT  8722.5 47432.5 8787.5 46547.5 ;
      RECT  8532.5 46547.5 8597.5 46412.5 ;
      RECT  8722.5 46547.5 8787.5 46412.5 ;
      RECT  8722.5 46547.5 8787.5 46412.5 ;
      RECT  8532.5 46547.5 8597.5 46412.5 ;
      RECT  8532.5 47432.5 8597.5 47297.5 ;
      RECT  8722.5 47432.5 8787.5 47297.5 ;
      RECT  8722.5 47432.5 8787.5 47297.5 ;
      RECT  8532.5 47432.5 8597.5 47297.5 ;
      RECT  8892.5 46457.5 8957.5 46322.5 ;
      RECT  8892.5 47432.5 8957.5 47297.5 ;
      RECT  8590.0 46990.0 8655.0 46855.0 ;
      RECT  8590.0 46990.0 8655.0 46855.0 ;
      RECT  8755.0 46955.0 8820.0 46890.0 ;
      RECT  8465.0 46237.5 9025.0 46172.5 ;
      RECT  8465.0 47582.5 9025.0 47517.5 ;
      RECT  8892.5 48710.0 8957.5 48895.0 ;
      RECT  8892.5 47550.0 8957.5 47735.0 ;
      RECT  8532.5 47667.5 8597.5 47517.5 ;
      RECT  8532.5 48552.5 8597.5 48927.5 ;
      RECT  8722.5 47667.5 8787.5 48552.5 ;
      RECT  8532.5 48552.5 8597.5 48687.5 ;
      RECT  8722.5 48552.5 8787.5 48687.5 ;
      RECT  8722.5 48552.5 8787.5 48687.5 ;
      RECT  8532.5 48552.5 8597.5 48687.5 ;
      RECT  8532.5 47667.5 8597.5 47802.5 ;
      RECT  8722.5 47667.5 8787.5 47802.5 ;
      RECT  8722.5 47667.5 8787.5 47802.5 ;
      RECT  8532.5 47667.5 8597.5 47802.5 ;
      RECT  8892.5 48642.5 8957.5 48777.5 ;
      RECT  8892.5 47667.5 8957.5 47802.5 ;
      RECT  8590.0 48110.0 8655.0 48245.0 ;
      RECT  8590.0 48110.0 8655.0 48245.0 ;
      RECT  8755.0 48145.0 8820.0 48210.0 ;
      RECT  8465.0 48862.5 9025.0 48927.5 ;
      RECT  8465.0 47517.5 9025.0 47582.5 ;
      RECT  8892.5 49080.0 8957.5 48895.0 ;
      RECT  8892.5 50240.0 8957.5 50055.0 ;
      RECT  8532.5 50122.5 8597.5 50272.5 ;
      RECT  8532.5 49237.5 8597.5 48862.5 ;
      RECT  8722.5 50122.5 8787.5 49237.5 ;
      RECT  8532.5 49237.5 8597.5 49102.5 ;
      RECT  8722.5 49237.5 8787.5 49102.5 ;
      RECT  8722.5 49237.5 8787.5 49102.5 ;
      RECT  8532.5 49237.5 8597.5 49102.5 ;
      RECT  8532.5 50122.5 8597.5 49987.5 ;
      RECT  8722.5 50122.5 8787.5 49987.5 ;
      RECT  8722.5 50122.5 8787.5 49987.5 ;
      RECT  8532.5 50122.5 8597.5 49987.5 ;
      RECT  8892.5 49147.5 8957.5 49012.5 ;
      RECT  8892.5 50122.5 8957.5 49987.5 ;
      RECT  8590.0 49680.0 8655.0 49545.0 ;
      RECT  8590.0 49680.0 8655.0 49545.0 ;
      RECT  8755.0 49645.0 8820.0 49580.0 ;
      RECT  8465.0 48927.5 9025.0 48862.5 ;
      RECT  8465.0 50272.5 9025.0 50207.5 ;
      RECT  8892.5 51400.0 8957.5 51585.0 ;
      RECT  8892.5 50240.0 8957.5 50425.0 ;
      RECT  8532.5 50357.5 8597.5 50207.5 ;
      RECT  8532.5 51242.5 8597.5 51617.5 ;
      RECT  8722.5 50357.5 8787.5 51242.5 ;
      RECT  8532.5 51242.5 8597.5 51377.5 ;
      RECT  8722.5 51242.5 8787.5 51377.5 ;
      RECT  8722.5 51242.5 8787.5 51377.5 ;
      RECT  8532.5 51242.5 8597.5 51377.5 ;
      RECT  8532.5 50357.5 8597.5 50492.5 ;
      RECT  8722.5 50357.5 8787.5 50492.5 ;
      RECT  8722.5 50357.5 8787.5 50492.5 ;
      RECT  8532.5 50357.5 8597.5 50492.5 ;
      RECT  8892.5 51332.5 8957.5 51467.5 ;
      RECT  8892.5 50357.5 8957.5 50492.5 ;
      RECT  8590.0 50800.0 8655.0 50935.0 ;
      RECT  8590.0 50800.0 8655.0 50935.0 ;
      RECT  8755.0 50835.0 8820.0 50900.0 ;
      RECT  8465.0 51552.5 9025.0 51617.5 ;
      RECT  8465.0 50207.5 9025.0 50272.5 ;
      RECT  8892.5 51770.0 8957.5 51585.0 ;
      RECT  8892.5 52930.0 8957.5 52745.0 ;
      RECT  8532.5 52812.5 8597.5 52962.5 ;
      RECT  8532.5 51927.5 8597.5 51552.5 ;
      RECT  8722.5 52812.5 8787.5 51927.5 ;
      RECT  8532.5 51927.5 8597.5 51792.5 ;
      RECT  8722.5 51927.5 8787.5 51792.5 ;
      RECT  8722.5 51927.5 8787.5 51792.5 ;
      RECT  8532.5 51927.5 8597.5 51792.5 ;
      RECT  8532.5 52812.5 8597.5 52677.5 ;
      RECT  8722.5 52812.5 8787.5 52677.5 ;
      RECT  8722.5 52812.5 8787.5 52677.5 ;
      RECT  8532.5 52812.5 8597.5 52677.5 ;
      RECT  8892.5 51837.5 8957.5 51702.5 ;
      RECT  8892.5 52812.5 8957.5 52677.5 ;
      RECT  8590.0 52370.0 8655.0 52235.0 ;
      RECT  8590.0 52370.0 8655.0 52235.0 ;
      RECT  8755.0 52335.0 8820.0 52270.0 ;
      RECT  8465.0 51617.5 9025.0 51552.5 ;
      RECT  8465.0 52962.5 9025.0 52897.5 ;
      RECT  8892.5 54090.0 8957.5 54275.0 ;
      RECT  8892.5 52930.0 8957.5 53115.0 ;
      RECT  8532.5 53047.5 8597.5 52897.5 ;
      RECT  8532.5 53932.5 8597.5 54307.5 ;
      RECT  8722.5 53047.5 8787.5 53932.5 ;
      RECT  8532.5 53932.5 8597.5 54067.5 ;
      RECT  8722.5 53932.5 8787.5 54067.5 ;
      RECT  8722.5 53932.5 8787.5 54067.5 ;
      RECT  8532.5 53932.5 8597.5 54067.5 ;
      RECT  8532.5 53047.5 8597.5 53182.5 ;
      RECT  8722.5 53047.5 8787.5 53182.5 ;
      RECT  8722.5 53047.5 8787.5 53182.5 ;
      RECT  8532.5 53047.5 8597.5 53182.5 ;
      RECT  8892.5 54022.5 8957.5 54157.5 ;
      RECT  8892.5 53047.5 8957.5 53182.5 ;
      RECT  8590.0 53490.0 8655.0 53625.0 ;
      RECT  8590.0 53490.0 8655.0 53625.0 ;
      RECT  8755.0 53525.0 8820.0 53590.0 ;
      RECT  8465.0 54242.5 9025.0 54307.5 ;
      RECT  8465.0 52897.5 9025.0 52962.5 ;
      RECT  8892.5 54460.0 8957.5 54275.0 ;
      RECT  8892.5 55620.0 8957.5 55435.0 ;
      RECT  8532.5 55502.5 8597.5 55652.5 ;
      RECT  8532.5 54617.5 8597.5 54242.5 ;
      RECT  8722.5 55502.5 8787.5 54617.5 ;
      RECT  8532.5 54617.5 8597.5 54482.5 ;
      RECT  8722.5 54617.5 8787.5 54482.5 ;
      RECT  8722.5 54617.5 8787.5 54482.5 ;
      RECT  8532.5 54617.5 8597.5 54482.5 ;
      RECT  8532.5 55502.5 8597.5 55367.5 ;
      RECT  8722.5 55502.5 8787.5 55367.5 ;
      RECT  8722.5 55502.5 8787.5 55367.5 ;
      RECT  8532.5 55502.5 8597.5 55367.5 ;
      RECT  8892.5 54527.5 8957.5 54392.5 ;
      RECT  8892.5 55502.5 8957.5 55367.5 ;
      RECT  8590.0 55060.0 8655.0 54925.0 ;
      RECT  8590.0 55060.0 8655.0 54925.0 ;
      RECT  8755.0 55025.0 8820.0 54960.0 ;
      RECT  8465.0 54307.5 9025.0 54242.5 ;
      RECT  8465.0 55652.5 9025.0 55587.5 ;
      RECT  8892.5 56780.0 8957.5 56965.0 ;
      RECT  8892.5 55620.0 8957.5 55805.0 ;
      RECT  8532.5 55737.5 8597.5 55587.5 ;
      RECT  8532.5 56622.5 8597.5 56997.5 ;
      RECT  8722.5 55737.5 8787.5 56622.5 ;
      RECT  8532.5 56622.5 8597.5 56757.5 ;
      RECT  8722.5 56622.5 8787.5 56757.5 ;
      RECT  8722.5 56622.5 8787.5 56757.5 ;
      RECT  8532.5 56622.5 8597.5 56757.5 ;
      RECT  8532.5 55737.5 8597.5 55872.5 ;
      RECT  8722.5 55737.5 8787.5 55872.5 ;
      RECT  8722.5 55737.5 8787.5 55872.5 ;
      RECT  8532.5 55737.5 8597.5 55872.5 ;
      RECT  8892.5 56712.5 8957.5 56847.5 ;
      RECT  8892.5 55737.5 8957.5 55872.5 ;
      RECT  8590.0 56180.0 8655.0 56315.0 ;
      RECT  8590.0 56180.0 8655.0 56315.0 ;
      RECT  8755.0 56215.0 8820.0 56280.0 ;
      RECT  8465.0 56932.5 9025.0 56997.5 ;
      RECT  8465.0 55587.5 9025.0 55652.5 ;
      RECT  8892.5 57150.0 8957.5 56965.0 ;
      RECT  8892.5 58310.0 8957.5 58125.0 ;
      RECT  8532.5 58192.5 8597.5 58342.5 ;
      RECT  8532.5 57307.5 8597.5 56932.5 ;
      RECT  8722.5 58192.5 8787.5 57307.5 ;
      RECT  8532.5 57307.5 8597.5 57172.5 ;
      RECT  8722.5 57307.5 8787.5 57172.5 ;
      RECT  8722.5 57307.5 8787.5 57172.5 ;
      RECT  8532.5 57307.5 8597.5 57172.5 ;
      RECT  8532.5 58192.5 8597.5 58057.5 ;
      RECT  8722.5 58192.5 8787.5 58057.5 ;
      RECT  8722.5 58192.5 8787.5 58057.5 ;
      RECT  8532.5 58192.5 8597.5 58057.5 ;
      RECT  8892.5 57217.5 8957.5 57082.5 ;
      RECT  8892.5 58192.5 8957.5 58057.5 ;
      RECT  8590.0 57750.0 8655.0 57615.0 ;
      RECT  8590.0 57750.0 8655.0 57615.0 ;
      RECT  8755.0 57715.0 8820.0 57650.0 ;
      RECT  8465.0 56997.5 9025.0 56932.5 ;
      RECT  8465.0 58342.5 9025.0 58277.5 ;
      RECT  8892.5 59470.0 8957.5 59655.0 ;
      RECT  8892.5 58310.0 8957.5 58495.0 ;
      RECT  8532.5 58427.5 8597.5 58277.5 ;
      RECT  8532.5 59312.5 8597.5 59687.5 ;
      RECT  8722.5 58427.5 8787.5 59312.5 ;
      RECT  8532.5 59312.5 8597.5 59447.5 ;
      RECT  8722.5 59312.5 8787.5 59447.5 ;
      RECT  8722.5 59312.5 8787.5 59447.5 ;
      RECT  8532.5 59312.5 8597.5 59447.5 ;
      RECT  8532.5 58427.5 8597.5 58562.5 ;
      RECT  8722.5 58427.5 8787.5 58562.5 ;
      RECT  8722.5 58427.5 8787.5 58562.5 ;
      RECT  8532.5 58427.5 8597.5 58562.5 ;
      RECT  8892.5 59402.5 8957.5 59537.5 ;
      RECT  8892.5 58427.5 8957.5 58562.5 ;
      RECT  8590.0 58870.0 8655.0 59005.0 ;
      RECT  8590.0 58870.0 8655.0 59005.0 ;
      RECT  8755.0 58905.0 8820.0 58970.0 ;
      RECT  8465.0 59622.5 9025.0 59687.5 ;
      RECT  8465.0 58277.5 9025.0 58342.5 ;
      RECT  8892.5 59840.0 8957.5 59655.0 ;
      RECT  8892.5 61000.0 8957.5 60815.0 ;
      RECT  8532.5 60882.5 8597.5 61032.5 ;
      RECT  8532.5 59997.5 8597.5 59622.5 ;
      RECT  8722.5 60882.5 8787.5 59997.5 ;
      RECT  8532.5 59997.5 8597.5 59862.5 ;
      RECT  8722.5 59997.5 8787.5 59862.5 ;
      RECT  8722.5 59997.5 8787.5 59862.5 ;
      RECT  8532.5 59997.5 8597.5 59862.5 ;
      RECT  8532.5 60882.5 8597.5 60747.5 ;
      RECT  8722.5 60882.5 8787.5 60747.5 ;
      RECT  8722.5 60882.5 8787.5 60747.5 ;
      RECT  8532.5 60882.5 8597.5 60747.5 ;
      RECT  8892.5 59907.5 8957.5 59772.5 ;
      RECT  8892.5 60882.5 8957.5 60747.5 ;
      RECT  8590.0 60440.0 8655.0 60305.0 ;
      RECT  8590.0 60440.0 8655.0 60305.0 ;
      RECT  8755.0 60405.0 8820.0 60340.0 ;
      RECT  8465.0 59687.5 9025.0 59622.5 ;
      RECT  8465.0 61032.5 9025.0 60967.5 ;
      RECT  8892.5 62160.0 8957.5 62345.0 ;
      RECT  8892.5 61000.0 8957.5 61185.0 ;
      RECT  8532.5 61117.5 8597.5 60967.5 ;
      RECT  8532.5 62002.5 8597.5 62377.5 ;
      RECT  8722.5 61117.5 8787.5 62002.5 ;
      RECT  8532.5 62002.5 8597.5 62137.5 ;
      RECT  8722.5 62002.5 8787.5 62137.5 ;
      RECT  8722.5 62002.5 8787.5 62137.5 ;
      RECT  8532.5 62002.5 8597.5 62137.5 ;
      RECT  8532.5 61117.5 8597.5 61252.5 ;
      RECT  8722.5 61117.5 8787.5 61252.5 ;
      RECT  8722.5 61117.5 8787.5 61252.5 ;
      RECT  8532.5 61117.5 8597.5 61252.5 ;
      RECT  8892.5 62092.5 8957.5 62227.5 ;
      RECT  8892.5 61117.5 8957.5 61252.5 ;
      RECT  8590.0 61560.0 8655.0 61695.0 ;
      RECT  8590.0 61560.0 8655.0 61695.0 ;
      RECT  8755.0 61595.0 8820.0 61660.0 ;
      RECT  8465.0 62312.5 9025.0 62377.5 ;
      RECT  8465.0 60967.5 9025.0 61032.5 ;
      RECT  8892.5 62530.0 8957.5 62345.0 ;
      RECT  8892.5 63690.0 8957.5 63505.0 ;
      RECT  8532.5 63572.5 8597.5 63722.5 ;
      RECT  8532.5 62687.5 8597.5 62312.5 ;
      RECT  8722.5 63572.5 8787.5 62687.5 ;
      RECT  8532.5 62687.5 8597.5 62552.5 ;
      RECT  8722.5 62687.5 8787.5 62552.5 ;
      RECT  8722.5 62687.5 8787.5 62552.5 ;
      RECT  8532.5 62687.5 8597.5 62552.5 ;
      RECT  8532.5 63572.5 8597.5 63437.5 ;
      RECT  8722.5 63572.5 8787.5 63437.5 ;
      RECT  8722.5 63572.5 8787.5 63437.5 ;
      RECT  8532.5 63572.5 8597.5 63437.5 ;
      RECT  8892.5 62597.5 8957.5 62462.5 ;
      RECT  8892.5 63572.5 8957.5 63437.5 ;
      RECT  8590.0 63130.0 8655.0 62995.0 ;
      RECT  8590.0 63130.0 8655.0 62995.0 ;
      RECT  8755.0 63095.0 8820.0 63030.0 ;
      RECT  8465.0 62377.5 9025.0 62312.5 ;
      RECT  8465.0 63722.5 9025.0 63657.5 ;
      RECT  8892.5 64850.0 8957.5 65035.0 ;
      RECT  8892.5 63690.0 8957.5 63875.0 ;
      RECT  8532.5 63807.5 8597.5 63657.5 ;
      RECT  8532.5 64692.5 8597.5 65067.5 ;
      RECT  8722.5 63807.5 8787.5 64692.5 ;
      RECT  8532.5 64692.5 8597.5 64827.5 ;
      RECT  8722.5 64692.5 8787.5 64827.5 ;
      RECT  8722.5 64692.5 8787.5 64827.5 ;
      RECT  8532.5 64692.5 8597.5 64827.5 ;
      RECT  8532.5 63807.5 8597.5 63942.5 ;
      RECT  8722.5 63807.5 8787.5 63942.5 ;
      RECT  8722.5 63807.5 8787.5 63942.5 ;
      RECT  8532.5 63807.5 8597.5 63942.5 ;
      RECT  8892.5 64782.5 8957.5 64917.5 ;
      RECT  8892.5 63807.5 8957.5 63942.5 ;
      RECT  8590.0 64250.0 8655.0 64385.0 ;
      RECT  8590.0 64250.0 8655.0 64385.0 ;
      RECT  8755.0 64285.0 8820.0 64350.0 ;
      RECT  8465.0 65002.5 9025.0 65067.5 ;
      RECT  8465.0 63657.5 9025.0 63722.5 ;
      RECT  8892.5 65220.0 8957.5 65035.0 ;
      RECT  8892.5 66380.0 8957.5 66195.0 ;
      RECT  8532.5 66262.5 8597.5 66412.5 ;
      RECT  8532.5 65377.5 8597.5 65002.5 ;
      RECT  8722.5 66262.5 8787.5 65377.5 ;
      RECT  8532.5 65377.5 8597.5 65242.5 ;
      RECT  8722.5 65377.5 8787.5 65242.5 ;
      RECT  8722.5 65377.5 8787.5 65242.5 ;
      RECT  8532.5 65377.5 8597.5 65242.5 ;
      RECT  8532.5 66262.5 8597.5 66127.5 ;
      RECT  8722.5 66262.5 8787.5 66127.5 ;
      RECT  8722.5 66262.5 8787.5 66127.5 ;
      RECT  8532.5 66262.5 8597.5 66127.5 ;
      RECT  8892.5 65287.5 8957.5 65152.5 ;
      RECT  8892.5 66262.5 8957.5 66127.5 ;
      RECT  8590.0 65820.0 8655.0 65685.0 ;
      RECT  8590.0 65820.0 8655.0 65685.0 ;
      RECT  8755.0 65785.0 8820.0 65720.0 ;
      RECT  8465.0 65067.5 9025.0 65002.5 ;
      RECT  8465.0 66412.5 9025.0 66347.5 ;
      RECT  8892.5 67540.0 8957.5 67725.0 ;
      RECT  8892.5 66380.0 8957.5 66565.0 ;
      RECT  8532.5 66497.5 8597.5 66347.5 ;
      RECT  8532.5 67382.5 8597.5 67757.5 ;
      RECT  8722.5 66497.5 8787.5 67382.5 ;
      RECT  8532.5 67382.5 8597.5 67517.5 ;
      RECT  8722.5 67382.5 8787.5 67517.5 ;
      RECT  8722.5 67382.5 8787.5 67517.5 ;
      RECT  8532.5 67382.5 8597.5 67517.5 ;
      RECT  8532.5 66497.5 8597.5 66632.5 ;
      RECT  8722.5 66497.5 8787.5 66632.5 ;
      RECT  8722.5 66497.5 8787.5 66632.5 ;
      RECT  8532.5 66497.5 8597.5 66632.5 ;
      RECT  8892.5 67472.5 8957.5 67607.5 ;
      RECT  8892.5 66497.5 8957.5 66632.5 ;
      RECT  8590.0 66940.0 8655.0 67075.0 ;
      RECT  8590.0 66940.0 8655.0 67075.0 ;
      RECT  8755.0 66975.0 8820.0 67040.0 ;
      RECT  8465.0 67692.5 9025.0 67757.5 ;
      RECT  8465.0 66347.5 9025.0 66412.5 ;
      RECT  8892.5 67910.0 8957.5 67725.0 ;
      RECT  8892.5 69070.0 8957.5 68885.0 ;
      RECT  8532.5 68952.5 8597.5 69102.5 ;
      RECT  8532.5 68067.5 8597.5 67692.5 ;
      RECT  8722.5 68952.5 8787.5 68067.5 ;
      RECT  8532.5 68067.5 8597.5 67932.5 ;
      RECT  8722.5 68067.5 8787.5 67932.5 ;
      RECT  8722.5 68067.5 8787.5 67932.5 ;
      RECT  8532.5 68067.5 8597.5 67932.5 ;
      RECT  8532.5 68952.5 8597.5 68817.5 ;
      RECT  8722.5 68952.5 8787.5 68817.5 ;
      RECT  8722.5 68952.5 8787.5 68817.5 ;
      RECT  8532.5 68952.5 8597.5 68817.5 ;
      RECT  8892.5 67977.5 8957.5 67842.5 ;
      RECT  8892.5 68952.5 8957.5 68817.5 ;
      RECT  8590.0 68510.0 8655.0 68375.0 ;
      RECT  8590.0 68510.0 8655.0 68375.0 ;
      RECT  8755.0 68475.0 8820.0 68410.0 ;
      RECT  8465.0 67757.5 9025.0 67692.5 ;
      RECT  8465.0 69102.5 9025.0 69037.5 ;
      RECT  8892.5 70230.0 8957.5 70415.0 ;
      RECT  8892.5 69070.0 8957.5 69255.0 ;
      RECT  8532.5 69187.5 8597.5 69037.5 ;
      RECT  8532.5 70072.5 8597.5 70447.5 ;
      RECT  8722.5 69187.5 8787.5 70072.5 ;
      RECT  8532.5 70072.5 8597.5 70207.5 ;
      RECT  8722.5 70072.5 8787.5 70207.5 ;
      RECT  8722.5 70072.5 8787.5 70207.5 ;
      RECT  8532.5 70072.5 8597.5 70207.5 ;
      RECT  8532.5 69187.5 8597.5 69322.5 ;
      RECT  8722.5 69187.5 8787.5 69322.5 ;
      RECT  8722.5 69187.5 8787.5 69322.5 ;
      RECT  8532.5 69187.5 8597.5 69322.5 ;
      RECT  8892.5 70162.5 8957.5 70297.5 ;
      RECT  8892.5 69187.5 8957.5 69322.5 ;
      RECT  8590.0 69630.0 8655.0 69765.0 ;
      RECT  8590.0 69630.0 8655.0 69765.0 ;
      RECT  8755.0 69665.0 8820.0 69730.0 ;
      RECT  8465.0 70382.5 9025.0 70447.5 ;
      RECT  8465.0 69037.5 9025.0 69102.5 ;
      RECT  8892.5 70600.0 8957.5 70415.0 ;
      RECT  8892.5 71760.0 8957.5 71575.0 ;
      RECT  8532.5 71642.5 8597.5 71792.5 ;
      RECT  8532.5 70757.5 8597.5 70382.5 ;
      RECT  8722.5 71642.5 8787.5 70757.5 ;
      RECT  8532.5 70757.5 8597.5 70622.5 ;
      RECT  8722.5 70757.5 8787.5 70622.5 ;
      RECT  8722.5 70757.5 8787.5 70622.5 ;
      RECT  8532.5 70757.5 8597.5 70622.5 ;
      RECT  8532.5 71642.5 8597.5 71507.5 ;
      RECT  8722.5 71642.5 8787.5 71507.5 ;
      RECT  8722.5 71642.5 8787.5 71507.5 ;
      RECT  8532.5 71642.5 8597.5 71507.5 ;
      RECT  8892.5 70667.5 8957.5 70532.5 ;
      RECT  8892.5 71642.5 8957.5 71507.5 ;
      RECT  8590.0 71200.0 8655.0 71065.0 ;
      RECT  8590.0 71200.0 8655.0 71065.0 ;
      RECT  8755.0 71165.0 8820.0 71100.0 ;
      RECT  8465.0 70447.5 9025.0 70382.5 ;
      RECT  8465.0 71792.5 9025.0 71727.5 ;
      RECT  8892.5 72920.0 8957.5 73105.0 ;
      RECT  8892.5 71760.0 8957.5 71945.0 ;
      RECT  8532.5 71877.5 8597.5 71727.5 ;
      RECT  8532.5 72762.5 8597.5 73137.5 ;
      RECT  8722.5 71877.5 8787.5 72762.5 ;
      RECT  8532.5 72762.5 8597.5 72897.5 ;
      RECT  8722.5 72762.5 8787.5 72897.5 ;
      RECT  8722.5 72762.5 8787.5 72897.5 ;
      RECT  8532.5 72762.5 8597.5 72897.5 ;
      RECT  8532.5 71877.5 8597.5 72012.5 ;
      RECT  8722.5 71877.5 8787.5 72012.5 ;
      RECT  8722.5 71877.5 8787.5 72012.5 ;
      RECT  8532.5 71877.5 8597.5 72012.5 ;
      RECT  8892.5 72852.5 8957.5 72987.5 ;
      RECT  8892.5 71877.5 8957.5 72012.5 ;
      RECT  8590.0 72320.0 8655.0 72455.0 ;
      RECT  8590.0 72320.0 8655.0 72455.0 ;
      RECT  8755.0 72355.0 8820.0 72420.0 ;
      RECT  8465.0 73072.5 9025.0 73137.5 ;
      RECT  8465.0 71727.5 9025.0 71792.5 ;
      RECT  8892.5 73290.0 8957.5 73105.0 ;
      RECT  8892.5 74450.0 8957.5 74265.0 ;
      RECT  8532.5 74332.5 8597.5 74482.5 ;
      RECT  8532.5 73447.5 8597.5 73072.5 ;
      RECT  8722.5 74332.5 8787.5 73447.5 ;
      RECT  8532.5 73447.5 8597.5 73312.5 ;
      RECT  8722.5 73447.5 8787.5 73312.5 ;
      RECT  8722.5 73447.5 8787.5 73312.5 ;
      RECT  8532.5 73447.5 8597.5 73312.5 ;
      RECT  8532.5 74332.5 8597.5 74197.5 ;
      RECT  8722.5 74332.5 8787.5 74197.5 ;
      RECT  8722.5 74332.5 8787.5 74197.5 ;
      RECT  8532.5 74332.5 8597.5 74197.5 ;
      RECT  8892.5 73357.5 8957.5 73222.5 ;
      RECT  8892.5 74332.5 8957.5 74197.5 ;
      RECT  8590.0 73890.0 8655.0 73755.0 ;
      RECT  8590.0 73890.0 8655.0 73755.0 ;
      RECT  8755.0 73855.0 8820.0 73790.0 ;
      RECT  8465.0 73137.5 9025.0 73072.5 ;
      RECT  8465.0 74482.5 9025.0 74417.5 ;
      RECT  8892.5 75610.0 8957.5 75795.0 ;
      RECT  8892.5 74450.0 8957.5 74635.0 ;
      RECT  8532.5 74567.5 8597.5 74417.5 ;
      RECT  8532.5 75452.5 8597.5 75827.5 ;
      RECT  8722.5 74567.5 8787.5 75452.5 ;
      RECT  8532.5 75452.5 8597.5 75587.5 ;
      RECT  8722.5 75452.5 8787.5 75587.5 ;
      RECT  8722.5 75452.5 8787.5 75587.5 ;
      RECT  8532.5 75452.5 8597.5 75587.5 ;
      RECT  8532.5 74567.5 8597.5 74702.5 ;
      RECT  8722.5 74567.5 8787.5 74702.5 ;
      RECT  8722.5 74567.5 8787.5 74702.5 ;
      RECT  8532.5 74567.5 8597.5 74702.5 ;
      RECT  8892.5 75542.5 8957.5 75677.5 ;
      RECT  8892.5 74567.5 8957.5 74702.5 ;
      RECT  8590.0 75010.0 8655.0 75145.0 ;
      RECT  8590.0 75010.0 8655.0 75145.0 ;
      RECT  8755.0 75045.0 8820.0 75110.0 ;
      RECT  8465.0 75762.5 9025.0 75827.5 ;
      RECT  8465.0 74417.5 9025.0 74482.5 ;
      RECT  8892.5 75980.0 8957.5 75795.0 ;
      RECT  8892.5 77140.0 8957.5 76955.0 ;
      RECT  8532.5 77022.5 8597.5 77172.5 ;
      RECT  8532.5 76137.5 8597.5 75762.5 ;
      RECT  8722.5 77022.5 8787.5 76137.5 ;
      RECT  8532.5 76137.5 8597.5 76002.5 ;
      RECT  8722.5 76137.5 8787.5 76002.5 ;
      RECT  8722.5 76137.5 8787.5 76002.5 ;
      RECT  8532.5 76137.5 8597.5 76002.5 ;
      RECT  8532.5 77022.5 8597.5 76887.5 ;
      RECT  8722.5 77022.5 8787.5 76887.5 ;
      RECT  8722.5 77022.5 8787.5 76887.5 ;
      RECT  8532.5 77022.5 8597.5 76887.5 ;
      RECT  8892.5 76047.5 8957.5 75912.5 ;
      RECT  8892.5 77022.5 8957.5 76887.5 ;
      RECT  8590.0 76580.0 8655.0 76445.0 ;
      RECT  8590.0 76580.0 8655.0 76445.0 ;
      RECT  8755.0 76545.0 8820.0 76480.0 ;
      RECT  8465.0 75827.5 9025.0 75762.5 ;
      RECT  8465.0 77172.5 9025.0 77107.5 ;
      RECT  8892.5 78300.0 8957.5 78485.0 ;
      RECT  8892.5 77140.0 8957.5 77325.0 ;
      RECT  8532.5 77257.5 8597.5 77107.5 ;
      RECT  8532.5 78142.5 8597.5 78517.5 ;
      RECT  8722.5 77257.5 8787.5 78142.5 ;
      RECT  8532.5 78142.5 8597.5 78277.5 ;
      RECT  8722.5 78142.5 8787.5 78277.5 ;
      RECT  8722.5 78142.5 8787.5 78277.5 ;
      RECT  8532.5 78142.5 8597.5 78277.5 ;
      RECT  8532.5 77257.5 8597.5 77392.5 ;
      RECT  8722.5 77257.5 8787.5 77392.5 ;
      RECT  8722.5 77257.5 8787.5 77392.5 ;
      RECT  8532.5 77257.5 8597.5 77392.5 ;
      RECT  8892.5 78232.5 8957.5 78367.5 ;
      RECT  8892.5 77257.5 8957.5 77392.5 ;
      RECT  8590.0 77700.0 8655.0 77835.0 ;
      RECT  8590.0 77700.0 8655.0 77835.0 ;
      RECT  8755.0 77735.0 8820.0 77800.0 ;
      RECT  8465.0 78452.5 9025.0 78517.5 ;
      RECT  8465.0 77107.5 9025.0 77172.5 ;
      RECT  8892.5 78670.0 8957.5 78485.0 ;
      RECT  8892.5 79830.0 8957.5 79645.0 ;
      RECT  8532.5 79712.5 8597.5 79862.5 ;
      RECT  8532.5 78827.5 8597.5 78452.5 ;
      RECT  8722.5 79712.5 8787.5 78827.5 ;
      RECT  8532.5 78827.5 8597.5 78692.5 ;
      RECT  8722.5 78827.5 8787.5 78692.5 ;
      RECT  8722.5 78827.5 8787.5 78692.5 ;
      RECT  8532.5 78827.5 8597.5 78692.5 ;
      RECT  8532.5 79712.5 8597.5 79577.5 ;
      RECT  8722.5 79712.5 8787.5 79577.5 ;
      RECT  8722.5 79712.5 8787.5 79577.5 ;
      RECT  8532.5 79712.5 8597.5 79577.5 ;
      RECT  8892.5 78737.5 8957.5 78602.5 ;
      RECT  8892.5 79712.5 8957.5 79577.5 ;
      RECT  8590.0 79270.0 8655.0 79135.0 ;
      RECT  8590.0 79270.0 8655.0 79135.0 ;
      RECT  8755.0 79235.0 8820.0 79170.0 ;
      RECT  8465.0 78517.5 9025.0 78452.5 ;
      RECT  8465.0 79862.5 9025.0 79797.5 ;
      RECT  8892.5 80990.0 8957.5 81175.0 ;
      RECT  8892.5 79830.0 8957.5 80015.0 ;
      RECT  8532.5 79947.5 8597.5 79797.5 ;
      RECT  8532.5 80832.5 8597.5 81207.5 ;
      RECT  8722.5 79947.5 8787.5 80832.5 ;
      RECT  8532.5 80832.5 8597.5 80967.5 ;
      RECT  8722.5 80832.5 8787.5 80967.5 ;
      RECT  8722.5 80832.5 8787.5 80967.5 ;
      RECT  8532.5 80832.5 8597.5 80967.5 ;
      RECT  8532.5 79947.5 8597.5 80082.5 ;
      RECT  8722.5 79947.5 8787.5 80082.5 ;
      RECT  8722.5 79947.5 8787.5 80082.5 ;
      RECT  8532.5 79947.5 8597.5 80082.5 ;
      RECT  8892.5 80922.5 8957.5 81057.5 ;
      RECT  8892.5 79947.5 8957.5 80082.5 ;
      RECT  8590.0 80390.0 8655.0 80525.0 ;
      RECT  8590.0 80390.0 8655.0 80525.0 ;
      RECT  8755.0 80425.0 8820.0 80490.0 ;
      RECT  8465.0 81142.5 9025.0 81207.5 ;
      RECT  8465.0 79797.5 9025.0 79862.5 ;
      RECT  8892.5 81360.0 8957.5 81175.0 ;
      RECT  8892.5 82520.0 8957.5 82335.0 ;
      RECT  8532.5 82402.5 8597.5 82552.5 ;
      RECT  8532.5 81517.5 8597.5 81142.5 ;
      RECT  8722.5 82402.5 8787.5 81517.5 ;
      RECT  8532.5 81517.5 8597.5 81382.5 ;
      RECT  8722.5 81517.5 8787.5 81382.5 ;
      RECT  8722.5 81517.5 8787.5 81382.5 ;
      RECT  8532.5 81517.5 8597.5 81382.5 ;
      RECT  8532.5 82402.5 8597.5 82267.5 ;
      RECT  8722.5 82402.5 8787.5 82267.5 ;
      RECT  8722.5 82402.5 8787.5 82267.5 ;
      RECT  8532.5 82402.5 8597.5 82267.5 ;
      RECT  8892.5 81427.5 8957.5 81292.5 ;
      RECT  8892.5 82402.5 8957.5 82267.5 ;
      RECT  8590.0 81960.0 8655.0 81825.0 ;
      RECT  8590.0 81960.0 8655.0 81825.0 ;
      RECT  8755.0 81925.0 8820.0 81860.0 ;
      RECT  8465.0 81207.5 9025.0 81142.5 ;
      RECT  8465.0 82552.5 9025.0 82487.5 ;
      RECT  8892.5 83680.0 8957.5 83865.0 ;
      RECT  8892.5 82520.0 8957.5 82705.0 ;
      RECT  8532.5 82637.5 8597.5 82487.5 ;
      RECT  8532.5 83522.5 8597.5 83897.5 ;
      RECT  8722.5 82637.5 8787.5 83522.5 ;
      RECT  8532.5 83522.5 8597.5 83657.5 ;
      RECT  8722.5 83522.5 8787.5 83657.5 ;
      RECT  8722.5 83522.5 8787.5 83657.5 ;
      RECT  8532.5 83522.5 8597.5 83657.5 ;
      RECT  8532.5 82637.5 8597.5 82772.5 ;
      RECT  8722.5 82637.5 8787.5 82772.5 ;
      RECT  8722.5 82637.5 8787.5 82772.5 ;
      RECT  8532.5 82637.5 8597.5 82772.5 ;
      RECT  8892.5 83612.5 8957.5 83747.5 ;
      RECT  8892.5 82637.5 8957.5 82772.5 ;
      RECT  8590.0 83080.0 8655.0 83215.0 ;
      RECT  8590.0 83080.0 8655.0 83215.0 ;
      RECT  8755.0 83115.0 8820.0 83180.0 ;
      RECT  8465.0 83832.5 9025.0 83897.5 ;
      RECT  8465.0 82487.5 9025.0 82552.5 ;
      RECT  8892.5 84050.0 8957.5 83865.0 ;
      RECT  8892.5 85210.0 8957.5 85025.0 ;
      RECT  8532.5 85092.5 8597.5 85242.5 ;
      RECT  8532.5 84207.5 8597.5 83832.5 ;
      RECT  8722.5 85092.5 8787.5 84207.5 ;
      RECT  8532.5 84207.5 8597.5 84072.5 ;
      RECT  8722.5 84207.5 8787.5 84072.5 ;
      RECT  8722.5 84207.5 8787.5 84072.5 ;
      RECT  8532.5 84207.5 8597.5 84072.5 ;
      RECT  8532.5 85092.5 8597.5 84957.5 ;
      RECT  8722.5 85092.5 8787.5 84957.5 ;
      RECT  8722.5 85092.5 8787.5 84957.5 ;
      RECT  8532.5 85092.5 8597.5 84957.5 ;
      RECT  8892.5 84117.5 8957.5 83982.5 ;
      RECT  8892.5 85092.5 8957.5 84957.5 ;
      RECT  8590.0 84650.0 8655.0 84515.0 ;
      RECT  8590.0 84650.0 8655.0 84515.0 ;
      RECT  8755.0 84615.0 8820.0 84550.0 ;
      RECT  8465.0 83897.5 9025.0 83832.5 ;
      RECT  8465.0 85242.5 9025.0 85177.5 ;
      RECT  8892.5 86370.0 8957.5 86555.0 ;
      RECT  8892.5 85210.0 8957.5 85395.0 ;
      RECT  8532.5 85327.5 8597.5 85177.5 ;
      RECT  8532.5 86212.5 8597.5 86587.5 ;
      RECT  8722.5 85327.5 8787.5 86212.5 ;
      RECT  8532.5 86212.5 8597.5 86347.5 ;
      RECT  8722.5 86212.5 8787.5 86347.5 ;
      RECT  8722.5 86212.5 8787.5 86347.5 ;
      RECT  8532.5 86212.5 8597.5 86347.5 ;
      RECT  8532.5 85327.5 8597.5 85462.5 ;
      RECT  8722.5 85327.5 8787.5 85462.5 ;
      RECT  8722.5 85327.5 8787.5 85462.5 ;
      RECT  8532.5 85327.5 8597.5 85462.5 ;
      RECT  8892.5 86302.5 8957.5 86437.5 ;
      RECT  8892.5 85327.5 8957.5 85462.5 ;
      RECT  8590.0 85770.0 8655.0 85905.0 ;
      RECT  8590.0 85770.0 8655.0 85905.0 ;
      RECT  8755.0 85805.0 8820.0 85870.0 ;
      RECT  8465.0 86522.5 9025.0 86587.5 ;
      RECT  8465.0 85177.5 9025.0 85242.5 ;
      RECT  8892.5 86740.0 8957.5 86555.0 ;
      RECT  8892.5 87900.0 8957.5 87715.0 ;
      RECT  8532.5 87782.5 8597.5 87932.5 ;
      RECT  8532.5 86897.5 8597.5 86522.5 ;
      RECT  8722.5 87782.5 8787.5 86897.5 ;
      RECT  8532.5 86897.5 8597.5 86762.5 ;
      RECT  8722.5 86897.5 8787.5 86762.5 ;
      RECT  8722.5 86897.5 8787.5 86762.5 ;
      RECT  8532.5 86897.5 8597.5 86762.5 ;
      RECT  8532.5 87782.5 8597.5 87647.5 ;
      RECT  8722.5 87782.5 8787.5 87647.5 ;
      RECT  8722.5 87782.5 8787.5 87647.5 ;
      RECT  8532.5 87782.5 8597.5 87647.5 ;
      RECT  8892.5 86807.5 8957.5 86672.5 ;
      RECT  8892.5 87782.5 8957.5 87647.5 ;
      RECT  8590.0 87340.0 8655.0 87205.0 ;
      RECT  8590.0 87340.0 8655.0 87205.0 ;
      RECT  8755.0 87305.0 8820.0 87240.0 ;
      RECT  8465.0 86587.5 9025.0 86522.5 ;
      RECT  8465.0 87932.5 9025.0 87867.5 ;
      RECT  8892.5 89060.0 8957.5 89245.0 ;
      RECT  8892.5 87900.0 8957.5 88085.0 ;
      RECT  8532.5 88017.5 8597.5 87867.5 ;
      RECT  8532.5 88902.5 8597.5 89277.5 ;
      RECT  8722.5 88017.5 8787.5 88902.5 ;
      RECT  8532.5 88902.5 8597.5 89037.5 ;
      RECT  8722.5 88902.5 8787.5 89037.5 ;
      RECT  8722.5 88902.5 8787.5 89037.5 ;
      RECT  8532.5 88902.5 8597.5 89037.5 ;
      RECT  8532.5 88017.5 8597.5 88152.5 ;
      RECT  8722.5 88017.5 8787.5 88152.5 ;
      RECT  8722.5 88017.5 8787.5 88152.5 ;
      RECT  8532.5 88017.5 8597.5 88152.5 ;
      RECT  8892.5 88992.5 8957.5 89127.5 ;
      RECT  8892.5 88017.5 8957.5 88152.5 ;
      RECT  8590.0 88460.0 8655.0 88595.0 ;
      RECT  8590.0 88460.0 8655.0 88595.0 ;
      RECT  8755.0 88495.0 8820.0 88560.0 ;
      RECT  8465.0 89212.5 9025.0 89277.5 ;
      RECT  8465.0 87867.5 9025.0 87932.5 ;
      RECT  8892.5 89430.0 8957.5 89245.0 ;
      RECT  8892.5 90590.0 8957.5 90405.0 ;
      RECT  8532.5 90472.5 8597.5 90622.5 ;
      RECT  8532.5 89587.5 8597.5 89212.5 ;
      RECT  8722.5 90472.5 8787.5 89587.5 ;
      RECT  8532.5 89587.5 8597.5 89452.5 ;
      RECT  8722.5 89587.5 8787.5 89452.5 ;
      RECT  8722.5 89587.5 8787.5 89452.5 ;
      RECT  8532.5 89587.5 8597.5 89452.5 ;
      RECT  8532.5 90472.5 8597.5 90337.5 ;
      RECT  8722.5 90472.5 8787.5 90337.5 ;
      RECT  8722.5 90472.5 8787.5 90337.5 ;
      RECT  8532.5 90472.5 8597.5 90337.5 ;
      RECT  8892.5 89497.5 8957.5 89362.5 ;
      RECT  8892.5 90472.5 8957.5 90337.5 ;
      RECT  8590.0 90030.0 8655.0 89895.0 ;
      RECT  8590.0 90030.0 8655.0 89895.0 ;
      RECT  8755.0 89995.0 8820.0 89930.0 ;
      RECT  8465.0 89277.5 9025.0 89212.5 ;
      RECT  8465.0 90622.5 9025.0 90557.5 ;
      RECT  8892.5 91750.0 8957.5 91935.0 ;
      RECT  8892.5 90590.0 8957.5 90775.0 ;
      RECT  8532.5 90707.5 8597.5 90557.5 ;
      RECT  8532.5 91592.5 8597.5 91967.5 ;
      RECT  8722.5 90707.5 8787.5 91592.5 ;
      RECT  8532.5 91592.5 8597.5 91727.5 ;
      RECT  8722.5 91592.5 8787.5 91727.5 ;
      RECT  8722.5 91592.5 8787.5 91727.5 ;
      RECT  8532.5 91592.5 8597.5 91727.5 ;
      RECT  8532.5 90707.5 8597.5 90842.5 ;
      RECT  8722.5 90707.5 8787.5 90842.5 ;
      RECT  8722.5 90707.5 8787.5 90842.5 ;
      RECT  8532.5 90707.5 8597.5 90842.5 ;
      RECT  8892.5 91682.5 8957.5 91817.5 ;
      RECT  8892.5 90707.5 8957.5 90842.5 ;
      RECT  8590.0 91150.0 8655.0 91285.0 ;
      RECT  8590.0 91150.0 8655.0 91285.0 ;
      RECT  8755.0 91185.0 8820.0 91250.0 ;
      RECT  8465.0 91902.5 9025.0 91967.5 ;
      RECT  8465.0 90557.5 9025.0 90622.5 ;
      RECT  8892.5 92120.0 8957.5 91935.0 ;
      RECT  8892.5 93280.0 8957.5 93095.0 ;
      RECT  8532.5 93162.5 8597.5 93312.5 ;
      RECT  8532.5 92277.5 8597.5 91902.5 ;
      RECT  8722.5 93162.5 8787.5 92277.5 ;
      RECT  8532.5 92277.5 8597.5 92142.5 ;
      RECT  8722.5 92277.5 8787.5 92142.5 ;
      RECT  8722.5 92277.5 8787.5 92142.5 ;
      RECT  8532.5 92277.5 8597.5 92142.5 ;
      RECT  8532.5 93162.5 8597.5 93027.5 ;
      RECT  8722.5 93162.5 8787.5 93027.5 ;
      RECT  8722.5 93162.5 8787.5 93027.5 ;
      RECT  8532.5 93162.5 8597.5 93027.5 ;
      RECT  8892.5 92187.5 8957.5 92052.5 ;
      RECT  8892.5 93162.5 8957.5 93027.5 ;
      RECT  8590.0 92720.0 8655.0 92585.0 ;
      RECT  8590.0 92720.0 8655.0 92585.0 ;
      RECT  8755.0 92685.0 8820.0 92620.0 ;
      RECT  8465.0 91967.5 9025.0 91902.5 ;
      RECT  8465.0 93312.5 9025.0 93247.5 ;
      RECT  8892.5 94440.0 8957.5 94625.0 ;
      RECT  8892.5 93280.0 8957.5 93465.0 ;
      RECT  8532.5 93397.5 8597.5 93247.5 ;
      RECT  8532.5 94282.5 8597.5 94657.5 ;
      RECT  8722.5 93397.5 8787.5 94282.5 ;
      RECT  8532.5 94282.5 8597.5 94417.5 ;
      RECT  8722.5 94282.5 8787.5 94417.5 ;
      RECT  8722.5 94282.5 8787.5 94417.5 ;
      RECT  8532.5 94282.5 8597.5 94417.5 ;
      RECT  8532.5 93397.5 8597.5 93532.5 ;
      RECT  8722.5 93397.5 8787.5 93532.5 ;
      RECT  8722.5 93397.5 8787.5 93532.5 ;
      RECT  8532.5 93397.5 8597.5 93532.5 ;
      RECT  8892.5 94372.5 8957.5 94507.5 ;
      RECT  8892.5 93397.5 8957.5 93532.5 ;
      RECT  8590.0 93840.0 8655.0 93975.0 ;
      RECT  8590.0 93840.0 8655.0 93975.0 ;
      RECT  8755.0 93875.0 8820.0 93940.0 ;
      RECT  8465.0 94592.5 9025.0 94657.5 ;
      RECT  8465.0 93247.5 9025.0 93312.5 ;
      RECT  8892.5 94810.0 8957.5 94625.0 ;
      RECT  8892.5 95970.0 8957.5 95785.0 ;
      RECT  8532.5 95852.5 8597.5 96002.5 ;
      RECT  8532.5 94967.5 8597.5 94592.5 ;
      RECT  8722.5 95852.5 8787.5 94967.5 ;
      RECT  8532.5 94967.5 8597.5 94832.5 ;
      RECT  8722.5 94967.5 8787.5 94832.5 ;
      RECT  8722.5 94967.5 8787.5 94832.5 ;
      RECT  8532.5 94967.5 8597.5 94832.5 ;
      RECT  8532.5 95852.5 8597.5 95717.5 ;
      RECT  8722.5 95852.5 8787.5 95717.5 ;
      RECT  8722.5 95852.5 8787.5 95717.5 ;
      RECT  8532.5 95852.5 8597.5 95717.5 ;
      RECT  8892.5 94877.5 8957.5 94742.5 ;
      RECT  8892.5 95852.5 8957.5 95717.5 ;
      RECT  8590.0 95410.0 8655.0 95275.0 ;
      RECT  8590.0 95410.0 8655.0 95275.0 ;
      RECT  8755.0 95375.0 8820.0 95310.0 ;
      RECT  8465.0 94657.5 9025.0 94592.5 ;
      RECT  8465.0 96002.5 9025.0 95937.5 ;
      RECT  8892.5 97130.0 8957.5 97315.0 ;
      RECT  8892.5 95970.0 8957.5 96155.0 ;
      RECT  8532.5 96087.5 8597.5 95937.5 ;
      RECT  8532.5 96972.5 8597.5 97347.5 ;
      RECT  8722.5 96087.5 8787.5 96972.5 ;
      RECT  8532.5 96972.5 8597.5 97107.5 ;
      RECT  8722.5 96972.5 8787.5 97107.5 ;
      RECT  8722.5 96972.5 8787.5 97107.5 ;
      RECT  8532.5 96972.5 8597.5 97107.5 ;
      RECT  8532.5 96087.5 8597.5 96222.5 ;
      RECT  8722.5 96087.5 8787.5 96222.5 ;
      RECT  8722.5 96087.5 8787.5 96222.5 ;
      RECT  8532.5 96087.5 8597.5 96222.5 ;
      RECT  8892.5 97062.5 8957.5 97197.5 ;
      RECT  8892.5 96087.5 8957.5 96222.5 ;
      RECT  8590.0 96530.0 8655.0 96665.0 ;
      RECT  8590.0 96530.0 8655.0 96665.0 ;
      RECT  8755.0 96565.0 8820.0 96630.0 ;
      RECT  8465.0 97282.5 9025.0 97347.5 ;
      RECT  8465.0 95937.5 9025.0 96002.5 ;
      RECT  8892.5 97500.0 8957.5 97315.0 ;
      RECT  8892.5 98660.0 8957.5 98475.0 ;
      RECT  8532.5 98542.5 8597.5 98692.5 ;
      RECT  8532.5 97657.5 8597.5 97282.5 ;
      RECT  8722.5 98542.5 8787.5 97657.5 ;
      RECT  8532.5 97657.5 8597.5 97522.5 ;
      RECT  8722.5 97657.5 8787.5 97522.5 ;
      RECT  8722.5 97657.5 8787.5 97522.5 ;
      RECT  8532.5 97657.5 8597.5 97522.5 ;
      RECT  8532.5 98542.5 8597.5 98407.5 ;
      RECT  8722.5 98542.5 8787.5 98407.5 ;
      RECT  8722.5 98542.5 8787.5 98407.5 ;
      RECT  8532.5 98542.5 8597.5 98407.5 ;
      RECT  8892.5 97567.5 8957.5 97432.5 ;
      RECT  8892.5 98542.5 8957.5 98407.5 ;
      RECT  8590.0 98100.0 8655.0 97965.0 ;
      RECT  8590.0 98100.0 8655.0 97965.0 ;
      RECT  8755.0 98065.0 8820.0 98000.0 ;
      RECT  8465.0 97347.5 9025.0 97282.5 ;
      RECT  8465.0 98692.5 9025.0 98627.5 ;
      RECT  8892.5 99820.0 8957.5 100005.0 ;
      RECT  8892.5 98660.0 8957.5 98845.0 ;
      RECT  8532.5 98777.5 8597.5 98627.5 ;
      RECT  8532.5 99662.5 8597.5 100037.5 ;
      RECT  8722.5 98777.5 8787.5 99662.5 ;
      RECT  8532.5 99662.5 8597.5 99797.5 ;
      RECT  8722.5 99662.5 8787.5 99797.5 ;
      RECT  8722.5 99662.5 8787.5 99797.5 ;
      RECT  8532.5 99662.5 8597.5 99797.5 ;
      RECT  8532.5 98777.5 8597.5 98912.5 ;
      RECT  8722.5 98777.5 8787.5 98912.5 ;
      RECT  8722.5 98777.5 8787.5 98912.5 ;
      RECT  8532.5 98777.5 8597.5 98912.5 ;
      RECT  8892.5 99752.5 8957.5 99887.5 ;
      RECT  8892.5 98777.5 8957.5 98912.5 ;
      RECT  8590.0 99220.0 8655.0 99355.0 ;
      RECT  8590.0 99220.0 8655.0 99355.0 ;
      RECT  8755.0 99255.0 8820.0 99320.0 ;
      RECT  8465.0 99972.5 9025.0 100037.5 ;
      RECT  8465.0 98627.5 9025.0 98692.5 ;
      RECT  8892.5 100190.0 8957.5 100005.0 ;
      RECT  8892.5 101350.0 8957.5 101165.0 ;
      RECT  8532.5 101232.5 8597.5 101382.5 ;
      RECT  8532.5 100347.5 8597.5 99972.5 ;
      RECT  8722.5 101232.5 8787.5 100347.5 ;
      RECT  8532.5 100347.5 8597.5 100212.5 ;
      RECT  8722.5 100347.5 8787.5 100212.5 ;
      RECT  8722.5 100347.5 8787.5 100212.5 ;
      RECT  8532.5 100347.5 8597.5 100212.5 ;
      RECT  8532.5 101232.5 8597.5 101097.5 ;
      RECT  8722.5 101232.5 8787.5 101097.5 ;
      RECT  8722.5 101232.5 8787.5 101097.5 ;
      RECT  8532.5 101232.5 8597.5 101097.5 ;
      RECT  8892.5 100257.5 8957.5 100122.5 ;
      RECT  8892.5 101232.5 8957.5 101097.5 ;
      RECT  8590.0 100790.0 8655.0 100655.0 ;
      RECT  8590.0 100790.0 8655.0 100655.0 ;
      RECT  8755.0 100755.0 8820.0 100690.0 ;
      RECT  8465.0 100037.5 9025.0 99972.5 ;
      RECT  8465.0 101382.5 9025.0 101317.5 ;
      RECT  8892.5 102510.0 8957.5 102695.0 ;
      RECT  8892.5 101350.0 8957.5 101535.0 ;
      RECT  8532.5 101467.5 8597.5 101317.5 ;
      RECT  8532.5 102352.5 8597.5 102727.5 ;
      RECT  8722.5 101467.5 8787.5 102352.5 ;
      RECT  8532.5 102352.5 8597.5 102487.5 ;
      RECT  8722.5 102352.5 8787.5 102487.5 ;
      RECT  8722.5 102352.5 8787.5 102487.5 ;
      RECT  8532.5 102352.5 8597.5 102487.5 ;
      RECT  8532.5 101467.5 8597.5 101602.5 ;
      RECT  8722.5 101467.5 8787.5 101602.5 ;
      RECT  8722.5 101467.5 8787.5 101602.5 ;
      RECT  8532.5 101467.5 8597.5 101602.5 ;
      RECT  8892.5 102442.5 8957.5 102577.5 ;
      RECT  8892.5 101467.5 8957.5 101602.5 ;
      RECT  8590.0 101910.0 8655.0 102045.0 ;
      RECT  8590.0 101910.0 8655.0 102045.0 ;
      RECT  8755.0 101945.0 8820.0 102010.0 ;
      RECT  8465.0 102662.5 9025.0 102727.5 ;
      RECT  8465.0 101317.5 9025.0 101382.5 ;
      RECT  8892.5 102880.0 8957.5 102695.0 ;
      RECT  8892.5 104040.0 8957.5 103855.0 ;
      RECT  8532.5 103922.5 8597.5 104072.5 ;
      RECT  8532.5 103037.5 8597.5 102662.5 ;
      RECT  8722.5 103922.5 8787.5 103037.5 ;
      RECT  8532.5 103037.5 8597.5 102902.5 ;
      RECT  8722.5 103037.5 8787.5 102902.5 ;
      RECT  8722.5 103037.5 8787.5 102902.5 ;
      RECT  8532.5 103037.5 8597.5 102902.5 ;
      RECT  8532.5 103922.5 8597.5 103787.5 ;
      RECT  8722.5 103922.5 8787.5 103787.5 ;
      RECT  8722.5 103922.5 8787.5 103787.5 ;
      RECT  8532.5 103922.5 8597.5 103787.5 ;
      RECT  8892.5 102947.5 8957.5 102812.5 ;
      RECT  8892.5 103922.5 8957.5 103787.5 ;
      RECT  8590.0 103480.0 8655.0 103345.0 ;
      RECT  8590.0 103480.0 8655.0 103345.0 ;
      RECT  8755.0 103445.0 8820.0 103380.0 ;
      RECT  8465.0 102727.5 9025.0 102662.5 ;
      RECT  8465.0 104072.5 9025.0 104007.5 ;
      RECT  8892.5 105200.0 8957.5 105385.0 ;
      RECT  8892.5 104040.0 8957.5 104225.0 ;
      RECT  8532.5 104157.5 8597.5 104007.5 ;
      RECT  8532.5 105042.5 8597.5 105417.5 ;
      RECT  8722.5 104157.5 8787.5 105042.5 ;
      RECT  8532.5 105042.5 8597.5 105177.5 ;
      RECT  8722.5 105042.5 8787.5 105177.5 ;
      RECT  8722.5 105042.5 8787.5 105177.5 ;
      RECT  8532.5 105042.5 8597.5 105177.5 ;
      RECT  8532.5 104157.5 8597.5 104292.5 ;
      RECT  8722.5 104157.5 8787.5 104292.5 ;
      RECT  8722.5 104157.5 8787.5 104292.5 ;
      RECT  8532.5 104157.5 8597.5 104292.5 ;
      RECT  8892.5 105132.5 8957.5 105267.5 ;
      RECT  8892.5 104157.5 8957.5 104292.5 ;
      RECT  8590.0 104600.0 8655.0 104735.0 ;
      RECT  8590.0 104600.0 8655.0 104735.0 ;
      RECT  8755.0 104635.0 8820.0 104700.0 ;
      RECT  8465.0 105352.5 9025.0 105417.5 ;
      RECT  8465.0 104007.5 9025.0 104072.5 ;
      RECT  8892.5 105570.0 8957.5 105385.0 ;
      RECT  8892.5 106730.0 8957.5 106545.0 ;
      RECT  8532.5 106612.5 8597.5 106762.5 ;
      RECT  8532.5 105727.5 8597.5 105352.5 ;
      RECT  8722.5 106612.5 8787.5 105727.5 ;
      RECT  8532.5 105727.5 8597.5 105592.5 ;
      RECT  8722.5 105727.5 8787.5 105592.5 ;
      RECT  8722.5 105727.5 8787.5 105592.5 ;
      RECT  8532.5 105727.5 8597.5 105592.5 ;
      RECT  8532.5 106612.5 8597.5 106477.5 ;
      RECT  8722.5 106612.5 8787.5 106477.5 ;
      RECT  8722.5 106612.5 8787.5 106477.5 ;
      RECT  8532.5 106612.5 8597.5 106477.5 ;
      RECT  8892.5 105637.5 8957.5 105502.5 ;
      RECT  8892.5 106612.5 8957.5 106477.5 ;
      RECT  8590.0 106170.0 8655.0 106035.0 ;
      RECT  8590.0 106170.0 8655.0 106035.0 ;
      RECT  8755.0 106135.0 8820.0 106070.0 ;
      RECT  8465.0 105417.5 9025.0 105352.5 ;
      RECT  8465.0 106762.5 9025.0 106697.5 ;
      RECT  8892.5 107890.0 8957.5 108075.0 ;
      RECT  8892.5 106730.0 8957.5 106915.0 ;
      RECT  8532.5 106847.5 8597.5 106697.5 ;
      RECT  8532.5 107732.5 8597.5 108107.5 ;
      RECT  8722.5 106847.5 8787.5 107732.5 ;
      RECT  8532.5 107732.5 8597.5 107867.5 ;
      RECT  8722.5 107732.5 8787.5 107867.5 ;
      RECT  8722.5 107732.5 8787.5 107867.5 ;
      RECT  8532.5 107732.5 8597.5 107867.5 ;
      RECT  8532.5 106847.5 8597.5 106982.5 ;
      RECT  8722.5 106847.5 8787.5 106982.5 ;
      RECT  8722.5 106847.5 8787.5 106982.5 ;
      RECT  8532.5 106847.5 8597.5 106982.5 ;
      RECT  8892.5 107822.5 8957.5 107957.5 ;
      RECT  8892.5 106847.5 8957.5 106982.5 ;
      RECT  8590.0 107290.0 8655.0 107425.0 ;
      RECT  8590.0 107290.0 8655.0 107425.0 ;
      RECT  8755.0 107325.0 8820.0 107390.0 ;
      RECT  8465.0 108042.5 9025.0 108107.5 ;
      RECT  8465.0 106697.5 9025.0 106762.5 ;
      RECT  8892.5 108260.0 8957.5 108075.0 ;
      RECT  8892.5 109420.0 8957.5 109235.0 ;
      RECT  8532.5 109302.5 8597.5 109452.5 ;
      RECT  8532.5 108417.5 8597.5 108042.5 ;
      RECT  8722.5 109302.5 8787.5 108417.5 ;
      RECT  8532.5 108417.5 8597.5 108282.5 ;
      RECT  8722.5 108417.5 8787.5 108282.5 ;
      RECT  8722.5 108417.5 8787.5 108282.5 ;
      RECT  8532.5 108417.5 8597.5 108282.5 ;
      RECT  8532.5 109302.5 8597.5 109167.5 ;
      RECT  8722.5 109302.5 8787.5 109167.5 ;
      RECT  8722.5 109302.5 8787.5 109167.5 ;
      RECT  8532.5 109302.5 8597.5 109167.5 ;
      RECT  8892.5 108327.5 8957.5 108192.5 ;
      RECT  8892.5 109302.5 8957.5 109167.5 ;
      RECT  8590.0 108860.0 8655.0 108725.0 ;
      RECT  8590.0 108860.0 8655.0 108725.0 ;
      RECT  8755.0 108825.0 8820.0 108760.0 ;
      RECT  8465.0 108107.5 9025.0 108042.5 ;
      RECT  8465.0 109452.5 9025.0 109387.5 ;
      RECT  8892.5 110580.0 8957.5 110765.0 ;
      RECT  8892.5 109420.0 8957.5 109605.0 ;
      RECT  8532.5 109537.5 8597.5 109387.5 ;
      RECT  8532.5 110422.5 8597.5 110797.5 ;
      RECT  8722.5 109537.5 8787.5 110422.5 ;
      RECT  8532.5 110422.5 8597.5 110557.5 ;
      RECT  8722.5 110422.5 8787.5 110557.5 ;
      RECT  8722.5 110422.5 8787.5 110557.5 ;
      RECT  8532.5 110422.5 8597.5 110557.5 ;
      RECT  8532.5 109537.5 8597.5 109672.5 ;
      RECT  8722.5 109537.5 8787.5 109672.5 ;
      RECT  8722.5 109537.5 8787.5 109672.5 ;
      RECT  8532.5 109537.5 8597.5 109672.5 ;
      RECT  8892.5 110512.5 8957.5 110647.5 ;
      RECT  8892.5 109537.5 8957.5 109672.5 ;
      RECT  8590.0 109980.0 8655.0 110115.0 ;
      RECT  8590.0 109980.0 8655.0 110115.0 ;
      RECT  8755.0 110015.0 8820.0 110080.0 ;
      RECT  8465.0 110732.5 9025.0 110797.5 ;
      RECT  8465.0 109387.5 9025.0 109452.5 ;
      RECT  8892.5 110950.0 8957.5 110765.0 ;
      RECT  8892.5 112110.0 8957.5 111925.0 ;
      RECT  8532.5 111992.5 8597.5 112142.5 ;
      RECT  8532.5 111107.5 8597.5 110732.5 ;
      RECT  8722.5 111992.5 8787.5 111107.5 ;
      RECT  8532.5 111107.5 8597.5 110972.5 ;
      RECT  8722.5 111107.5 8787.5 110972.5 ;
      RECT  8722.5 111107.5 8787.5 110972.5 ;
      RECT  8532.5 111107.5 8597.5 110972.5 ;
      RECT  8532.5 111992.5 8597.5 111857.5 ;
      RECT  8722.5 111992.5 8787.5 111857.5 ;
      RECT  8722.5 111992.5 8787.5 111857.5 ;
      RECT  8532.5 111992.5 8597.5 111857.5 ;
      RECT  8892.5 111017.5 8957.5 110882.5 ;
      RECT  8892.5 111992.5 8957.5 111857.5 ;
      RECT  8590.0 111550.0 8655.0 111415.0 ;
      RECT  8590.0 111550.0 8655.0 111415.0 ;
      RECT  8755.0 111515.0 8820.0 111450.0 ;
      RECT  8465.0 110797.5 9025.0 110732.5 ;
      RECT  8465.0 112142.5 9025.0 112077.5 ;
      RECT  8892.5 113270.0 8957.5 113455.0 ;
      RECT  8892.5 112110.0 8957.5 112295.0 ;
      RECT  8532.5 112227.5 8597.5 112077.5 ;
      RECT  8532.5 113112.5 8597.5 113487.5 ;
      RECT  8722.5 112227.5 8787.5 113112.5 ;
      RECT  8532.5 113112.5 8597.5 113247.5 ;
      RECT  8722.5 113112.5 8787.5 113247.5 ;
      RECT  8722.5 113112.5 8787.5 113247.5 ;
      RECT  8532.5 113112.5 8597.5 113247.5 ;
      RECT  8532.5 112227.5 8597.5 112362.5 ;
      RECT  8722.5 112227.5 8787.5 112362.5 ;
      RECT  8722.5 112227.5 8787.5 112362.5 ;
      RECT  8532.5 112227.5 8597.5 112362.5 ;
      RECT  8892.5 113202.5 8957.5 113337.5 ;
      RECT  8892.5 112227.5 8957.5 112362.5 ;
      RECT  8590.0 112670.0 8655.0 112805.0 ;
      RECT  8590.0 112670.0 8655.0 112805.0 ;
      RECT  8755.0 112705.0 8820.0 112770.0 ;
      RECT  8465.0 113422.5 9025.0 113487.5 ;
      RECT  8465.0 112077.5 9025.0 112142.5 ;
      RECT  8892.5 113640.0 8957.5 113455.0 ;
      RECT  8892.5 114800.0 8957.5 114615.0 ;
      RECT  8532.5 114682.5 8597.5 114832.5 ;
      RECT  8532.5 113797.5 8597.5 113422.5 ;
      RECT  8722.5 114682.5 8787.5 113797.5 ;
      RECT  8532.5 113797.5 8597.5 113662.5 ;
      RECT  8722.5 113797.5 8787.5 113662.5 ;
      RECT  8722.5 113797.5 8787.5 113662.5 ;
      RECT  8532.5 113797.5 8597.5 113662.5 ;
      RECT  8532.5 114682.5 8597.5 114547.5 ;
      RECT  8722.5 114682.5 8787.5 114547.5 ;
      RECT  8722.5 114682.5 8787.5 114547.5 ;
      RECT  8532.5 114682.5 8597.5 114547.5 ;
      RECT  8892.5 113707.5 8957.5 113572.5 ;
      RECT  8892.5 114682.5 8957.5 114547.5 ;
      RECT  8590.0 114240.0 8655.0 114105.0 ;
      RECT  8590.0 114240.0 8655.0 114105.0 ;
      RECT  8755.0 114205.0 8820.0 114140.0 ;
      RECT  8465.0 113487.5 9025.0 113422.5 ;
      RECT  8465.0 114832.5 9025.0 114767.5 ;
      RECT  8892.5 115960.0 8957.5 116145.0 ;
      RECT  8892.5 114800.0 8957.5 114985.0 ;
      RECT  8532.5 114917.5 8597.5 114767.5 ;
      RECT  8532.5 115802.5 8597.5 116177.5 ;
      RECT  8722.5 114917.5 8787.5 115802.5 ;
      RECT  8532.5 115802.5 8597.5 115937.5 ;
      RECT  8722.5 115802.5 8787.5 115937.5 ;
      RECT  8722.5 115802.5 8787.5 115937.5 ;
      RECT  8532.5 115802.5 8597.5 115937.5 ;
      RECT  8532.5 114917.5 8597.5 115052.5 ;
      RECT  8722.5 114917.5 8787.5 115052.5 ;
      RECT  8722.5 114917.5 8787.5 115052.5 ;
      RECT  8532.5 114917.5 8597.5 115052.5 ;
      RECT  8892.5 115892.5 8957.5 116027.5 ;
      RECT  8892.5 114917.5 8957.5 115052.5 ;
      RECT  8590.0 115360.0 8655.0 115495.0 ;
      RECT  8590.0 115360.0 8655.0 115495.0 ;
      RECT  8755.0 115395.0 8820.0 115460.0 ;
      RECT  8465.0 116112.5 9025.0 116177.5 ;
      RECT  8465.0 114767.5 9025.0 114832.5 ;
      RECT  8892.5 116330.0 8957.5 116145.0 ;
      RECT  8892.5 117490.0 8957.5 117305.0 ;
      RECT  8532.5 117372.5 8597.5 117522.5 ;
      RECT  8532.5 116487.5 8597.5 116112.5 ;
      RECT  8722.5 117372.5 8787.5 116487.5 ;
      RECT  8532.5 116487.5 8597.5 116352.5 ;
      RECT  8722.5 116487.5 8787.5 116352.5 ;
      RECT  8722.5 116487.5 8787.5 116352.5 ;
      RECT  8532.5 116487.5 8597.5 116352.5 ;
      RECT  8532.5 117372.5 8597.5 117237.5 ;
      RECT  8722.5 117372.5 8787.5 117237.5 ;
      RECT  8722.5 117372.5 8787.5 117237.5 ;
      RECT  8532.5 117372.5 8597.5 117237.5 ;
      RECT  8892.5 116397.5 8957.5 116262.5 ;
      RECT  8892.5 117372.5 8957.5 117237.5 ;
      RECT  8590.0 116930.0 8655.0 116795.0 ;
      RECT  8590.0 116930.0 8655.0 116795.0 ;
      RECT  8755.0 116895.0 8820.0 116830.0 ;
      RECT  8465.0 116177.5 9025.0 116112.5 ;
      RECT  8465.0 117522.5 9025.0 117457.5 ;
      RECT  8892.5 118650.0 8957.5 118835.0 ;
      RECT  8892.5 117490.0 8957.5 117675.0 ;
      RECT  8532.5 117607.5 8597.5 117457.5 ;
      RECT  8532.5 118492.5 8597.5 118867.5 ;
      RECT  8722.5 117607.5 8787.5 118492.5 ;
      RECT  8532.5 118492.5 8597.5 118627.5 ;
      RECT  8722.5 118492.5 8787.5 118627.5 ;
      RECT  8722.5 118492.5 8787.5 118627.5 ;
      RECT  8532.5 118492.5 8597.5 118627.5 ;
      RECT  8532.5 117607.5 8597.5 117742.5 ;
      RECT  8722.5 117607.5 8787.5 117742.5 ;
      RECT  8722.5 117607.5 8787.5 117742.5 ;
      RECT  8532.5 117607.5 8597.5 117742.5 ;
      RECT  8892.5 118582.5 8957.5 118717.5 ;
      RECT  8892.5 117607.5 8957.5 117742.5 ;
      RECT  8590.0 118050.0 8655.0 118185.0 ;
      RECT  8590.0 118050.0 8655.0 118185.0 ;
      RECT  8755.0 118085.0 8820.0 118150.0 ;
      RECT  8465.0 118802.5 9025.0 118867.5 ;
      RECT  8465.0 117457.5 9025.0 117522.5 ;
      RECT  8892.5 119020.0 8957.5 118835.0 ;
      RECT  8892.5 120180.0 8957.5 119995.0 ;
      RECT  8532.5 120062.5 8597.5 120212.5 ;
      RECT  8532.5 119177.5 8597.5 118802.5 ;
      RECT  8722.5 120062.5 8787.5 119177.5 ;
      RECT  8532.5 119177.5 8597.5 119042.5 ;
      RECT  8722.5 119177.5 8787.5 119042.5 ;
      RECT  8722.5 119177.5 8787.5 119042.5 ;
      RECT  8532.5 119177.5 8597.5 119042.5 ;
      RECT  8532.5 120062.5 8597.5 119927.5 ;
      RECT  8722.5 120062.5 8787.5 119927.5 ;
      RECT  8722.5 120062.5 8787.5 119927.5 ;
      RECT  8532.5 120062.5 8597.5 119927.5 ;
      RECT  8892.5 119087.5 8957.5 118952.5 ;
      RECT  8892.5 120062.5 8957.5 119927.5 ;
      RECT  8590.0 119620.0 8655.0 119485.0 ;
      RECT  8590.0 119620.0 8655.0 119485.0 ;
      RECT  8755.0 119585.0 8820.0 119520.0 ;
      RECT  8465.0 118867.5 9025.0 118802.5 ;
      RECT  8465.0 120212.5 9025.0 120147.5 ;
      RECT  8892.5 121340.0 8957.5 121525.0 ;
      RECT  8892.5 120180.0 8957.5 120365.0 ;
      RECT  8532.5 120297.5 8597.5 120147.5 ;
      RECT  8532.5 121182.5 8597.5 121557.5 ;
      RECT  8722.5 120297.5 8787.5 121182.5 ;
      RECT  8532.5 121182.5 8597.5 121317.5 ;
      RECT  8722.5 121182.5 8787.5 121317.5 ;
      RECT  8722.5 121182.5 8787.5 121317.5 ;
      RECT  8532.5 121182.5 8597.5 121317.5 ;
      RECT  8532.5 120297.5 8597.5 120432.5 ;
      RECT  8722.5 120297.5 8787.5 120432.5 ;
      RECT  8722.5 120297.5 8787.5 120432.5 ;
      RECT  8532.5 120297.5 8597.5 120432.5 ;
      RECT  8892.5 121272.5 8957.5 121407.5 ;
      RECT  8892.5 120297.5 8957.5 120432.5 ;
      RECT  8590.0 120740.0 8655.0 120875.0 ;
      RECT  8590.0 120740.0 8655.0 120875.0 ;
      RECT  8755.0 120775.0 8820.0 120840.0 ;
      RECT  8465.0 121492.5 9025.0 121557.5 ;
      RECT  8465.0 120147.5 9025.0 120212.5 ;
      RECT  8892.5 121710.0 8957.5 121525.0 ;
      RECT  8892.5 122870.0 8957.5 122685.0 ;
      RECT  8532.5 122752.5 8597.5 122902.5 ;
      RECT  8532.5 121867.5 8597.5 121492.5 ;
      RECT  8722.5 122752.5 8787.5 121867.5 ;
      RECT  8532.5 121867.5 8597.5 121732.5 ;
      RECT  8722.5 121867.5 8787.5 121732.5 ;
      RECT  8722.5 121867.5 8787.5 121732.5 ;
      RECT  8532.5 121867.5 8597.5 121732.5 ;
      RECT  8532.5 122752.5 8597.5 122617.5 ;
      RECT  8722.5 122752.5 8787.5 122617.5 ;
      RECT  8722.5 122752.5 8787.5 122617.5 ;
      RECT  8532.5 122752.5 8597.5 122617.5 ;
      RECT  8892.5 121777.5 8957.5 121642.5 ;
      RECT  8892.5 122752.5 8957.5 122617.5 ;
      RECT  8590.0 122310.0 8655.0 122175.0 ;
      RECT  8590.0 122310.0 8655.0 122175.0 ;
      RECT  8755.0 122275.0 8820.0 122210.0 ;
      RECT  8465.0 121557.5 9025.0 121492.5 ;
      RECT  8465.0 122902.5 9025.0 122837.5 ;
      RECT  8892.5 124030.0 8957.5 124215.0 ;
      RECT  8892.5 122870.0 8957.5 123055.0 ;
      RECT  8532.5 122987.5 8597.5 122837.5 ;
      RECT  8532.5 123872.5 8597.5 124247.5 ;
      RECT  8722.5 122987.5 8787.5 123872.5 ;
      RECT  8532.5 123872.5 8597.5 124007.5 ;
      RECT  8722.5 123872.5 8787.5 124007.5 ;
      RECT  8722.5 123872.5 8787.5 124007.5 ;
      RECT  8532.5 123872.5 8597.5 124007.5 ;
      RECT  8532.5 122987.5 8597.5 123122.5 ;
      RECT  8722.5 122987.5 8787.5 123122.5 ;
      RECT  8722.5 122987.5 8787.5 123122.5 ;
      RECT  8532.5 122987.5 8597.5 123122.5 ;
      RECT  8892.5 123962.5 8957.5 124097.5 ;
      RECT  8892.5 122987.5 8957.5 123122.5 ;
      RECT  8590.0 123430.0 8655.0 123565.0 ;
      RECT  8590.0 123430.0 8655.0 123565.0 ;
      RECT  8755.0 123465.0 8820.0 123530.0 ;
      RECT  8465.0 124182.5 9025.0 124247.5 ;
      RECT  8465.0 122837.5 9025.0 122902.5 ;
      RECT  8892.5 124400.0 8957.5 124215.0 ;
      RECT  8892.5 125560.0 8957.5 125375.0 ;
      RECT  8532.5 125442.5 8597.5 125592.5 ;
      RECT  8532.5 124557.5 8597.5 124182.5 ;
      RECT  8722.5 125442.5 8787.5 124557.5 ;
      RECT  8532.5 124557.5 8597.5 124422.5 ;
      RECT  8722.5 124557.5 8787.5 124422.5 ;
      RECT  8722.5 124557.5 8787.5 124422.5 ;
      RECT  8532.5 124557.5 8597.5 124422.5 ;
      RECT  8532.5 125442.5 8597.5 125307.5 ;
      RECT  8722.5 125442.5 8787.5 125307.5 ;
      RECT  8722.5 125442.5 8787.5 125307.5 ;
      RECT  8532.5 125442.5 8597.5 125307.5 ;
      RECT  8892.5 124467.5 8957.5 124332.5 ;
      RECT  8892.5 125442.5 8957.5 125307.5 ;
      RECT  8590.0 125000.0 8655.0 124865.0 ;
      RECT  8590.0 125000.0 8655.0 124865.0 ;
      RECT  8755.0 124965.0 8820.0 124900.0 ;
      RECT  8465.0 124247.5 9025.0 124182.5 ;
      RECT  8465.0 125592.5 9025.0 125527.5 ;
      RECT  8892.5 126720.0 8957.5 126905.0 ;
      RECT  8892.5 125560.0 8957.5 125745.0 ;
      RECT  8532.5 125677.5 8597.5 125527.5 ;
      RECT  8532.5 126562.5 8597.5 126937.5 ;
      RECT  8722.5 125677.5 8787.5 126562.5 ;
      RECT  8532.5 126562.5 8597.5 126697.5 ;
      RECT  8722.5 126562.5 8787.5 126697.5 ;
      RECT  8722.5 126562.5 8787.5 126697.5 ;
      RECT  8532.5 126562.5 8597.5 126697.5 ;
      RECT  8532.5 125677.5 8597.5 125812.5 ;
      RECT  8722.5 125677.5 8787.5 125812.5 ;
      RECT  8722.5 125677.5 8787.5 125812.5 ;
      RECT  8532.5 125677.5 8597.5 125812.5 ;
      RECT  8892.5 126652.5 8957.5 126787.5 ;
      RECT  8892.5 125677.5 8957.5 125812.5 ;
      RECT  8590.0 126120.0 8655.0 126255.0 ;
      RECT  8590.0 126120.0 8655.0 126255.0 ;
      RECT  8755.0 126155.0 8820.0 126220.0 ;
      RECT  8465.0 126872.5 9025.0 126937.5 ;
      RECT  8465.0 125527.5 9025.0 125592.5 ;
      RECT  8892.5 127090.0 8957.5 126905.0 ;
      RECT  8892.5 128250.0 8957.5 128065.0 ;
      RECT  8532.5 128132.5 8597.5 128282.5 ;
      RECT  8532.5 127247.5 8597.5 126872.5 ;
      RECT  8722.5 128132.5 8787.5 127247.5 ;
      RECT  8532.5 127247.5 8597.5 127112.5 ;
      RECT  8722.5 127247.5 8787.5 127112.5 ;
      RECT  8722.5 127247.5 8787.5 127112.5 ;
      RECT  8532.5 127247.5 8597.5 127112.5 ;
      RECT  8532.5 128132.5 8597.5 127997.5 ;
      RECT  8722.5 128132.5 8787.5 127997.5 ;
      RECT  8722.5 128132.5 8787.5 127997.5 ;
      RECT  8532.5 128132.5 8597.5 127997.5 ;
      RECT  8892.5 127157.5 8957.5 127022.5 ;
      RECT  8892.5 128132.5 8957.5 127997.5 ;
      RECT  8590.0 127690.0 8655.0 127555.0 ;
      RECT  8590.0 127690.0 8655.0 127555.0 ;
      RECT  8755.0 127655.0 8820.0 127590.0 ;
      RECT  8465.0 126937.5 9025.0 126872.5 ;
      RECT  8465.0 128282.5 9025.0 128217.5 ;
      RECT  8892.5 129410.0 8957.5 129595.0 ;
      RECT  8892.5 128250.0 8957.5 128435.0 ;
      RECT  8532.5 128367.5 8597.5 128217.5 ;
      RECT  8532.5 129252.5 8597.5 129627.5 ;
      RECT  8722.5 128367.5 8787.5 129252.5 ;
      RECT  8532.5 129252.5 8597.5 129387.5 ;
      RECT  8722.5 129252.5 8787.5 129387.5 ;
      RECT  8722.5 129252.5 8787.5 129387.5 ;
      RECT  8532.5 129252.5 8597.5 129387.5 ;
      RECT  8532.5 128367.5 8597.5 128502.5 ;
      RECT  8722.5 128367.5 8787.5 128502.5 ;
      RECT  8722.5 128367.5 8787.5 128502.5 ;
      RECT  8532.5 128367.5 8597.5 128502.5 ;
      RECT  8892.5 129342.5 8957.5 129477.5 ;
      RECT  8892.5 128367.5 8957.5 128502.5 ;
      RECT  8590.0 128810.0 8655.0 128945.0 ;
      RECT  8590.0 128810.0 8655.0 128945.0 ;
      RECT  8755.0 128845.0 8820.0 128910.0 ;
      RECT  8465.0 129562.5 9025.0 129627.5 ;
      RECT  8465.0 128217.5 9025.0 128282.5 ;
      RECT  8892.5 129780.0 8957.5 129595.0 ;
      RECT  8892.5 130940.0 8957.5 130755.0 ;
      RECT  8532.5 130822.5 8597.5 130972.5 ;
      RECT  8532.5 129937.5 8597.5 129562.5 ;
      RECT  8722.5 130822.5 8787.5 129937.5 ;
      RECT  8532.5 129937.5 8597.5 129802.5 ;
      RECT  8722.5 129937.5 8787.5 129802.5 ;
      RECT  8722.5 129937.5 8787.5 129802.5 ;
      RECT  8532.5 129937.5 8597.5 129802.5 ;
      RECT  8532.5 130822.5 8597.5 130687.5 ;
      RECT  8722.5 130822.5 8787.5 130687.5 ;
      RECT  8722.5 130822.5 8787.5 130687.5 ;
      RECT  8532.5 130822.5 8597.5 130687.5 ;
      RECT  8892.5 129847.5 8957.5 129712.5 ;
      RECT  8892.5 130822.5 8957.5 130687.5 ;
      RECT  8590.0 130380.0 8655.0 130245.0 ;
      RECT  8590.0 130380.0 8655.0 130245.0 ;
      RECT  8755.0 130345.0 8820.0 130280.0 ;
      RECT  8465.0 129627.5 9025.0 129562.5 ;
      RECT  8465.0 130972.5 9025.0 130907.5 ;
      RECT  8892.5 132100.0 8957.5 132285.0 ;
      RECT  8892.5 130940.0 8957.5 131125.0 ;
      RECT  8532.5 131057.5 8597.5 130907.5 ;
      RECT  8532.5 131942.5 8597.5 132317.5 ;
      RECT  8722.5 131057.5 8787.5 131942.5 ;
      RECT  8532.5 131942.5 8597.5 132077.5 ;
      RECT  8722.5 131942.5 8787.5 132077.5 ;
      RECT  8722.5 131942.5 8787.5 132077.5 ;
      RECT  8532.5 131942.5 8597.5 132077.5 ;
      RECT  8532.5 131057.5 8597.5 131192.5 ;
      RECT  8722.5 131057.5 8787.5 131192.5 ;
      RECT  8722.5 131057.5 8787.5 131192.5 ;
      RECT  8532.5 131057.5 8597.5 131192.5 ;
      RECT  8892.5 132032.5 8957.5 132167.5 ;
      RECT  8892.5 131057.5 8957.5 131192.5 ;
      RECT  8590.0 131500.0 8655.0 131635.0 ;
      RECT  8590.0 131500.0 8655.0 131635.0 ;
      RECT  8755.0 131535.0 8820.0 131600.0 ;
      RECT  8465.0 132252.5 9025.0 132317.5 ;
      RECT  8465.0 130907.5 9025.0 130972.5 ;
      RECT  8892.5 132470.0 8957.5 132285.0 ;
      RECT  8892.5 133630.0 8957.5 133445.0 ;
      RECT  8532.5 133512.5 8597.5 133662.5 ;
      RECT  8532.5 132627.5 8597.5 132252.5 ;
      RECT  8722.5 133512.5 8787.5 132627.5 ;
      RECT  8532.5 132627.5 8597.5 132492.5 ;
      RECT  8722.5 132627.5 8787.5 132492.5 ;
      RECT  8722.5 132627.5 8787.5 132492.5 ;
      RECT  8532.5 132627.5 8597.5 132492.5 ;
      RECT  8532.5 133512.5 8597.5 133377.5 ;
      RECT  8722.5 133512.5 8787.5 133377.5 ;
      RECT  8722.5 133512.5 8787.5 133377.5 ;
      RECT  8532.5 133512.5 8597.5 133377.5 ;
      RECT  8892.5 132537.5 8957.5 132402.5 ;
      RECT  8892.5 133512.5 8957.5 133377.5 ;
      RECT  8590.0 133070.0 8655.0 132935.0 ;
      RECT  8590.0 133070.0 8655.0 132935.0 ;
      RECT  8755.0 133035.0 8820.0 132970.0 ;
      RECT  8465.0 132317.5 9025.0 132252.5 ;
      RECT  8465.0 133662.5 9025.0 133597.5 ;
      RECT  8892.5 134790.0 8957.5 134975.0 ;
      RECT  8892.5 133630.0 8957.5 133815.0 ;
      RECT  8532.5 133747.5 8597.5 133597.5 ;
      RECT  8532.5 134632.5 8597.5 135007.5 ;
      RECT  8722.5 133747.5 8787.5 134632.5 ;
      RECT  8532.5 134632.5 8597.5 134767.5 ;
      RECT  8722.5 134632.5 8787.5 134767.5 ;
      RECT  8722.5 134632.5 8787.5 134767.5 ;
      RECT  8532.5 134632.5 8597.5 134767.5 ;
      RECT  8532.5 133747.5 8597.5 133882.5 ;
      RECT  8722.5 133747.5 8787.5 133882.5 ;
      RECT  8722.5 133747.5 8787.5 133882.5 ;
      RECT  8532.5 133747.5 8597.5 133882.5 ;
      RECT  8892.5 134722.5 8957.5 134857.5 ;
      RECT  8892.5 133747.5 8957.5 133882.5 ;
      RECT  8590.0 134190.0 8655.0 134325.0 ;
      RECT  8590.0 134190.0 8655.0 134325.0 ;
      RECT  8755.0 134225.0 8820.0 134290.0 ;
      RECT  8465.0 134942.5 9025.0 135007.5 ;
      RECT  8465.0 133597.5 9025.0 133662.5 ;
      RECT  8892.5 135160.0 8957.5 134975.0 ;
      RECT  8892.5 136320.0 8957.5 136135.0 ;
      RECT  8532.5 136202.5 8597.5 136352.5 ;
      RECT  8532.5 135317.5 8597.5 134942.5 ;
      RECT  8722.5 136202.5 8787.5 135317.5 ;
      RECT  8532.5 135317.5 8597.5 135182.5 ;
      RECT  8722.5 135317.5 8787.5 135182.5 ;
      RECT  8722.5 135317.5 8787.5 135182.5 ;
      RECT  8532.5 135317.5 8597.5 135182.5 ;
      RECT  8532.5 136202.5 8597.5 136067.5 ;
      RECT  8722.5 136202.5 8787.5 136067.5 ;
      RECT  8722.5 136202.5 8787.5 136067.5 ;
      RECT  8532.5 136202.5 8597.5 136067.5 ;
      RECT  8892.5 135227.5 8957.5 135092.5 ;
      RECT  8892.5 136202.5 8957.5 136067.5 ;
      RECT  8590.0 135760.0 8655.0 135625.0 ;
      RECT  8590.0 135760.0 8655.0 135625.0 ;
      RECT  8755.0 135725.0 8820.0 135660.0 ;
      RECT  8465.0 135007.5 9025.0 134942.5 ;
      RECT  8465.0 136352.5 9025.0 136287.5 ;
      RECT  8892.5 137480.0 8957.5 137665.0 ;
      RECT  8892.5 136320.0 8957.5 136505.0 ;
      RECT  8532.5 136437.5 8597.5 136287.5 ;
      RECT  8532.5 137322.5 8597.5 137697.5 ;
      RECT  8722.5 136437.5 8787.5 137322.5 ;
      RECT  8532.5 137322.5 8597.5 137457.5 ;
      RECT  8722.5 137322.5 8787.5 137457.5 ;
      RECT  8722.5 137322.5 8787.5 137457.5 ;
      RECT  8532.5 137322.5 8597.5 137457.5 ;
      RECT  8532.5 136437.5 8597.5 136572.5 ;
      RECT  8722.5 136437.5 8787.5 136572.5 ;
      RECT  8722.5 136437.5 8787.5 136572.5 ;
      RECT  8532.5 136437.5 8597.5 136572.5 ;
      RECT  8892.5 137412.5 8957.5 137547.5 ;
      RECT  8892.5 136437.5 8957.5 136572.5 ;
      RECT  8590.0 136880.0 8655.0 137015.0 ;
      RECT  8590.0 136880.0 8655.0 137015.0 ;
      RECT  8755.0 136915.0 8820.0 136980.0 ;
      RECT  8465.0 137632.5 9025.0 137697.5 ;
      RECT  8465.0 136287.5 9025.0 136352.5 ;
      RECT  8892.5 137850.0 8957.5 137665.0 ;
      RECT  8892.5 139010.0 8957.5 138825.0 ;
      RECT  8532.5 138892.5 8597.5 139042.5 ;
      RECT  8532.5 138007.5 8597.5 137632.5 ;
      RECT  8722.5 138892.5 8787.5 138007.5 ;
      RECT  8532.5 138007.5 8597.5 137872.5 ;
      RECT  8722.5 138007.5 8787.5 137872.5 ;
      RECT  8722.5 138007.5 8787.5 137872.5 ;
      RECT  8532.5 138007.5 8597.5 137872.5 ;
      RECT  8532.5 138892.5 8597.5 138757.5 ;
      RECT  8722.5 138892.5 8787.5 138757.5 ;
      RECT  8722.5 138892.5 8787.5 138757.5 ;
      RECT  8532.5 138892.5 8597.5 138757.5 ;
      RECT  8892.5 137917.5 8957.5 137782.5 ;
      RECT  8892.5 138892.5 8957.5 138757.5 ;
      RECT  8590.0 138450.0 8655.0 138315.0 ;
      RECT  8590.0 138450.0 8655.0 138315.0 ;
      RECT  8755.0 138415.0 8820.0 138350.0 ;
      RECT  8465.0 137697.5 9025.0 137632.5 ;
      RECT  8465.0 139042.5 9025.0 138977.5 ;
      RECT  8892.5 140170.0 8957.5 140355.0 ;
      RECT  8892.5 139010.0 8957.5 139195.0 ;
      RECT  8532.5 139127.5 8597.5 138977.5 ;
      RECT  8532.5 140012.5 8597.5 140387.5 ;
      RECT  8722.5 139127.5 8787.5 140012.5 ;
      RECT  8532.5 140012.5 8597.5 140147.5 ;
      RECT  8722.5 140012.5 8787.5 140147.5 ;
      RECT  8722.5 140012.5 8787.5 140147.5 ;
      RECT  8532.5 140012.5 8597.5 140147.5 ;
      RECT  8532.5 139127.5 8597.5 139262.5 ;
      RECT  8722.5 139127.5 8787.5 139262.5 ;
      RECT  8722.5 139127.5 8787.5 139262.5 ;
      RECT  8532.5 139127.5 8597.5 139262.5 ;
      RECT  8892.5 140102.5 8957.5 140237.5 ;
      RECT  8892.5 139127.5 8957.5 139262.5 ;
      RECT  8590.0 139570.0 8655.0 139705.0 ;
      RECT  8590.0 139570.0 8655.0 139705.0 ;
      RECT  8755.0 139605.0 8820.0 139670.0 ;
      RECT  8465.0 140322.5 9025.0 140387.5 ;
      RECT  8465.0 138977.5 9025.0 139042.5 ;
      RECT  8892.5 140540.0 8957.5 140355.0 ;
      RECT  8892.5 141700.0 8957.5 141515.0 ;
      RECT  8532.5 141582.5 8597.5 141732.5 ;
      RECT  8532.5 140697.5 8597.5 140322.5 ;
      RECT  8722.5 141582.5 8787.5 140697.5 ;
      RECT  8532.5 140697.5 8597.5 140562.5 ;
      RECT  8722.5 140697.5 8787.5 140562.5 ;
      RECT  8722.5 140697.5 8787.5 140562.5 ;
      RECT  8532.5 140697.5 8597.5 140562.5 ;
      RECT  8532.5 141582.5 8597.5 141447.5 ;
      RECT  8722.5 141582.5 8787.5 141447.5 ;
      RECT  8722.5 141582.5 8787.5 141447.5 ;
      RECT  8532.5 141582.5 8597.5 141447.5 ;
      RECT  8892.5 140607.5 8957.5 140472.5 ;
      RECT  8892.5 141582.5 8957.5 141447.5 ;
      RECT  8590.0 141140.0 8655.0 141005.0 ;
      RECT  8590.0 141140.0 8655.0 141005.0 ;
      RECT  8755.0 141105.0 8820.0 141040.0 ;
      RECT  8465.0 140387.5 9025.0 140322.5 ;
      RECT  8465.0 141732.5 9025.0 141667.5 ;
      RECT  8892.5 142860.0 8957.5 143045.0 ;
      RECT  8892.5 141700.0 8957.5 141885.0 ;
      RECT  8532.5 141817.5 8597.5 141667.5 ;
      RECT  8532.5 142702.5 8597.5 143077.5 ;
      RECT  8722.5 141817.5 8787.5 142702.5 ;
      RECT  8532.5 142702.5 8597.5 142837.5 ;
      RECT  8722.5 142702.5 8787.5 142837.5 ;
      RECT  8722.5 142702.5 8787.5 142837.5 ;
      RECT  8532.5 142702.5 8597.5 142837.5 ;
      RECT  8532.5 141817.5 8597.5 141952.5 ;
      RECT  8722.5 141817.5 8787.5 141952.5 ;
      RECT  8722.5 141817.5 8787.5 141952.5 ;
      RECT  8532.5 141817.5 8597.5 141952.5 ;
      RECT  8892.5 142792.5 8957.5 142927.5 ;
      RECT  8892.5 141817.5 8957.5 141952.5 ;
      RECT  8590.0 142260.0 8655.0 142395.0 ;
      RECT  8590.0 142260.0 8655.0 142395.0 ;
      RECT  8755.0 142295.0 8820.0 142360.0 ;
      RECT  8465.0 143012.5 9025.0 143077.5 ;
      RECT  8465.0 141667.5 9025.0 141732.5 ;
      RECT  8892.5 143230.0 8957.5 143045.0 ;
      RECT  8892.5 144390.0 8957.5 144205.0 ;
      RECT  8532.5 144272.5 8597.5 144422.5 ;
      RECT  8532.5 143387.5 8597.5 143012.5 ;
      RECT  8722.5 144272.5 8787.5 143387.5 ;
      RECT  8532.5 143387.5 8597.5 143252.5 ;
      RECT  8722.5 143387.5 8787.5 143252.5 ;
      RECT  8722.5 143387.5 8787.5 143252.5 ;
      RECT  8532.5 143387.5 8597.5 143252.5 ;
      RECT  8532.5 144272.5 8597.5 144137.5 ;
      RECT  8722.5 144272.5 8787.5 144137.5 ;
      RECT  8722.5 144272.5 8787.5 144137.5 ;
      RECT  8532.5 144272.5 8597.5 144137.5 ;
      RECT  8892.5 143297.5 8957.5 143162.5 ;
      RECT  8892.5 144272.5 8957.5 144137.5 ;
      RECT  8590.0 143830.0 8655.0 143695.0 ;
      RECT  8590.0 143830.0 8655.0 143695.0 ;
      RECT  8755.0 143795.0 8820.0 143730.0 ;
      RECT  8465.0 143077.5 9025.0 143012.5 ;
      RECT  8465.0 144422.5 9025.0 144357.5 ;
      RECT  8892.5 145550.0 8957.5 145735.0 ;
      RECT  8892.5 144390.0 8957.5 144575.0 ;
      RECT  8532.5 144507.5 8597.5 144357.5 ;
      RECT  8532.5 145392.5 8597.5 145767.5 ;
      RECT  8722.5 144507.5 8787.5 145392.5 ;
      RECT  8532.5 145392.5 8597.5 145527.5 ;
      RECT  8722.5 145392.5 8787.5 145527.5 ;
      RECT  8722.5 145392.5 8787.5 145527.5 ;
      RECT  8532.5 145392.5 8597.5 145527.5 ;
      RECT  8532.5 144507.5 8597.5 144642.5 ;
      RECT  8722.5 144507.5 8787.5 144642.5 ;
      RECT  8722.5 144507.5 8787.5 144642.5 ;
      RECT  8532.5 144507.5 8597.5 144642.5 ;
      RECT  8892.5 145482.5 8957.5 145617.5 ;
      RECT  8892.5 144507.5 8957.5 144642.5 ;
      RECT  8590.0 144950.0 8655.0 145085.0 ;
      RECT  8590.0 144950.0 8655.0 145085.0 ;
      RECT  8755.0 144985.0 8820.0 145050.0 ;
      RECT  8465.0 145702.5 9025.0 145767.5 ;
      RECT  8465.0 144357.5 9025.0 144422.5 ;
      RECT  8892.5 145920.0 8957.5 145735.0 ;
      RECT  8892.5 147080.0 8957.5 146895.0 ;
      RECT  8532.5 146962.5 8597.5 147112.5 ;
      RECT  8532.5 146077.5 8597.5 145702.5 ;
      RECT  8722.5 146962.5 8787.5 146077.5 ;
      RECT  8532.5 146077.5 8597.5 145942.5 ;
      RECT  8722.5 146077.5 8787.5 145942.5 ;
      RECT  8722.5 146077.5 8787.5 145942.5 ;
      RECT  8532.5 146077.5 8597.5 145942.5 ;
      RECT  8532.5 146962.5 8597.5 146827.5 ;
      RECT  8722.5 146962.5 8787.5 146827.5 ;
      RECT  8722.5 146962.5 8787.5 146827.5 ;
      RECT  8532.5 146962.5 8597.5 146827.5 ;
      RECT  8892.5 145987.5 8957.5 145852.5 ;
      RECT  8892.5 146962.5 8957.5 146827.5 ;
      RECT  8590.0 146520.0 8655.0 146385.0 ;
      RECT  8590.0 146520.0 8655.0 146385.0 ;
      RECT  8755.0 146485.0 8820.0 146420.0 ;
      RECT  8465.0 145767.5 9025.0 145702.5 ;
      RECT  8465.0 147112.5 9025.0 147047.5 ;
      RECT  8892.5 148240.0 8957.5 148425.0 ;
      RECT  8892.5 147080.0 8957.5 147265.0 ;
      RECT  8532.5 147197.5 8597.5 147047.5 ;
      RECT  8532.5 148082.5 8597.5 148457.5 ;
      RECT  8722.5 147197.5 8787.5 148082.5 ;
      RECT  8532.5 148082.5 8597.5 148217.5 ;
      RECT  8722.5 148082.5 8787.5 148217.5 ;
      RECT  8722.5 148082.5 8787.5 148217.5 ;
      RECT  8532.5 148082.5 8597.5 148217.5 ;
      RECT  8532.5 147197.5 8597.5 147332.5 ;
      RECT  8722.5 147197.5 8787.5 147332.5 ;
      RECT  8722.5 147197.5 8787.5 147332.5 ;
      RECT  8532.5 147197.5 8597.5 147332.5 ;
      RECT  8892.5 148172.5 8957.5 148307.5 ;
      RECT  8892.5 147197.5 8957.5 147332.5 ;
      RECT  8590.0 147640.0 8655.0 147775.0 ;
      RECT  8590.0 147640.0 8655.0 147775.0 ;
      RECT  8755.0 147675.0 8820.0 147740.0 ;
      RECT  8465.0 148392.5 9025.0 148457.5 ;
      RECT  8465.0 147047.5 9025.0 147112.5 ;
      RECT  8892.5 148610.0 8957.5 148425.0 ;
      RECT  8892.5 149770.0 8957.5 149585.0 ;
      RECT  8532.5 149652.5 8597.5 149802.5 ;
      RECT  8532.5 148767.5 8597.5 148392.5 ;
      RECT  8722.5 149652.5 8787.5 148767.5 ;
      RECT  8532.5 148767.5 8597.5 148632.5 ;
      RECT  8722.5 148767.5 8787.5 148632.5 ;
      RECT  8722.5 148767.5 8787.5 148632.5 ;
      RECT  8532.5 148767.5 8597.5 148632.5 ;
      RECT  8532.5 149652.5 8597.5 149517.5 ;
      RECT  8722.5 149652.5 8787.5 149517.5 ;
      RECT  8722.5 149652.5 8787.5 149517.5 ;
      RECT  8532.5 149652.5 8597.5 149517.5 ;
      RECT  8892.5 148677.5 8957.5 148542.5 ;
      RECT  8892.5 149652.5 8957.5 149517.5 ;
      RECT  8590.0 149210.0 8655.0 149075.0 ;
      RECT  8590.0 149210.0 8655.0 149075.0 ;
      RECT  8755.0 149175.0 8820.0 149110.0 ;
      RECT  8465.0 148457.5 9025.0 148392.5 ;
      RECT  8465.0 149802.5 9025.0 149737.5 ;
      RECT  8892.5 150930.0 8957.5 151115.0 ;
      RECT  8892.5 149770.0 8957.5 149955.0 ;
      RECT  8532.5 149887.5 8597.5 149737.5 ;
      RECT  8532.5 150772.5 8597.5 151147.5 ;
      RECT  8722.5 149887.5 8787.5 150772.5 ;
      RECT  8532.5 150772.5 8597.5 150907.5 ;
      RECT  8722.5 150772.5 8787.5 150907.5 ;
      RECT  8722.5 150772.5 8787.5 150907.5 ;
      RECT  8532.5 150772.5 8597.5 150907.5 ;
      RECT  8532.5 149887.5 8597.5 150022.5 ;
      RECT  8722.5 149887.5 8787.5 150022.5 ;
      RECT  8722.5 149887.5 8787.5 150022.5 ;
      RECT  8532.5 149887.5 8597.5 150022.5 ;
      RECT  8892.5 150862.5 8957.5 150997.5 ;
      RECT  8892.5 149887.5 8957.5 150022.5 ;
      RECT  8590.0 150330.0 8655.0 150465.0 ;
      RECT  8590.0 150330.0 8655.0 150465.0 ;
      RECT  8755.0 150365.0 8820.0 150430.0 ;
      RECT  8465.0 151082.5 9025.0 151147.5 ;
      RECT  8465.0 149737.5 9025.0 149802.5 ;
      RECT  8892.5 151300.0 8957.5 151115.0 ;
      RECT  8892.5 152460.0 8957.5 152275.0 ;
      RECT  8532.5 152342.5 8597.5 152492.5 ;
      RECT  8532.5 151457.5 8597.5 151082.5 ;
      RECT  8722.5 152342.5 8787.5 151457.5 ;
      RECT  8532.5 151457.5 8597.5 151322.5 ;
      RECT  8722.5 151457.5 8787.5 151322.5 ;
      RECT  8722.5 151457.5 8787.5 151322.5 ;
      RECT  8532.5 151457.5 8597.5 151322.5 ;
      RECT  8532.5 152342.5 8597.5 152207.5 ;
      RECT  8722.5 152342.5 8787.5 152207.5 ;
      RECT  8722.5 152342.5 8787.5 152207.5 ;
      RECT  8532.5 152342.5 8597.5 152207.5 ;
      RECT  8892.5 151367.5 8957.5 151232.5 ;
      RECT  8892.5 152342.5 8957.5 152207.5 ;
      RECT  8590.0 151900.0 8655.0 151765.0 ;
      RECT  8590.0 151900.0 8655.0 151765.0 ;
      RECT  8755.0 151865.0 8820.0 151800.0 ;
      RECT  8465.0 151147.5 9025.0 151082.5 ;
      RECT  8465.0 152492.5 9025.0 152427.5 ;
      RECT  8892.5 153620.0 8957.5 153805.0 ;
      RECT  8892.5 152460.0 8957.5 152645.0 ;
      RECT  8532.5 152577.5 8597.5 152427.5 ;
      RECT  8532.5 153462.5 8597.5 153837.5 ;
      RECT  8722.5 152577.5 8787.5 153462.5 ;
      RECT  8532.5 153462.5 8597.5 153597.5 ;
      RECT  8722.5 153462.5 8787.5 153597.5 ;
      RECT  8722.5 153462.5 8787.5 153597.5 ;
      RECT  8532.5 153462.5 8597.5 153597.5 ;
      RECT  8532.5 152577.5 8597.5 152712.5 ;
      RECT  8722.5 152577.5 8787.5 152712.5 ;
      RECT  8722.5 152577.5 8787.5 152712.5 ;
      RECT  8532.5 152577.5 8597.5 152712.5 ;
      RECT  8892.5 153552.5 8957.5 153687.5 ;
      RECT  8892.5 152577.5 8957.5 152712.5 ;
      RECT  8590.0 153020.0 8655.0 153155.0 ;
      RECT  8590.0 153020.0 8655.0 153155.0 ;
      RECT  8755.0 153055.0 8820.0 153120.0 ;
      RECT  8465.0 153772.5 9025.0 153837.5 ;
      RECT  8465.0 152427.5 9025.0 152492.5 ;
      RECT  8892.5 153990.0 8957.5 153805.0 ;
      RECT  8892.5 155150.0 8957.5 154965.0 ;
      RECT  8532.5 155032.5 8597.5 155182.5 ;
      RECT  8532.5 154147.5 8597.5 153772.5 ;
      RECT  8722.5 155032.5 8787.5 154147.5 ;
      RECT  8532.5 154147.5 8597.5 154012.5 ;
      RECT  8722.5 154147.5 8787.5 154012.5 ;
      RECT  8722.5 154147.5 8787.5 154012.5 ;
      RECT  8532.5 154147.5 8597.5 154012.5 ;
      RECT  8532.5 155032.5 8597.5 154897.5 ;
      RECT  8722.5 155032.5 8787.5 154897.5 ;
      RECT  8722.5 155032.5 8787.5 154897.5 ;
      RECT  8532.5 155032.5 8597.5 154897.5 ;
      RECT  8892.5 154057.5 8957.5 153922.5 ;
      RECT  8892.5 155032.5 8957.5 154897.5 ;
      RECT  8590.0 154590.0 8655.0 154455.0 ;
      RECT  8590.0 154590.0 8655.0 154455.0 ;
      RECT  8755.0 154555.0 8820.0 154490.0 ;
      RECT  8465.0 153837.5 9025.0 153772.5 ;
      RECT  8465.0 155182.5 9025.0 155117.5 ;
      RECT  8892.5 156310.0 8957.5 156495.0 ;
      RECT  8892.5 155150.0 8957.5 155335.0 ;
      RECT  8532.5 155267.5 8597.5 155117.5 ;
      RECT  8532.5 156152.5 8597.5 156527.5 ;
      RECT  8722.5 155267.5 8787.5 156152.5 ;
      RECT  8532.5 156152.5 8597.5 156287.5 ;
      RECT  8722.5 156152.5 8787.5 156287.5 ;
      RECT  8722.5 156152.5 8787.5 156287.5 ;
      RECT  8532.5 156152.5 8597.5 156287.5 ;
      RECT  8532.5 155267.5 8597.5 155402.5 ;
      RECT  8722.5 155267.5 8787.5 155402.5 ;
      RECT  8722.5 155267.5 8787.5 155402.5 ;
      RECT  8532.5 155267.5 8597.5 155402.5 ;
      RECT  8892.5 156242.5 8957.5 156377.5 ;
      RECT  8892.5 155267.5 8957.5 155402.5 ;
      RECT  8590.0 155710.0 8655.0 155845.0 ;
      RECT  8590.0 155710.0 8655.0 155845.0 ;
      RECT  8755.0 155745.0 8820.0 155810.0 ;
      RECT  8465.0 156462.5 9025.0 156527.5 ;
      RECT  8465.0 155117.5 9025.0 155182.5 ;
      RECT  8892.5 156680.0 8957.5 156495.0 ;
      RECT  8892.5 157840.0 8957.5 157655.0 ;
      RECT  8532.5 157722.5 8597.5 157872.5 ;
      RECT  8532.5 156837.5 8597.5 156462.5 ;
      RECT  8722.5 157722.5 8787.5 156837.5 ;
      RECT  8532.5 156837.5 8597.5 156702.5 ;
      RECT  8722.5 156837.5 8787.5 156702.5 ;
      RECT  8722.5 156837.5 8787.5 156702.5 ;
      RECT  8532.5 156837.5 8597.5 156702.5 ;
      RECT  8532.5 157722.5 8597.5 157587.5 ;
      RECT  8722.5 157722.5 8787.5 157587.5 ;
      RECT  8722.5 157722.5 8787.5 157587.5 ;
      RECT  8532.5 157722.5 8597.5 157587.5 ;
      RECT  8892.5 156747.5 8957.5 156612.5 ;
      RECT  8892.5 157722.5 8957.5 157587.5 ;
      RECT  8590.0 157280.0 8655.0 157145.0 ;
      RECT  8590.0 157280.0 8655.0 157145.0 ;
      RECT  8755.0 157245.0 8820.0 157180.0 ;
      RECT  8465.0 156527.5 9025.0 156462.5 ;
      RECT  8465.0 157872.5 9025.0 157807.5 ;
      RECT  8892.5 159000.0 8957.5 159185.0 ;
      RECT  8892.5 157840.0 8957.5 158025.0 ;
      RECT  8532.5 157957.5 8597.5 157807.5 ;
      RECT  8532.5 158842.5 8597.5 159217.5 ;
      RECT  8722.5 157957.5 8787.5 158842.5 ;
      RECT  8532.5 158842.5 8597.5 158977.5 ;
      RECT  8722.5 158842.5 8787.5 158977.5 ;
      RECT  8722.5 158842.5 8787.5 158977.5 ;
      RECT  8532.5 158842.5 8597.5 158977.5 ;
      RECT  8532.5 157957.5 8597.5 158092.5 ;
      RECT  8722.5 157957.5 8787.5 158092.5 ;
      RECT  8722.5 157957.5 8787.5 158092.5 ;
      RECT  8532.5 157957.5 8597.5 158092.5 ;
      RECT  8892.5 158932.5 8957.5 159067.5 ;
      RECT  8892.5 157957.5 8957.5 158092.5 ;
      RECT  8590.0 158400.0 8655.0 158535.0 ;
      RECT  8590.0 158400.0 8655.0 158535.0 ;
      RECT  8755.0 158435.0 8820.0 158500.0 ;
      RECT  8465.0 159152.5 9025.0 159217.5 ;
      RECT  8465.0 157807.5 9025.0 157872.5 ;
      RECT  8892.5 159370.0 8957.5 159185.0 ;
      RECT  8892.5 160530.0 8957.5 160345.0 ;
      RECT  8532.5 160412.5 8597.5 160562.5 ;
      RECT  8532.5 159527.5 8597.5 159152.5 ;
      RECT  8722.5 160412.5 8787.5 159527.5 ;
      RECT  8532.5 159527.5 8597.5 159392.5 ;
      RECT  8722.5 159527.5 8787.5 159392.5 ;
      RECT  8722.5 159527.5 8787.5 159392.5 ;
      RECT  8532.5 159527.5 8597.5 159392.5 ;
      RECT  8532.5 160412.5 8597.5 160277.5 ;
      RECT  8722.5 160412.5 8787.5 160277.5 ;
      RECT  8722.5 160412.5 8787.5 160277.5 ;
      RECT  8532.5 160412.5 8597.5 160277.5 ;
      RECT  8892.5 159437.5 8957.5 159302.5 ;
      RECT  8892.5 160412.5 8957.5 160277.5 ;
      RECT  8590.0 159970.0 8655.0 159835.0 ;
      RECT  8590.0 159970.0 8655.0 159835.0 ;
      RECT  8755.0 159935.0 8820.0 159870.0 ;
      RECT  8465.0 159217.5 9025.0 159152.5 ;
      RECT  8465.0 160562.5 9025.0 160497.5 ;
      RECT  8892.5 161690.0 8957.5 161875.0 ;
      RECT  8892.5 160530.0 8957.5 160715.0 ;
      RECT  8532.5 160647.5 8597.5 160497.5 ;
      RECT  8532.5 161532.5 8597.5 161907.5 ;
      RECT  8722.5 160647.5 8787.5 161532.5 ;
      RECT  8532.5 161532.5 8597.5 161667.5 ;
      RECT  8722.5 161532.5 8787.5 161667.5 ;
      RECT  8722.5 161532.5 8787.5 161667.5 ;
      RECT  8532.5 161532.5 8597.5 161667.5 ;
      RECT  8532.5 160647.5 8597.5 160782.5 ;
      RECT  8722.5 160647.5 8787.5 160782.5 ;
      RECT  8722.5 160647.5 8787.5 160782.5 ;
      RECT  8532.5 160647.5 8597.5 160782.5 ;
      RECT  8892.5 161622.5 8957.5 161757.5 ;
      RECT  8892.5 160647.5 8957.5 160782.5 ;
      RECT  8590.0 161090.0 8655.0 161225.0 ;
      RECT  8590.0 161090.0 8655.0 161225.0 ;
      RECT  8755.0 161125.0 8820.0 161190.0 ;
      RECT  8465.0 161842.5 9025.0 161907.5 ;
      RECT  8465.0 160497.5 9025.0 160562.5 ;
      RECT  8892.5 162060.0 8957.5 161875.0 ;
      RECT  8892.5 163220.0 8957.5 163035.0 ;
      RECT  8532.5 163102.5 8597.5 163252.5 ;
      RECT  8532.5 162217.5 8597.5 161842.5 ;
      RECT  8722.5 163102.5 8787.5 162217.5 ;
      RECT  8532.5 162217.5 8597.5 162082.5 ;
      RECT  8722.5 162217.5 8787.5 162082.5 ;
      RECT  8722.5 162217.5 8787.5 162082.5 ;
      RECT  8532.5 162217.5 8597.5 162082.5 ;
      RECT  8532.5 163102.5 8597.5 162967.5 ;
      RECT  8722.5 163102.5 8787.5 162967.5 ;
      RECT  8722.5 163102.5 8787.5 162967.5 ;
      RECT  8532.5 163102.5 8597.5 162967.5 ;
      RECT  8892.5 162127.5 8957.5 161992.5 ;
      RECT  8892.5 163102.5 8957.5 162967.5 ;
      RECT  8590.0 162660.0 8655.0 162525.0 ;
      RECT  8590.0 162660.0 8655.0 162525.0 ;
      RECT  8755.0 162625.0 8820.0 162560.0 ;
      RECT  8465.0 161907.5 9025.0 161842.5 ;
      RECT  8465.0 163252.5 9025.0 163187.5 ;
      RECT  8892.5 164380.0 8957.5 164565.0 ;
      RECT  8892.5 163220.0 8957.5 163405.0 ;
      RECT  8532.5 163337.5 8597.5 163187.5 ;
      RECT  8532.5 164222.5 8597.5 164597.5 ;
      RECT  8722.5 163337.5 8787.5 164222.5 ;
      RECT  8532.5 164222.5 8597.5 164357.5 ;
      RECT  8722.5 164222.5 8787.5 164357.5 ;
      RECT  8722.5 164222.5 8787.5 164357.5 ;
      RECT  8532.5 164222.5 8597.5 164357.5 ;
      RECT  8532.5 163337.5 8597.5 163472.5 ;
      RECT  8722.5 163337.5 8787.5 163472.5 ;
      RECT  8722.5 163337.5 8787.5 163472.5 ;
      RECT  8532.5 163337.5 8597.5 163472.5 ;
      RECT  8892.5 164312.5 8957.5 164447.5 ;
      RECT  8892.5 163337.5 8957.5 163472.5 ;
      RECT  8590.0 163780.0 8655.0 163915.0 ;
      RECT  8590.0 163780.0 8655.0 163915.0 ;
      RECT  8755.0 163815.0 8820.0 163880.0 ;
      RECT  8465.0 164532.5 9025.0 164597.5 ;
      RECT  8465.0 163187.5 9025.0 163252.5 ;
      RECT  8892.5 164750.0 8957.5 164565.0 ;
      RECT  8892.5 165910.0 8957.5 165725.0 ;
      RECT  8532.5 165792.5 8597.5 165942.5 ;
      RECT  8532.5 164907.5 8597.5 164532.5 ;
      RECT  8722.5 165792.5 8787.5 164907.5 ;
      RECT  8532.5 164907.5 8597.5 164772.5 ;
      RECT  8722.5 164907.5 8787.5 164772.5 ;
      RECT  8722.5 164907.5 8787.5 164772.5 ;
      RECT  8532.5 164907.5 8597.5 164772.5 ;
      RECT  8532.5 165792.5 8597.5 165657.5 ;
      RECT  8722.5 165792.5 8787.5 165657.5 ;
      RECT  8722.5 165792.5 8787.5 165657.5 ;
      RECT  8532.5 165792.5 8597.5 165657.5 ;
      RECT  8892.5 164817.5 8957.5 164682.5 ;
      RECT  8892.5 165792.5 8957.5 165657.5 ;
      RECT  8590.0 165350.0 8655.0 165215.0 ;
      RECT  8590.0 165350.0 8655.0 165215.0 ;
      RECT  8755.0 165315.0 8820.0 165250.0 ;
      RECT  8465.0 164597.5 9025.0 164532.5 ;
      RECT  8465.0 165942.5 9025.0 165877.5 ;
      RECT  8892.5 167070.0 8957.5 167255.0 ;
      RECT  8892.5 165910.0 8957.5 166095.0 ;
      RECT  8532.5 166027.5 8597.5 165877.5 ;
      RECT  8532.5 166912.5 8597.5 167287.5 ;
      RECT  8722.5 166027.5 8787.5 166912.5 ;
      RECT  8532.5 166912.5 8597.5 167047.5 ;
      RECT  8722.5 166912.5 8787.5 167047.5 ;
      RECT  8722.5 166912.5 8787.5 167047.5 ;
      RECT  8532.5 166912.5 8597.5 167047.5 ;
      RECT  8532.5 166027.5 8597.5 166162.5 ;
      RECT  8722.5 166027.5 8787.5 166162.5 ;
      RECT  8722.5 166027.5 8787.5 166162.5 ;
      RECT  8532.5 166027.5 8597.5 166162.5 ;
      RECT  8892.5 167002.5 8957.5 167137.5 ;
      RECT  8892.5 166027.5 8957.5 166162.5 ;
      RECT  8590.0 166470.0 8655.0 166605.0 ;
      RECT  8590.0 166470.0 8655.0 166605.0 ;
      RECT  8755.0 166505.0 8820.0 166570.0 ;
      RECT  8465.0 167222.5 9025.0 167287.5 ;
      RECT  8465.0 165877.5 9025.0 165942.5 ;
      RECT  8892.5 167440.0 8957.5 167255.0 ;
      RECT  8892.5 168600.0 8957.5 168415.0 ;
      RECT  8532.5 168482.5 8597.5 168632.5 ;
      RECT  8532.5 167597.5 8597.5 167222.5 ;
      RECT  8722.5 168482.5 8787.5 167597.5 ;
      RECT  8532.5 167597.5 8597.5 167462.5 ;
      RECT  8722.5 167597.5 8787.5 167462.5 ;
      RECT  8722.5 167597.5 8787.5 167462.5 ;
      RECT  8532.5 167597.5 8597.5 167462.5 ;
      RECT  8532.5 168482.5 8597.5 168347.5 ;
      RECT  8722.5 168482.5 8787.5 168347.5 ;
      RECT  8722.5 168482.5 8787.5 168347.5 ;
      RECT  8532.5 168482.5 8597.5 168347.5 ;
      RECT  8892.5 167507.5 8957.5 167372.5 ;
      RECT  8892.5 168482.5 8957.5 168347.5 ;
      RECT  8590.0 168040.0 8655.0 167905.0 ;
      RECT  8590.0 168040.0 8655.0 167905.0 ;
      RECT  8755.0 168005.0 8820.0 167940.0 ;
      RECT  8465.0 167287.5 9025.0 167222.5 ;
      RECT  8465.0 168632.5 9025.0 168567.5 ;
      RECT  8892.5 169760.0 8957.5 169945.0 ;
      RECT  8892.5 168600.0 8957.5 168785.0 ;
      RECT  8532.5 168717.5 8597.5 168567.5 ;
      RECT  8532.5 169602.5 8597.5 169977.5 ;
      RECT  8722.5 168717.5 8787.5 169602.5 ;
      RECT  8532.5 169602.5 8597.5 169737.5 ;
      RECT  8722.5 169602.5 8787.5 169737.5 ;
      RECT  8722.5 169602.5 8787.5 169737.5 ;
      RECT  8532.5 169602.5 8597.5 169737.5 ;
      RECT  8532.5 168717.5 8597.5 168852.5 ;
      RECT  8722.5 168717.5 8787.5 168852.5 ;
      RECT  8722.5 168717.5 8787.5 168852.5 ;
      RECT  8532.5 168717.5 8597.5 168852.5 ;
      RECT  8892.5 169692.5 8957.5 169827.5 ;
      RECT  8892.5 168717.5 8957.5 168852.5 ;
      RECT  8590.0 169160.0 8655.0 169295.0 ;
      RECT  8590.0 169160.0 8655.0 169295.0 ;
      RECT  8755.0 169195.0 8820.0 169260.0 ;
      RECT  8465.0 169912.5 9025.0 169977.5 ;
      RECT  8465.0 168567.5 9025.0 168632.5 ;
      RECT  8892.5 170130.0 8957.5 169945.0 ;
      RECT  8892.5 171290.0 8957.5 171105.0 ;
      RECT  8532.5 171172.5 8597.5 171322.5 ;
      RECT  8532.5 170287.5 8597.5 169912.5 ;
      RECT  8722.5 171172.5 8787.5 170287.5 ;
      RECT  8532.5 170287.5 8597.5 170152.5 ;
      RECT  8722.5 170287.5 8787.5 170152.5 ;
      RECT  8722.5 170287.5 8787.5 170152.5 ;
      RECT  8532.5 170287.5 8597.5 170152.5 ;
      RECT  8532.5 171172.5 8597.5 171037.5 ;
      RECT  8722.5 171172.5 8787.5 171037.5 ;
      RECT  8722.5 171172.5 8787.5 171037.5 ;
      RECT  8532.5 171172.5 8597.5 171037.5 ;
      RECT  8892.5 170197.5 8957.5 170062.5 ;
      RECT  8892.5 171172.5 8957.5 171037.5 ;
      RECT  8590.0 170730.0 8655.0 170595.0 ;
      RECT  8590.0 170730.0 8655.0 170595.0 ;
      RECT  8755.0 170695.0 8820.0 170630.0 ;
      RECT  8465.0 169977.5 9025.0 169912.5 ;
      RECT  8465.0 171322.5 9025.0 171257.5 ;
      RECT  8892.5 172450.0 8957.5 172635.0 ;
      RECT  8892.5 171290.0 8957.5 171475.0 ;
      RECT  8532.5 171407.5 8597.5 171257.5 ;
      RECT  8532.5 172292.5 8597.5 172667.5 ;
      RECT  8722.5 171407.5 8787.5 172292.5 ;
      RECT  8532.5 172292.5 8597.5 172427.5 ;
      RECT  8722.5 172292.5 8787.5 172427.5 ;
      RECT  8722.5 172292.5 8787.5 172427.5 ;
      RECT  8532.5 172292.5 8597.5 172427.5 ;
      RECT  8532.5 171407.5 8597.5 171542.5 ;
      RECT  8722.5 171407.5 8787.5 171542.5 ;
      RECT  8722.5 171407.5 8787.5 171542.5 ;
      RECT  8532.5 171407.5 8597.5 171542.5 ;
      RECT  8892.5 172382.5 8957.5 172517.5 ;
      RECT  8892.5 171407.5 8957.5 171542.5 ;
      RECT  8590.0 171850.0 8655.0 171985.0 ;
      RECT  8590.0 171850.0 8655.0 171985.0 ;
      RECT  8755.0 171885.0 8820.0 171950.0 ;
      RECT  8465.0 172602.5 9025.0 172667.5 ;
      RECT  8465.0 171257.5 9025.0 171322.5 ;
      RECT  8892.5 172820.0 8957.5 172635.0 ;
      RECT  8892.5 173980.0 8957.5 173795.0 ;
      RECT  8532.5 173862.5 8597.5 174012.5 ;
      RECT  8532.5 172977.5 8597.5 172602.5 ;
      RECT  8722.5 173862.5 8787.5 172977.5 ;
      RECT  8532.5 172977.5 8597.5 172842.5 ;
      RECT  8722.5 172977.5 8787.5 172842.5 ;
      RECT  8722.5 172977.5 8787.5 172842.5 ;
      RECT  8532.5 172977.5 8597.5 172842.5 ;
      RECT  8532.5 173862.5 8597.5 173727.5 ;
      RECT  8722.5 173862.5 8787.5 173727.5 ;
      RECT  8722.5 173862.5 8787.5 173727.5 ;
      RECT  8532.5 173862.5 8597.5 173727.5 ;
      RECT  8892.5 172887.5 8957.5 172752.5 ;
      RECT  8892.5 173862.5 8957.5 173727.5 ;
      RECT  8590.0 173420.0 8655.0 173285.0 ;
      RECT  8590.0 173420.0 8655.0 173285.0 ;
      RECT  8755.0 173385.0 8820.0 173320.0 ;
      RECT  8465.0 172667.5 9025.0 172602.5 ;
      RECT  8465.0 174012.5 9025.0 173947.5 ;
      RECT  8892.5 175140.0 8957.5 175325.0 ;
      RECT  8892.5 173980.0 8957.5 174165.0 ;
      RECT  8532.5 174097.5 8597.5 173947.5 ;
      RECT  8532.5 174982.5 8597.5 175357.5 ;
      RECT  8722.5 174097.5 8787.5 174982.5 ;
      RECT  8532.5 174982.5 8597.5 175117.5 ;
      RECT  8722.5 174982.5 8787.5 175117.5 ;
      RECT  8722.5 174982.5 8787.5 175117.5 ;
      RECT  8532.5 174982.5 8597.5 175117.5 ;
      RECT  8532.5 174097.5 8597.5 174232.5 ;
      RECT  8722.5 174097.5 8787.5 174232.5 ;
      RECT  8722.5 174097.5 8787.5 174232.5 ;
      RECT  8532.5 174097.5 8597.5 174232.5 ;
      RECT  8892.5 175072.5 8957.5 175207.5 ;
      RECT  8892.5 174097.5 8957.5 174232.5 ;
      RECT  8590.0 174540.0 8655.0 174675.0 ;
      RECT  8590.0 174540.0 8655.0 174675.0 ;
      RECT  8755.0 174575.0 8820.0 174640.0 ;
      RECT  8465.0 175292.5 9025.0 175357.5 ;
      RECT  8465.0 173947.5 9025.0 174012.5 ;
      RECT  8892.5 175510.0 8957.5 175325.0 ;
      RECT  8892.5 176670.0 8957.5 176485.0 ;
      RECT  8532.5 176552.5 8597.5 176702.5 ;
      RECT  8532.5 175667.5 8597.5 175292.5 ;
      RECT  8722.5 176552.5 8787.5 175667.5 ;
      RECT  8532.5 175667.5 8597.5 175532.5 ;
      RECT  8722.5 175667.5 8787.5 175532.5 ;
      RECT  8722.5 175667.5 8787.5 175532.5 ;
      RECT  8532.5 175667.5 8597.5 175532.5 ;
      RECT  8532.5 176552.5 8597.5 176417.5 ;
      RECT  8722.5 176552.5 8787.5 176417.5 ;
      RECT  8722.5 176552.5 8787.5 176417.5 ;
      RECT  8532.5 176552.5 8597.5 176417.5 ;
      RECT  8892.5 175577.5 8957.5 175442.5 ;
      RECT  8892.5 176552.5 8957.5 176417.5 ;
      RECT  8590.0 176110.0 8655.0 175975.0 ;
      RECT  8590.0 176110.0 8655.0 175975.0 ;
      RECT  8755.0 176075.0 8820.0 176010.0 ;
      RECT  8465.0 175357.5 9025.0 175292.5 ;
      RECT  8465.0 176702.5 9025.0 176637.5 ;
      RECT  8892.5 177830.0 8957.5 178015.0 ;
      RECT  8892.5 176670.0 8957.5 176855.0 ;
      RECT  8532.5 176787.5 8597.5 176637.5 ;
      RECT  8532.5 177672.5 8597.5 178047.5 ;
      RECT  8722.5 176787.5 8787.5 177672.5 ;
      RECT  8532.5 177672.5 8597.5 177807.5 ;
      RECT  8722.5 177672.5 8787.5 177807.5 ;
      RECT  8722.5 177672.5 8787.5 177807.5 ;
      RECT  8532.5 177672.5 8597.5 177807.5 ;
      RECT  8532.5 176787.5 8597.5 176922.5 ;
      RECT  8722.5 176787.5 8787.5 176922.5 ;
      RECT  8722.5 176787.5 8787.5 176922.5 ;
      RECT  8532.5 176787.5 8597.5 176922.5 ;
      RECT  8892.5 177762.5 8957.5 177897.5 ;
      RECT  8892.5 176787.5 8957.5 176922.5 ;
      RECT  8590.0 177230.0 8655.0 177365.0 ;
      RECT  8590.0 177230.0 8655.0 177365.0 ;
      RECT  8755.0 177265.0 8820.0 177330.0 ;
      RECT  8465.0 177982.5 9025.0 178047.5 ;
      RECT  8465.0 176637.5 9025.0 176702.5 ;
      RECT  8892.5 178200.0 8957.5 178015.0 ;
      RECT  8892.5 179360.0 8957.5 179175.0 ;
      RECT  8532.5 179242.5 8597.5 179392.5 ;
      RECT  8532.5 178357.5 8597.5 177982.5 ;
      RECT  8722.5 179242.5 8787.5 178357.5 ;
      RECT  8532.5 178357.5 8597.5 178222.5 ;
      RECT  8722.5 178357.5 8787.5 178222.5 ;
      RECT  8722.5 178357.5 8787.5 178222.5 ;
      RECT  8532.5 178357.5 8597.5 178222.5 ;
      RECT  8532.5 179242.5 8597.5 179107.5 ;
      RECT  8722.5 179242.5 8787.5 179107.5 ;
      RECT  8722.5 179242.5 8787.5 179107.5 ;
      RECT  8532.5 179242.5 8597.5 179107.5 ;
      RECT  8892.5 178267.5 8957.5 178132.5 ;
      RECT  8892.5 179242.5 8957.5 179107.5 ;
      RECT  8590.0 178800.0 8655.0 178665.0 ;
      RECT  8590.0 178800.0 8655.0 178665.0 ;
      RECT  8755.0 178765.0 8820.0 178700.0 ;
      RECT  8465.0 178047.5 9025.0 177982.5 ;
      RECT  8465.0 179392.5 9025.0 179327.5 ;
      RECT  8892.5 180520.0 8957.5 180705.0 ;
      RECT  8892.5 179360.0 8957.5 179545.0 ;
      RECT  8532.5 179477.5 8597.5 179327.5 ;
      RECT  8532.5 180362.5 8597.5 180737.5 ;
      RECT  8722.5 179477.5 8787.5 180362.5 ;
      RECT  8532.5 180362.5 8597.5 180497.5 ;
      RECT  8722.5 180362.5 8787.5 180497.5 ;
      RECT  8722.5 180362.5 8787.5 180497.5 ;
      RECT  8532.5 180362.5 8597.5 180497.5 ;
      RECT  8532.5 179477.5 8597.5 179612.5 ;
      RECT  8722.5 179477.5 8787.5 179612.5 ;
      RECT  8722.5 179477.5 8787.5 179612.5 ;
      RECT  8532.5 179477.5 8597.5 179612.5 ;
      RECT  8892.5 180452.5 8957.5 180587.5 ;
      RECT  8892.5 179477.5 8957.5 179612.5 ;
      RECT  8590.0 179920.0 8655.0 180055.0 ;
      RECT  8590.0 179920.0 8655.0 180055.0 ;
      RECT  8755.0 179955.0 8820.0 180020.0 ;
      RECT  8465.0 180672.5 9025.0 180737.5 ;
      RECT  8465.0 179327.5 9025.0 179392.5 ;
      RECT  8892.5 180890.0 8957.5 180705.0 ;
      RECT  8892.5 182050.0 8957.5 181865.0 ;
      RECT  8532.5 181932.5 8597.5 182082.5 ;
      RECT  8532.5 181047.5 8597.5 180672.5 ;
      RECT  8722.5 181932.5 8787.5 181047.5 ;
      RECT  8532.5 181047.5 8597.5 180912.5 ;
      RECT  8722.5 181047.5 8787.5 180912.5 ;
      RECT  8722.5 181047.5 8787.5 180912.5 ;
      RECT  8532.5 181047.5 8597.5 180912.5 ;
      RECT  8532.5 181932.5 8597.5 181797.5 ;
      RECT  8722.5 181932.5 8787.5 181797.5 ;
      RECT  8722.5 181932.5 8787.5 181797.5 ;
      RECT  8532.5 181932.5 8597.5 181797.5 ;
      RECT  8892.5 180957.5 8957.5 180822.5 ;
      RECT  8892.5 181932.5 8957.5 181797.5 ;
      RECT  8590.0 181490.0 8655.0 181355.0 ;
      RECT  8590.0 181490.0 8655.0 181355.0 ;
      RECT  8755.0 181455.0 8820.0 181390.0 ;
      RECT  8465.0 180737.5 9025.0 180672.5 ;
      RECT  8465.0 182082.5 9025.0 182017.5 ;
      RECT  8892.5 183210.0 8957.5 183395.0 ;
      RECT  8892.5 182050.0 8957.5 182235.0 ;
      RECT  8532.5 182167.5 8597.5 182017.5 ;
      RECT  8532.5 183052.5 8597.5 183427.5 ;
      RECT  8722.5 182167.5 8787.5 183052.5 ;
      RECT  8532.5 183052.5 8597.5 183187.5 ;
      RECT  8722.5 183052.5 8787.5 183187.5 ;
      RECT  8722.5 183052.5 8787.5 183187.5 ;
      RECT  8532.5 183052.5 8597.5 183187.5 ;
      RECT  8532.5 182167.5 8597.5 182302.5 ;
      RECT  8722.5 182167.5 8787.5 182302.5 ;
      RECT  8722.5 182167.5 8787.5 182302.5 ;
      RECT  8532.5 182167.5 8597.5 182302.5 ;
      RECT  8892.5 183142.5 8957.5 183277.5 ;
      RECT  8892.5 182167.5 8957.5 182302.5 ;
      RECT  8590.0 182610.0 8655.0 182745.0 ;
      RECT  8590.0 182610.0 8655.0 182745.0 ;
      RECT  8755.0 182645.0 8820.0 182710.0 ;
      RECT  8465.0 183362.5 9025.0 183427.5 ;
      RECT  8465.0 182017.5 9025.0 182082.5 ;
      RECT  8892.5 183580.0 8957.5 183395.0 ;
      RECT  8892.5 184740.0 8957.5 184555.0 ;
      RECT  8532.5 184622.5 8597.5 184772.5 ;
      RECT  8532.5 183737.5 8597.5 183362.5 ;
      RECT  8722.5 184622.5 8787.5 183737.5 ;
      RECT  8532.5 183737.5 8597.5 183602.5 ;
      RECT  8722.5 183737.5 8787.5 183602.5 ;
      RECT  8722.5 183737.5 8787.5 183602.5 ;
      RECT  8532.5 183737.5 8597.5 183602.5 ;
      RECT  8532.5 184622.5 8597.5 184487.5 ;
      RECT  8722.5 184622.5 8787.5 184487.5 ;
      RECT  8722.5 184622.5 8787.5 184487.5 ;
      RECT  8532.5 184622.5 8597.5 184487.5 ;
      RECT  8892.5 183647.5 8957.5 183512.5 ;
      RECT  8892.5 184622.5 8957.5 184487.5 ;
      RECT  8590.0 184180.0 8655.0 184045.0 ;
      RECT  8590.0 184180.0 8655.0 184045.0 ;
      RECT  8755.0 184145.0 8820.0 184080.0 ;
      RECT  8465.0 183427.5 9025.0 183362.5 ;
      RECT  8465.0 184772.5 9025.0 184707.5 ;
      RECT  8892.5 185900.0 8957.5 186085.0 ;
      RECT  8892.5 184740.0 8957.5 184925.0 ;
      RECT  8532.5 184857.5 8597.5 184707.5 ;
      RECT  8532.5 185742.5 8597.5 186117.5 ;
      RECT  8722.5 184857.5 8787.5 185742.5 ;
      RECT  8532.5 185742.5 8597.5 185877.5 ;
      RECT  8722.5 185742.5 8787.5 185877.5 ;
      RECT  8722.5 185742.5 8787.5 185877.5 ;
      RECT  8532.5 185742.5 8597.5 185877.5 ;
      RECT  8532.5 184857.5 8597.5 184992.5 ;
      RECT  8722.5 184857.5 8787.5 184992.5 ;
      RECT  8722.5 184857.5 8787.5 184992.5 ;
      RECT  8532.5 184857.5 8597.5 184992.5 ;
      RECT  8892.5 185832.5 8957.5 185967.5 ;
      RECT  8892.5 184857.5 8957.5 184992.5 ;
      RECT  8590.0 185300.0 8655.0 185435.0 ;
      RECT  8590.0 185300.0 8655.0 185435.0 ;
      RECT  8755.0 185335.0 8820.0 185400.0 ;
      RECT  8465.0 186052.5 9025.0 186117.5 ;
      RECT  8465.0 184707.5 9025.0 184772.5 ;
      RECT  8892.5 186270.0 8957.5 186085.0 ;
      RECT  8892.5 187430.0 8957.5 187245.0 ;
      RECT  8532.5 187312.5 8597.5 187462.5 ;
      RECT  8532.5 186427.5 8597.5 186052.5 ;
      RECT  8722.5 187312.5 8787.5 186427.5 ;
      RECT  8532.5 186427.5 8597.5 186292.5 ;
      RECT  8722.5 186427.5 8787.5 186292.5 ;
      RECT  8722.5 186427.5 8787.5 186292.5 ;
      RECT  8532.5 186427.5 8597.5 186292.5 ;
      RECT  8532.5 187312.5 8597.5 187177.5 ;
      RECT  8722.5 187312.5 8787.5 187177.5 ;
      RECT  8722.5 187312.5 8787.5 187177.5 ;
      RECT  8532.5 187312.5 8597.5 187177.5 ;
      RECT  8892.5 186337.5 8957.5 186202.5 ;
      RECT  8892.5 187312.5 8957.5 187177.5 ;
      RECT  8590.0 186870.0 8655.0 186735.0 ;
      RECT  8590.0 186870.0 8655.0 186735.0 ;
      RECT  8755.0 186835.0 8820.0 186770.0 ;
      RECT  8465.0 186117.5 9025.0 186052.5 ;
      RECT  8465.0 187462.5 9025.0 187397.5 ;
      RECT  8892.5 188590.0 8957.5 188775.0 ;
      RECT  8892.5 187430.0 8957.5 187615.0 ;
      RECT  8532.5 187547.5 8597.5 187397.5 ;
      RECT  8532.5 188432.5 8597.5 188807.5 ;
      RECT  8722.5 187547.5 8787.5 188432.5 ;
      RECT  8532.5 188432.5 8597.5 188567.5 ;
      RECT  8722.5 188432.5 8787.5 188567.5 ;
      RECT  8722.5 188432.5 8787.5 188567.5 ;
      RECT  8532.5 188432.5 8597.5 188567.5 ;
      RECT  8532.5 187547.5 8597.5 187682.5 ;
      RECT  8722.5 187547.5 8787.5 187682.5 ;
      RECT  8722.5 187547.5 8787.5 187682.5 ;
      RECT  8532.5 187547.5 8597.5 187682.5 ;
      RECT  8892.5 188522.5 8957.5 188657.5 ;
      RECT  8892.5 187547.5 8957.5 187682.5 ;
      RECT  8590.0 187990.0 8655.0 188125.0 ;
      RECT  8590.0 187990.0 8655.0 188125.0 ;
      RECT  8755.0 188025.0 8820.0 188090.0 ;
      RECT  8465.0 188742.5 9025.0 188807.5 ;
      RECT  8465.0 187397.5 9025.0 187462.5 ;
      RECT  8892.5 188960.0 8957.5 188775.0 ;
      RECT  8892.5 190120.0 8957.5 189935.0 ;
      RECT  8532.5 190002.5 8597.5 190152.5 ;
      RECT  8532.5 189117.5 8597.5 188742.5 ;
      RECT  8722.5 190002.5 8787.5 189117.5 ;
      RECT  8532.5 189117.5 8597.5 188982.5 ;
      RECT  8722.5 189117.5 8787.5 188982.5 ;
      RECT  8722.5 189117.5 8787.5 188982.5 ;
      RECT  8532.5 189117.5 8597.5 188982.5 ;
      RECT  8532.5 190002.5 8597.5 189867.5 ;
      RECT  8722.5 190002.5 8787.5 189867.5 ;
      RECT  8722.5 190002.5 8787.5 189867.5 ;
      RECT  8532.5 190002.5 8597.5 189867.5 ;
      RECT  8892.5 189027.5 8957.5 188892.5 ;
      RECT  8892.5 190002.5 8957.5 189867.5 ;
      RECT  8590.0 189560.0 8655.0 189425.0 ;
      RECT  8590.0 189560.0 8655.0 189425.0 ;
      RECT  8755.0 189525.0 8820.0 189460.0 ;
      RECT  8465.0 188807.5 9025.0 188742.5 ;
      RECT  8465.0 190152.5 9025.0 190087.5 ;
      RECT  8892.5 191280.0 8957.5 191465.0 ;
      RECT  8892.5 190120.0 8957.5 190305.0 ;
      RECT  8532.5 190237.5 8597.5 190087.5 ;
      RECT  8532.5 191122.5 8597.5 191497.5 ;
      RECT  8722.5 190237.5 8787.5 191122.5 ;
      RECT  8532.5 191122.5 8597.5 191257.5 ;
      RECT  8722.5 191122.5 8787.5 191257.5 ;
      RECT  8722.5 191122.5 8787.5 191257.5 ;
      RECT  8532.5 191122.5 8597.5 191257.5 ;
      RECT  8532.5 190237.5 8597.5 190372.5 ;
      RECT  8722.5 190237.5 8787.5 190372.5 ;
      RECT  8722.5 190237.5 8787.5 190372.5 ;
      RECT  8532.5 190237.5 8597.5 190372.5 ;
      RECT  8892.5 191212.5 8957.5 191347.5 ;
      RECT  8892.5 190237.5 8957.5 190372.5 ;
      RECT  8590.0 190680.0 8655.0 190815.0 ;
      RECT  8590.0 190680.0 8655.0 190815.0 ;
      RECT  8755.0 190715.0 8820.0 190780.0 ;
      RECT  8465.0 191432.5 9025.0 191497.5 ;
      RECT  8465.0 190087.5 9025.0 190152.5 ;
      RECT  8892.5 191650.0 8957.5 191465.0 ;
      RECT  8892.5 192810.0 8957.5 192625.0 ;
      RECT  8532.5 192692.5 8597.5 192842.5 ;
      RECT  8532.5 191807.5 8597.5 191432.5 ;
      RECT  8722.5 192692.5 8787.5 191807.5 ;
      RECT  8532.5 191807.5 8597.5 191672.5 ;
      RECT  8722.5 191807.5 8787.5 191672.5 ;
      RECT  8722.5 191807.5 8787.5 191672.5 ;
      RECT  8532.5 191807.5 8597.5 191672.5 ;
      RECT  8532.5 192692.5 8597.5 192557.5 ;
      RECT  8722.5 192692.5 8787.5 192557.5 ;
      RECT  8722.5 192692.5 8787.5 192557.5 ;
      RECT  8532.5 192692.5 8597.5 192557.5 ;
      RECT  8892.5 191717.5 8957.5 191582.5 ;
      RECT  8892.5 192692.5 8957.5 192557.5 ;
      RECT  8590.0 192250.0 8655.0 192115.0 ;
      RECT  8590.0 192250.0 8655.0 192115.0 ;
      RECT  8755.0 192215.0 8820.0 192150.0 ;
      RECT  8465.0 191497.5 9025.0 191432.5 ;
      RECT  8465.0 192842.5 9025.0 192777.5 ;
      RECT  8892.5 193970.0 8957.5 194155.0 ;
      RECT  8892.5 192810.0 8957.5 192995.0 ;
      RECT  8532.5 192927.5 8597.5 192777.5 ;
      RECT  8532.5 193812.5 8597.5 194187.5 ;
      RECT  8722.5 192927.5 8787.5 193812.5 ;
      RECT  8532.5 193812.5 8597.5 193947.5 ;
      RECT  8722.5 193812.5 8787.5 193947.5 ;
      RECT  8722.5 193812.5 8787.5 193947.5 ;
      RECT  8532.5 193812.5 8597.5 193947.5 ;
      RECT  8532.5 192927.5 8597.5 193062.5 ;
      RECT  8722.5 192927.5 8787.5 193062.5 ;
      RECT  8722.5 192927.5 8787.5 193062.5 ;
      RECT  8532.5 192927.5 8597.5 193062.5 ;
      RECT  8892.5 193902.5 8957.5 194037.5 ;
      RECT  8892.5 192927.5 8957.5 193062.5 ;
      RECT  8590.0 193370.0 8655.0 193505.0 ;
      RECT  8590.0 193370.0 8655.0 193505.0 ;
      RECT  8755.0 193405.0 8820.0 193470.0 ;
      RECT  8465.0 194122.5 9025.0 194187.5 ;
      RECT  8465.0 192777.5 9025.0 192842.5 ;
      RECT  8892.5 194340.0 8957.5 194155.0 ;
      RECT  8892.5 195500.0 8957.5 195315.0 ;
      RECT  8532.5 195382.5 8597.5 195532.5 ;
      RECT  8532.5 194497.5 8597.5 194122.5 ;
      RECT  8722.5 195382.5 8787.5 194497.5 ;
      RECT  8532.5 194497.5 8597.5 194362.5 ;
      RECT  8722.5 194497.5 8787.5 194362.5 ;
      RECT  8722.5 194497.5 8787.5 194362.5 ;
      RECT  8532.5 194497.5 8597.5 194362.5 ;
      RECT  8532.5 195382.5 8597.5 195247.5 ;
      RECT  8722.5 195382.5 8787.5 195247.5 ;
      RECT  8722.5 195382.5 8787.5 195247.5 ;
      RECT  8532.5 195382.5 8597.5 195247.5 ;
      RECT  8892.5 194407.5 8957.5 194272.5 ;
      RECT  8892.5 195382.5 8957.5 195247.5 ;
      RECT  8590.0 194940.0 8655.0 194805.0 ;
      RECT  8590.0 194940.0 8655.0 194805.0 ;
      RECT  8755.0 194905.0 8820.0 194840.0 ;
      RECT  8465.0 194187.5 9025.0 194122.5 ;
      RECT  8465.0 195532.5 9025.0 195467.5 ;
      RECT  8892.5 196660.0 8957.5 196845.0 ;
      RECT  8892.5 195500.0 8957.5 195685.0 ;
      RECT  8532.5 195617.5 8597.5 195467.5 ;
      RECT  8532.5 196502.5 8597.5 196877.5 ;
      RECT  8722.5 195617.5 8787.5 196502.5 ;
      RECT  8532.5 196502.5 8597.5 196637.5 ;
      RECT  8722.5 196502.5 8787.5 196637.5 ;
      RECT  8722.5 196502.5 8787.5 196637.5 ;
      RECT  8532.5 196502.5 8597.5 196637.5 ;
      RECT  8532.5 195617.5 8597.5 195752.5 ;
      RECT  8722.5 195617.5 8787.5 195752.5 ;
      RECT  8722.5 195617.5 8787.5 195752.5 ;
      RECT  8532.5 195617.5 8597.5 195752.5 ;
      RECT  8892.5 196592.5 8957.5 196727.5 ;
      RECT  8892.5 195617.5 8957.5 195752.5 ;
      RECT  8590.0 196060.0 8655.0 196195.0 ;
      RECT  8590.0 196060.0 8655.0 196195.0 ;
      RECT  8755.0 196095.0 8820.0 196160.0 ;
      RECT  8465.0 196812.5 9025.0 196877.5 ;
      RECT  8465.0 195467.5 9025.0 195532.5 ;
      RECT  8892.5 197030.0 8957.5 196845.0 ;
      RECT  8892.5 198190.0 8957.5 198005.0 ;
      RECT  8532.5 198072.5 8597.5 198222.5 ;
      RECT  8532.5 197187.5 8597.5 196812.5 ;
      RECT  8722.5 198072.5 8787.5 197187.5 ;
      RECT  8532.5 197187.5 8597.5 197052.5 ;
      RECT  8722.5 197187.5 8787.5 197052.5 ;
      RECT  8722.5 197187.5 8787.5 197052.5 ;
      RECT  8532.5 197187.5 8597.5 197052.5 ;
      RECT  8532.5 198072.5 8597.5 197937.5 ;
      RECT  8722.5 198072.5 8787.5 197937.5 ;
      RECT  8722.5 198072.5 8787.5 197937.5 ;
      RECT  8532.5 198072.5 8597.5 197937.5 ;
      RECT  8892.5 197097.5 8957.5 196962.5 ;
      RECT  8892.5 198072.5 8957.5 197937.5 ;
      RECT  8590.0 197630.0 8655.0 197495.0 ;
      RECT  8590.0 197630.0 8655.0 197495.0 ;
      RECT  8755.0 197595.0 8820.0 197530.0 ;
      RECT  8465.0 196877.5 9025.0 196812.5 ;
      RECT  8465.0 198222.5 9025.0 198157.5 ;
      RECT  8892.5 199350.0 8957.5 199535.0 ;
      RECT  8892.5 198190.0 8957.5 198375.0 ;
      RECT  8532.5 198307.5 8597.5 198157.5 ;
      RECT  8532.5 199192.5 8597.5 199567.5 ;
      RECT  8722.5 198307.5 8787.5 199192.5 ;
      RECT  8532.5 199192.5 8597.5 199327.5 ;
      RECT  8722.5 199192.5 8787.5 199327.5 ;
      RECT  8722.5 199192.5 8787.5 199327.5 ;
      RECT  8532.5 199192.5 8597.5 199327.5 ;
      RECT  8532.5 198307.5 8597.5 198442.5 ;
      RECT  8722.5 198307.5 8787.5 198442.5 ;
      RECT  8722.5 198307.5 8787.5 198442.5 ;
      RECT  8532.5 198307.5 8597.5 198442.5 ;
      RECT  8892.5 199282.5 8957.5 199417.5 ;
      RECT  8892.5 198307.5 8957.5 198442.5 ;
      RECT  8590.0 198750.0 8655.0 198885.0 ;
      RECT  8590.0 198750.0 8655.0 198885.0 ;
      RECT  8755.0 198785.0 8820.0 198850.0 ;
      RECT  8465.0 199502.5 9025.0 199567.5 ;
      RECT  8465.0 198157.5 9025.0 198222.5 ;
      RECT  8892.5 199720.0 8957.5 199535.0 ;
      RECT  8892.5 200880.0 8957.5 200695.0 ;
      RECT  8532.5 200762.5 8597.5 200912.5 ;
      RECT  8532.5 199877.5 8597.5 199502.5 ;
      RECT  8722.5 200762.5 8787.5 199877.5 ;
      RECT  8532.5 199877.5 8597.5 199742.5 ;
      RECT  8722.5 199877.5 8787.5 199742.5 ;
      RECT  8722.5 199877.5 8787.5 199742.5 ;
      RECT  8532.5 199877.5 8597.5 199742.5 ;
      RECT  8532.5 200762.5 8597.5 200627.5 ;
      RECT  8722.5 200762.5 8787.5 200627.5 ;
      RECT  8722.5 200762.5 8787.5 200627.5 ;
      RECT  8532.5 200762.5 8597.5 200627.5 ;
      RECT  8892.5 199787.5 8957.5 199652.5 ;
      RECT  8892.5 200762.5 8957.5 200627.5 ;
      RECT  8590.0 200320.0 8655.0 200185.0 ;
      RECT  8590.0 200320.0 8655.0 200185.0 ;
      RECT  8755.0 200285.0 8820.0 200220.0 ;
      RECT  8465.0 199567.5 9025.0 199502.5 ;
      RECT  8465.0 200912.5 9025.0 200847.5 ;
      RECT  8892.5 202040.0 8957.5 202225.0 ;
      RECT  8892.5 200880.0 8957.5 201065.0 ;
      RECT  8532.5 200997.5 8597.5 200847.5 ;
      RECT  8532.5 201882.5 8597.5 202257.5 ;
      RECT  8722.5 200997.5 8787.5 201882.5 ;
      RECT  8532.5 201882.5 8597.5 202017.5 ;
      RECT  8722.5 201882.5 8787.5 202017.5 ;
      RECT  8722.5 201882.5 8787.5 202017.5 ;
      RECT  8532.5 201882.5 8597.5 202017.5 ;
      RECT  8532.5 200997.5 8597.5 201132.5 ;
      RECT  8722.5 200997.5 8787.5 201132.5 ;
      RECT  8722.5 200997.5 8787.5 201132.5 ;
      RECT  8532.5 200997.5 8597.5 201132.5 ;
      RECT  8892.5 201972.5 8957.5 202107.5 ;
      RECT  8892.5 200997.5 8957.5 201132.5 ;
      RECT  8590.0 201440.0 8655.0 201575.0 ;
      RECT  8590.0 201440.0 8655.0 201575.0 ;
      RECT  8755.0 201475.0 8820.0 201540.0 ;
      RECT  8465.0 202192.5 9025.0 202257.5 ;
      RECT  8465.0 200847.5 9025.0 200912.5 ;
      RECT  8892.5 202410.0 8957.5 202225.0 ;
      RECT  8892.5 203570.0 8957.5 203385.0 ;
      RECT  8532.5 203452.5 8597.5 203602.5 ;
      RECT  8532.5 202567.5 8597.5 202192.5 ;
      RECT  8722.5 203452.5 8787.5 202567.5 ;
      RECT  8532.5 202567.5 8597.5 202432.5 ;
      RECT  8722.5 202567.5 8787.5 202432.5 ;
      RECT  8722.5 202567.5 8787.5 202432.5 ;
      RECT  8532.5 202567.5 8597.5 202432.5 ;
      RECT  8532.5 203452.5 8597.5 203317.5 ;
      RECT  8722.5 203452.5 8787.5 203317.5 ;
      RECT  8722.5 203452.5 8787.5 203317.5 ;
      RECT  8532.5 203452.5 8597.5 203317.5 ;
      RECT  8892.5 202477.5 8957.5 202342.5 ;
      RECT  8892.5 203452.5 8957.5 203317.5 ;
      RECT  8590.0 203010.0 8655.0 202875.0 ;
      RECT  8590.0 203010.0 8655.0 202875.0 ;
      RECT  8755.0 202975.0 8820.0 202910.0 ;
      RECT  8465.0 202257.5 9025.0 202192.5 ;
      RECT  8465.0 203602.5 9025.0 203537.5 ;
      RECT  8892.5 204730.0 8957.5 204915.0 ;
      RECT  8892.5 203570.0 8957.5 203755.0 ;
      RECT  8532.5 203687.5 8597.5 203537.5 ;
      RECT  8532.5 204572.5 8597.5 204947.5 ;
      RECT  8722.5 203687.5 8787.5 204572.5 ;
      RECT  8532.5 204572.5 8597.5 204707.5 ;
      RECT  8722.5 204572.5 8787.5 204707.5 ;
      RECT  8722.5 204572.5 8787.5 204707.5 ;
      RECT  8532.5 204572.5 8597.5 204707.5 ;
      RECT  8532.5 203687.5 8597.5 203822.5 ;
      RECT  8722.5 203687.5 8787.5 203822.5 ;
      RECT  8722.5 203687.5 8787.5 203822.5 ;
      RECT  8532.5 203687.5 8597.5 203822.5 ;
      RECT  8892.5 204662.5 8957.5 204797.5 ;
      RECT  8892.5 203687.5 8957.5 203822.5 ;
      RECT  8590.0 204130.0 8655.0 204265.0 ;
      RECT  8590.0 204130.0 8655.0 204265.0 ;
      RECT  8755.0 204165.0 8820.0 204230.0 ;
      RECT  8465.0 204882.5 9025.0 204947.5 ;
      RECT  8465.0 203537.5 9025.0 203602.5 ;
      RECT  8892.5 205100.0 8957.5 204915.0 ;
      RECT  8892.5 206260.0 8957.5 206075.0 ;
      RECT  8532.5 206142.5 8597.5 206292.5 ;
      RECT  8532.5 205257.5 8597.5 204882.5 ;
      RECT  8722.5 206142.5 8787.5 205257.5 ;
      RECT  8532.5 205257.5 8597.5 205122.5 ;
      RECT  8722.5 205257.5 8787.5 205122.5 ;
      RECT  8722.5 205257.5 8787.5 205122.5 ;
      RECT  8532.5 205257.5 8597.5 205122.5 ;
      RECT  8532.5 206142.5 8597.5 206007.5 ;
      RECT  8722.5 206142.5 8787.5 206007.5 ;
      RECT  8722.5 206142.5 8787.5 206007.5 ;
      RECT  8532.5 206142.5 8597.5 206007.5 ;
      RECT  8892.5 205167.5 8957.5 205032.5 ;
      RECT  8892.5 206142.5 8957.5 206007.5 ;
      RECT  8590.0 205700.0 8655.0 205565.0 ;
      RECT  8590.0 205700.0 8655.0 205565.0 ;
      RECT  8755.0 205665.0 8820.0 205600.0 ;
      RECT  8465.0 204947.5 9025.0 204882.5 ;
      RECT  8465.0 206292.5 9025.0 206227.5 ;
      RECT  4757.5 13175.0 4622.5 13240.0 ;
      RECT  4932.5 14610.0 4797.5 14675.0 ;
      RECT  5107.5 15865.0 4972.5 15930.0 ;
      RECT  5282.5 17300.0 5147.5 17365.0 ;
      RECT  5457.5 18555.0 5322.5 18620.0 ;
      RECT  5632.5 19990.0 5497.5 20055.0 ;
      RECT  5807.5 21245.0 5672.5 21310.0 ;
      RECT  5982.5 22680.0 5847.5 22745.0 ;
      RECT  6157.5 23935.0 6022.5 24000.0 ;
      RECT  6332.5 25370.0 6197.5 25435.0 ;
      RECT  6507.5 26625.0 6372.5 26690.0 ;
      RECT  6682.5 28060.0 6547.5 28125.0 ;
      RECT  6857.5 29315.0 6722.5 29380.0 ;
      RECT  7032.5 30750.0 6897.5 30815.0 ;
      RECT  7207.5 32005.0 7072.5 32070.0 ;
      RECT  7382.5 33440.0 7247.5 33505.0 ;
      RECT  4757.5 34755.0 4622.5 34820.0 ;
      RECT  5457.5 34615.0 5322.5 34680.0 ;
      RECT  6157.5 34475.0 6022.5 34540.0 ;
      RECT  4757.5 36070.0 4622.5 36135.0 ;
      RECT  5457.5 36210.0 5322.5 36275.0 ;
      RECT  6332.5 36350.0 6197.5 36415.0 ;
      RECT  4757.5 37445.0 4622.5 37510.0 ;
      RECT  5457.5 37305.0 5322.5 37370.0 ;
      RECT  6507.5 37165.0 6372.5 37230.0 ;
      RECT  4757.5 38760.0 4622.5 38825.0 ;
      RECT  5457.5 38900.0 5322.5 38965.0 ;
      RECT  6682.5 39040.0 6547.5 39105.0 ;
      RECT  4757.5 40135.0 4622.5 40200.0 ;
      RECT  5457.5 39995.0 5322.5 40060.0 ;
      RECT  6857.5 39855.0 6722.5 39920.0 ;
      RECT  4757.5 41450.0 4622.5 41515.0 ;
      RECT  5457.5 41590.0 5322.5 41655.0 ;
      RECT  7032.5 41730.0 6897.5 41795.0 ;
      RECT  4757.5 42825.0 4622.5 42890.0 ;
      RECT  5457.5 42685.0 5322.5 42750.0 ;
      RECT  7207.5 42545.0 7072.5 42610.0 ;
      RECT  4757.5 44140.0 4622.5 44205.0 ;
      RECT  5457.5 44280.0 5322.5 44345.0 ;
      RECT  7382.5 44420.0 7247.5 44485.0 ;
      RECT  4757.5 45515.0 4622.5 45580.0 ;
      RECT  5632.5 45375.0 5497.5 45440.0 ;
      RECT  6157.5 45235.0 6022.5 45300.0 ;
      RECT  4757.5 46830.0 4622.5 46895.0 ;
      RECT  5632.5 46970.0 5497.5 47035.0 ;
      RECT  6332.5 47110.0 6197.5 47175.0 ;
      RECT  4757.5 48205.0 4622.5 48270.0 ;
      RECT  5632.5 48065.0 5497.5 48130.0 ;
      RECT  6507.5 47925.0 6372.5 47990.0 ;
      RECT  4757.5 49520.0 4622.5 49585.0 ;
      RECT  5632.5 49660.0 5497.5 49725.0 ;
      RECT  6682.5 49800.0 6547.5 49865.0 ;
      RECT  4757.5 50895.0 4622.5 50960.0 ;
      RECT  5632.5 50755.0 5497.5 50820.0 ;
      RECT  6857.5 50615.0 6722.5 50680.0 ;
      RECT  4757.5 52210.0 4622.5 52275.0 ;
      RECT  5632.5 52350.0 5497.5 52415.0 ;
      RECT  7032.5 52490.0 6897.5 52555.0 ;
      RECT  4757.5 53585.0 4622.5 53650.0 ;
      RECT  5632.5 53445.0 5497.5 53510.0 ;
      RECT  7207.5 53305.0 7072.5 53370.0 ;
      RECT  4757.5 54900.0 4622.5 54965.0 ;
      RECT  5632.5 55040.0 5497.5 55105.0 ;
      RECT  7382.5 55180.0 7247.5 55245.0 ;
      RECT  4757.5 56275.0 4622.5 56340.0 ;
      RECT  5807.5 56135.0 5672.5 56200.0 ;
      RECT  6157.5 55995.0 6022.5 56060.0 ;
      RECT  4757.5 57590.0 4622.5 57655.0 ;
      RECT  5807.5 57730.0 5672.5 57795.0 ;
      RECT  6332.5 57870.0 6197.5 57935.0 ;
      RECT  4757.5 58965.0 4622.5 59030.0 ;
      RECT  5807.5 58825.0 5672.5 58890.0 ;
      RECT  6507.5 58685.0 6372.5 58750.0 ;
      RECT  4757.5 60280.0 4622.5 60345.0 ;
      RECT  5807.5 60420.0 5672.5 60485.0 ;
      RECT  6682.5 60560.0 6547.5 60625.0 ;
      RECT  4757.5 61655.0 4622.5 61720.0 ;
      RECT  5807.5 61515.0 5672.5 61580.0 ;
      RECT  6857.5 61375.0 6722.5 61440.0 ;
      RECT  4757.5 62970.0 4622.5 63035.0 ;
      RECT  5807.5 63110.0 5672.5 63175.0 ;
      RECT  7032.5 63250.0 6897.5 63315.0 ;
      RECT  4757.5 64345.0 4622.5 64410.0 ;
      RECT  5807.5 64205.0 5672.5 64270.0 ;
      RECT  7207.5 64065.0 7072.5 64130.0 ;
      RECT  4757.5 65660.0 4622.5 65725.0 ;
      RECT  5807.5 65800.0 5672.5 65865.0 ;
      RECT  7382.5 65940.0 7247.5 66005.0 ;
      RECT  4757.5 67035.0 4622.5 67100.0 ;
      RECT  5982.5 66895.0 5847.5 66960.0 ;
      RECT  6157.5 66755.0 6022.5 66820.0 ;
      RECT  4757.5 68350.0 4622.5 68415.0 ;
      RECT  5982.5 68490.0 5847.5 68555.0 ;
      RECT  6332.5 68630.0 6197.5 68695.0 ;
      RECT  4757.5 69725.0 4622.5 69790.0 ;
      RECT  5982.5 69585.0 5847.5 69650.0 ;
      RECT  6507.5 69445.0 6372.5 69510.0 ;
      RECT  4757.5 71040.0 4622.5 71105.0 ;
      RECT  5982.5 71180.0 5847.5 71245.0 ;
      RECT  6682.5 71320.0 6547.5 71385.0 ;
      RECT  4757.5 72415.0 4622.5 72480.0 ;
      RECT  5982.5 72275.0 5847.5 72340.0 ;
      RECT  6857.5 72135.0 6722.5 72200.0 ;
      RECT  4757.5 73730.0 4622.5 73795.0 ;
      RECT  5982.5 73870.0 5847.5 73935.0 ;
      RECT  7032.5 74010.0 6897.5 74075.0 ;
      RECT  4757.5 75105.0 4622.5 75170.0 ;
      RECT  5982.5 74965.0 5847.5 75030.0 ;
      RECT  7207.5 74825.0 7072.5 74890.0 ;
      RECT  4757.5 76420.0 4622.5 76485.0 ;
      RECT  5982.5 76560.0 5847.5 76625.0 ;
      RECT  7382.5 76700.0 7247.5 76765.0 ;
      RECT  4932.5 77795.0 4797.5 77860.0 ;
      RECT  5457.5 77655.0 5322.5 77720.0 ;
      RECT  6157.5 77515.0 6022.5 77580.0 ;
      RECT  4932.5 79110.0 4797.5 79175.0 ;
      RECT  5457.5 79250.0 5322.5 79315.0 ;
      RECT  6332.5 79390.0 6197.5 79455.0 ;
      RECT  4932.5 80485.0 4797.5 80550.0 ;
      RECT  5457.5 80345.0 5322.5 80410.0 ;
      RECT  6507.5 80205.0 6372.5 80270.0 ;
      RECT  4932.5 81800.0 4797.5 81865.0 ;
      RECT  5457.5 81940.0 5322.5 82005.0 ;
      RECT  6682.5 82080.0 6547.5 82145.0 ;
      RECT  4932.5 83175.0 4797.5 83240.0 ;
      RECT  5457.5 83035.0 5322.5 83100.0 ;
      RECT  6857.5 82895.0 6722.5 82960.0 ;
      RECT  4932.5 84490.0 4797.5 84555.0 ;
      RECT  5457.5 84630.0 5322.5 84695.0 ;
      RECT  7032.5 84770.0 6897.5 84835.0 ;
      RECT  4932.5 85865.0 4797.5 85930.0 ;
      RECT  5457.5 85725.0 5322.5 85790.0 ;
      RECT  7207.5 85585.0 7072.5 85650.0 ;
      RECT  4932.5 87180.0 4797.5 87245.0 ;
      RECT  5457.5 87320.0 5322.5 87385.0 ;
      RECT  7382.5 87460.0 7247.5 87525.0 ;
      RECT  4932.5 88555.0 4797.5 88620.0 ;
      RECT  5632.5 88415.0 5497.5 88480.0 ;
      RECT  6157.5 88275.0 6022.5 88340.0 ;
      RECT  4932.5 89870.0 4797.5 89935.0 ;
      RECT  5632.5 90010.0 5497.5 90075.0 ;
      RECT  6332.5 90150.0 6197.5 90215.0 ;
      RECT  4932.5 91245.0 4797.5 91310.0 ;
      RECT  5632.5 91105.0 5497.5 91170.0 ;
      RECT  6507.5 90965.0 6372.5 91030.0 ;
      RECT  4932.5 92560.0 4797.5 92625.0 ;
      RECT  5632.5 92700.0 5497.5 92765.0 ;
      RECT  6682.5 92840.0 6547.5 92905.0 ;
      RECT  4932.5 93935.0 4797.5 94000.0 ;
      RECT  5632.5 93795.0 5497.5 93860.0 ;
      RECT  6857.5 93655.0 6722.5 93720.0 ;
      RECT  4932.5 95250.0 4797.5 95315.0 ;
      RECT  5632.5 95390.0 5497.5 95455.0 ;
      RECT  7032.5 95530.0 6897.5 95595.0 ;
      RECT  4932.5 96625.0 4797.5 96690.0 ;
      RECT  5632.5 96485.0 5497.5 96550.0 ;
      RECT  7207.5 96345.0 7072.5 96410.0 ;
      RECT  4932.5 97940.0 4797.5 98005.0 ;
      RECT  5632.5 98080.0 5497.5 98145.0 ;
      RECT  7382.5 98220.0 7247.5 98285.0 ;
      RECT  4932.5 99315.0 4797.5 99380.0 ;
      RECT  5807.5 99175.0 5672.5 99240.0 ;
      RECT  6157.5 99035.0 6022.5 99100.0 ;
      RECT  4932.5 100630.0 4797.5 100695.0 ;
      RECT  5807.5 100770.0 5672.5 100835.0 ;
      RECT  6332.5 100910.0 6197.5 100975.0 ;
      RECT  4932.5 102005.0 4797.5 102070.0 ;
      RECT  5807.5 101865.0 5672.5 101930.0 ;
      RECT  6507.5 101725.0 6372.5 101790.0 ;
      RECT  4932.5 103320.0 4797.5 103385.0 ;
      RECT  5807.5 103460.0 5672.5 103525.0 ;
      RECT  6682.5 103600.0 6547.5 103665.0 ;
      RECT  4932.5 104695.0 4797.5 104760.0 ;
      RECT  5807.5 104555.0 5672.5 104620.0 ;
      RECT  6857.5 104415.0 6722.5 104480.0 ;
      RECT  4932.5 106010.0 4797.5 106075.0 ;
      RECT  5807.5 106150.0 5672.5 106215.0 ;
      RECT  7032.5 106290.0 6897.5 106355.0 ;
      RECT  4932.5 107385.0 4797.5 107450.0 ;
      RECT  5807.5 107245.0 5672.5 107310.0 ;
      RECT  7207.5 107105.0 7072.5 107170.0 ;
      RECT  4932.5 108700.0 4797.5 108765.0 ;
      RECT  5807.5 108840.0 5672.5 108905.0 ;
      RECT  7382.5 108980.0 7247.5 109045.0 ;
      RECT  4932.5 110075.0 4797.5 110140.0 ;
      RECT  5982.5 109935.0 5847.5 110000.0 ;
      RECT  6157.5 109795.0 6022.5 109860.0 ;
      RECT  4932.5 111390.0 4797.5 111455.0 ;
      RECT  5982.5 111530.0 5847.5 111595.0 ;
      RECT  6332.5 111670.0 6197.5 111735.0 ;
      RECT  4932.5 112765.0 4797.5 112830.0 ;
      RECT  5982.5 112625.0 5847.5 112690.0 ;
      RECT  6507.5 112485.0 6372.5 112550.0 ;
      RECT  4932.5 114080.0 4797.5 114145.0 ;
      RECT  5982.5 114220.0 5847.5 114285.0 ;
      RECT  6682.5 114360.0 6547.5 114425.0 ;
      RECT  4932.5 115455.0 4797.5 115520.0 ;
      RECT  5982.5 115315.0 5847.5 115380.0 ;
      RECT  6857.5 115175.0 6722.5 115240.0 ;
      RECT  4932.5 116770.0 4797.5 116835.0 ;
      RECT  5982.5 116910.0 5847.5 116975.0 ;
      RECT  7032.5 117050.0 6897.5 117115.0 ;
      RECT  4932.5 118145.0 4797.5 118210.0 ;
      RECT  5982.5 118005.0 5847.5 118070.0 ;
      RECT  7207.5 117865.0 7072.5 117930.0 ;
      RECT  4932.5 119460.0 4797.5 119525.0 ;
      RECT  5982.5 119600.0 5847.5 119665.0 ;
      RECT  7382.5 119740.0 7247.5 119805.0 ;
      RECT  5107.5 120835.0 4972.5 120900.0 ;
      RECT  5457.5 120695.0 5322.5 120760.0 ;
      RECT  6157.5 120555.0 6022.5 120620.0 ;
      RECT  5107.5 122150.0 4972.5 122215.0 ;
      RECT  5457.5 122290.0 5322.5 122355.0 ;
      RECT  6332.5 122430.0 6197.5 122495.0 ;
      RECT  5107.5 123525.0 4972.5 123590.0 ;
      RECT  5457.5 123385.0 5322.5 123450.0 ;
      RECT  6507.5 123245.0 6372.5 123310.0 ;
      RECT  5107.5 124840.0 4972.5 124905.0 ;
      RECT  5457.5 124980.0 5322.5 125045.0 ;
      RECT  6682.5 125120.0 6547.5 125185.0 ;
      RECT  5107.5 126215.0 4972.5 126280.0 ;
      RECT  5457.5 126075.0 5322.5 126140.0 ;
      RECT  6857.5 125935.0 6722.5 126000.0 ;
      RECT  5107.5 127530.0 4972.5 127595.0 ;
      RECT  5457.5 127670.0 5322.5 127735.0 ;
      RECT  7032.5 127810.0 6897.5 127875.0 ;
      RECT  5107.5 128905.0 4972.5 128970.0 ;
      RECT  5457.5 128765.0 5322.5 128830.0 ;
      RECT  7207.5 128625.0 7072.5 128690.0 ;
      RECT  5107.5 130220.0 4972.5 130285.0 ;
      RECT  5457.5 130360.0 5322.5 130425.0 ;
      RECT  7382.5 130500.0 7247.5 130565.0 ;
      RECT  5107.5 131595.0 4972.5 131660.0 ;
      RECT  5632.5 131455.0 5497.5 131520.0 ;
      RECT  6157.5 131315.0 6022.5 131380.0 ;
      RECT  5107.5 132910.0 4972.5 132975.0 ;
      RECT  5632.5 133050.0 5497.5 133115.0 ;
      RECT  6332.5 133190.0 6197.5 133255.0 ;
      RECT  5107.5 134285.0 4972.5 134350.0 ;
      RECT  5632.5 134145.0 5497.5 134210.0 ;
      RECT  6507.5 134005.0 6372.5 134070.0 ;
      RECT  5107.5 135600.0 4972.5 135665.0 ;
      RECT  5632.5 135740.0 5497.5 135805.0 ;
      RECT  6682.5 135880.0 6547.5 135945.0 ;
      RECT  5107.5 136975.0 4972.5 137040.0 ;
      RECT  5632.5 136835.0 5497.5 136900.0 ;
      RECT  6857.5 136695.0 6722.5 136760.0 ;
      RECT  5107.5 138290.0 4972.5 138355.0 ;
      RECT  5632.5 138430.0 5497.5 138495.0 ;
      RECT  7032.5 138570.0 6897.5 138635.0 ;
      RECT  5107.5 139665.0 4972.5 139730.0 ;
      RECT  5632.5 139525.0 5497.5 139590.0 ;
      RECT  7207.5 139385.0 7072.5 139450.0 ;
      RECT  5107.5 140980.0 4972.5 141045.0 ;
      RECT  5632.5 141120.0 5497.5 141185.0 ;
      RECT  7382.5 141260.0 7247.5 141325.0 ;
      RECT  5107.5 142355.0 4972.5 142420.0 ;
      RECT  5807.5 142215.0 5672.5 142280.0 ;
      RECT  6157.5 142075.0 6022.5 142140.0 ;
      RECT  5107.5 143670.0 4972.5 143735.0 ;
      RECT  5807.5 143810.0 5672.5 143875.0 ;
      RECT  6332.5 143950.0 6197.5 144015.0 ;
      RECT  5107.5 145045.0 4972.5 145110.0 ;
      RECT  5807.5 144905.0 5672.5 144970.0 ;
      RECT  6507.5 144765.0 6372.5 144830.0 ;
      RECT  5107.5 146360.0 4972.5 146425.0 ;
      RECT  5807.5 146500.0 5672.5 146565.0 ;
      RECT  6682.5 146640.0 6547.5 146705.0 ;
      RECT  5107.5 147735.0 4972.5 147800.0 ;
      RECT  5807.5 147595.0 5672.5 147660.0 ;
      RECT  6857.5 147455.0 6722.5 147520.0 ;
      RECT  5107.5 149050.0 4972.5 149115.0 ;
      RECT  5807.5 149190.0 5672.5 149255.0 ;
      RECT  7032.5 149330.0 6897.5 149395.0 ;
      RECT  5107.5 150425.0 4972.5 150490.0 ;
      RECT  5807.5 150285.0 5672.5 150350.0 ;
      RECT  7207.5 150145.0 7072.5 150210.0 ;
      RECT  5107.5 151740.0 4972.5 151805.0 ;
      RECT  5807.5 151880.0 5672.5 151945.0 ;
      RECT  7382.5 152020.0 7247.5 152085.0 ;
      RECT  5107.5 153115.0 4972.5 153180.0 ;
      RECT  5982.5 152975.0 5847.5 153040.0 ;
      RECT  6157.5 152835.0 6022.5 152900.0 ;
      RECT  5107.5 154430.0 4972.5 154495.0 ;
      RECT  5982.5 154570.0 5847.5 154635.0 ;
      RECT  6332.5 154710.0 6197.5 154775.0 ;
      RECT  5107.5 155805.0 4972.5 155870.0 ;
      RECT  5982.5 155665.0 5847.5 155730.0 ;
      RECT  6507.5 155525.0 6372.5 155590.0 ;
      RECT  5107.5 157120.0 4972.5 157185.0 ;
      RECT  5982.5 157260.0 5847.5 157325.0 ;
      RECT  6682.5 157400.0 6547.5 157465.0 ;
      RECT  5107.5 158495.0 4972.5 158560.0 ;
      RECT  5982.5 158355.0 5847.5 158420.0 ;
      RECT  6857.5 158215.0 6722.5 158280.0 ;
      RECT  5107.5 159810.0 4972.5 159875.0 ;
      RECT  5982.5 159950.0 5847.5 160015.0 ;
      RECT  7032.5 160090.0 6897.5 160155.0 ;
      RECT  5107.5 161185.0 4972.5 161250.0 ;
      RECT  5982.5 161045.0 5847.5 161110.0 ;
      RECT  7207.5 160905.0 7072.5 160970.0 ;
      RECT  5107.5 162500.0 4972.5 162565.0 ;
      RECT  5982.5 162640.0 5847.5 162705.0 ;
      RECT  7382.5 162780.0 7247.5 162845.0 ;
      RECT  5282.5 163875.0 5147.5 163940.0 ;
      RECT  5457.5 163735.0 5322.5 163800.0 ;
      RECT  6157.5 163595.0 6022.5 163660.0 ;
      RECT  5282.5 165190.0 5147.5 165255.0 ;
      RECT  5457.5 165330.0 5322.5 165395.0 ;
      RECT  6332.5 165470.0 6197.5 165535.0 ;
      RECT  5282.5 166565.0 5147.5 166630.0 ;
      RECT  5457.5 166425.0 5322.5 166490.0 ;
      RECT  6507.5 166285.0 6372.5 166350.0 ;
      RECT  5282.5 167880.0 5147.5 167945.0 ;
      RECT  5457.5 168020.0 5322.5 168085.0 ;
      RECT  6682.5 168160.0 6547.5 168225.0 ;
      RECT  5282.5 169255.0 5147.5 169320.0 ;
      RECT  5457.5 169115.0 5322.5 169180.0 ;
      RECT  6857.5 168975.0 6722.5 169040.0 ;
      RECT  5282.5 170570.0 5147.5 170635.0 ;
      RECT  5457.5 170710.0 5322.5 170775.0 ;
      RECT  7032.5 170850.0 6897.5 170915.0 ;
      RECT  5282.5 171945.0 5147.5 172010.0 ;
      RECT  5457.5 171805.0 5322.5 171870.0 ;
      RECT  7207.5 171665.0 7072.5 171730.0 ;
      RECT  5282.5 173260.0 5147.5 173325.0 ;
      RECT  5457.5 173400.0 5322.5 173465.0 ;
      RECT  7382.5 173540.0 7247.5 173605.0 ;
      RECT  5282.5 174635.0 5147.5 174700.0 ;
      RECT  5632.5 174495.0 5497.5 174560.0 ;
      RECT  6157.5 174355.0 6022.5 174420.0 ;
      RECT  5282.5 175950.0 5147.5 176015.0 ;
      RECT  5632.5 176090.0 5497.5 176155.0 ;
      RECT  6332.5 176230.0 6197.5 176295.0 ;
      RECT  5282.5 177325.0 5147.5 177390.0 ;
      RECT  5632.5 177185.0 5497.5 177250.0 ;
      RECT  6507.5 177045.0 6372.5 177110.0 ;
      RECT  5282.5 178640.0 5147.5 178705.0 ;
      RECT  5632.5 178780.0 5497.5 178845.0 ;
      RECT  6682.5 178920.0 6547.5 178985.0 ;
      RECT  5282.5 180015.0 5147.5 180080.0 ;
      RECT  5632.5 179875.0 5497.5 179940.0 ;
      RECT  6857.5 179735.0 6722.5 179800.0 ;
      RECT  5282.5 181330.0 5147.5 181395.0 ;
      RECT  5632.5 181470.0 5497.5 181535.0 ;
      RECT  7032.5 181610.0 6897.5 181675.0 ;
      RECT  5282.5 182705.0 5147.5 182770.0 ;
      RECT  5632.5 182565.0 5497.5 182630.0 ;
      RECT  7207.5 182425.0 7072.5 182490.0 ;
      RECT  5282.5 184020.0 5147.5 184085.0 ;
      RECT  5632.5 184160.0 5497.5 184225.0 ;
      RECT  7382.5 184300.0 7247.5 184365.0 ;
      RECT  5282.5 185395.0 5147.5 185460.0 ;
      RECT  5807.5 185255.0 5672.5 185320.0 ;
      RECT  6157.5 185115.0 6022.5 185180.0 ;
      RECT  5282.5 186710.0 5147.5 186775.0 ;
      RECT  5807.5 186850.0 5672.5 186915.0 ;
      RECT  6332.5 186990.0 6197.5 187055.0 ;
      RECT  5282.5 188085.0 5147.5 188150.0 ;
      RECT  5807.5 187945.0 5672.5 188010.0 ;
      RECT  6507.5 187805.0 6372.5 187870.0 ;
      RECT  5282.5 189400.0 5147.5 189465.0 ;
      RECT  5807.5 189540.0 5672.5 189605.0 ;
      RECT  6682.5 189680.0 6547.5 189745.0 ;
      RECT  5282.5 190775.0 5147.5 190840.0 ;
      RECT  5807.5 190635.0 5672.5 190700.0 ;
      RECT  6857.5 190495.0 6722.5 190560.0 ;
      RECT  5282.5 192090.0 5147.5 192155.0 ;
      RECT  5807.5 192230.0 5672.5 192295.0 ;
      RECT  7032.5 192370.0 6897.5 192435.0 ;
      RECT  5282.5 193465.0 5147.5 193530.0 ;
      RECT  5807.5 193325.0 5672.5 193390.0 ;
      RECT  7207.5 193185.0 7072.5 193250.0 ;
      RECT  5282.5 194780.0 5147.5 194845.0 ;
      RECT  5807.5 194920.0 5672.5 194985.0 ;
      RECT  7382.5 195060.0 7247.5 195125.0 ;
      RECT  5282.5 196155.0 5147.5 196220.0 ;
      RECT  5982.5 196015.0 5847.5 196080.0 ;
      RECT  6157.5 195875.0 6022.5 195940.0 ;
      RECT  5282.5 197470.0 5147.5 197535.0 ;
      RECT  5982.5 197610.0 5847.5 197675.0 ;
      RECT  6332.5 197750.0 6197.5 197815.0 ;
      RECT  5282.5 198845.0 5147.5 198910.0 ;
      RECT  5982.5 198705.0 5847.5 198770.0 ;
      RECT  6507.5 198565.0 6372.5 198630.0 ;
      RECT  5282.5 200160.0 5147.5 200225.0 ;
      RECT  5982.5 200300.0 5847.5 200365.0 ;
      RECT  6682.5 200440.0 6547.5 200505.0 ;
      RECT  5282.5 201535.0 5147.5 201600.0 ;
      RECT  5982.5 201395.0 5847.5 201460.0 ;
      RECT  6857.5 201255.0 6722.5 201320.0 ;
      RECT  5282.5 202850.0 5147.5 202915.0 ;
      RECT  5982.5 202990.0 5847.5 203055.0 ;
      RECT  7032.5 203130.0 6897.5 203195.0 ;
      RECT  5282.5 204225.0 5147.5 204290.0 ;
      RECT  5982.5 204085.0 5847.5 204150.0 ;
      RECT  7207.5 203945.0 7072.5 204010.0 ;
      RECT  5282.5 205540.0 5147.5 205605.0 ;
      RECT  5982.5 205680.0 5847.5 205745.0 ;
      RECT  7382.5 205820.0 7247.5 205885.0 ;
      RECT  8755.0 34695.0 8820.0 34760.0 ;
      RECT  8755.0 36130.0 8820.0 36195.0 ;
      RECT  8755.0 37385.0 8820.0 37450.0 ;
      RECT  8755.0 38820.0 8820.0 38885.0 ;
      RECT  8755.0 40075.0 8820.0 40140.0 ;
      RECT  8755.0 41510.0 8820.0 41575.0 ;
      RECT  8755.0 42765.0 8820.0 42830.0 ;
      RECT  8755.0 44200.0 8820.0 44265.0 ;
      RECT  8755.0 45455.0 8820.0 45520.0 ;
      RECT  8755.0 46890.0 8820.0 46955.0 ;
      RECT  8755.0 48145.0 8820.0 48210.0 ;
      RECT  8755.0 49580.0 8820.0 49645.0 ;
      RECT  8755.0 50835.0 8820.0 50900.0 ;
      RECT  8755.0 52270.0 8820.0 52335.0 ;
      RECT  8755.0 53525.0 8820.0 53590.0 ;
      RECT  8755.0 54960.0 8820.0 55025.0 ;
      RECT  8755.0 56215.0 8820.0 56280.0 ;
      RECT  8755.0 57650.0 8820.0 57715.0 ;
      RECT  8755.0 58905.0 8820.0 58970.0 ;
      RECT  8755.0 60340.0 8820.0 60405.0 ;
      RECT  8755.0 61595.0 8820.0 61660.0 ;
      RECT  8755.0 63030.0 8820.0 63095.0 ;
      RECT  8755.0 64285.0 8820.0 64350.0 ;
      RECT  8755.0 65720.0 8820.0 65785.0 ;
      RECT  8755.0 66975.0 8820.0 67040.0 ;
      RECT  8755.0 68410.0 8820.0 68475.0 ;
      RECT  8755.0 69665.0 8820.0 69730.0 ;
      RECT  8755.0 71100.0 8820.0 71165.0 ;
      RECT  8755.0 72355.0 8820.0 72420.0 ;
      RECT  8755.0 73790.0 8820.0 73855.0 ;
      RECT  8755.0 75045.0 8820.0 75110.0 ;
      RECT  8755.0 76480.0 8820.0 76545.0 ;
      RECT  8755.0 77735.0 8820.0 77800.0 ;
      RECT  8755.0 79170.0 8820.0 79235.0 ;
      RECT  8755.0 80425.0 8820.0 80490.0 ;
      RECT  8755.0 81860.0 8820.0 81925.0 ;
      RECT  8755.0 83115.0 8820.0 83180.0 ;
      RECT  8755.0 84550.0 8820.0 84615.0 ;
      RECT  8755.0 85805.0 8820.0 85870.0 ;
      RECT  8755.0 87240.0 8820.0 87305.0 ;
      RECT  8755.0 88495.0 8820.0 88560.0 ;
      RECT  8755.0 89930.0 8820.0 89995.0 ;
      RECT  8755.0 91185.0 8820.0 91250.0 ;
      RECT  8755.0 92620.0 8820.0 92685.0 ;
      RECT  8755.0 93875.0 8820.0 93940.0 ;
      RECT  8755.0 95310.0 8820.0 95375.0 ;
      RECT  8755.0 96565.0 8820.0 96630.0 ;
      RECT  8755.0 98000.0 8820.0 98065.0 ;
      RECT  8755.0 99255.0 8820.0 99320.0 ;
      RECT  8755.0 100690.0 8820.0 100755.0 ;
      RECT  8755.0 101945.0 8820.0 102010.0 ;
      RECT  8755.0 103380.0 8820.0 103445.0 ;
      RECT  8755.0 104635.0 8820.0 104700.0 ;
      RECT  8755.0 106070.0 8820.0 106135.0 ;
      RECT  8755.0 107325.0 8820.0 107390.0 ;
      RECT  8755.0 108760.0 8820.0 108825.0 ;
      RECT  8755.0 110015.0 8820.0 110080.0 ;
      RECT  8755.0 111450.0 8820.0 111515.0 ;
      RECT  8755.0 112705.0 8820.0 112770.0 ;
      RECT  8755.0 114140.0 8820.0 114205.0 ;
      RECT  8755.0 115395.0 8820.0 115460.0 ;
      RECT  8755.0 116830.0 8820.0 116895.0 ;
      RECT  8755.0 118085.0 8820.0 118150.0 ;
      RECT  8755.0 119520.0 8820.0 119585.0 ;
      RECT  8755.0 120775.0 8820.0 120840.0 ;
      RECT  8755.0 122210.0 8820.0 122275.0 ;
      RECT  8755.0 123465.0 8820.0 123530.0 ;
      RECT  8755.0 124900.0 8820.0 124965.0 ;
      RECT  8755.0 126155.0 8820.0 126220.0 ;
      RECT  8755.0 127590.0 8820.0 127655.0 ;
      RECT  8755.0 128845.0 8820.0 128910.0 ;
      RECT  8755.0 130280.0 8820.0 130345.0 ;
      RECT  8755.0 131535.0 8820.0 131600.0 ;
      RECT  8755.0 132970.0 8820.0 133035.0 ;
      RECT  8755.0 134225.0 8820.0 134290.0 ;
      RECT  8755.0 135660.0 8820.0 135725.0 ;
      RECT  8755.0 136915.0 8820.0 136980.0 ;
      RECT  8755.0 138350.0 8820.0 138415.0 ;
      RECT  8755.0 139605.0 8820.0 139670.0 ;
      RECT  8755.0 141040.0 8820.0 141105.0 ;
      RECT  8755.0 142295.0 8820.0 142360.0 ;
      RECT  8755.0 143730.0 8820.0 143795.0 ;
      RECT  8755.0 144985.0 8820.0 145050.0 ;
      RECT  8755.0 146420.0 8820.0 146485.0 ;
      RECT  8755.0 147675.0 8820.0 147740.0 ;
      RECT  8755.0 149110.0 8820.0 149175.0 ;
      RECT  8755.0 150365.0 8820.0 150430.0 ;
      RECT  8755.0 151800.0 8820.0 151865.0 ;
      RECT  8755.0 153055.0 8820.0 153120.0 ;
      RECT  8755.0 154490.0 8820.0 154555.0 ;
      RECT  8755.0 155745.0 8820.0 155810.0 ;
      RECT  8755.0 157180.0 8820.0 157245.0 ;
      RECT  8755.0 158435.0 8820.0 158500.0 ;
      RECT  8755.0 159870.0 8820.0 159935.0 ;
      RECT  8755.0 161125.0 8820.0 161190.0 ;
      RECT  8755.0 162560.0 8820.0 162625.0 ;
      RECT  8755.0 163815.0 8820.0 163880.0 ;
      RECT  8755.0 165250.0 8820.0 165315.0 ;
      RECT  8755.0 166505.0 8820.0 166570.0 ;
      RECT  8755.0 167940.0 8820.0 168005.0 ;
      RECT  8755.0 169195.0 8820.0 169260.0 ;
      RECT  8755.0 170630.0 8820.0 170695.0 ;
      RECT  8755.0 171885.0 8820.0 171950.0 ;
      RECT  8755.0 173320.0 8820.0 173385.0 ;
      RECT  8755.0 174575.0 8820.0 174640.0 ;
      RECT  8755.0 176010.0 8820.0 176075.0 ;
      RECT  8755.0 177265.0 8820.0 177330.0 ;
      RECT  8755.0 178700.0 8820.0 178765.0 ;
      RECT  8755.0 179955.0 8820.0 180020.0 ;
      RECT  8755.0 181390.0 8820.0 181455.0 ;
      RECT  8755.0 182645.0 8820.0 182710.0 ;
      RECT  8755.0 184080.0 8820.0 184145.0 ;
      RECT  8755.0 185335.0 8820.0 185400.0 ;
      RECT  8755.0 186770.0 8820.0 186835.0 ;
      RECT  8755.0 188025.0 8820.0 188090.0 ;
      RECT  8755.0 189460.0 8820.0 189525.0 ;
      RECT  8755.0 190715.0 8820.0 190780.0 ;
      RECT  8755.0 192150.0 8820.0 192215.0 ;
      RECT  8755.0 193405.0 8820.0 193470.0 ;
      RECT  8755.0 194840.0 8820.0 194905.0 ;
      RECT  8755.0 196095.0 8820.0 196160.0 ;
      RECT  8755.0 197530.0 8820.0 197595.0 ;
      RECT  8755.0 198785.0 8820.0 198850.0 ;
      RECT  8755.0 200220.0 8820.0 200285.0 ;
      RECT  8755.0 201475.0 8820.0 201540.0 ;
      RECT  8755.0 202910.0 8820.0 202975.0 ;
      RECT  8755.0 204165.0 8820.0 204230.0 ;
      RECT  8755.0 205600.0 8820.0 205665.0 ;
      RECT  4655.0 13892.5 12335.0 13957.5 ;
      RECT  4655.0 16582.5 12335.0 16647.5 ;
      RECT  4655.0 19272.5 12335.0 19337.5 ;
      RECT  4655.0 21962.5 12335.0 22027.5 ;
      RECT  4655.0 24652.5 12335.0 24717.5 ;
      RECT  4655.0 27342.5 12335.0 27407.5 ;
      RECT  4655.0 30032.5 12335.0 30097.5 ;
      RECT  4655.0 32722.5 12335.0 32787.5 ;
      RECT  4655.0 35412.5 12335.0 35477.5 ;
      RECT  4655.0 38102.5 12335.0 38167.5 ;
      RECT  4655.0 40792.5 12335.0 40857.5 ;
      RECT  4655.0 43482.5 12335.0 43547.5 ;
      RECT  4655.0 46172.5 12335.0 46237.5 ;
      RECT  4655.0 48862.5 12335.0 48927.5 ;
      RECT  4655.0 51552.5 12335.0 51617.5 ;
      RECT  4655.0 54242.5 12335.0 54307.5 ;
      RECT  4655.0 56932.5 12335.0 56997.5 ;
      RECT  4655.0 59622.5 12335.0 59687.5 ;
      RECT  4655.0 62312.5 12335.0 62377.5 ;
      RECT  4655.0 65002.5 12335.0 65067.5 ;
      RECT  4655.0 67692.5 12335.0 67757.5 ;
      RECT  4655.0 70382.5 12335.0 70447.5 ;
      RECT  4655.0 73072.5 12335.0 73137.5 ;
      RECT  4655.0 75762.5 12335.0 75827.5 ;
      RECT  4655.0 78452.5 12335.0 78517.5 ;
      RECT  4655.0 81142.5 12335.0 81207.5 ;
      RECT  4655.0 83832.5 12335.0 83897.5 ;
      RECT  4655.0 86522.5 12335.0 86587.5 ;
      RECT  4655.0 89212.5 12335.0 89277.5 ;
      RECT  4655.0 91902.5 12335.0 91967.5 ;
      RECT  4655.0 94592.5 12335.0 94657.5 ;
      RECT  4655.0 97282.5 12335.0 97347.5 ;
      RECT  4655.0 99972.5 12335.0 100037.5 ;
      RECT  4655.0 102662.5 12335.0 102727.5 ;
      RECT  4655.0 105352.5 12335.0 105417.5 ;
      RECT  4655.0 108042.5 12335.0 108107.5 ;
      RECT  4655.0 110732.5 12335.0 110797.5 ;
      RECT  4655.0 113422.5 12335.0 113487.5 ;
      RECT  4655.0 116112.5 12335.0 116177.5 ;
      RECT  4655.0 118802.5 12335.0 118867.5 ;
      RECT  4655.0 121492.5 12335.0 121557.5 ;
      RECT  4655.0 124182.5 12335.0 124247.5 ;
      RECT  4655.0 126872.5 12335.0 126937.5 ;
      RECT  4655.0 129562.5 12335.0 129627.5 ;
      RECT  4655.0 132252.5 12335.0 132317.5 ;
      RECT  4655.0 134942.5 12335.0 135007.5 ;
      RECT  4655.0 137632.5 12335.0 137697.5 ;
      RECT  4655.0 140322.5 12335.0 140387.5 ;
      RECT  4655.0 143012.5 12335.0 143077.5 ;
      RECT  4655.0 145702.5 12335.0 145767.5 ;
      RECT  4655.0 148392.5 12335.0 148457.5 ;
      RECT  4655.0 151082.5 12335.0 151147.5 ;
      RECT  4655.0 153772.5 12335.0 153837.5 ;
      RECT  4655.0 156462.5 12335.0 156527.5 ;
      RECT  4655.0 159152.5 12335.0 159217.5 ;
      RECT  4655.0 161842.5 12335.0 161907.5 ;
      RECT  4655.0 164532.5 12335.0 164597.5 ;
      RECT  4655.0 167222.5 12335.0 167287.5 ;
      RECT  4655.0 169912.5 12335.0 169977.5 ;
      RECT  4655.0 172602.5 12335.0 172667.5 ;
      RECT  4655.0 175292.5 12335.0 175357.5 ;
      RECT  4655.0 177982.5 12335.0 178047.5 ;
      RECT  4655.0 180672.5 12335.0 180737.5 ;
      RECT  4655.0 183362.5 12335.0 183427.5 ;
      RECT  4655.0 186052.5 12335.0 186117.5 ;
      RECT  4655.0 188742.5 12335.0 188807.5 ;
      RECT  4655.0 191432.5 12335.0 191497.5 ;
      RECT  4655.0 194122.5 12335.0 194187.5 ;
      RECT  4655.0 196812.5 12335.0 196877.5 ;
      RECT  4655.0 199502.5 12335.0 199567.5 ;
      RECT  4655.0 202192.5 12335.0 202257.5 ;
      RECT  4655.0 204882.5 12335.0 204947.5 ;
      RECT  4655.0 12547.5 12335.0 12612.5 ;
      RECT  4655.0 15237.5 12335.0 15302.5 ;
      RECT  4655.0 17927.5 12335.0 17992.5 ;
      RECT  4655.0 20617.5 12335.0 20682.5 ;
      RECT  4655.0 23307.5 12335.0 23372.5 ;
      RECT  4655.0 25997.5 12335.0 26062.5 ;
      RECT  4655.0 28687.5 12335.0 28752.5 ;
      RECT  4655.0 31377.5 12335.0 31442.5 ;
      RECT  4655.0 34067.5 12335.0 34132.5 ;
      RECT  4655.0 36757.5 12335.0 36822.5 ;
      RECT  4655.0 39447.5 12335.0 39512.5 ;
      RECT  4655.0 42137.5 12335.0 42202.5 ;
      RECT  4655.0 44827.5 12335.0 44892.5 ;
      RECT  4655.0 47517.5 12335.0 47582.5 ;
      RECT  4655.0 50207.5 12335.0 50272.5 ;
      RECT  4655.0 52897.5 12335.0 52962.5 ;
      RECT  4655.0 55587.5 12335.0 55652.5 ;
      RECT  4655.0 58277.5 12335.0 58342.5 ;
      RECT  4655.0 60967.5 12335.0 61032.5 ;
      RECT  4655.0 63657.5 12335.0 63722.5 ;
      RECT  4655.0 66347.5 12335.0 66412.5 ;
      RECT  4655.0 69037.5 12335.0 69102.5 ;
      RECT  4655.0 71727.5 12335.0 71792.5 ;
      RECT  4655.0 74417.5 12335.0 74482.5 ;
      RECT  4655.0 77107.5 12335.0 77172.5 ;
      RECT  4655.0 79797.5 12335.0 79862.5 ;
      RECT  4655.0 82487.5 12335.0 82552.5 ;
      RECT  4655.0 85177.5 12335.0 85242.5 ;
      RECT  4655.0 87867.5 12335.0 87932.5 ;
      RECT  4655.0 90557.5 12335.0 90622.5 ;
      RECT  4655.0 93247.5 12335.0 93312.5 ;
      RECT  4655.0 95937.5 12335.0 96002.5 ;
      RECT  4655.0 98627.5 12335.0 98692.5 ;
      RECT  4655.0 101317.5 12335.0 101382.5 ;
      RECT  4655.0 104007.5 12335.0 104072.5 ;
      RECT  4655.0 106697.5 12335.0 106762.5 ;
      RECT  4655.0 109387.5 12335.0 109452.5 ;
      RECT  4655.0 112077.5 12335.0 112142.5 ;
      RECT  4655.0 114767.5 12335.0 114832.5 ;
      RECT  4655.0 117457.5 12335.0 117522.5 ;
      RECT  4655.0 120147.5 12335.0 120212.5 ;
      RECT  4655.0 122837.5 12335.0 122902.5 ;
      RECT  4655.0 125527.5 12335.0 125592.5 ;
      RECT  4655.0 128217.5 12335.0 128282.5 ;
      RECT  4655.0 130907.5 12335.0 130972.5 ;
      RECT  4655.0 133597.5 12335.0 133662.5 ;
      RECT  4655.0 136287.5 12335.0 136352.5 ;
      RECT  4655.0 138977.5 12335.0 139042.5 ;
      RECT  4655.0 141667.5 12335.0 141732.5 ;
      RECT  4655.0 144357.5 12335.0 144422.5 ;
      RECT  4655.0 147047.5 12335.0 147112.5 ;
      RECT  4655.0 149737.5 12335.0 149802.5 ;
      RECT  4655.0 152427.5 12335.0 152492.5 ;
      RECT  4655.0 155117.5 12335.0 155182.5 ;
      RECT  4655.0 157807.5 12335.0 157872.5 ;
      RECT  4655.0 160497.5 12335.0 160562.5 ;
      RECT  4655.0 163187.5 12335.0 163252.5 ;
      RECT  4655.0 165877.5 12335.0 165942.5 ;
      RECT  4655.0 168567.5 12335.0 168632.5 ;
      RECT  4655.0 171257.5 12335.0 171322.5 ;
      RECT  4655.0 173947.5 12335.0 174012.5 ;
      RECT  4655.0 176637.5 12335.0 176702.5 ;
      RECT  4655.0 179327.5 12335.0 179392.5 ;
      RECT  4655.0 182017.5 12335.0 182082.5 ;
      RECT  4655.0 184707.5 12335.0 184772.5 ;
      RECT  4655.0 187397.5 12335.0 187462.5 ;
      RECT  4655.0 190087.5 12335.0 190152.5 ;
      RECT  4655.0 192777.5 12335.0 192842.5 ;
      RECT  4655.0 195467.5 12335.0 195532.5 ;
      RECT  4655.0 198157.5 12335.0 198222.5 ;
      RECT  4655.0 200847.5 12335.0 200912.5 ;
      RECT  4655.0 203537.5 12335.0 203602.5 ;
      RECT  4655.0 206227.5 12335.0 206292.5 ;
      RECT  9255.0 34695.0 9605.0 34760.0 ;
      RECT  9770.0 34707.5 9835.0 34772.5 ;
      RECT  9770.0 34695.0 9835.0 34760.0 ;
      RECT  9770.0 34740.0 9835.0 34760.0 ;
      RECT  9802.5 34707.5 10100.0 34772.5 ;
      RECT  10100.0 34707.5 10235.0 34772.5 ;
      RECT  10805.0 34707.5 10870.0 34772.5 ;
      RECT  10805.0 34695.0 10870.0 34760.0 ;
      RECT  10587.5 34707.5 10837.5 34772.5 ;
      RECT  10805.0 34727.5 10870.0 34740.0 ;
      RECT  10837.5 34695.0 11085.0 34760.0 ;
      RECT  9255.0 36130.0 9605.0 36195.0 ;
      RECT  9770.0 36117.5 9835.0 36182.5 ;
      RECT  9770.0 36130.0 9835.0 36195.0 ;
      RECT  9770.0 36150.0 9835.0 36195.0 ;
      RECT  9802.5 36117.5 10100.0 36182.5 ;
      RECT  10100.0 36117.5 10235.0 36182.5 ;
      RECT  10805.0 36117.5 10870.0 36182.5 ;
      RECT  10805.0 36130.0 10870.0 36195.0 ;
      RECT  10587.5 36117.5 10837.5 36182.5 ;
      RECT  10805.0 36150.0 10870.0 36162.5 ;
      RECT  10837.5 36130.0 11085.0 36195.0 ;
      RECT  9255.0 37385.0 9605.0 37450.0 ;
      RECT  9770.0 37397.5 9835.0 37462.5 ;
      RECT  9770.0 37385.0 9835.0 37450.0 ;
      RECT  9770.0 37430.0 9835.0 37450.0 ;
      RECT  9802.5 37397.5 10100.0 37462.5 ;
      RECT  10100.0 37397.5 10235.0 37462.5 ;
      RECT  10805.0 37397.5 10870.0 37462.5 ;
      RECT  10805.0 37385.0 10870.0 37450.0 ;
      RECT  10587.5 37397.5 10837.5 37462.5 ;
      RECT  10805.0 37417.5 10870.0 37430.0 ;
      RECT  10837.5 37385.0 11085.0 37450.0 ;
      RECT  9255.0 38820.0 9605.0 38885.0 ;
      RECT  9770.0 38807.5 9835.0 38872.5 ;
      RECT  9770.0 38820.0 9835.0 38885.0 ;
      RECT  9770.0 38840.0 9835.0 38885.0 ;
      RECT  9802.5 38807.5 10100.0 38872.5 ;
      RECT  10100.0 38807.5 10235.0 38872.5 ;
      RECT  10805.0 38807.5 10870.0 38872.5 ;
      RECT  10805.0 38820.0 10870.0 38885.0 ;
      RECT  10587.5 38807.5 10837.5 38872.5 ;
      RECT  10805.0 38840.0 10870.0 38852.5 ;
      RECT  10837.5 38820.0 11085.0 38885.0 ;
      RECT  9255.0 40075.0 9605.0 40140.0 ;
      RECT  9770.0 40087.5 9835.0 40152.5 ;
      RECT  9770.0 40075.0 9835.0 40140.0 ;
      RECT  9770.0 40120.0 9835.0 40140.0 ;
      RECT  9802.5 40087.5 10100.0 40152.5 ;
      RECT  10100.0 40087.5 10235.0 40152.5 ;
      RECT  10805.0 40087.5 10870.0 40152.5 ;
      RECT  10805.0 40075.0 10870.0 40140.0 ;
      RECT  10587.5 40087.5 10837.5 40152.5 ;
      RECT  10805.0 40107.5 10870.0 40120.0 ;
      RECT  10837.5 40075.0 11085.0 40140.0 ;
      RECT  9255.0 41510.0 9605.0 41575.0 ;
      RECT  9770.0 41497.5 9835.0 41562.5 ;
      RECT  9770.0 41510.0 9835.0 41575.0 ;
      RECT  9770.0 41530.0 9835.0 41575.0 ;
      RECT  9802.5 41497.5 10100.0 41562.5 ;
      RECT  10100.0 41497.5 10235.0 41562.5 ;
      RECT  10805.0 41497.5 10870.0 41562.5 ;
      RECT  10805.0 41510.0 10870.0 41575.0 ;
      RECT  10587.5 41497.5 10837.5 41562.5 ;
      RECT  10805.0 41530.0 10870.0 41542.5 ;
      RECT  10837.5 41510.0 11085.0 41575.0 ;
      RECT  9255.0 42765.0 9605.0 42830.0 ;
      RECT  9770.0 42777.5 9835.0 42842.5 ;
      RECT  9770.0 42765.0 9835.0 42830.0 ;
      RECT  9770.0 42810.0 9835.0 42830.0 ;
      RECT  9802.5 42777.5 10100.0 42842.5 ;
      RECT  10100.0 42777.5 10235.0 42842.5 ;
      RECT  10805.0 42777.5 10870.0 42842.5 ;
      RECT  10805.0 42765.0 10870.0 42830.0 ;
      RECT  10587.5 42777.5 10837.5 42842.5 ;
      RECT  10805.0 42797.5 10870.0 42810.0 ;
      RECT  10837.5 42765.0 11085.0 42830.0 ;
      RECT  9255.0 44200.0 9605.0 44265.0 ;
      RECT  9770.0 44187.5 9835.0 44252.5 ;
      RECT  9770.0 44200.0 9835.0 44265.0 ;
      RECT  9770.0 44220.0 9835.0 44265.0 ;
      RECT  9802.5 44187.5 10100.0 44252.5 ;
      RECT  10100.0 44187.5 10235.0 44252.5 ;
      RECT  10805.0 44187.5 10870.0 44252.5 ;
      RECT  10805.0 44200.0 10870.0 44265.0 ;
      RECT  10587.5 44187.5 10837.5 44252.5 ;
      RECT  10805.0 44220.0 10870.0 44232.5 ;
      RECT  10837.5 44200.0 11085.0 44265.0 ;
      RECT  9255.0 45455.0 9605.0 45520.0 ;
      RECT  9770.0 45467.5 9835.0 45532.5 ;
      RECT  9770.0 45455.0 9835.0 45520.0 ;
      RECT  9770.0 45500.0 9835.0 45520.0 ;
      RECT  9802.5 45467.5 10100.0 45532.5 ;
      RECT  10100.0 45467.5 10235.0 45532.5 ;
      RECT  10805.0 45467.5 10870.0 45532.5 ;
      RECT  10805.0 45455.0 10870.0 45520.0 ;
      RECT  10587.5 45467.5 10837.5 45532.5 ;
      RECT  10805.0 45487.5 10870.0 45500.0 ;
      RECT  10837.5 45455.0 11085.0 45520.0 ;
      RECT  9255.0 46890.0 9605.0 46955.0 ;
      RECT  9770.0 46877.5 9835.0 46942.5 ;
      RECT  9770.0 46890.0 9835.0 46955.0 ;
      RECT  9770.0 46910.0 9835.0 46955.0 ;
      RECT  9802.5 46877.5 10100.0 46942.5 ;
      RECT  10100.0 46877.5 10235.0 46942.5 ;
      RECT  10805.0 46877.5 10870.0 46942.5 ;
      RECT  10805.0 46890.0 10870.0 46955.0 ;
      RECT  10587.5 46877.5 10837.5 46942.5 ;
      RECT  10805.0 46910.0 10870.0 46922.5 ;
      RECT  10837.5 46890.0 11085.0 46955.0 ;
      RECT  9255.0 48145.0 9605.0 48210.0 ;
      RECT  9770.0 48157.5 9835.0 48222.5 ;
      RECT  9770.0 48145.0 9835.0 48210.0 ;
      RECT  9770.0 48190.0 9835.0 48210.0 ;
      RECT  9802.5 48157.5 10100.0 48222.5 ;
      RECT  10100.0 48157.5 10235.0 48222.5 ;
      RECT  10805.0 48157.5 10870.0 48222.5 ;
      RECT  10805.0 48145.0 10870.0 48210.0 ;
      RECT  10587.5 48157.5 10837.5 48222.5 ;
      RECT  10805.0 48177.5 10870.0 48190.0 ;
      RECT  10837.5 48145.0 11085.0 48210.0 ;
      RECT  9255.0 49580.0 9605.0 49645.0 ;
      RECT  9770.0 49567.5 9835.0 49632.5 ;
      RECT  9770.0 49580.0 9835.0 49645.0 ;
      RECT  9770.0 49600.0 9835.0 49645.0 ;
      RECT  9802.5 49567.5 10100.0 49632.5 ;
      RECT  10100.0 49567.5 10235.0 49632.5 ;
      RECT  10805.0 49567.5 10870.0 49632.5 ;
      RECT  10805.0 49580.0 10870.0 49645.0 ;
      RECT  10587.5 49567.5 10837.5 49632.5 ;
      RECT  10805.0 49600.0 10870.0 49612.5 ;
      RECT  10837.5 49580.0 11085.0 49645.0 ;
      RECT  9255.0 50835.0 9605.0 50900.0 ;
      RECT  9770.0 50847.5 9835.0 50912.5 ;
      RECT  9770.0 50835.0 9835.0 50900.0 ;
      RECT  9770.0 50880.0 9835.0 50900.0 ;
      RECT  9802.5 50847.5 10100.0 50912.5 ;
      RECT  10100.0 50847.5 10235.0 50912.5 ;
      RECT  10805.0 50847.5 10870.0 50912.5 ;
      RECT  10805.0 50835.0 10870.0 50900.0 ;
      RECT  10587.5 50847.5 10837.5 50912.5 ;
      RECT  10805.0 50867.5 10870.0 50880.0 ;
      RECT  10837.5 50835.0 11085.0 50900.0 ;
      RECT  9255.0 52270.0 9605.0 52335.0 ;
      RECT  9770.0 52257.5 9835.0 52322.5 ;
      RECT  9770.0 52270.0 9835.0 52335.0 ;
      RECT  9770.0 52290.0 9835.0 52335.0 ;
      RECT  9802.5 52257.5 10100.0 52322.5 ;
      RECT  10100.0 52257.5 10235.0 52322.5 ;
      RECT  10805.0 52257.5 10870.0 52322.5 ;
      RECT  10805.0 52270.0 10870.0 52335.0 ;
      RECT  10587.5 52257.5 10837.5 52322.5 ;
      RECT  10805.0 52290.0 10870.0 52302.5 ;
      RECT  10837.5 52270.0 11085.0 52335.0 ;
      RECT  9255.0 53525.0 9605.0 53590.0 ;
      RECT  9770.0 53537.5 9835.0 53602.5 ;
      RECT  9770.0 53525.0 9835.0 53590.0 ;
      RECT  9770.0 53570.0 9835.0 53590.0 ;
      RECT  9802.5 53537.5 10100.0 53602.5 ;
      RECT  10100.0 53537.5 10235.0 53602.5 ;
      RECT  10805.0 53537.5 10870.0 53602.5 ;
      RECT  10805.0 53525.0 10870.0 53590.0 ;
      RECT  10587.5 53537.5 10837.5 53602.5 ;
      RECT  10805.0 53557.5 10870.0 53570.0 ;
      RECT  10837.5 53525.0 11085.0 53590.0 ;
      RECT  9255.0 54960.0 9605.0 55025.0 ;
      RECT  9770.0 54947.5 9835.0 55012.5 ;
      RECT  9770.0 54960.0 9835.0 55025.0 ;
      RECT  9770.0 54980.0 9835.0 55025.0 ;
      RECT  9802.5 54947.5 10100.0 55012.5 ;
      RECT  10100.0 54947.5 10235.0 55012.5 ;
      RECT  10805.0 54947.5 10870.0 55012.5 ;
      RECT  10805.0 54960.0 10870.0 55025.0 ;
      RECT  10587.5 54947.5 10837.5 55012.5 ;
      RECT  10805.0 54980.0 10870.0 54992.5 ;
      RECT  10837.5 54960.0 11085.0 55025.0 ;
      RECT  9255.0 56215.0 9605.0 56280.0 ;
      RECT  9770.0 56227.5 9835.0 56292.5 ;
      RECT  9770.0 56215.0 9835.0 56280.0 ;
      RECT  9770.0 56260.0 9835.0 56280.0 ;
      RECT  9802.5 56227.5 10100.0 56292.5 ;
      RECT  10100.0 56227.5 10235.0 56292.5 ;
      RECT  10805.0 56227.5 10870.0 56292.5 ;
      RECT  10805.0 56215.0 10870.0 56280.0 ;
      RECT  10587.5 56227.5 10837.5 56292.5 ;
      RECT  10805.0 56247.5 10870.0 56260.0 ;
      RECT  10837.5 56215.0 11085.0 56280.0 ;
      RECT  9255.0 57650.0 9605.0 57715.0 ;
      RECT  9770.0 57637.5 9835.0 57702.5 ;
      RECT  9770.0 57650.0 9835.0 57715.0 ;
      RECT  9770.0 57670.0 9835.0 57715.0 ;
      RECT  9802.5 57637.5 10100.0 57702.5 ;
      RECT  10100.0 57637.5 10235.0 57702.5 ;
      RECT  10805.0 57637.5 10870.0 57702.5 ;
      RECT  10805.0 57650.0 10870.0 57715.0 ;
      RECT  10587.5 57637.5 10837.5 57702.5 ;
      RECT  10805.0 57670.0 10870.0 57682.5 ;
      RECT  10837.5 57650.0 11085.0 57715.0 ;
      RECT  9255.0 58905.0 9605.0 58970.0 ;
      RECT  9770.0 58917.5 9835.0 58982.5 ;
      RECT  9770.0 58905.0 9835.0 58970.0 ;
      RECT  9770.0 58950.0 9835.0 58970.0 ;
      RECT  9802.5 58917.5 10100.0 58982.5 ;
      RECT  10100.0 58917.5 10235.0 58982.5 ;
      RECT  10805.0 58917.5 10870.0 58982.5 ;
      RECT  10805.0 58905.0 10870.0 58970.0 ;
      RECT  10587.5 58917.5 10837.5 58982.5 ;
      RECT  10805.0 58937.5 10870.0 58950.0 ;
      RECT  10837.5 58905.0 11085.0 58970.0 ;
      RECT  9255.0 60340.0 9605.0 60405.0 ;
      RECT  9770.0 60327.5 9835.0 60392.5 ;
      RECT  9770.0 60340.0 9835.0 60405.0 ;
      RECT  9770.0 60360.0 9835.0 60405.0 ;
      RECT  9802.5 60327.5 10100.0 60392.5 ;
      RECT  10100.0 60327.5 10235.0 60392.5 ;
      RECT  10805.0 60327.5 10870.0 60392.5 ;
      RECT  10805.0 60340.0 10870.0 60405.0 ;
      RECT  10587.5 60327.5 10837.5 60392.5 ;
      RECT  10805.0 60360.0 10870.0 60372.5 ;
      RECT  10837.5 60340.0 11085.0 60405.0 ;
      RECT  9255.0 61595.0 9605.0 61660.0 ;
      RECT  9770.0 61607.5 9835.0 61672.5 ;
      RECT  9770.0 61595.0 9835.0 61660.0 ;
      RECT  9770.0 61640.0 9835.0 61660.0 ;
      RECT  9802.5 61607.5 10100.0 61672.5 ;
      RECT  10100.0 61607.5 10235.0 61672.5 ;
      RECT  10805.0 61607.5 10870.0 61672.5 ;
      RECT  10805.0 61595.0 10870.0 61660.0 ;
      RECT  10587.5 61607.5 10837.5 61672.5 ;
      RECT  10805.0 61627.5 10870.0 61640.0 ;
      RECT  10837.5 61595.0 11085.0 61660.0 ;
      RECT  9255.0 63030.0 9605.0 63095.0 ;
      RECT  9770.0 63017.5 9835.0 63082.5 ;
      RECT  9770.0 63030.0 9835.0 63095.0 ;
      RECT  9770.0 63050.0 9835.0 63095.0 ;
      RECT  9802.5 63017.5 10100.0 63082.5 ;
      RECT  10100.0 63017.5 10235.0 63082.5 ;
      RECT  10805.0 63017.5 10870.0 63082.5 ;
      RECT  10805.0 63030.0 10870.0 63095.0 ;
      RECT  10587.5 63017.5 10837.5 63082.5 ;
      RECT  10805.0 63050.0 10870.0 63062.5 ;
      RECT  10837.5 63030.0 11085.0 63095.0 ;
      RECT  9255.0 64285.0 9605.0 64350.0 ;
      RECT  9770.0 64297.5 9835.0 64362.5 ;
      RECT  9770.0 64285.0 9835.0 64350.0 ;
      RECT  9770.0 64330.0 9835.0 64350.0 ;
      RECT  9802.5 64297.5 10100.0 64362.5 ;
      RECT  10100.0 64297.5 10235.0 64362.5 ;
      RECT  10805.0 64297.5 10870.0 64362.5 ;
      RECT  10805.0 64285.0 10870.0 64350.0 ;
      RECT  10587.5 64297.5 10837.5 64362.5 ;
      RECT  10805.0 64317.5 10870.0 64330.0 ;
      RECT  10837.5 64285.0 11085.0 64350.0 ;
      RECT  9255.0 65720.0 9605.0 65785.0 ;
      RECT  9770.0 65707.5 9835.0 65772.5 ;
      RECT  9770.0 65720.0 9835.0 65785.0 ;
      RECT  9770.0 65740.0 9835.0 65785.0 ;
      RECT  9802.5 65707.5 10100.0 65772.5 ;
      RECT  10100.0 65707.5 10235.0 65772.5 ;
      RECT  10805.0 65707.5 10870.0 65772.5 ;
      RECT  10805.0 65720.0 10870.0 65785.0 ;
      RECT  10587.5 65707.5 10837.5 65772.5 ;
      RECT  10805.0 65740.0 10870.0 65752.5 ;
      RECT  10837.5 65720.0 11085.0 65785.0 ;
      RECT  9255.0 66975.0 9605.0 67040.0 ;
      RECT  9770.0 66987.5 9835.0 67052.5 ;
      RECT  9770.0 66975.0 9835.0 67040.0 ;
      RECT  9770.0 67020.0 9835.0 67040.0 ;
      RECT  9802.5 66987.5 10100.0 67052.5 ;
      RECT  10100.0 66987.5 10235.0 67052.5 ;
      RECT  10805.0 66987.5 10870.0 67052.5 ;
      RECT  10805.0 66975.0 10870.0 67040.0 ;
      RECT  10587.5 66987.5 10837.5 67052.5 ;
      RECT  10805.0 67007.5 10870.0 67020.0 ;
      RECT  10837.5 66975.0 11085.0 67040.0 ;
      RECT  9255.0 68410.0 9605.0 68475.0 ;
      RECT  9770.0 68397.5 9835.0 68462.5 ;
      RECT  9770.0 68410.0 9835.0 68475.0 ;
      RECT  9770.0 68430.0 9835.0 68475.0 ;
      RECT  9802.5 68397.5 10100.0 68462.5 ;
      RECT  10100.0 68397.5 10235.0 68462.5 ;
      RECT  10805.0 68397.5 10870.0 68462.5 ;
      RECT  10805.0 68410.0 10870.0 68475.0 ;
      RECT  10587.5 68397.5 10837.5 68462.5 ;
      RECT  10805.0 68430.0 10870.0 68442.5 ;
      RECT  10837.5 68410.0 11085.0 68475.0 ;
      RECT  9255.0 69665.0 9605.0 69730.0 ;
      RECT  9770.0 69677.5 9835.0 69742.5 ;
      RECT  9770.0 69665.0 9835.0 69730.0 ;
      RECT  9770.0 69710.0 9835.0 69730.0 ;
      RECT  9802.5 69677.5 10100.0 69742.5 ;
      RECT  10100.0 69677.5 10235.0 69742.5 ;
      RECT  10805.0 69677.5 10870.0 69742.5 ;
      RECT  10805.0 69665.0 10870.0 69730.0 ;
      RECT  10587.5 69677.5 10837.5 69742.5 ;
      RECT  10805.0 69697.5 10870.0 69710.0 ;
      RECT  10837.5 69665.0 11085.0 69730.0 ;
      RECT  9255.0 71100.0 9605.0 71165.0 ;
      RECT  9770.0 71087.5 9835.0 71152.5 ;
      RECT  9770.0 71100.0 9835.0 71165.0 ;
      RECT  9770.0 71120.0 9835.0 71165.0 ;
      RECT  9802.5 71087.5 10100.0 71152.5 ;
      RECT  10100.0 71087.5 10235.0 71152.5 ;
      RECT  10805.0 71087.5 10870.0 71152.5 ;
      RECT  10805.0 71100.0 10870.0 71165.0 ;
      RECT  10587.5 71087.5 10837.5 71152.5 ;
      RECT  10805.0 71120.0 10870.0 71132.5 ;
      RECT  10837.5 71100.0 11085.0 71165.0 ;
      RECT  9255.0 72355.0 9605.0 72420.0 ;
      RECT  9770.0 72367.5 9835.0 72432.5 ;
      RECT  9770.0 72355.0 9835.0 72420.0 ;
      RECT  9770.0 72400.0 9835.0 72420.0 ;
      RECT  9802.5 72367.5 10100.0 72432.5 ;
      RECT  10100.0 72367.5 10235.0 72432.5 ;
      RECT  10805.0 72367.5 10870.0 72432.5 ;
      RECT  10805.0 72355.0 10870.0 72420.0 ;
      RECT  10587.5 72367.5 10837.5 72432.5 ;
      RECT  10805.0 72387.5 10870.0 72400.0 ;
      RECT  10837.5 72355.0 11085.0 72420.0 ;
      RECT  9255.0 73790.0 9605.0 73855.0 ;
      RECT  9770.0 73777.5 9835.0 73842.5 ;
      RECT  9770.0 73790.0 9835.0 73855.0 ;
      RECT  9770.0 73810.0 9835.0 73855.0 ;
      RECT  9802.5 73777.5 10100.0 73842.5 ;
      RECT  10100.0 73777.5 10235.0 73842.5 ;
      RECT  10805.0 73777.5 10870.0 73842.5 ;
      RECT  10805.0 73790.0 10870.0 73855.0 ;
      RECT  10587.5 73777.5 10837.5 73842.5 ;
      RECT  10805.0 73810.0 10870.0 73822.5 ;
      RECT  10837.5 73790.0 11085.0 73855.0 ;
      RECT  9255.0 75045.0 9605.0 75110.0 ;
      RECT  9770.0 75057.5 9835.0 75122.5 ;
      RECT  9770.0 75045.0 9835.0 75110.0 ;
      RECT  9770.0 75090.0 9835.0 75110.0 ;
      RECT  9802.5 75057.5 10100.0 75122.5 ;
      RECT  10100.0 75057.5 10235.0 75122.5 ;
      RECT  10805.0 75057.5 10870.0 75122.5 ;
      RECT  10805.0 75045.0 10870.0 75110.0 ;
      RECT  10587.5 75057.5 10837.5 75122.5 ;
      RECT  10805.0 75077.5 10870.0 75090.0 ;
      RECT  10837.5 75045.0 11085.0 75110.0 ;
      RECT  9255.0 76480.0 9605.0 76545.0 ;
      RECT  9770.0 76467.5 9835.0 76532.5 ;
      RECT  9770.0 76480.0 9835.0 76545.0 ;
      RECT  9770.0 76500.0 9835.0 76545.0 ;
      RECT  9802.5 76467.5 10100.0 76532.5 ;
      RECT  10100.0 76467.5 10235.0 76532.5 ;
      RECT  10805.0 76467.5 10870.0 76532.5 ;
      RECT  10805.0 76480.0 10870.0 76545.0 ;
      RECT  10587.5 76467.5 10837.5 76532.5 ;
      RECT  10805.0 76500.0 10870.0 76512.5 ;
      RECT  10837.5 76480.0 11085.0 76545.0 ;
      RECT  9255.0 77735.0 9605.0 77800.0 ;
      RECT  9770.0 77747.5 9835.0 77812.5 ;
      RECT  9770.0 77735.0 9835.0 77800.0 ;
      RECT  9770.0 77780.0 9835.0 77800.0 ;
      RECT  9802.5 77747.5 10100.0 77812.5 ;
      RECT  10100.0 77747.5 10235.0 77812.5 ;
      RECT  10805.0 77747.5 10870.0 77812.5 ;
      RECT  10805.0 77735.0 10870.0 77800.0 ;
      RECT  10587.5 77747.5 10837.5 77812.5 ;
      RECT  10805.0 77767.5 10870.0 77780.0 ;
      RECT  10837.5 77735.0 11085.0 77800.0 ;
      RECT  9255.0 79170.0 9605.0 79235.0 ;
      RECT  9770.0 79157.5 9835.0 79222.5 ;
      RECT  9770.0 79170.0 9835.0 79235.0 ;
      RECT  9770.0 79190.0 9835.0 79235.0 ;
      RECT  9802.5 79157.5 10100.0 79222.5 ;
      RECT  10100.0 79157.5 10235.0 79222.5 ;
      RECT  10805.0 79157.5 10870.0 79222.5 ;
      RECT  10805.0 79170.0 10870.0 79235.0 ;
      RECT  10587.5 79157.5 10837.5 79222.5 ;
      RECT  10805.0 79190.0 10870.0 79202.5 ;
      RECT  10837.5 79170.0 11085.0 79235.0 ;
      RECT  9255.0 80425.0 9605.0 80490.0 ;
      RECT  9770.0 80437.5 9835.0 80502.5 ;
      RECT  9770.0 80425.0 9835.0 80490.0 ;
      RECT  9770.0 80470.0 9835.0 80490.0 ;
      RECT  9802.5 80437.5 10100.0 80502.5 ;
      RECT  10100.0 80437.5 10235.0 80502.5 ;
      RECT  10805.0 80437.5 10870.0 80502.5 ;
      RECT  10805.0 80425.0 10870.0 80490.0 ;
      RECT  10587.5 80437.5 10837.5 80502.5 ;
      RECT  10805.0 80457.5 10870.0 80470.0 ;
      RECT  10837.5 80425.0 11085.0 80490.0 ;
      RECT  9255.0 81860.0 9605.0 81925.0 ;
      RECT  9770.0 81847.5 9835.0 81912.5 ;
      RECT  9770.0 81860.0 9835.0 81925.0 ;
      RECT  9770.0 81880.0 9835.0 81925.0 ;
      RECT  9802.5 81847.5 10100.0 81912.5 ;
      RECT  10100.0 81847.5 10235.0 81912.5 ;
      RECT  10805.0 81847.5 10870.0 81912.5 ;
      RECT  10805.0 81860.0 10870.0 81925.0 ;
      RECT  10587.5 81847.5 10837.5 81912.5 ;
      RECT  10805.0 81880.0 10870.0 81892.5 ;
      RECT  10837.5 81860.0 11085.0 81925.0 ;
      RECT  9255.0 83115.0 9605.0 83180.0 ;
      RECT  9770.0 83127.5 9835.0 83192.5 ;
      RECT  9770.0 83115.0 9835.0 83180.0 ;
      RECT  9770.0 83160.0 9835.0 83180.0 ;
      RECT  9802.5 83127.5 10100.0 83192.5 ;
      RECT  10100.0 83127.5 10235.0 83192.5 ;
      RECT  10805.0 83127.5 10870.0 83192.5 ;
      RECT  10805.0 83115.0 10870.0 83180.0 ;
      RECT  10587.5 83127.5 10837.5 83192.5 ;
      RECT  10805.0 83147.5 10870.0 83160.0 ;
      RECT  10837.5 83115.0 11085.0 83180.0 ;
      RECT  9255.0 84550.0 9605.0 84615.0 ;
      RECT  9770.0 84537.5 9835.0 84602.5 ;
      RECT  9770.0 84550.0 9835.0 84615.0 ;
      RECT  9770.0 84570.0 9835.0 84615.0 ;
      RECT  9802.5 84537.5 10100.0 84602.5 ;
      RECT  10100.0 84537.5 10235.0 84602.5 ;
      RECT  10805.0 84537.5 10870.0 84602.5 ;
      RECT  10805.0 84550.0 10870.0 84615.0 ;
      RECT  10587.5 84537.5 10837.5 84602.5 ;
      RECT  10805.0 84570.0 10870.0 84582.5 ;
      RECT  10837.5 84550.0 11085.0 84615.0 ;
      RECT  9255.0 85805.0 9605.0 85870.0 ;
      RECT  9770.0 85817.5 9835.0 85882.5 ;
      RECT  9770.0 85805.0 9835.0 85870.0 ;
      RECT  9770.0 85850.0 9835.0 85870.0 ;
      RECT  9802.5 85817.5 10100.0 85882.5 ;
      RECT  10100.0 85817.5 10235.0 85882.5 ;
      RECT  10805.0 85817.5 10870.0 85882.5 ;
      RECT  10805.0 85805.0 10870.0 85870.0 ;
      RECT  10587.5 85817.5 10837.5 85882.5 ;
      RECT  10805.0 85837.5 10870.0 85850.0 ;
      RECT  10837.5 85805.0 11085.0 85870.0 ;
      RECT  9255.0 87240.0 9605.0 87305.0 ;
      RECT  9770.0 87227.5 9835.0 87292.5 ;
      RECT  9770.0 87240.0 9835.0 87305.0 ;
      RECT  9770.0 87260.0 9835.0 87305.0 ;
      RECT  9802.5 87227.5 10100.0 87292.5 ;
      RECT  10100.0 87227.5 10235.0 87292.5 ;
      RECT  10805.0 87227.5 10870.0 87292.5 ;
      RECT  10805.0 87240.0 10870.0 87305.0 ;
      RECT  10587.5 87227.5 10837.5 87292.5 ;
      RECT  10805.0 87260.0 10870.0 87272.5 ;
      RECT  10837.5 87240.0 11085.0 87305.0 ;
      RECT  9255.0 88495.0 9605.0 88560.0 ;
      RECT  9770.0 88507.5 9835.0 88572.5 ;
      RECT  9770.0 88495.0 9835.0 88560.0 ;
      RECT  9770.0 88540.0 9835.0 88560.0 ;
      RECT  9802.5 88507.5 10100.0 88572.5 ;
      RECT  10100.0 88507.5 10235.0 88572.5 ;
      RECT  10805.0 88507.5 10870.0 88572.5 ;
      RECT  10805.0 88495.0 10870.0 88560.0 ;
      RECT  10587.5 88507.5 10837.5 88572.5 ;
      RECT  10805.0 88527.5 10870.0 88540.0 ;
      RECT  10837.5 88495.0 11085.0 88560.0 ;
      RECT  9255.0 89930.0 9605.0 89995.0 ;
      RECT  9770.0 89917.5 9835.0 89982.5 ;
      RECT  9770.0 89930.0 9835.0 89995.0 ;
      RECT  9770.0 89950.0 9835.0 89995.0 ;
      RECT  9802.5 89917.5 10100.0 89982.5 ;
      RECT  10100.0 89917.5 10235.0 89982.5 ;
      RECT  10805.0 89917.5 10870.0 89982.5 ;
      RECT  10805.0 89930.0 10870.0 89995.0 ;
      RECT  10587.5 89917.5 10837.5 89982.5 ;
      RECT  10805.0 89950.0 10870.0 89962.5 ;
      RECT  10837.5 89930.0 11085.0 89995.0 ;
      RECT  9255.0 91185.0 9605.0 91250.0 ;
      RECT  9770.0 91197.5 9835.0 91262.5 ;
      RECT  9770.0 91185.0 9835.0 91250.0 ;
      RECT  9770.0 91230.0 9835.0 91250.0 ;
      RECT  9802.5 91197.5 10100.0 91262.5 ;
      RECT  10100.0 91197.5 10235.0 91262.5 ;
      RECT  10805.0 91197.5 10870.0 91262.5 ;
      RECT  10805.0 91185.0 10870.0 91250.0 ;
      RECT  10587.5 91197.5 10837.5 91262.5 ;
      RECT  10805.0 91217.5 10870.0 91230.0 ;
      RECT  10837.5 91185.0 11085.0 91250.0 ;
      RECT  9255.0 92620.0 9605.0 92685.0 ;
      RECT  9770.0 92607.5 9835.0 92672.5 ;
      RECT  9770.0 92620.0 9835.0 92685.0 ;
      RECT  9770.0 92640.0 9835.0 92685.0 ;
      RECT  9802.5 92607.5 10100.0 92672.5 ;
      RECT  10100.0 92607.5 10235.0 92672.5 ;
      RECT  10805.0 92607.5 10870.0 92672.5 ;
      RECT  10805.0 92620.0 10870.0 92685.0 ;
      RECT  10587.5 92607.5 10837.5 92672.5 ;
      RECT  10805.0 92640.0 10870.0 92652.5 ;
      RECT  10837.5 92620.0 11085.0 92685.0 ;
      RECT  9255.0 93875.0 9605.0 93940.0 ;
      RECT  9770.0 93887.5 9835.0 93952.5 ;
      RECT  9770.0 93875.0 9835.0 93940.0 ;
      RECT  9770.0 93920.0 9835.0 93940.0 ;
      RECT  9802.5 93887.5 10100.0 93952.5 ;
      RECT  10100.0 93887.5 10235.0 93952.5 ;
      RECT  10805.0 93887.5 10870.0 93952.5 ;
      RECT  10805.0 93875.0 10870.0 93940.0 ;
      RECT  10587.5 93887.5 10837.5 93952.5 ;
      RECT  10805.0 93907.5 10870.0 93920.0 ;
      RECT  10837.5 93875.0 11085.0 93940.0 ;
      RECT  9255.0 95310.0 9605.0 95375.0 ;
      RECT  9770.0 95297.5 9835.0 95362.5 ;
      RECT  9770.0 95310.0 9835.0 95375.0 ;
      RECT  9770.0 95330.0 9835.0 95375.0 ;
      RECT  9802.5 95297.5 10100.0 95362.5 ;
      RECT  10100.0 95297.5 10235.0 95362.5 ;
      RECT  10805.0 95297.5 10870.0 95362.5 ;
      RECT  10805.0 95310.0 10870.0 95375.0 ;
      RECT  10587.5 95297.5 10837.5 95362.5 ;
      RECT  10805.0 95330.0 10870.0 95342.5 ;
      RECT  10837.5 95310.0 11085.0 95375.0 ;
      RECT  9255.0 96565.0 9605.0 96630.0 ;
      RECT  9770.0 96577.5 9835.0 96642.5 ;
      RECT  9770.0 96565.0 9835.0 96630.0 ;
      RECT  9770.0 96610.0 9835.0 96630.0 ;
      RECT  9802.5 96577.5 10100.0 96642.5 ;
      RECT  10100.0 96577.5 10235.0 96642.5 ;
      RECT  10805.0 96577.5 10870.0 96642.5 ;
      RECT  10805.0 96565.0 10870.0 96630.0 ;
      RECT  10587.5 96577.5 10837.5 96642.5 ;
      RECT  10805.0 96597.5 10870.0 96610.0 ;
      RECT  10837.5 96565.0 11085.0 96630.0 ;
      RECT  9255.0 98000.0 9605.0 98065.0 ;
      RECT  9770.0 97987.5 9835.0 98052.5 ;
      RECT  9770.0 98000.0 9835.0 98065.0 ;
      RECT  9770.0 98020.0 9835.0 98065.0 ;
      RECT  9802.5 97987.5 10100.0 98052.5 ;
      RECT  10100.0 97987.5 10235.0 98052.5 ;
      RECT  10805.0 97987.5 10870.0 98052.5 ;
      RECT  10805.0 98000.0 10870.0 98065.0 ;
      RECT  10587.5 97987.5 10837.5 98052.5 ;
      RECT  10805.0 98020.0 10870.0 98032.5 ;
      RECT  10837.5 98000.0 11085.0 98065.0 ;
      RECT  9255.0 99255.0 9605.0 99320.0 ;
      RECT  9770.0 99267.5 9835.0 99332.5 ;
      RECT  9770.0 99255.0 9835.0 99320.0 ;
      RECT  9770.0 99300.0 9835.0 99320.0 ;
      RECT  9802.5 99267.5 10100.0 99332.5 ;
      RECT  10100.0 99267.5 10235.0 99332.5 ;
      RECT  10805.0 99267.5 10870.0 99332.5 ;
      RECT  10805.0 99255.0 10870.0 99320.0 ;
      RECT  10587.5 99267.5 10837.5 99332.5 ;
      RECT  10805.0 99287.5 10870.0 99300.0 ;
      RECT  10837.5 99255.0 11085.0 99320.0 ;
      RECT  9255.0 100690.0 9605.0 100755.0 ;
      RECT  9770.0 100677.5 9835.0 100742.5 ;
      RECT  9770.0 100690.0 9835.0 100755.0 ;
      RECT  9770.0 100710.0 9835.0 100755.0 ;
      RECT  9802.5 100677.5 10100.0 100742.5 ;
      RECT  10100.0 100677.5 10235.0 100742.5 ;
      RECT  10805.0 100677.5 10870.0 100742.5 ;
      RECT  10805.0 100690.0 10870.0 100755.0 ;
      RECT  10587.5 100677.5 10837.5 100742.5 ;
      RECT  10805.0 100710.0 10870.0 100722.5 ;
      RECT  10837.5 100690.0 11085.0 100755.0 ;
      RECT  9255.0 101945.0 9605.0 102010.0 ;
      RECT  9770.0 101957.5 9835.0 102022.5 ;
      RECT  9770.0 101945.0 9835.0 102010.0 ;
      RECT  9770.0 101990.0 9835.0 102010.0 ;
      RECT  9802.5 101957.5 10100.0 102022.5 ;
      RECT  10100.0 101957.5 10235.0 102022.5 ;
      RECT  10805.0 101957.5 10870.0 102022.5 ;
      RECT  10805.0 101945.0 10870.0 102010.0 ;
      RECT  10587.5 101957.5 10837.5 102022.5 ;
      RECT  10805.0 101977.5 10870.0 101990.0 ;
      RECT  10837.5 101945.0 11085.0 102010.0 ;
      RECT  9255.0 103380.0 9605.0 103445.0 ;
      RECT  9770.0 103367.5 9835.0 103432.5 ;
      RECT  9770.0 103380.0 9835.0 103445.0 ;
      RECT  9770.0 103400.0 9835.0 103445.0 ;
      RECT  9802.5 103367.5 10100.0 103432.5 ;
      RECT  10100.0 103367.5 10235.0 103432.5 ;
      RECT  10805.0 103367.5 10870.0 103432.5 ;
      RECT  10805.0 103380.0 10870.0 103445.0 ;
      RECT  10587.5 103367.5 10837.5 103432.5 ;
      RECT  10805.0 103400.0 10870.0 103412.5 ;
      RECT  10837.5 103380.0 11085.0 103445.0 ;
      RECT  9255.0 104635.0 9605.0 104700.0 ;
      RECT  9770.0 104647.5 9835.0 104712.5 ;
      RECT  9770.0 104635.0 9835.0 104700.0 ;
      RECT  9770.0 104680.0 9835.0 104700.0 ;
      RECT  9802.5 104647.5 10100.0 104712.5 ;
      RECT  10100.0 104647.5 10235.0 104712.5 ;
      RECT  10805.0 104647.5 10870.0 104712.5 ;
      RECT  10805.0 104635.0 10870.0 104700.0 ;
      RECT  10587.5 104647.5 10837.5 104712.5 ;
      RECT  10805.0 104667.5 10870.0 104680.0 ;
      RECT  10837.5 104635.0 11085.0 104700.0 ;
      RECT  9255.0 106070.0 9605.0 106135.0 ;
      RECT  9770.0 106057.5 9835.0 106122.5 ;
      RECT  9770.0 106070.0 9835.0 106135.0 ;
      RECT  9770.0 106090.0 9835.0 106135.0 ;
      RECT  9802.5 106057.5 10100.0 106122.5 ;
      RECT  10100.0 106057.5 10235.0 106122.5 ;
      RECT  10805.0 106057.5 10870.0 106122.5 ;
      RECT  10805.0 106070.0 10870.0 106135.0 ;
      RECT  10587.5 106057.5 10837.5 106122.5 ;
      RECT  10805.0 106090.0 10870.0 106102.5 ;
      RECT  10837.5 106070.0 11085.0 106135.0 ;
      RECT  9255.0 107325.0 9605.0 107390.0 ;
      RECT  9770.0 107337.5 9835.0 107402.5 ;
      RECT  9770.0 107325.0 9835.0 107390.0 ;
      RECT  9770.0 107370.0 9835.0 107390.0 ;
      RECT  9802.5 107337.5 10100.0 107402.5 ;
      RECT  10100.0 107337.5 10235.0 107402.5 ;
      RECT  10805.0 107337.5 10870.0 107402.5 ;
      RECT  10805.0 107325.0 10870.0 107390.0 ;
      RECT  10587.5 107337.5 10837.5 107402.5 ;
      RECT  10805.0 107357.5 10870.0 107370.0 ;
      RECT  10837.5 107325.0 11085.0 107390.0 ;
      RECT  9255.0 108760.0 9605.0 108825.0 ;
      RECT  9770.0 108747.5 9835.0 108812.5 ;
      RECT  9770.0 108760.0 9835.0 108825.0 ;
      RECT  9770.0 108780.0 9835.0 108825.0 ;
      RECT  9802.5 108747.5 10100.0 108812.5 ;
      RECT  10100.0 108747.5 10235.0 108812.5 ;
      RECT  10805.0 108747.5 10870.0 108812.5 ;
      RECT  10805.0 108760.0 10870.0 108825.0 ;
      RECT  10587.5 108747.5 10837.5 108812.5 ;
      RECT  10805.0 108780.0 10870.0 108792.5 ;
      RECT  10837.5 108760.0 11085.0 108825.0 ;
      RECT  9255.0 110015.0 9605.0 110080.0 ;
      RECT  9770.0 110027.5 9835.0 110092.5 ;
      RECT  9770.0 110015.0 9835.0 110080.0 ;
      RECT  9770.0 110060.0 9835.0 110080.0 ;
      RECT  9802.5 110027.5 10100.0 110092.5 ;
      RECT  10100.0 110027.5 10235.0 110092.5 ;
      RECT  10805.0 110027.5 10870.0 110092.5 ;
      RECT  10805.0 110015.0 10870.0 110080.0 ;
      RECT  10587.5 110027.5 10837.5 110092.5 ;
      RECT  10805.0 110047.5 10870.0 110060.0 ;
      RECT  10837.5 110015.0 11085.0 110080.0 ;
      RECT  9255.0 111450.0 9605.0 111515.0 ;
      RECT  9770.0 111437.5 9835.0 111502.5 ;
      RECT  9770.0 111450.0 9835.0 111515.0 ;
      RECT  9770.0 111470.0 9835.0 111515.0 ;
      RECT  9802.5 111437.5 10100.0 111502.5 ;
      RECT  10100.0 111437.5 10235.0 111502.5 ;
      RECT  10805.0 111437.5 10870.0 111502.5 ;
      RECT  10805.0 111450.0 10870.0 111515.0 ;
      RECT  10587.5 111437.5 10837.5 111502.5 ;
      RECT  10805.0 111470.0 10870.0 111482.5 ;
      RECT  10837.5 111450.0 11085.0 111515.0 ;
      RECT  9255.0 112705.0 9605.0 112770.0 ;
      RECT  9770.0 112717.5 9835.0 112782.5 ;
      RECT  9770.0 112705.0 9835.0 112770.0 ;
      RECT  9770.0 112750.0 9835.0 112770.0 ;
      RECT  9802.5 112717.5 10100.0 112782.5 ;
      RECT  10100.0 112717.5 10235.0 112782.5 ;
      RECT  10805.0 112717.5 10870.0 112782.5 ;
      RECT  10805.0 112705.0 10870.0 112770.0 ;
      RECT  10587.5 112717.5 10837.5 112782.5 ;
      RECT  10805.0 112737.5 10870.0 112750.0 ;
      RECT  10837.5 112705.0 11085.0 112770.0 ;
      RECT  9255.0 114140.0 9605.0 114205.0 ;
      RECT  9770.0 114127.5 9835.0 114192.5 ;
      RECT  9770.0 114140.0 9835.0 114205.0 ;
      RECT  9770.0 114160.0 9835.0 114205.0 ;
      RECT  9802.5 114127.5 10100.0 114192.5 ;
      RECT  10100.0 114127.5 10235.0 114192.5 ;
      RECT  10805.0 114127.5 10870.0 114192.5 ;
      RECT  10805.0 114140.0 10870.0 114205.0 ;
      RECT  10587.5 114127.5 10837.5 114192.5 ;
      RECT  10805.0 114160.0 10870.0 114172.5 ;
      RECT  10837.5 114140.0 11085.0 114205.0 ;
      RECT  9255.0 115395.0 9605.0 115460.0 ;
      RECT  9770.0 115407.5 9835.0 115472.5 ;
      RECT  9770.0 115395.0 9835.0 115460.0 ;
      RECT  9770.0 115440.0 9835.0 115460.0 ;
      RECT  9802.5 115407.5 10100.0 115472.5 ;
      RECT  10100.0 115407.5 10235.0 115472.5 ;
      RECT  10805.0 115407.5 10870.0 115472.5 ;
      RECT  10805.0 115395.0 10870.0 115460.0 ;
      RECT  10587.5 115407.5 10837.5 115472.5 ;
      RECT  10805.0 115427.5 10870.0 115440.0 ;
      RECT  10837.5 115395.0 11085.0 115460.0 ;
      RECT  9255.0 116830.0 9605.0 116895.0 ;
      RECT  9770.0 116817.5 9835.0 116882.5 ;
      RECT  9770.0 116830.0 9835.0 116895.0 ;
      RECT  9770.0 116850.0 9835.0 116895.0 ;
      RECT  9802.5 116817.5 10100.0 116882.5 ;
      RECT  10100.0 116817.5 10235.0 116882.5 ;
      RECT  10805.0 116817.5 10870.0 116882.5 ;
      RECT  10805.0 116830.0 10870.0 116895.0 ;
      RECT  10587.5 116817.5 10837.5 116882.5 ;
      RECT  10805.0 116850.0 10870.0 116862.5 ;
      RECT  10837.5 116830.0 11085.0 116895.0 ;
      RECT  9255.0 118085.0 9605.0 118150.0 ;
      RECT  9770.0 118097.5 9835.0 118162.5 ;
      RECT  9770.0 118085.0 9835.0 118150.0 ;
      RECT  9770.0 118130.0 9835.0 118150.0 ;
      RECT  9802.5 118097.5 10100.0 118162.5 ;
      RECT  10100.0 118097.5 10235.0 118162.5 ;
      RECT  10805.0 118097.5 10870.0 118162.5 ;
      RECT  10805.0 118085.0 10870.0 118150.0 ;
      RECT  10587.5 118097.5 10837.5 118162.5 ;
      RECT  10805.0 118117.5 10870.0 118130.0 ;
      RECT  10837.5 118085.0 11085.0 118150.0 ;
      RECT  9255.0 119520.0 9605.0 119585.0 ;
      RECT  9770.0 119507.5 9835.0 119572.5 ;
      RECT  9770.0 119520.0 9835.0 119585.0 ;
      RECT  9770.0 119540.0 9835.0 119585.0 ;
      RECT  9802.5 119507.5 10100.0 119572.5 ;
      RECT  10100.0 119507.5 10235.0 119572.5 ;
      RECT  10805.0 119507.5 10870.0 119572.5 ;
      RECT  10805.0 119520.0 10870.0 119585.0 ;
      RECT  10587.5 119507.5 10837.5 119572.5 ;
      RECT  10805.0 119540.0 10870.0 119552.5 ;
      RECT  10837.5 119520.0 11085.0 119585.0 ;
      RECT  9255.0 120775.0 9605.0 120840.0 ;
      RECT  9770.0 120787.5 9835.0 120852.5 ;
      RECT  9770.0 120775.0 9835.0 120840.0 ;
      RECT  9770.0 120820.0 9835.0 120840.0 ;
      RECT  9802.5 120787.5 10100.0 120852.5 ;
      RECT  10100.0 120787.5 10235.0 120852.5 ;
      RECT  10805.0 120787.5 10870.0 120852.5 ;
      RECT  10805.0 120775.0 10870.0 120840.0 ;
      RECT  10587.5 120787.5 10837.5 120852.5 ;
      RECT  10805.0 120807.5 10870.0 120820.0 ;
      RECT  10837.5 120775.0 11085.0 120840.0 ;
      RECT  9255.0 122210.0 9605.0 122275.0 ;
      RECT  9770.0 122197.5 9835.0 122262.5 ;
      RECT  9770.0 122210.0 9835.0 122275.0 ;
      RECT  9770.0 122230.0 9835.0 122275.0 ;
      RECT  9802.5 122197.5 10100.0 122262.5 ;
      RECT  10100.0 122197.5 10235.0 122262.5 ;
      RECT  10805.0 122197.5 10870.0 122262.5 ;
      RECT  10805.0 122210.0 10870.0 122275.0 ;
      RECT  10587.5 122197.5 10837.5 122262.5 ;
      RECT  10805.0 122230.0 10870.0 122242.5 ;
      RECT  10837.5 122210.0 11085.0 122275.0 ;
      RECT  9255.0 123465.0 9605.0 123530.0 ;
      RECT  9770.0 123477.5 9835.0 123542.5 ;
      RECT  9770.0 123465.0 9835.0 123530.0 ;
      RECT  9770.0 123510.0 9835.0 123530.0 ;
      RECT  9802.5 123477.5 10100.0 123542.5 ;
      RECT  10100.0 123477.5 10235.0 123542.5 ;
      RECT  10805.0 123477.5 10870.0 123542.5 ;
      RECT  10805.0 123465.0 10870.0 123530.0 ;
      RECT  10587.5 123477.5 10837.5 123542.5 ;
      RECT  10805.0 123497.5 10870.0 123510.0 ;
      RECT  10837.5 123465.0 11085.0 123530.0 ;
      RECT  9255.0 124900.0 9605.0 124965.0 ;
      RECT  9770.0 124887.5 9835.0 124952.5 ;
      RECT  9770.0 124900.0 9835.0 124965.0 ;
      RECT  9770.0 124920.0 9835.0 124965.0 ;
      RECT  9802.5 124887.5 10100.0 124952.5 ;
      RECT  10100.0 124887.5 10235.0 124952.5 ;
      RECT  10805.0 124887.5 10870.0 124952.5 ;
      RECT  10805.0 124900.0 10870.0 124965.0 ;
      RECT  10587.5 124887.5 10837.5 124952.5 ;
      RECT  10805.0 124920.0 10870.0 124932.5 ;
      RECT  10837.5 124900.0 11085.0 124965.0 ;
      RECT  9255.0 126155.0 9605.0 126220.0 ;
      RECT  9770.0 126167.5 9835.0 126232.5 ;
      RECT  9770.0 126155.0 9835.0 126220.0 ;
      RECT  9770.0 126200.0 9835.0 126220.0 ;
      RECT  9802.5 126167.5 10100.0 126232.5 ;
      RECT  10100.0 126167.5 10235.0 126232.5 ;
      RECT  10805.0 126167.5 10870.0 126232.5 ;
      RECT  10805.0 126155.0 10870.0 126220.0 ;
      RECT  10587.5 126167.5 10837.5 126232.5 ;
      RECT  10805.0 126187.5 10870.0 126200.0 ;
      RECT  10837.5 126155.0 11085.0 126220.0 ;
      RECT  9255.0 127590.0 9605.0 127655.0 ;
      RECT  9770.0 127577.5 9835.0 127642.5 ;
      RECT  9770.0 127590.0 9835.0 127655.0 ;
      RECT  9770.0 127610.0 9835.0 127655.0 ;
      RECT  9802.5 127577.5 10100.0 127642.5 ;
      RECT  10100.0 127577.5 10235.0 127642.5 ;
      RECT  10805.0 127577.5 10870.0 127642.5 ;
      RECT  10805.0 127590.0 10870.0 127655.0 ;
      RECT  10587.5 127577.5 10837.5 127642.5 ;
      RECT  10805.0 127610.0 10870.0 127622.5 ;
      RECT  10837.5 127590.0 11085.0 127655.0 ;
      RECT  9255.0 128845.0 9605.0 128910.0 ;
      RECT  9770.0 128857.5 9835.0 128922.5 ;
      RECT  9770.0 128845.0 9835.0 128910.0 ;
      RECT  9770.0 128890.0 9835.0 128910.0 ;
      RECT  9802.5 128857.5 10100.0 128922.5 ;
      RECT  10100.0 128857.5 10235.0 128922.5 ;
      RECT  10805.0 128857.5 10870.0 128922.5 ;
      RECT  10805.0 128845.0 10870.0 128910.0 ;
      RECT  10587.5 128857.5 10837.5 128922.5 ;
      RECT  10805.0 128877.5 10870.0 128890.0 ;
      RECT  10837.5 128845.0 11085.0 128910.0 ;
      RECT  9255.0 130280.0 9605.0 130345.0 ;
      RECT  9770.0 130267.5 9835.0 130332.5 ;
      RECT  9770.0 130280.0 9835.0 130345.0 ;
      RECT  9770.0 130300.0 9835.0 130345.0 ;
      RECT  9802.5 130267.5 10100.0 130332.5 ;
      RECT  10100.0 130267.5 10235.0 130332.5 ;
      RECT  10805.0 130267.5 10870.0 130332.5 ;
      RECT  10805.0 130280.0 10870.0 130345.0 ;
      RECT  10587.5 130267.5 10837.5 130332.5 ;
      RECT  10805.0 130300.0 10870.0 130312.5 ;
      RECT  10837.5 130280.0 11085.0 130345.0 ;
      RECT  9255.0 131535.0 9605.0 131600.0 ;
      RECT  9770.0 131547.5 9835.0 131612.5 ;
      RECT  9770.0 131535.0 9835.0 131600.0 ;
      RECT  9770.0 131580.0 9835.0 131600.0 ;
      RECT  9802.5 131547.5 10100.0 131612.5 ;
      RECT  10100.0 131547.5 10235.0 131612.5 ;
      RECT  10805.0 131547.5 10870.0 131612.5 ;
      RECT  10805.0 131535.0 10870.0 131600.0 ;
      RECT  10587.5 131547.5 10837.5 131612.5 ;
      RECT  10805.0 131567.5 10870.0 131580.0 ;
      RECT  10837.5 131535.0 11085.0 131600.0 ;
      RECT  9255.0 132970.0 9605.0 133035.0 ;
      RECT  9770.0 132957.5 9835.0 133022.5 ;
      RECT  9770.0 132970.0 9835.0 133035.0 ;
      RECT  9770.0 132990.0 9835.0 133035.0 ;
      RECT  9802.5 132957.5 10100.0 133022.5 ;
      RECT  10100.0 132957.5 10235.0 133022.5 ;
      RECT  10805.0 132957.5 10870.0 133022.5 ;
      RECT  10805.0 132970.0 10870.0 133035.0 ;
      RECT  10587.5 132957.5 10837.5 133022.5 ;
      RECT  10805.0 132990.0 10870.0 133002.5 ;
      RECT  10837.5 132970.0 11085.0 133035.0 ;
      RECT  9255.0 134225.0 9605.0 134290.0 ;
      RECT  9770.0 134237.5 9835.0 134302.5 ;
      RECT  9770.0 134225.0 9835.0 134290.0 ;
      RECT  9770.0 134270.0 9835.0 134290.0 ;
      RECT  9802.5 134237.5 10100.0 134302.5 ;
      RECT  10100.0 134237.5 10235.0 134302.5 ;
      RECT  10805.0 134237.5 10870.0 134302.5 ;
      RECT  10805.0 134225.0 10870.0 134290.0 ;
      RECT  10587.5 134237.5 10837.5 134302.5 ;
      RECT  10805.0 134257.5 10870.0 134270.0 ;
      RECT  10837.5 134225.0 11085.0 134290.0 ;
      RECT  9255.0 135660.0 9605.0 135725.0 ;
      RECT  9770.0 135647.5 9835.0 135712.5 ;
      RECT  9770.0 135660.0 9835.0 135725.0 ;
      RECT  9770.0 135680.0 9835.0 135725.0 ;
      RECT  9802.5 135647.5 10100.0 135712.5 ;
      RECT  10100.0 135647.5 10235.0 135712.5 ;
      RECT  10805.0 135647.5 10870.0 135712.5 ;
      RECT  10805.0 135660.0 10870.0 135725.0 ;
      RECT  10587.5 135647.5 10837.5 135712.5 ;
      RECT  10805.0 135680.0 10870.0 135692.5 ;
      RECT  10837.5 135660.0 11085.0 135725.0 ;
      RECT  9255.0 136915.0 9605.0 136980.0 ;
      RECT  9770.0 136927.5 9835.0 136992.5 ;
      RECT  9770.0 136915.0 9835.0 136980.0 ;
      RECT  9770.0 136960.0 9835.0 136980.0 ;
      RECT  9802.5 136927.5 10100.0 136992.5 ;
      RECT  10100.0 136927.5 10235.0 136992.5 ;
      RECT  10805.0 136927.5 10870.0 136992.5 ;
      RECT  10805.0 136915.0 10870.0 136980.0 ;
      RECT  10587.5 136927.5 10837.5 136992.5 ;
      RECT  10805.0 136947.5 10870.0 136960.0 ;
      RECT  10837.5 136915.0 11085.0 136980.0 ;
      RECT  9255.0 138350.0 9605.0 138415.0 ;
      RECT  9770.0 138337.5 9835.0 138402.5 ;
      RECT  9770.0 138350.0 9835.0 138415.0 ;
      RECT  9770.0 138370.0 9835.0 138415.0 ;
      RECT  9802.5 138337.5 10100.0 138402.5 ;
      RECT  10100.0 138337.5 10235.0 138402.5 ;
      RECT  10805.0 138337.5 10870.0 138402.5 ;
      RECT  10805.0 138350.0 10870.0 138415.0 ;
      RECT  10587.5 138337.5 10837.5 138402.5 ;
      RECT  10805.0 138370.0 10870.0 138382.5 ;
      RECT  10837.5 138350.0 11085.0 138415.0 ;
      RECT  9255.0 139605.0 9605.0 139670.0 ;
      RECT  9770.0 139617.5 9835.0 139682.5 ;
      RECT  9770.0 139605.0 9835.0 139670.0 ;
      RECT  9770.0 139650.0 9835.0 139670.0 ;
      RECT  9802.5 139617.5 10100.0 139682.5 ;
      RECT  10100.0 139617.5 10235.0 139682.5 ;
      RECT  10805.0 139617.5 10870.0 139682.5 ;
      RECT  10805.0 139605.0 10870.0 139670.0 ;
      RECT  10587.5 139617.5 10837.5 139682.5 ;
      RECT  10805.0 139637.5 10870.0 139650.0 ;
      RECT  10837.5 139605.0 11085.0 139670.0 ;
      RECT  9255.0 141040.0 9605.0 141105.0 ;
      RECT  9770.0 141027.5 9835.0 141092.5 ;
      RECT  9770.0 141040.0 9835.0 141105.0 ;
      RECT  9770.0 141060.0 9835.0 141105.0 ;
      RECT  9802.5 141027.5 10100.0 141092.5 ;
      RECT  10100.0 141027.5 10235.0 141092.5 ;
      RECT  10805.0 141027.5 10870.0 141092.5 ;
      RECT  10805.0 141040.0 10870.0 141105.0 ;
      RECT  10587.5 141027.5 10837.5 141092.5 ;
      RECT  10805.0 141060.0 10870.0 141072.5 ;
      RECT  10837.5 141040.0 11085.0 141105.0 ;
      RECT  9255.0 142295.0 9605.0 142360.0 ;
      RECT  9770.0 142307.5 9835.0 142372.5 ;
      RECT  9770.0 142295.0 9835.0 142360.0 ;
      RECT  9770.0 142340.0 9835.0 142360.0 ;
      RECT  9802.5 142307.5 10100.0 142372.5 ;
      RECT  10100.0 142307.5 10235.0 142372.5 ;
      RECT  10805.0 142307.5 10870.0 142372.5 ;
      RECT  10805.0 142295.0 10870.0 142360.0 ;
      RECT  10587.5 142307.5 10837.5 142372.5 ;
      RECT  10805.0 142327.5 10870.0 142340.0 ;
      RECT  10837.5 142295.0 11085.0 142360.0 ;
      RECT  9255.0 143730.0 9605.0 143795.0 ;
      RECT  9770.0 143717.5 9835.0 143782.5 ;
      RECT  9770.0 143730.0 9835.0 143795.0 ;
      RECT  9770.0 143750.0 9835.0 143795.0 ;
      RECT  9802.5 143717.5 10100.0 143782.5 ;
      RECT  10100.0 143717.5 10235.0 143782.5 ;
      RECT  10805.0 143717.5 10870.0 143782.5 ;
      RECT  10805.0 143730.0 10870.0 143795.0 ;
      RECT  10587.5 143717.5 10837.5 143782.5 ;
      RECT  10805.0 143750.0 10870.0 143762.5 ;
      RECT  10837.5 143730.0 11085.0 143795.0 ;
      RECT  9255.0 144985.0 9605.0 145050.0 ;
      RECT  9770.0 144997.5 9835.0 145062.5 ;
      RECT  9770.0 144985.0 9835.0 145050.0 ;
      RECT  9770.0 145030.0 9835.0 145050.0 ;
      RECT  9802.5 144997.5 10100.0 145062.5 ;
      RECT  10100.0 144997.5 10235.0 145062.5 ;
      RECT  10805.0 144997.5 10870.0 145062.5 ;
      RECT  10805.0 144985.0 10870.0 145050.0 ;
      RECT  10587.5 144997.5 10837.5 145062.5 ;
      RECT  10805.0 145017.5 10870.0 145030.0 ;
      RECT  10837.5 144985.0 11085.0 145050.0 ;
      RECT  9255.0 146420.0 9605.0 146485.0 ;
      RECT  9770.0 146407.5 9835.0 146472.5 ;
      RECT  9770.0 146420.0 9835.0 146485.0 ;
      RECT  9770.0 146440.0 9835.0 146485.0 ;
      RECT  9802.5 146407.5 10100.0 146472.5 ;
      RECT  10100.0 146407.5 10235.0 146472.5 ;
      RECT  10805.0 146407.5 10870.0 146472.5 ;
      RECT  10805.0 146420.0 10870.0 146485.0 ;
      RECT  10587.5 146407.5 10837.5 146472.5 ;
      RECT  10805.0 146440.0 10870.0 146452.5 ;
      RECT  10837.5 146420.0 11085.0 146485.0 ;
      RECT  9255.0 147675.0 9605.0 147740.0 ;
      RECT  9770.0 147687.5 9835.0 147752.5 ;
      RECT  9770.0 147675.0 9835.0 147740.0 ;
      RECT  9770.0 147720.0 9835.0 147740.0 ;
      RECT  9802.5 147687.5 10100.0 147752.5 ;
      RECT  10100.0 147687.5 10235.0 147752.5 ;
      RECT  10805.0 147687.5 10870.0 147752.5 ;
      RECT  10805.0 147675.0 10870.0 147740.0 ;
      RECT  10587.5 147687.5 10837.5 147752.5 ;
      RECT  10805.0 147707.5 10870.0 147720.0 ;
      RECT  10837.5 147675.0 11085.0 147740.0 ;
      RECT  9255.0 149110.0 9605.0 149175.0 ;
      RECT  9770.0 149097.5 9835.0 149162.5 ;
      RECT  9770.0 149110.0 9835.0 149175.0 ;
      RECT  9770.0 149130.0 9835.0 149175.0 ;
      RECT  9802.5 149097.5 10100.0 149162.5 ;
      RECT  10100.0 149097.5 10235.0 149162.5 ;
      RECT  10805.0 149097.5 10870.0 149162.5 ;
      RECT  10805.0 149110.0 10870.0 149175.0 ;
      RECT  10587.5 149097.5 10837.5 149162.5 ;
      RECT  10805.0 149130.0 10870.0 149142.5 ;
      RECT  10837.5 149110.0 11085.0 149175.0 ;
      RECT  9255.0 150365.0 9605.0 150430.0 ;
      RECT  9770.0 150377.5 9835.0 150442.5 ;
      RECT  9770.0 150365.0 9835.0 150430.0 ;
      RECT  9770.0 150410.0 9835.0 150430.0 ;
      RECT  9802.5 150377.5 10100.0 150442.5 ;
      RECT  10100.0 150377.5 10235.0 150442.5 ;
      RECT  10805.0 150377.5 10870.0 150442.5 ;
      RECT  10805.0 150365.0 10870.0 150430.0 ;
      RECT  10587.5 150377.5 10837.5 150442.5 ;
      RECT  10805.0 150397.5 10870.0 150410.0 ;
      RECT  10837.5 150365.0 11085.0 150430.0 ;
      RECT  9255.0 151800.0 9605.0 151865.0 ;
      RECT  9770.0 151787.5 9835.0 151852.5 ;
      RECT  9770.0 151800.0 9835.0 151865.0 ;
      RECT  9770.0 151820.0 9835.0 151865.0 ;
      RECT  9802.5 151787.5 10100.0 151852.5 ;
      RECT  10100.0 151787.5 10235.0 151852.5 ;
      RECT  10805.0 151787.5 10870.0 151852.5 ;
      RECT  10805.0 151800.0 10870.0 151865.0 ;
      RECT  10587.5 151787.5 10837.5 151852.5 ;
      RECT  10805.0 151820.0 10870.0 151832.5 ;
      RECT  10837.5 151800.0 11085.0 151865.0 ;
      RECT  9255.0 153055.0 9605.0 153120.0 ;
      RECT  9770.0 153067.5 9835.0 153132.5 ;
      RECT  9770.0 153055.0 9835.0 153120.0 ;
      RECT  9770.0 153100.0 9835.0 153120.0 ;
      RECT  9802.5 153067.5 10100.0 153132.5 ;
      RECT  10100.0 153067.5 10235.0 153132.5 ;
      RECT  10805.0 153067.5 10870.0 153132.5 ;
      RECT  10805.0 153055.0 10870.0 153120.0 ;
      RECT  10587.5 153067.5 10837.5 153132.5 ;
      RECT  10805.0 153087.5 10870.0 153100.0 ;
      RECT  10837.5 153055.0 11085.0 153120.0 ;
      RECT  9255.0 154490.0 9605.0 154555.0 ;
      RECT  9770.0 154477.5 9835.0 154542.5 ;
      RECT  9770.0 154490.0 9835.0 154555.0 ;
      RECT  9770.0 154510.0 9835.0 154555.0 ;
      RECT  9802.5 154477.5 10100.0 154542.5 ;
      RECT  10100.0 154477.5 10235.0 154542.5 ;
      RECT  10805.0 154477.5 10870.0 154542.5 ;
      RECT  10805.0 154490.0 10870.0 154555.0 ;
      RECT  10587.5 154477.5 10837.5 154542.5 ;
      RECT  10805.0 154510.0 10870.0 154522.5 ;
      RECT  10837.5 154490.0 11085.0 154555.0 ;
      RECT  9255.0 155745.0 9605.0 155810.0 ;
      RECT  9770.0 155757.5 9835.0 155822.5 ;
      RECT  9770.0 155745.0 9835.0 155810.0 ;
      RECT  9770.0 155790.0 9835.0 155810.0 ;
      RECT  9802.5 155757.5 10100.0 155822.5 ;
      RECT  10100.0 155757.5 10235.0 155822.5 ;
      RECT  10805.0 155757.5 10870.0 155822.5 ;
      RECT  10805.0 155745.0 10870.0 155810.0 ;
      RECT  10587.5 155757.5 10837.5 155822.5 ;
      RECT  10805.0 155777.5 10870.0 155790.0 ;
      RECT  10837.5 155745.0 11085.0 155810.0 ;
      RECT  9255.0 157180.0 9605.0 157245.0 ;
      RECT  9770.0 157167.5 9835.0 157232.5 ;
      RECT  9770.0 157180.0 9835.0 157245.0 ;
      RECT  9770.0 157200.0 9835.0 157245.0 ;
      RECT  9802.5 157167.5 10100.0 157232.5 ;
      RECT  10100.0 157167.5 10235.0 157232.5 ;
      RECT  10805.0 157167.5 10870.0 157232.5 ;
      RECT  10805.0 157180.0 10870.0 157245.0 ;
      RECT  10587.5 157167.5 10837.5 157232.5 ;
      RECT  10805.0 157200.0 10870.0 157212.5 ;
      RECT  10837.5 157180.0 11085.0 157245.0 ;
      RECT  9255.0 158435.0 9605.0 158500.0 ;
      RECT  9770.0 158447.5 9835.0 158512.5 ;
      RECT  9770.0 158435.0 9835.0 158500.0 ;
      RECT  9770.0 158480.0 9835.0 158500.0 ;
      RECT  9802.5 158447.5 10100.0 158512.5 ;
      RECT  10100.0 158447.5 10235.0 158512.5 ;
      RECT  10805.0 158447.5 10870.0 158512.5 ;
      RECT  10805.0 158435.0 10870.0 158500.0 ;
      RECT  10587.5 158447.5 10837.5 158512.5 ;
      RECT  10805.0 158467.5 10870.0 158480.0 ;
      RECT  10837.5 158435.0 11085.0 158500.0 ;
      RECT  9255.0 159870.0 9605.0 159935.0 ;
      RECT  9770.0 159857.5 9835.0 159922.5 ;
      RECT  9770.0 159870.0 9835.0 159935.0 ;
      RECT  9770.0 159890.0 9835.0 159935.0 ;
      RECT  9802.5 159857.5 10100.0 159922.5 ;
      RECT  10100.0 159857.5 10235.0 159922.5 ;
      RECT  10805.0 159857.5 10870.0 159922.5 ;
      RECT  10805.0 159870.0 10870.0 159935.0 ;
      RECT  10587.5 159857.5 10837.5 159922.5 ;
      RECT  10805.0 159890.0 10870.0 159902.5 ;
      RECT  10837.5 159870.0 11085.0 159935.0 ;
      RECT  9255.0 161125.0 9605.0 161190.0 ;
      RECT  9770.0 161137.5 9835.0 161202.5 ;
      RECT  9770.0 161125.0 9835.0 161190.0 ;
      RECT  9770.0 161170.0 9835.0 161190.0 ;
      RECT  9802.5 161137.5 10100.0 161202.5 ;
      RECT  10100.0 161137.5 10235.0 161202.5 ;
      RECT  10805.0 161137.5 10870.0 161202.5 ;
      RECT  10805.0 161125.0 10870.0 161190.0 ;
      RECT  10587.5 161137.5 10837.5 161202.5 ;
      RECT  10805.0 161157.5 10870.0 161170.0 ;
      RECT  10837.5 161125.0 11085.0 161190.0 ;
      RECT  9255.0 162560.0 9605.0 162625.0 ;
      RECT  9770.0 162547.5 9835.0 162612.5 ;
      RECT  9770.0 162560.0 9835.0 162625.0 ;
      RECT  9770.0 162580.0 9835.0 162625.0 ;
      RECT  9802.5 162547.5 10100.0 162612.5 ;
      RECT  10100.0 162547.5 10235.0 162612.5 ;
      RECT  10805.0 162547.5 10870.0 162612.5 ;
      RECT  10805.0 162560.0 10870.0 162625.0 ;
      RECT  10587.5 162547.5 10837.5 162612.5 ;
      RECT  10805.0 162580.0 10870.0 162592.5 ;
      RECT  10837.5 162560.0 11085.0 162625.0 ;
      RECT  9255.0 163815.0 9605.0 163880.0 ;
      RECT  9770.0 163827.5 9835.0 163892.5 ;
      RECT  9770.0 163815.0 9835.0 163880.0 ;
      RECT  9770.0 163860.0 9835.0 163880.0 ;
      RECT  9802.5 163827.5 10100.0 163892.5 ;
      RECT  10100.0 163827.5 10235.0 163892.5 ;
      RECT  10805.0 163827.5 10870.0 163892.5 ;
      RECT  10805.0 163815.0 10870.0 163880.0 ;
      RECT  10587.5 163827.5 10837.5 163892.5 ;
      RECT  10805.0 163847.5 10870.0 163860.0 ;
      RECT  10837.5 163815.0 11085.0 163880.0 ;
      RECT  9255.0 165250.0 9605.0 165315.0 ;
      RECT  9770.0 165237.5 9835.0 165302.5 ;
      RECT  9770.0 165250.0 9835.0 165315.0 ;
      RECT  9770.0 165270.0 9835.0 165315.0 ;
      RECT  9802.5 165237.5 10100.0 165302.5 ;
      RECT  10100.0 165237.5 10235.0 165302.5 ;
      RECT  10805.0 165237.5 10870.0 165302.5 ;
      RECT  10805.0 165250.0 10870.0 165315.0 ;
      RECT  10587.5 165237.5 10837.5 165302.5 ;
      RECT  10805.0 165270.0 10870.0 165282.5 ;
      RECT  10837.5 165250.0 11085.0 165315.0 ;
      RECT  9255.0 166505.0 9605.0 166570.0 ;
      RECT  9770.0 166517.5 9835.0 166582.5 ;
      RECT  9770.0 166505.0 9835.0 166570.0 ;
      RECT  9770.0 166550.0 9835.0 166570.0 ;
      RECT  9802.5 166517.5 10100.0 166582.5 ;
      RECT  10100.0 166517.5 10235.0 166582.5 ;
      RECT  10805.0 166517.5 10870.0 166582.5 ;
      RECT  10805.0 166505.0 10870.0 166570.0 ;
      RECT  10587.5 166517.5 10837.5 166582.5 ;
      RECT  10805.0 166537.5 10870.0 166550.0 ;
      RECT  10837.5 166505.0 11085.0 166570.0 ;
      RECT  9255.0 167940.0 9605.0 168005.0 ;
      RECT  9770.0 167927.5 9835.0 167992.5 ;
      RECT  9770.0 167940.0 9835.0 168005.0 ;
      RECT  9770.0 167960.0 9835.0 168005.0 ;
      RECT  9802.5 167927.5 10100.0 167992.5 ;
      RECT  10100.0 167927.5 10235.0 167992.5 ;
      RECT  10805.0 167927.5 10870.0 167992.5 ;
      RECT  10805.0 167940.0 10870.0 168005.0 ;
      RECT  10587.5 167927.5 10837.5 167992.5 ;
      RECT  10805.0 167960.0 10870.0 167972.5 ;
      RECT  10837.5 167940.0 11085.0 168005.0 ;
      RECT  9255.0 169195.0 9605.0 169260.0 ;
      RECT  9770.0 169207.5 9835.0 169272.5 ;
      RECT  9770.0 169195.0 9835.0 169260.0 ;
      RECT  9770.0 169240.0 9835.0 169260.0 ;
      RECT  9802.5 169207.5 10100.0 169272.5 ;
      RECT  10100.0 169207.5 10235.0 169272.5 ;
      RECT  10805.0 169207.5 10870.0 169272.5 ;
      RECT  10805.0 169195.0 10870.0 169260.0 ;
      RECT  10587.5 169207.5 10837.5 169272.5 ;
      RECT  10805.0 169227.5 10870.0 169240.0 ;
      RECT  10837.5 169195.0 11085.0 169260.0 ;
      RECT  9255.0 170630.0 9605.0 170695.0 ;
      RECT  9770.0 170617.5 9835.0 170682.5 ;
      RECT  9770.0 170630.0 9835.0 170695.0 ;
      RECT  9770.0 170650.0 9835.0 170695.0 ;
      RECT  9802.5 170617.5 10100.0 170682.5 ;
      RECT  10100.0 170617.5 10235.0 170682.5 ;
      RECT  10805.0 170617.5 10870.0 170682.5 ;
      RECT  10805.0 170630.0 10870.0 170695.0 ;
      RECT  10587.5 170617.5 10837.5 170682.5 ;
      RECT  10805.0 170650.0 10870.0 170662.5 ;
      RECT  10837.5 170630.0 11085.0 170695.0 ;
      RECT  9255.0 171885.0 9605.0 171950.0 ;
      RECT  9770.0 171897.5 9835.0 171962.5 ;
      RECT  9770.0 171885.0 9835.0 171950.0 ;
      RECT  9770.0 171930.0 9835.0 171950.0 ;
      RECT  9802.5 171897.5 10100.0 171962.5 ;
      RECT  10100.0 171897.5 10235.0 171962.5 ;
      RECT  10805.0 171897.5 10870.0 171962.5 ;
      RECT  10805.0 171885.0 10870.0 171950.0 ;
      RECT  10587.5 171897.5 10837.5 171962.5 ;
      RECT  10805.0 171917.5 10870.0 171930.0 ;
      RECT  10837.5 171885.0 11085.0 171950.0 ;
      RECT  9255.0 173320.0 9605.0 173385.0 ;
      RECT  9770.0 173307.5 9835.0 173372.5 ;
      RECT  9770.0 173320.0 9835.0 173385.0 ;
      RECT  9770.0 173340.0 9835.0 173385.0 ;
      RECT  9802.5 173307.5 10100.0 173372.5 ;
      RECT  10100.0 173307.5 10235.0 173372.5 ;
      RECT  10805.0 173307.5 10870.0 173372.5 ;
      RECT  10805.0 173320.0 10870.0 173385.0 ;
      RECT  10587.5 173307.5 10837.5 173372.5 ;
      RECT  10805.0 173340.0 10870.0 173352.5 ;
      RECT  10837.5 173320.0 11085.0 173385.0 ;
      RECT  9255.0 174575.0 9605.0 174640.0 ;
      RECT  9770.0 174587.5 9835.0 174652.5 ;
      RECT  9770.0 174575.0 9835.0 174640.0 ;
      RECT  9770.0 174620.0 9835.0 174640.0 ;
      RECT  9802.5 174587.5 10100.0 174652.5 ;
      RECT  10100.0 174587.5 10235.0 174652.5 ;
      RECT  10805.0 174587.5 10870.0 174652.5 ;
      RECT  10805.0 174575.0 10870.0 174640.0 ;
      RECT  10587.5 174587.5 10837.5 174652.5 ;
      RECT  10805.0 174607.5 10870.0 174620.0 ;
      RECT  10837.5 174575.0 11085.0 174640.0 ;
      RECT  9255.0 176010.0 9605.0 176075.0 ;
      RECT  9770.0 175997.5 9835.0 176062.5 ;
      RECT  9770.0 176010.0 9835.0 176075.0 ;
      RECT  9770.0 176030.0 9835.0 176075.0 ;
      RECT  9802.5 175997.5 10100.0 176062.5 ;
      RECT  10100.0 175997.5 10235.0 176062.5 ;
      RECT  10805.0 175997.5 10870.0 176062.5 ;
      RECT  10805.0 176010.0 10870.0 176075.0 ;
      RECT  10587.5 175997.5 10837.5 176062.5 ;
      RECT  10805.0 176030.0 10870.0 176042.5 ;
      RECT  10837.5 176010.0 11085.0 176075.0 ;
      RECT  9255.0 177265.0 9605.0 177330.0 ;
      RECT  9770.0 177277.5 9835.0 177342.5 ;
      RECT  9770.0 177265.0 9835.0 177330.0 ;
      RECT  9770.0 177310.0 9835.0 177330.0 ;
      RECT  9802.5 177277.5 10100.0 177342.5 ;
      RECT  10100.0 177277.5 10235.0 177342.5 ;
      RECT  10805.0 177277.5 10870.0 177342.5 ;
      RECT  10805.0 177265.0 10870.0 177330.0 ;
      RECT  10587.5 177277.5 10837.5 177342.5 ;
      RECT  10805.0 177297.5 10870.0 177310.0 ;
      RECT  10837.5 177265.0 11085.0 177330.0 ;
      RECT  9255.0 178700.0 9605.0 178765.0 ;
      RECT  9770.0 178687.5 9835.0 178752.5 ;
      RECT  9770.0 178700.0 9835.0 178765.0 ;
      RECT  9770.0 178720.0 9835.0 178765.0 ;
      RECT  9802.5 178687.5 10100.0 178752.5 ;
      RECT  10100.0 178687.5 10235.0 178752.5 ;
      RECT  10805.0 178687.5 10870.0 178752.5 ;
      RECT  10805.0 178700.0 10870.0 178765.0 ;
      RECT  10587.5 178687.5 10837.5 178752.5 ;
      RECT  10805.0 178720.0 10870.0 178732.5 ;
      RECT  10837.5 178700.0 11085.0 178765.0 ;
      RECT  9255.0 179955.0 9605.0 180020.0 ;
      RECT  9770.0 179967.5 9835.0 180032.5 ;
      RECT  9770.0 179955.0 9835.0 180020.0 ;
      RECT  9770.0 180000.0 9835.0 180020.0 ;
      RECT  9802.5 179967.5 10100.0 180032.5 ;
      RECT  10100.0 179967.5 10235.0 180032.5 ;
      RECT  10805.0 179967.5 10870.0 180032.5 ;
      RECT  10805.0 179955.0 10870.0 180020.0 ;
      RECT  10587.5 179967.5 10837.5 180032.5 ;
      RECT  10805.0 179987.5 10870.0 180000.0 ;
      RECT  10837.5 179955.0 11085.0 180020.0 ;
      RECT  9255.0 181390.0 9605.0 181455.0 ;
      RECT  9770.0 181377.5 9835.0 181442.5 ;
      RECT  9770.0 181390.0 9835.0 181455.0 ;
      RECT  9770.0 181410.0 9835.0 181455.0 ;
      RECT  9802.5 181377.5 10100.0 181442.5 ;
      RECT  10100.0 181377.5 10235.0 181442.5 ;
      RECT  10805.0 181377.5 10870.0 181442.5 ;
      RECT  10805.0 181390.0 10870.0 181455.0 ;
      RECT  10587.5 181377.5 10837.5 181442.5 ;
      RECT  10805.0 181410.0 10870.0 181422.5 ;
      RECT  10837.5 181390.0 11085.0 181455.0 ;
      RECT  9255.0 182645.0 9605.0 182710.0 ;
      RECT  9770.0 182657.5 9835.0 182722.5 ;
      RECT  9770.0 182645.0 9835.0 182710.0 ;
      RECT  9770.0 182690.0 9835.0 182710.0 ;
      RECT  9802.5 182657.5 10100.0 182722.5 ;
      RECT  10100.0 182657.5 10235.0 182722.5 ;
      RECT  10805.0 182657.5 10870.0 182722.5 ;
      RECT  10805.0 182645.0 10870.0 182710.0 ;
      RECT  10587.5 182657.5 10837.5 182722.5 ;
      RECT  10805.0 182677.5 10870.0 182690.0 ;
      RECT  10837.5 182645.0 11085.0 182710.0 ;
      RECT  9255.0 184080.0 9605.0 184145.0 ;
      RECT  9770.0 184067.5 9835.0 184132.5 ;
      RECT  9770.0 184080.0 9835.0 184145.0 ;
      RECT  9770.0 184100.0 9835.0 184145.0 ;
      RECT  9802.5 184067.5 10100.0 184132.5 ;
      RECT  10100.0 184067.5 10235.0 184132.5 ;
      RECT  10805.0 184067.5 10870.0 184132.5 ;
      RECT  10805.0 184080.0 10870.0 184145.0 ;
      RECT  10587.5 184067.5 10837.5 184132.5 ;
      RECT  10805.0 184100.0 10870.0 184112.5 ;
      RECT  10837.5 184080.0 11085.0 184145.0 ;
      RECT  9255.0 185335.0 9605.0 185400.0 ;
      RECT  9770.0 185347.5 9835.0 185412.5 ;
      RECT  9770.0 185335.0 9835.0 185400.0 ;
      RECT  9770.0 185380.0 9835.0 185400.0 ;
      RECT  9802.5 185347.5 10100.0 185412.5 ;
      RECT  10100.0 185347.5 10235.0 185412.5 ;
      RECT  10805.0 185347.5 10870.0 185412.5 ;
      RECT  10805.0 185335.0 10870.0 185400.0 ;
      RECT  10587.5 185347.5 10837.5 185412.5 ;
      RECT  10805.0 185367.5 10870.0 185380.0 ;
      RECT  10837.5 185335.0 11085.0 185400.0 ;
      RECT  9255.0 186770.0 9605.0 186835.0 ;
      RECT  9770.0 186757.5 9835.0 186822.5 ;
      RECT  9770.0 186770.0 9835.0 186835.0 ;
      RECT  9770.0 186790.0 9835.0 186835.0 ;
      RECT  9802.5 186757.5 10100.0 186822.5 ;
      RECT  10100.0 186757.5 10235.0 186822.5 ;
      RECT  10805.0 186757.5 10870.0 186822.5 ;
      RECT  10805.0 186770.0 10870.0 186835.0 ;
      RECT  10587.5 186757.5 10837.5 186822.5 ;
      RECT  10805.0 186790.0 10870.0 186802.5 ;
      RECT  10837.5 186770.0 11085.0 186835.0 ;
      RECT  9255.0 188025.0 9605.0 188090.0 ;
      RECT  9770.0 188037.5 9835.0 188102.5 ;
      RECT  9770.0 188025.0 9835.0 188090.0 ;
      RECT  9770.0 188070.0 9835.0 188090.0 ;
      RECT  9802.5 188037.5 10100.0 188102.5 ;
      RECT  10100.0 188037.5 10235.0 188102.5 ;
      RECT  10805.0 188037.5 10870.0 188102.5 ;
      RECT  10805.0 188025.0 10870.0 188090.0 ;
      RECT  10587.5 188037.5 10837.5 188102.5 ;
      RECT  10805.0 188057.5 10870.0 188070.0 ;
      RECT  10837.5 188025.0 11085.0 188090.0 ;
      RECT  9255.0 189460.0 9605.0 189525.0 ;
      RECT  9770.0 189447.5 9835.0 189512.5 ;
      RECT  9770.0 189460.0 9835.0 189525.0 ;
      RECT  9770.0 189480.0 9835.0 189525.0 ;
      RECT  9802.5 189447.5 10100.0 189512.5 ;
      RECT  10100.0 189447.5 10235.0 189512.5 ;
      RECT  10805.0 189447.5 10870.0 189512.5 ;
      RECT  10805.0 189460.0 10870.0 189525.0 ;
      RECT  10587.5 189447.5 10837.5 189512.5 ;
      RECT  10805.0 189480.0 10870.0 189492.5 ;
      RECT  10837.5 189460.0 11085.0 189525.0 ;
      RECT  9255.0 190715.0 9605.0 190780.0 ;
      RECT  9770.0 190727.5 9835.0 190792.5 ;
      RECT  9770.0 190715.0 9835.0 190780.0 ;
      RECT  9770.0 190760.0 9835.0 190780.0 ;
      RECT  9802.5 190727.5 10100.0 190792.5 ;
      RECT  10100.0 190727.5 10235.0 190792.5 ;
      RECT  10805.0 190727.5 10870.0 190792.5 ;
      RECT  10805.0 190715.0 10870.0 190780.0 ;
      RECT  10587.5 190727.5 10837.5 190792.5 ;
      RECT  10805.0 190747.5 10870.0 190760.0 ;
      RECT  10837.5 190715.0 11085.0 190780.0 ;
      RECT  9255.0 192150.0 9605.0 192215.0 ;
      RECT  9770.0 192137.5 9835.0 192202.5 ;
      RECT  9770.0 192150.0 9835.0 192215.0 ;
      RECT  9770.0 192170.0 9835.0 192215.0 ;
      RECT  9802.5 192137.5 10100.0 192202.5 ;
      RECT  10100.0 192137.5 10235.0 192202.5 ;
      RECT  10805.0 192137.5 10870.0 192202.5 ;
      RECT  10805.0 192150.0 10870.0 192215.0 ;
      RECT  10587.5 192137.5 10837.5 192202.5 ;
      RECT  10805.0 192170.0 10870.0 192182.5 ;
      RECT  10837.5 192150.0 11085.0 192215.0 ;
      RECT  9255.0 193405.0 9605.0 193470.0 ;
      RECT  9770.0 193417.5 9835.0 193482.5 ;
      RECT  9770.0 193405.0 9835.0 193470.0 ;
      RECT  9770.0 193450.0 9835.0 193470.0 ;
      RECT  9802.5 193417.5 10100.0 193482.5 ;
      RECT  10100.0 193417.5 10235.0 193482.5 ;
      RECT  10805.0 193417.5 10870.0 193482.5 ;
      RECT  10805.0 193405.0 10870.0 193470.0 ;
      RECT  10587.5 193417.5 10837.5 193482.5 ;
      RECT  10805.0 193437.5 10870.0 193450.0 ;
      RECT  10837.5 193405.0 11085.0 193470.0 ;
      RECT  9255.0 194840.0 9605.0 194905.0 ;
      RECT  9770.0 194827.5 9835.0 194892.5 ;
      RECT  9770.0 194840.0 9835.0 194905.0 ;
      RECT  9770.0 194860.0 9835.0 194905.0 ;
      RECT  9802.5 194827.5 10100.0 194892.5 ;
      RECT  10100.0 194827.5 10235.0 194892.5 ;
      RECT  10805.0 194827.5 10870.0 194892.5 ;
      RECT  10805.0 194840.0 10870.0 194905.0 ;
      RECT  10587.5 194827.5 10837.5 194892.5 ;
      RECT  10805.0 194860.0 10870.0 194872.5 ;
      RECT  10837.5 194840.0 11085.0 194905.0 ;
      RECT  9255.0 196095.0 9605.0 196160.0 ;
      RECT  9770.0 196107.5 9835.0 196172.5 ;
      RECT  9770.0 196095.0 9835.0 196160.0 ;
      RECT  9770.0 196140.0 9835.0 196160.0 ;
      RECT  9802.5 196107.5 10100.0 196172.5 ;
      RECT  10100.0 196107.5 10235.0 196172.5 ;
      RECT  10805.0 196107.5 10870.0 196172.5 ;
      RECT  10805.0 196095.0 10870.0 196160.0 ;
      RECT  10587.5 196107.5 10837.5 196172.5 ;
      RECT  10805.0 196127.5 10870.0 196140.0 ;
      RECT  10837.5 196095.0 11085.0 196160.0 ;
      RECT  9255.0 197530.0 9605.0 197595.0 ;
      RECT  9770.0 197517.5 9835.0 197582.5 ;
      RECT  9770.0 197530.0 9835.0 197595.0 ;
      RECT  9770.0 197550.0 9835.0 197595.0 ;
      RECT  9802.5 197517.5 10100.0 197582.5 ;
      RECT  10100.0 197517.5 10235.0 197582.5 ;
      RECT  10805.0 197517.5 10870.0 197582.5 ;
      RECT  10805.0 197530.0 10870.0 197595.0 ;
      RECT  10587.5 197517.5 10837.5 197582.5 ;
      RECT  10805.0 197550.0 10870.0 197562.5 ;
      RECT  10837.5 197530.0 11085.0 197595.0 ;
      RECT  9255.0 198785.0 9605.0 198850.0 ;
      RECT  9770.0 198797.5 9835.0 198862.5 ;
      RECT  9770.0 198785.0 9835.0 198850.0 ;
      RECT  9770.0 198830.0 9835.0 198850.0 ;
      RECT  9802.5 198797.5 10100.0 198862.5 ;
      RECT  10100.0 198797.5 10235.0 198862.5 ;
      RECT  10805.0 198797.5 10870.0 198862.5 ;
      RECT  10805.0 198785.0 10870.0 198850.0 ;
      RECT  10587.5 198797.5 10837.5 198862.5 ;
      RECT  10805.0 198817.5 10870.0 198830.0 ;
      RECT  10837.5 198785.0 11085.0 198850.0 ;
      RECT  9255.0 200220.0 9605.0 200285.0 ;
      RECT  9770.0 200207.5 9835.0 200272.5 ;
      RECT  9770.0 200220.0 9835.0 200285.0 ;
      RECT  9770.0 200240.0 9835.0 200285.0 ;
      RECT  9802.5 200207.5 10100.0 200272.5 ;
      RECT  10100.0 200207.5 10235.0 200272.5 ;
      RECT  10805.0 200207.5 10870.0 200272.5 ;
      RECT  10805.0 200220.0 10870.0 200285.0 ;
      RECT  10587.5 200207.5 10837.5 200272.5 ;
      RECT  10805.0 200240.0 10870.0 200252.5 ;
      RECT  10837.5 200220.0 11085.0 200285.0 ;
      RECT  9255.0 201475.0 9605.0 201540.0 ;
      RECT  9770.0 201487.5 9835.0 201552.5 ;
      RECT  9770.0 201475.0 9835.0 201540.0 ;
      RECT  9770.0 201520.0 9835.0 201540.0 ;
      RECT  9802.5 201487.5 10100.0 201552.5 ;
      RECT  10100.0 201487.5 10235.0 201552.5 ;
      RECT  10805.0 201487.5 10870.0 201552.5 ;
      RECT  10805.0 201475.0 10870.0 201540.0 ;
      RECT  10587.5 201487.5 10837.5 201552.5 ;
      RECT  10805.0 201507.5 10870.0 201520.0 ;
      RECT  10837.5 201475.0 11085.0 201540.0 ;
      RECT  9255.0 202910.0 9605.0 202975.0 ;
      RECT  9770.0 202897.5 9835.0 202962.5 ;
      RECT  9770.0 202910.0 9835.0 202975.0 ;
      RECT  9770.0 202930.0 9835.0 202975.0 ;
      RECT  9802.5 202897.5 10100.0 202962.5 ;
      RECT  10100.0 202897.5 10235.0 202962.5 ;
      RECT  10805.0 202897.5 10870.0 202962.5 ;
      RECT  10805.0 202910.0 10870.0 202975.0 ;
      RECT  10587.5 202897.5 10837.5 202962.5 ;
      RECT  10805.0 202930.0 10870.0 202942.5 ;
      RECT  10837.5 202910.0 11085.0 202975.0 ;
      RECT  9255.0 204165.0 9605.0 204230.0 ;
      RECT  9770.0 204177.5 9835.0 204242.5 ;
      RECT  9770.0 204165.0 9835.0 204230.0 ;
      RECT  9770.0 204210.0 9835.0 204230.0 ;
      RECT  9802.5 204177.5 10100.0 204242.5 ;
      RECT  10100.0 204177.5 10235.0 204242.5 ;
      RECT  10805.0 204177.5 10870.0 204242.5 ;
      RECT  10805.0 204165.0 10870.0 204230.0 ;
      RECT  10587.5 204177.5 10837.5 204242.5 ;
      RECT  10805.0 204197.5 10870.0 204210.0 ;
      RECT  10837.5 204165.0 11085.0 204230.0 ;
      RECT  9255.0 205600.0 9605.0 205665.0 ;
      RECT  9770.0 205587.5 9835.0 205652.5 ;
      RECT  9770.0 205600.0 9835.0 205665.0 ;
      RECT  9770.0 205620.0 9835.0 205665.0 ;
      RECT  9802.5 205587.5 10100.0 205652.5 ;
      RECT  10100.0 205587.5 10235.0 205652.5 ;
      RECT  10805.0 205587.5 10870.0 205652.5 ;
      RECT  10805.0 205600.0 10870.0 205665.0 ;
      RECT  10587.5 205587.5 10837.5 205652.5 ;
      RECT  10805.0 205620.0 10870.0 205632.5 ;
      RECT  10837.5 205600.0 11085.0 205665.0 ;
      RECT  9907.5 35260.0 9972.5 35445.0 ;
      RECT  9907.5 34100.0 9972.5 34285.0 ;
      RECT  9547.5 34217.5 9612.5 34067.5 ;
      RECT  9547.5 35102.5 9612.5 35477.5 ;
      RECT  9737.5 34217.5 9802.5 35102.5 ;
      RECT  9547.5 35102.5 9612.5 35237.5 ;
      RECT  9737.5 35102.5 9802.5 35237.5 ;
      RECT  9737.5 35102.5 9802.5 35237.5 ;
      RECT  9547.5 35102.5 9612.5 35237.5 ;
      RECT  9547.5 34217.5 9612.5 34352.5 ;
      RECT  9737.5 34217.5 9802.5 34352.5 ;
      RECT  9737.5 34217.5 9802.5 34352.5 ;
      RECT  9547.5 34217.5 9612.5 34352.5 ;
      RECT  9907.5 35192.5 9972.5 35327.5 ;
      RECT  9907.5 34217.5 9972.5 34352.5 ;
      RECT  9605.0 34660.0 9670.0 34795.0 ;
      RECT  9605.0 34660.0 9670.0 34795.0 ;
      RECT  9770.0 34695.0 9835.0 34760.0 ;
      RECT  9480.0 35412.5 10040.0 35477.5 ;
      RECT  9480.0 34067.5 10040.0 34132.5 ;
      RECT  10107.5 34262.5 10172.5 34067.5 ;
      RECT  10107.5 35102.5 10172.5 35477.5 ;
      RECT  10487.5 35102.5 10552.5 35477.5 ;
      RECT  10657.5 35260.0 10722.5 35445.0 ;
      RECT  10657.5 34100.0 10722.5 34285.0 ;
      RECT  10107.5 35102.5 10172.5 35237.5 ;
      RECT  10297.5 35102.5 10362.5 35237.5 ;
      RECT  10297.5 35102.5 10362.5 35237.5 ;
      RECT  10107.5 35102.5 10172.5 35237.5 ;
      RECT  10297.5 35102.5 10362.5 35237.5 ;
      RECT  10487.5 35102.5 10552.5 35237.5 ;
      RECT  10487.5 35102.5 10552.5 35237.5 ;
      RECT  10297.5 35102.5 10362.5 35237.5 ;
      RECT  10107.5 34262.5 10172.5 34397.5 ;
      RECT  10297.5 34262.5 10362.5 34397.5 ;
      RECT  10297.5 34262.5 10362.5 34397.5 ;
      RECT  10107.5 34262.5 10172.5 34397.5 ;
      RECT  10297.5 34262.5 10362.5 34397.5 ;
      RECT  10487.5 34262.5 10552.5 34397.5 ;
      RECT  10487.5 34262.5 10552.5 34397.5 ;
      RECT  10297.5 34262.5 10362.5 34397.5 ;
      RECT  10657.5 35192.5 10722.5 35327.5 ;
      RECT  10657.5 34217.5 10722.5 34352.5 ;
      RECT  10492.5 34492.5 10357.5 34557.5 ;
      RECT  10235.0 34707.5 10100.0 34772.5 ;
      RECT  10297.5 35102.5 10362.5 35237.5 ;
      RECT  10487.5 34262.5 10552.5 34397.5 ;
      RECT  10587.5 34707.5 10452.5 34772.5 ;
      RECT  10100.0 34707.5 10235.0 34772.5 ;
      RECT  10357.5 34492.5 10492.5 34557.5 ;
      RECT  10452.5 34707.5 10587.5 34772.5 ;
      RECT  10040.0 35412.5 10960.0 35477.5 ;
      RECT  10040.0 34067.5 10960.0 34132.5 ;
      RECT  11387.5 35260.0 11452.5 35445.0 ;
      RECT  11387.5 34100.0 11452.5 34285.0 ;
      RECT  11027.5 34217.5 11092.5 34067.5 ;
      RECT  11027.5 35102.5 11092.5 35477.5 ;
      RECT  11217.5 34217.5 11282.5 35102.5 ;
      RECT  11027.5 35102.5 11092.5 35237.5 ;
      RECT  11217.5 35102.5 11282.5 35237.5 ;
      RECT  11217.5 35102.5 11282.5 35237.5 ;
      RECT  11027.5 35102.5 11092.5 35237.5 ;
      RECT  11027.5 34217.5 11092.5 34352.5 ;
      RECT  11217.5 34217.5 11282.5 34352.5 ;
      RECT  11217.5 34217.5 11282.5 34352.5 ;
      RECT  11027.5 34217.5 11092.5 34352.5 ;
      RECT  11387.5 35192.5 11452.5 35327.5 ;
      RECT  11387.5 34217.5 11452.5 34352.5 ;
      RECT  11085.0 34660.0 11150.0 34795.0 ;
      RECT  11085.0 34660.0 11150.0 34795.0 ;
      RECT  11250.0 34695.0 11315.0 34760.0 ;
      RECT  10960.0 35412.5 11520.0 35477.5 ;
      RECT  10960.0 34067.5 11520.0 34132.5 ;
      RECT  9222.5 34660.0 9287.5 34795.0 ;
      RECT  9362.5 34387.5 9427.5 34522.5 ;
      RECT  10357.5 34492.5 10222.5 34557.5 ;
      RECT  9907.5 35630.0 9972.5 35445.0 ;
      RECT  9907.5 36790.0 9972.5 36605.0 ;
      RECT  9547.5 36672.5 9612.5 36822.5 ;
      RECT  9547.5 35787.5 9612.5 35412.5 ;
      RECT  9737.5 36672.5 9802.5 35787.5 ;
      RECT  9547.5 35787.5 9612.5 35652.5 ;
      RECT  9737.5 35787.5 9802.5 35652.5 ;
      RECT  9737.5 35787.5 9802.5 35652.5 ;
      RECT  9547.5 35787.5 9612.5 35652.5 ;
      RECT  9547.5 36672.5 9612.5 36537.5 ;
      RECT  9737.5 36672.5 9802.5 36537.5 ;
      RECT  9737.5 36672.5 9802.5 36537.5 ;
      RECT  9547.5 36672.5 9612.5 36537.5 ;
      RECT  9907.5 35697.5 9972.5 35562.5 ;
      RECT  9907.5 36672.5 9972.5 36537.5 ;
      RECT  9605.0 36230.0 9670.0 36095.0 ;
      RECT  9605.0 36230.0 9670.0 36095.0 ;
      RECT  9770.0 36195.0 9835.0 36130.0 ;
      RECT  9480.0 35477.5 10040.0 35412.5 ;
      RECT  9480.0 36822.5 10040.0 36757.5 ;
      RECT  10107.5 36627.5 10172.5 36822.5 ;
      RECT  10107.5 35787.5 10172.5 35412.5 ;
      RECT  10487.5 35787.5 10552.5 35412.5 ;
      RECT  10657.5 35630.0 10722.5 35445.0 ;
      RECT  10657.5 36790.0 10722.5 36605.0 ;
      RECT  10107.5 35787.5 10172.5 35652.5 ;
      RECT  10297.5 35787.5 10362.5 35652.5 ;
      RECT  10297.5 35787.5 10362.5 35652.5 ;
      RECT  10107.5 35787.5 10172.5 35652.5 ;
      RECT  10297.5 35787.5 10362.5 35652.5 ;
      RECT  10487.5 35787.5 10552.5 35652.5 ;
      RECT  10487.5 35787.5 10552.5 35652.5 ;
      RECT  10297.5 35787.5 10362.5 35652.5 ;
      RECT  10107.5 36627.5 10172.5 36492.5 ;
      RECT  10297.5 36627.5 10362.5 36492.5 ;
      RECT  10297.5 36627.5 10362.5 36492.5 ;
      RECT  10107.5 36627.5 10172.5 36492.5 ;
      RECT  10297.5 36627.5 10362.5 36492.5 ;
      RECT  10487.5 36627.5 10552.5 36492.5 ;
      RECT  10487.5 36627.5 10552.5 36492.5 ;
      RECT  10297.5 36627.5 10362.5 36492.5 ;
      RECT  10657.5 35697.5 10722.5 35562.5 ;
      RECT  10657.5 36672.5 10722.5 36537.5 ;
      RECT  10492.5 36397.5 10357.5 36332.5 ;
      RECT  10235.0 36182.5 10100.0 36117.5 ;
      RECT  10297.5 35787.5 10362.5 35652.5 ;
      RECT  10487.5 36627.5 10552.5 36492.5 ;
      RECT  10587.5 36182.5 10452.5 36117.5 ;
      RECT  10100.0 36182.5 10235.0 36117.5 ;
      RECT  10357.5 36397.5 10492.5 36332.5 ;
      RECT  10452.5 36182.5 10587.5 36117.5 ;
      RECT  10040.0 35477.5 10960.0 35412.5 ;
      RECT  10040.0 36822.5 10960.0 36757.5 ;
      RECT  11387.5 35630.0 11452.5 35445.0 ;
      RECT  11387.5 36790.0 11452.5 36605.0 ;
      RECT  11027.5 36672.5 11092.5 36822.5 ;
      RECT  11027.5 35787.5 11092.5 35412.5 ;
      RECT  11217.5 36672.5 11282.5 35787.5 ;
      RECT  11027.5 35787.5 11092.5 35652.5 ;
      RECT  11217.5 35787.5 11282.5 35652.5 ;
      RECT  11217.5 35787.5 11282.5 35652.5 ;
      RECT  11027.5 35787.5 11092.5 35652.5 ;
      RECT  11027.5 36672.5 11092.5 36537.5 ;
      RECT  11217.5 36672.5 11282.5 36537.5 ;
      RECT  11217.5 36672.5 11282.5 36537.5 ;
      RECT  11027.5 36672.5 11092.5 36537.5 ;
      RECT  11387.5 35697.5 11452.5 35562.5 ;
      RECT  11387.5 36672.5 11452.5 36537.5 ;
      RECT  11085.0 36230.0 11150.0 36095.0 ;
      RECT  11085.0 36230.0 11150.0 36095.0 ;
      RECT  11250.0 36195.0 11315.0 36130.0 ;
      RECT  10960.0 35477.5 11520.0 35412.5 ;
      RECT  10960.0 36822.5 11520.0 36757.5 ;
      RECT  9222.5 36095.0 9287.5 36230.0 ;
      RECT  9362.5 36367.5 9427.5 36502.5 ;
      RECT  10357.5 36332.5 10222.5 36397.5 ;
      RECT  9907.5 37950.0 9972.5 38135.0 ;
      RECT  9907.5 36790.0 9972.5 36975.0 ;
      RECT  9547.5 36907.5 9612.5 36757.5 ;
      RECT  9547.5 37792.5 9612.5 38167.5 ;
      RECT  9737.5 36907.5 9802.5 37792.5 ;
      RECT  9547.5 37792.5 9612.5 37927.5 ;
      RECT  9737.5 37792.5 9802.5 37927.5 ;
      RECT  9737.5 37792.5 9802.5 37927.5 ;
      RECT  9547.5 37792.5 9612.5 37927.5 ;
      RECT  9547.5 36907.5 9612.5 37042.5 ;
      RECT  9737.5 36907.5 9802.5 37042.5 ;
      RECT  9737.5 36907.5 9802.5 37042.5 ;
      RECT  9547.5 36907.5 9612.5 37042.5 ;
      RECT  9907.5 37882.5 9972.5 38017.5 ;
      RECT  9907.5 36907.5 9972.5 37042.5 ;
      RECT  9605.0 37350.0 9670.0 37485.0 ;
      RECT  9605.0 37350.0 9670.0 37485.0 ;
      RECT  9770.0 37385.0 9835.0 37450.0 ;
      RECT  9480.0 38102.5 10040.0 38167.5 ;
      RECT  9480.0 36757.5 10040.0 36822.5 ;
      RECT  10107.5 36952.5 10172.5 36757.5 ;
      RECT  10107.5 37792.5 10172.5 38167.5 ;
      RECT  10487.5 37792.5 10552.5 38167.5 ;
      RECT  10657.5 37950.0 10722.5 38135.0 ;
      RECT  10657.5 36790.0 10722.5 36975.0 ;
      RECT  10107.5 37792.5 10172.5 37927.5 ;
      RECT  10297.5 37792.5 10362.5 37927.5 ;
      RECT  10297.5 37792.5 10362.5 37927.5 ;
      RECT  10107.5 37792.5 10172.5 37927.5 ;
      RECT  10297.5 37792.5 10362.5 37927.5 ;
      RECT  10487.5 37792.5 10552.5 37927.5 ;
      RECT  10487.5 37792.5 10552.5 37927.5 ;
      RECT  10297.5 37792.5 10362.5 37927.5 ;
      RECT  10107.5 36952.5 10172.5 37087.5 ;
      RECT  10297.5 36952.5 10362.5 37087.5 ;
      RECT  10297.5 36952.5 10362.5 37087.5 ;
      RECT  10107.5 36952.5 10172.5 37087.5 ;
      RECT  10297.5 36952.5 10362.5 37087.5 ;
      RECT  10487.5 36952.5 10552.5 37087.5 ;
      RECT  10487.5 36952.5 10552.5 37087.5 ;
      RECT  10297.5 36952.5 10362.5 37087.5 ;
      RECT  10657.5 37882.5 10722.5 38017.5 ;
      RECT  10657.5 36907.5 10722.5 37042.5 ;
      RECT  10492.5 37182.5 10357.5 37247.5 ;
      RECT  10235.0 37397.5 10100.0 37462.5 ;
      RECT  10297.5 37792.5 10362.5 37927.5 ;
      RECT  10487.5 36952.5 10552.5 37087.5 ;
      RECT  10587.5 37397.5 10452.5 37462.5 ;
      RECT  10100.0 37397.5 10235.0 37462.5 ;
      RECT  10357.5 37182.5 10492.5 37247.5 ;
      RECT  10452.5 37397.5 10587.5 37462.5 ;
      RECT  10040.0 38102.5 10960.0 38167.5 ;
      RECT  10040.0 36757.5 10960.0 36822.5 ;
      RECT  11387.5 37950.0 11452.5 38135.0 ;
      RECT  11387.5 36790.0 11452.5 36975.0 ;
      RECT  11027.5 36907.5 11092.5 36757.5 ;
      RECT  11027.5 37792.5 11092.5 38167.5 ;
      RECT  11217.5 36907.5 11282.5 37792.5 ;
      RECT  11027.5 37792.5 11092.5 37927.5 ;
      RECT  11217.5 37792.5 11282.5 37927.5 ;
      RECT  11217.5 37792.5 11282.5 37927.5 ;
      RECT  11027.5 37792.5 11092.5 37927.5 ;
      RECT  11027.5 36907.5 11092.5 37042.5 ;
      RECT  11217.5 36907.5 11282.5 37042.5 ;
      RECT  11217.5 36907.5 11282.5 37042.5 ;
      RECT  11027.5 36907.5 11092.5 37042.5 ;
      RECT  11387.5 37882.5 11452.5 38017.5 ;
      RECT  11387.5 36907.5 11452.5 37042.5 ;
      RECT  11085.0 37350.0 11150.0 37485.0 ;
      RECT  11085.0 37350.0 11150.0 37485.0 ;
      RECT  11250.0 37385.0 11315.0 37450.0 ;
      RECT  10960.0 38102.5 11520.0 38167.5 ;
      RECT  10960.0 36757.5 11520.0 36822.5 ;
      RECT  9222.5 37350.0 9287.5 37485.0 ;
      RECT  9362.5 37077.5 9427.5 37212.5 ;
      RECT  10357.5 37182.5 10222.5 37247.5 ;
      RECT  9907.5 38320.0 9972.5 38135.0 ;
      RECT  9907.5 39480.0 9972.5 39295.0 ;
      RECT  9547.5 39362.5 9612.5 39512.5 ;
      RECT  9547.5 38477.5 9612.5 38102.5 ;
      RECT  9737.5 39362.5 9802.5 38477.5 ;
      RECT  9547.5 38477.5 9612.5 38342.5 ;
      RECT  9737.5 38477.5 9802.5 38342.5 ;
      RECT  9737.5 38477.5 9802.5 38342.5 ;
      RECT  9547.5 38477.5 9612.5 38342.5 ;
      RECT  9547.5 39362.5 9612.5 39227.5 ;
      RECT  9737.5 39362.5 9802.5 39227.5 ;
      RECT  9737.5 39362.5 9802.5 39227.5 ;
      RECT  9547.5 39362.5 9612.5 39227.5 ;
      RECT  9907.5 38387.5 9972.5 38252.5 ;
      RECT  9907.5 39362.5 9972.5 39227.5 ;
      RECT  9605.0 38920.0 9670.0 38785.0 ;
      RECT  9605.0 38920.0 9670.0 38785.0 ;
      RECT  9770.0 38885.0 9835.0 38820.0 ;
      RECT  9480.0 38167.5 10040.0 38102.5 ;
      RECT  9480.0 39512.5 10040.0 39447.5 ;
      RECT  10107.5 39317.5 10172.5 39512.5 ;
      RECT  10107.5 38477.5 10172.5 38102.5 ;
      RECT  10487.5 38477.5 10552.5 38102.5 ;
      RECT  10657.5 38320.0 10722.5 38135.0 ;
      RECT  10657.5 39480.0 10722.5 39295.0 ;
      RECT  10107.5 38477.5 10172.5 38342.5 ;
      RECT  10297.5 38477.5 10362.5 38342.5 ;
      RECT  10297.5 38477.5 10362.5 38342.5 ;
      RECT  10107.5 38477.5 10172.5 38342.5 ;
      RECT  10297.5 38477.5 10362.5 38342.5 ;
      RECT  10487.5 38477.5 10552.5 38342.5 ;
      RECT  10487.5 38477.5 10552.5 38342.5 ;
      RECT  10297.5 38477.5 10362.5 38342.5 ;
      RECT  10107.5 39317.5 10172.5 39182.5 ;
      RECT  10297.5 39317.5 10362.5 39182.5 ;
      RECT  10297.5 39317.5 10362.5 39182.5 ;
      RECT  10107.5 39317.5 10172.5 39182.5 ;
      RECT  10297.5 39317.5 10362.5 39182.5 ;
      RECT  10487.5 39317.5 10552.5 39182.5 ;
      RECT  10487.5 39317.5 10552.5 39182.5 ;
      RECT  10297.5 39317.5 10362.5 39182.5 ;
      RECT  10657.5 38387.5 10722.5 38252.5 ;
      RECT  10657.5 39362.5 10722.5 39227.5 ;
      RECT  10492.5 39087.5 10357.5 39022.5 ;
      RECT  10235.0 38872.5 10100.0 38807.5 ;
      RECT  10297.5 38477.5 10362.5 38342.5 ;
      RECT  10487.5 39317.5 10552.5 39182.5 ;
      RECT  10587.5 38872.5 10452.5 38807.5 ;
      RECT  10100.0 38872.5 10235.0 38807.5 ;
      RECT  10357.5 39087.5 10492.5 39022.5 ;
      RECT  10452.5 38872.5 10587.5 38807.5 ;
      RECT  10040.0 38167.5 10960.0 38102.5 ;
      RECT  10040.0 39512.5 10960.0 39447.5 ;
      RECT  11387.5 38320.0 11452.5 38135.0 ;
      RECT  11387.5 39480.0 11452.5 39295.0 ;
      RECT  11027.5 39362.5 11092.5 39512.5 ;
      RECT  11027.5 38477.5 11092.5 38102.5 ;
      RECT  11217.5 39362.5 11282.5 38477.5 ;
      RECT  11027.5 38477.5 11092.5 38342.5 ;
      RECT  11217.5 38477.5 11282.5 38342.5 ;
      RECT  11217.5 38477.5 11282.5 38342.5 ;
      RECT  11027.5 38477.5 11092.5 38342.5 ;
      RECT  11027.5 39362.5 11092.5 39227.5 ;
      RECT  11217.5 39362.5 11282.5 39227.5 ;
      RECT  11217.5 39362.5 11282.5 39227.5 ;
      RECT  11027.5 39362.5 11092.5 39227.5 ;
      RECT  11387.5 38387.5 11452.5 38252.5 ;
      RECT  11387.5 39362.5 11452.5 39227.5 ;
      RECT  11085.0 38920.0 11150.0 38785.0 ;
      RECT  11085.0 38920.0 11150.0 38785.0 ;
      RECT  11250.0 38885.0 11315.0 38820.0 ;
      RECT  10960.0 38167.5 11520.0 38102.5 ;
      RECT  10960.0 39512.5 11520.0 39447.5 ;
      RECT  9222.5 38785.0 9287.5 38920.0 ;
      RECT  9362.5 39057.5 9427.5 39192.5 ;
      RECT  10357.5 39022.5 10222.5 39087.5 ;
      RECT  9907.5 40640.0 9972.5 40825.0 ;
      RECT  9907.5 39480.0 9972.5 39665.0 ;
      RECT  9547.5 39597.5 9612.5 39447.5 ;
      RECT  9547.5 40482.5 9612.5 40857.5 ;
      RECT  9737.5 39597.5 9802.5 40482.5 ;
      RECT  9547.5 40482.5 9612.5 40617.5 ;
      RECT  9737.5 40482.5 9802.5 40617.5 ;
      RECT  9737.5 40482.5 9802.5 40617.5 ;
      RECT  9547.5 40482.5 9612.5 40617.5 ;
      RECT  9547.5 39597.5 9612.5 39732.5 ;
      RECT  9737.5 39597.5 9802.5 39732.5 ;
      RECT  9737.5 39597.5 9802.5 39732.5 ;
      RECT  9547.5 39597.5 9612.5 39732.5 ;
      RECT  9907.5 40572.5 9972.5 40707.5 ;
      RECT  9907.5 39597.5 9972.5 39732.5 ;
      RECT  9605.0 40040.0 9670.0 40175.0 ;
      RECT  9605.0 40040.0 9670.0 40175.0 ;
      RECT  9770.0 40075.0 9835.0 40140.0 ;
      RECT  9480.0 40792.5 10040.0 40857.5 ;
      RECT  9480.0 39447.5 10040.0 39512.5 ;
      RECT  10107.5 39642.5 10172.5 39447.5 ;
      RECT  10107.5 40482.5 10172.5 40857.5 ;
      RECT  10487.5 40482.5 10552.5 40857.5 ;
      RECT  10657.5 40640.0 10722.5 40825.0 ;
      RECT  10657.5 39480.0 10722.5 39665.0 ;
      RECT  10107.5 40482.5 10172.5 40617.5 ;
      RECT  10297.5 40482.5 10362.5 40617.5 ;
      RECT  10297.5 40482.5 10362.5 40617.5 ;
      RECT  10107.5 40482.5 10172.5 40617.5 ;
      RECT  10297.5 40482.5 10362.5 40617.5 ;
      RECT  10487.5 40482.5 10552.5 40617.5 ;
      RECT  10487.5 40482.5 10552.5 40617.5 ;
      RECT  10297.5 40482.5 10362.5 40617.5 ;
      RECT  10107.5 39642.5 10172.5 39777.5 ;
      RECT  10297.5 39642.5 10362.5 39777.5 ;
      RECT  10297.5 39642.5 10362.5 39777.5 ;
      RECT  10107.5 39642.5 10172.5 39777.5 ;
      RECT  10297.5 39642.5 10362.5 39777.5 ;
      RECT  10487.5 39642.5 10552.5 39777.5 ;
      RECT  10487.5 39642.5 10552.5 39777.5 ;
      RECT  10297.5 39642.5 10362.5 39777.5 ;
      RECT  10657.5 40572.5 10722.5 40707.5 ;
      RECT  10657.5 39597.5 10722.5 39732.5 ;
      RECT  10492.5 39872.5 10357.5 39937.5 ;
      RECT  10235.0 40087.5 10100.0 40152.5 ;
      RECT  10297.5 40482.5 10362.5 40617.5 ;
      RECT  10487.5 39642.5 10552.5 39777.5 ;
      RECT  10587.5 40087.5 10452.5 40152.5 ;
      RECT  10100.0 40087.5 10235.0 40152.5 ;
      RECT  10357.5 39872.5 10492.5 39937.5 ;
      RECT  10452.5 40087.5 10587.5 40152.5 ;
      RECT  10040.0 40792.5 10960.0 40857.5 ;
      RECT  10040.0 39447.5 10960.0 39512.5 ;
      RECT  11387.5 40640.0 11452.5 40825.0 ;
      RECT  11387.5 39480.0 11452.5 39665.0 ;
      RECT  11027.5 39597.5 11092.5 39447.5 ;
      RECT  11027.5 40482.5 11092.5 40857.5 ;
      RECT  11217.5 39597.5 11282.5 40482.5 ;
      RECT  11027.5 40482.5 11092.5 40617.5 ;
      RECT  11217.5 40482.5 11282.5 40617.5 ;
      RECT  11217.5 40482.5 11282.5 40617.5 ;
      RECT  11027.5 40482.5 11092.5 40617.5 ;
      RECT  11027.5 39597.5 11092.5 39732.5 ;
      RECT  11217.5 39597.5 11282.5 39732.5 ;
      RECT  11217.5 39597.5 11282.5 39732.5 ;
      RECT  11027.5 39597.5 11092.5 39732.5 ;
      RECT  11387.5 40572.5 11452.5 40707.5 ;
      RECT  11387.5 39597.5 11452.5 39732.5 ;
      RECT  11085.0 40040.0 11150.0 40175.0 ;
      RECT  11085.0 40040.0 11150.0 40175.0 ;
      RECT  11250.0 40075.0 11315.0 40140.0 ;
      RECT  10960.0 40792.5 11520.0 40857.5 ;
      RECT  10960.0 39447.5 11520.0 39512.5 ;
      RECT  9222.5 40040.0 9287.5 40175.0 ;
      RECT  9362.5 39767.5 9427.5 39902.5 ;
      RECT  10357.5 39872.5 10222.5 39937.5 ;
      RECT  9907.5 41010.0 9972.5 40825.0 ;
      RECT  9907.5 42170.0 9972.5 41985.0 ;
      RECT  9547.5 42052.5 9612.5 42202.5 ;
      RECT  9547.5 41167.5 9612.5 40792.5 ;
      RECT  9737.5 42052.5 9802.5 41167.5 ;
      RECT  9547.5 41167.5 9612.5 41032.5 ;
      RECT  9737.5 41167.5 9802.5 41032.5 ;
      RECT  9737.5 41167.5 9802.5 41032.5 ;
      RECT  9547.5 41167.5 9612.5 41032.5 ;
      RECT  9547.5 42052.5 9612.5 41917.5 ;
      RECT  9737.5 42052.5 9802.5 41917.5 ;
      RECT  9737.5 42052.5 9802.5 41917.5 ;
      RECT  9547.5 42052.5 9612.5 41917.5 ;
      RECT  9907.5 41077.5 9972.5 40942.5 ;
      RECT  9907.5 42052.5 9972.5 41917.5 ;
      RECT  9605.0 41610.0 9670.0 41475.0 ;
      RECT  9605.0 41610.0 9670.0 41475.0 ;
      RECT  9770.0 41575.0 9835.0 41510.0 ;
      RECT  9480.0 40857.5 10040.0 40792.5 ;
      RECT  9480.0 42202.5 10040.0 42137.5 ;
      RECT  10107.5 42007.5 10172.5 42202.5 ;
      RECT  10107.5 41167.5 10172.5 40792.5 ;
      RECT  10487.5 41167.5 10552.5 40792.5 ;
      RECT  10657.5 41010.0 10722.5 40825.0 ;
      RECT  10657.5 42170.0 10722.5 41985.0 ;
      RECT  10107.5 41167.5 10172.5 41032.5 ;
      RECT  10297.5 41167.5 10362.5 41032.5 ;
      RECT  10297.5 41167.5 10362.5 41032.5 ;
      RECT  10107.5 41167.5 10172.5 41032.5 ;
      RECT  10297.5 41167.5 10362.5 41032.5 ;
      RECT  10487.5 41167.5 10552.5 41032.5 ;
      RECT  10487.5 41167.5 10552.5 41032.5 ;
      RECT  10297.5 41167.5 10362.5 41032.5 ;
      RECT  10107.5 42007.5 10172.5 41872.5 ;
      RECT  10297.5 42007.5 10362.5 41872.5 ;
      RECT  10297.5 42007.5 10362.5 41872.5 ;
      RECT  10107.5 42007.5 10172.5 41872.5 ;
      RECT  10297.5 42007.5 10362.5 41872.5 ;
      RECT  10487.5 42007.5 10552.5 41872.5 ;
      RECT  10487.5 42007.5 10552.5 41872.5 ;
      RECT  10297.5 42007.5 10362.5 41872.5 ;
      RECT  10657.5 41077.5 10722.5 40942.5 ;
      RECT  10657.5 42052.5 10722.5 41917.5 ;
      RECT  10492.5 41777.5 10357.5 41712.5 ;
      RECT  10235.0 41562.5 10100.0 41497.5 ;
      RECT  10297.5 41167.5 10362.5 41032.5 ;
      RECT  10487.5 42007.5 10552.5 41872.5 ;
      RECT  10587.5 41562.5 10452.5 41497.5 ;
      RECT  10100.0 41562.5 10235.0 41497.5 ;
      RECT  10357.5 41777.5 10492.5 41712.5 ;
      RECT  10452.5 41562.5 10587.5 41497.5 ;
      RECT  10040.0 40857.5 10960.0 40792.5 ;
      RECT  10040.0 42202.5 10960.0 42137.5 ;
      RECT  11387.5 41010.0 11452.5 40825.0 ;
      RECT  11387.5 42170.0 11452.5 41985.0 ;
      RECT  11027.5 42052.5 11092.5 42202.5 ;
      RECT  11027.5 41167.5 11092.5 40792.5 ;
      RECT  11217.5 42052.5 11282.5 41167.5 ;
      RECT  11027.5 41167.5 11092.5 41032.5 ;
      RECT  11217.5 41167.5 11282.5 41032.5 ;
      RECT  11217.5 41167.5 11282.5 41032.5 ;
      RECT  11027.5 41167.5 11092.5 41032.5 ;
      RECT  11027.5 42052.5 11092.5 41917.5 ;
      RECT  11217.5 42052.5 11282.5 41917.5 ;
      RECT  11217.5 42052.5 11282.5 41917.5 ;
      RECT  11027.5 42052.5 11092.5 41917.5 ;
      RECT  11387.5 41077.5 11452.5 40942.5 ;
      RECT  11387.5 42052.5 11452.5 41917.5 ;
      RECT  11085.0 41610.0 11150.0 41475.0 ;
      RECT  11085.0 41610.0 11150.0 41475.0 ;
      RECT  11250.0 41575.0 11315.0 41510.0 ;
      RECT  10960.0 40857.5 11520.0 40792.5 ;
      RECT  10960.0 42202.5 11520.0 42137.5 ;
      RECT  9222.5 41475.0 9287.5 41610.0 ;
      RECT  9362.5 41747.5 9427.5 41882.5 ;
      RECT  10357.5 41712.5 10222.5 41777.5 ;
      RECT  9907.5 43330.0 9972.5 43515.0 ;
      RECT  9907.5 42170.0 9972.5 42355.0 ;
      RECT  9547.5 42287.5 9612.5 42137.5 ;
      RECT  9547.5 43172.5 9612.5 43547.5 ;
      RECT  9737.5 42287.5 9802.5 43172.5 ;
      RECT  9547.5 43172.5 9612.5 43307.5 ;
      RECT  9737.5 43172.5 9802.5 43307.5 ;
      RECT  9737.5 43172.5 9802.5 43307.5 ;
      RECT  9547.5 43172.5 9612.5 43307.5 ;
      RECT  9547.5 42287.5 9612.5 42422.5 ;
      RECT  9737.5 42287.5 9802.5 42422.5 ;
      RECT  9737.5 42287.5 9802.5 42422.5 ;
      RECT  9547.5 42287.5 9612.5 42422.5 ;
      RECT  9907.5 43262.5 9972.5 43397.5 ;
      RECT  9907.5 42287.5 9972.5 42422.5 ;
      RECT  9605.0 42730.0 9670.0 42865.0 ;
      RECT  9605.0 42730.0 9670.0 42865.0 ;
      RECT  9770.0 42765.0 9835.0 42830.0 ;
      RECT  9480.0 43482.5 10040.0 43547.5 ;
      RECT  9480.0 42137.5 10040.0 42202.5 ;
      RECT  10107.5 42332.5 10172.5 42137.5 ;
      RECT  10107.5 43172.5 10172.5 43547.5 ;
      RECT  10487.5 43172.5 10552.5 43547.5 ;
      RECT  10657.5 43330.0 10722.5 43515.0 ;
      RECT  10657.5 42170.0 10722.5 42355.0 ;
      RECT  10107.5 43172.5 10172.5 43307.5 ;
      RECT  10297.5 43172.5 10362.5 43307.5 ;
      RECT  10297.5 43172.5 10362.5 43307.5 ;
      RECT  10107.5 43172.5 10172.5 43307.5 ;
      RECT  10297.5 43172.5 10362.5 43307.5 ;
      RECT  10487.5 43172.5 10552.5 43307.5 ;
      RECT  10487.5 43172.5 10552.5 43307.5 ;
      RECT  10297.5 43172.5 10362.5 43307.5 ;
      RECT  10107.5 42332.5 10172.5 42467.5 ;
      RECT  10297.5 42332.5 10362.5 42467.5 ;
      RECT  10297.5 42332.5 10362.5 42467.5 ;
      RECT  10107.5 42332.5 10172.5 42467.5 ;
      RECT  10297.5 42332.5 10362.5 42467.5 ;
      RECT  10487.5 42332.5 10552.5 42467.5 ;
      RECT  10487.5 42332.5 10552.5 42467.5 ;
      RECT  10297.5 42332.5 10362.5 42467.5 ;
      RECT  10657.5 43262.5 10722.5 43397.5 ;
      RECT  10657.5 42287.5 10722.5 42422.5 ;
      RECT  10492.5 42562.5 10357.5 42627.5 ;
      RECT  10235.0 42777.5 10100.0 42842.5 ;
      RECT  10297.5 43172.5 10362.5 43307.5 ;
      RECT  10487.5 42332.5 10552.5 42467.5 ;
      RECT  10587.5 42777.5 10452.5 42842.5 ;
      RECT  10100.0 42777.5 10235.0 42842.5 ;
      RECT  10357.5 42562.5 10492.5 42627.5 ;
      RECT  10452.5 42777.5 10587.5 42842.5 ;
      RECT  10040.0 43482.5 10960.0 43547.5 ;
      RECT  10040.0 42137.5 10960.0 42202.5 ;
      RECT  11387.5 43330.0 11452.5 43515.0 ;
      RECT  11387.5 42170.0 11452.5 42355.0 ;
      RECT  11027.5 42287.5 11092.5 42137.5 ;
      RECT  11027.5 43172.5 11092.5 43547.5 ;
      RECT  11217.5 42287.5 11282.5 43172.5 ;
      RECT  11027.5 43172.5 11092.5 43307.5 ;
      RECT  11217.5 43172.5 11282.5 43307.5 ;
      RECT  11217.5 43172.5 11282.5 43307.5 ;
      RECT  11027.5 43172.5 11092.5 43307.5 ;
      RECT  11027.5 42287.5 11092.5 42422.5 ;
      RECT  11217.5 42287.5 11282.5 42422.5 ;
      RECT  11217.5 42287.5 11282.5 42422.5 ;
      RECT  11027.5 42287.5 11092.5 42422.5 ;
      RECT  11387.5 43262.5 11452.5 43397.5 ;
      RECT  11387.5 42287.5 11452.5 42422.5 ;
      RECT  11085.0 42730.0 11150.0 42865.0 ;
      RECT  11085.0 42730.0 11150.0 42865.0 ;
      RECT  11250.0 42765.0 11315.0 42830.0 ;
      RECT  10960.0 43482.5 11520.0 43547.5 ;
      RECT  10960.0 42137.5 11520.0 42202.5 ;
      RECT  9222.5 42730.0 9287.5 42865.0 ;
      RECT  9362.5 42457.5 9427.5 42592.5 ;
      RECT  10357.5 42562.5 10222.5 42627.5 ;
      RECT  9907.5 43700.0 9972.5 43515.0 ;
      RECT  9907.5 44860.0 9972.5 44675.0 ;
      RECT  9547.5 44742.5 9612.5 44892.5 ;
      RECT  9547.5 43857.5 9612.5 43482.5 ;
      RECT  9737.5 44742.5 9802.5 43857.5 ;
      RECT  9547.5 43857.5 9612.5 43722.5 ;
      RECT  9737.5 43857.5 9802.5 43722.5 ;
      RECT  9737.5 43857.5 9802.5 43722.5 ;
      RECT  9547.5 43857.5 9612.5 43722.5 ;
      RECT  9547.5 44742.5 9612.5 44607.5 ;
      RECT  9737.5 44742.5 9802.5 44607.5 ;
      RECT  9737.5 44742.5 9802.5 44607.5 ;
      RECT  9547.5 44742.5 9612.5 44607.5 ;
      RECT  9907.5 43767.5 9972.5 43632.5 ;
      RECT  9907.5 44742.5 9972.5 44607.5 ;
      RECT  9605.0 44300.0 9670.0 44165.0 ;
      RECT  9605.0 44300.0 9670.0 44165.0 ;
      RECT  9770.0 44265.0 9835.0 44200.0 ;
      RECT  9480.0 43547.5 10040.0 43482.5 ;
      RECT  9480.0 44892.5 10040.0 44827.5 ;
      RECT  10107.5 44697.5 10172.5 44892.5 ;
      RECT  10107.5 43857.5 10172.5 43482.5 ;
      RECT  10487.5 43857.5 10552.5 43482.5 ;
      RECT  10657.5 43700.0 10722.5 43515.0 ;
      RECT  10657.5 44860.0 10722.5 44675.0 ;
      RECT  10107.5 43857.5 10172.5 43722.5 ;
      RECT  10297.5 43857.5 10362.5 43722.5 ;
      RECT  10297.5 43857.5 10362.5 43722.5 ;
      RECT  10107.5 43857.5 10172.5 43722.5 ;
      RECT  10297.5 43857.5 10362.5 43722.5 ;
      RECT  10487.5 43857.5 10552.5 43722.5 ;
      RECT  10487.5 43857.5 10552.5 43722.5 ;
      RECT  10297.5 43857.5 10362.5 43722.5 ;
      RECT  10107.5 44697.5 10172.5 44562.5 ;
      RECT  10297.5 44697.5 10362.5 44562.5 ;
      RECT  10297.5 44697.5 10362.5 44562.5 ;
      RECT  10107.5 44697.5 10172.5 44562.5 ;
      RECT  10297.5 44697.5 10362.5 44562.5 ;
      RECT  10487.5 44697.5 10552.5 44562.5 ;
      RECT  10487.5 44697.5 10552.5 44562.5 ;
      RECT  10297.5 44697.5 10362.5 44562.5 ;
      RECT  10657.5 43767.5 10722.5 43632.5 ;
      RECT  10657.5 44742.5 10722.5 44607.5 ;
      RECT  10492.5 44467.5 10357.5 44402.5 ;
      RECT  10235.0 44252.5 10100.0 44187.5 ;
      RECT  10297.5 43857.5 10362.5 43722.5 ;
      RECT  10487.5 44697.5 10552.5 44562.5 ;
      RECT  10587.5 44252.5 10452.5 44187.5 ;
      RECT  10100.0 44252.5 10235.0 44187.5 ;
      RECT  10357.5 44467.5 10492.5 44402.5 ;
      RECT  10452.5 44252.5 10587.5 44187.5 ;
      RECT  10040.0 43547.5 10960.0 43482.5 ;
      RECT  10040.0 44892.5 10960.0 44827.5 ;
      RECT  11387.5 43700.0 11452.5 43515.0 ;
      RECT  11387.5 44860.0 11452.5 44675.0 ;
      RECT  11027.5 44742.5 11092.5 44892.5 ;
      RECT  11027.5 43857.5 11092.5 43482.5 ;
      RECT  11217.5 44742.5 11282.5 43857.5 ;
      RECT  11027.5 43857.5 11092.5 43722.5 ;
      RECT  11217.5 43857.5 11282.5 43722.5 ;
      RECT  11217.5 43857.5 11282.5 43722.5 ;
      RECT  11027.5 43857.5 11092.5 43722.5 ;
      RECT  11027.5 44742.5 11092.5 44607.5 ;
      RECT  11217.5 44742.5 11282.5 44607.5 ;
      RECT  11217.5 44742.5 11282.5 44607.5 ;
      RECT  11027.5 44742.5 11092.5 44607.5 ;
      RECT  11387.5 43767.5 11452.5 43632.5 ;
      RECT  11387.5 44742.5 11452.5 44607.5 ;
      RECT  11085.0 44300.0 11150.0 44165.0 ;
      RECT  11085.0 44300.0 11150.0 44165.0 ;
      RECT  11250.0 44265.0 11315.0 44200.0 ;
      RECT  10960.0 43547.5 11520.0 43482.5 ;
      RECT  10960.0 44892.5 11520.0 44827.5 ;
      RECT  9222.5 44165.0 9287.5 44300.0 ;
      RECT  9362.5 44437.5 9427.5 44572.5 ;
      RECT  10357.5 44402.5 10222.5 44467.5 ;
      RECT  9907.5 46020.0 9972.5 46205.0 ;
      RECT  9907.5 44860.0 9972.5 45045.0 ;
      RECT  9547.5 44977.5 9612.5 44827.5 ;
      RECT  9547.5 45862.5 9612.5 46237.5 ;
      RECT  9737.5 44977.5 9802.5 45862.5 ;
      RECT  9547.5 45862.5 9612.5 45997.5 ;
      RECT  9737.5 45862.5 9802.5 45997.5 ;
      RECT  9737.5 45862.5 9802.5 45997.5 ;
      RECT  9547.5 45862.5 9612.5 45997.5 ;
      RECT  9547.5 44977.5 9612.5 45112.5 ;
      RECT  9737.5 44977.5 9802.5 45112.5 ;
      RECT  9737.5 44977.5 9802.5 45112.5 ;
      RECT  9547.5 44977.5 9612.5 45112.5 ;
      RECT  9907.5 45952.5 9972.5 46087.5 ;
      RECT  9907.5 44977.5 9972.5 45112.5 ;
      RECT  9605.0 45420.0 9670.0 45555.0 ;
      RECT  9605.0 45420.0 9670.0 45555.0 ;
      RECT  9770.0 45455.0 9835.0 45520.0 ;
      RECT  9480.0 46172.5 10040.0 46237.5 ;
      RECT  9480.0 44827.5 10040.0 44892.5 ;
      RECT  10107.5 45022.5 10172.5 44827.5 ;
      RECT  10107.5 45862.5 10172.5 46237.5 ;
      RECT  10487.5 45862.5 10552.5 46237.5 ;
      RECT  10657.5 46020.0 10722.5 46205.0 ;
      RECT  10657.5 44860.0 10722.5 45045.0 ;
      RECT  10107.5 45862.5 10172.5 45997.5 ;
      RECT  10297.5 45862.5 10362.5 45997.5 ;
      RECT  10297.5 45862.5 10362.5 45997.5 ;
      RECT  10107.5 45862.5 10172.5 45997.5 ;
      RECT  10297.5 45862.5 10362.5 45997.5 ;
      RECT  10487.5 45862.5 10552.5 45997.5 ;
      RECT  10487.5 45862.5 10552.5 45997.5 ;
      RECT  10297.5 45862.5 10362.5 45997.5 ;
      RECT  10107.5 45022.5 10172.5 45157.5 ;
      RECT  10297.5 45022.5 10362.5 45157.5 ;
      RECT  10297.5 45022.5 10362.5 45157.5 ;
      RECT  10107.5 45022.5 10172.5 45157.5 ;
      RECT  10297.5 45022.5 10362.5 45157.5 ;
      RECT  10487.5 45022.5 10552.5 45157.5 ;
      RECT  10487.5 45022.5 10552.5 45157.5 ;
      RECT  10297.5 45022.5 10362.5 45157.5 ;
      RECT  10657.5 45952.5 10722.5 46087.5 ;
      RECT  10657.5 44977.5 10722.5 45112.5 ;
      RECT  10492.5 45252.5 10357.5 45317.5 ;
      RECT  10235.0 45467.5 10100.0 45532.5 ;
      RECT  10297.5 45862.5 10362.5 45997.5 ;
      RECT  10487.5 45022.5 10552.5 45157.5 ;
      RECT  10587.5 45467.5 10452.5 45532.5 ;
      RECT  10100.0 45467.5 10235.0 45532.5 ;
      RECT  10357.5 45252.5 10492.5 45317.5 ;
      RECT  10452.5 45467.5 10587.5 45532.5 ;
      RECT  10040.0 46172.5 10960.0 46237.5 ;
      RECT  10040.0 44827.5 10960.0 44892.5 ;
      RECT  11387.5 46020.0 11452.5 46205.0 ;
      RECT  11387.5 44860.0 11452.5 45045.0 ;
      RECT  11027.5 44977.5 11092.5 44827.5 ;
      RECT  11027.5 45862.5 11092.5 46237.5 ;
      RECT  11217.5 44977.5 11282.5 45862.5 ;
      RECT  11027.5 45862.5 11092.5 45997.5 ;
      RECT  11217.5 45862.5 11282.5 45997.5 ;
      RECT  11217.5 45862.5 11282.5 45997.5 ;
      RECT  11027.5 45862.5 11092.5 45997.5 ;
      RECT  11027.5 44977.5 11092.5 45112.5 ;
      RECT  11217.5 44977.5 11282.5 45112.5 ;
      RECT  11217.5 44977.5 11282.5 45112.5 ;
      RECT  11027.5 44977.5 11092.5 45112.5 ;
      RECT  11387.5 45952.5 11452.5 46087.5 ;
      RECT  11387.5 44977.5 11452.5 45112.5 ;
      RECT  11085.0 45420.0 11150.0 45555.0 ;
      RECT  11085.0 45420.0 11150.0 45555.0 ;
      RECT  11250.0 45455.0 11315.0 45520.0 ;
      RECT  10960.0 46172.5 11520.0 46237.5 ;
      RECT  10960.0 44827.5 11520.0 44892.5 ;
      RECT  9222.5 45420.0 9287.5 45555.0 ;
      RECT  9362.5 45147.5 9427.5 45282.5 ;
      RECT  10357.5 45252.5 10222.5 45317.5 ;
      RECT  9907.5 46390.0 9972.5 46205.0 ;
      RECT  9907.5 47550.0 9972.5 47365.0 ;
      RECT  9547.5 47432.5 9612.5 47582.5 ;
      RECT  9547.5 46547.5 9612.5 46172.5 ;
      RECT  9737.5 47432.5 9802.5 46547.5 ;
      RECT  9547.5 46547.5 9612.5 46412.5 ;
      RECT  9737.5 46547.5 9802.5 46412.5 ;
      RECT  9737.5 46547.5 9802.5 46412.5 ;
      RECT  9547.5 46547.5 9612.5 46412.5 ;
      RECT  9547.5 47432.5 9612.5 47297.5 ;
      RECT  9737.5 47432.5 9802.5 47297.5 ;
      RECT  9737.5 47432.5 9802.5 47297.5 ;
      RECT  9547.5 47432.5 9612.5 47297.5 ;
      RECT  9907.5 46457.5 9972.5 46322.5 ;
      RECT  9907.5 47432.5 9972.5 47297.5 ;
      RECT  9605.0 46990.0 9670.0 46855.0 ;
      RECT  9605.0 46990.0 9670.0 46855.0 ;
      RECT  9770.0 46955.0 9835.0 46890.0 ;
      RECT  9480.0 46237.5 10040.0 46172.5 ;
      RECT  9480.0 47582.5 10040.0 47517.5 ;
      RECT  10107.5 47387.5 10172.5 47582.5 ;
      RECT  10107.5 46547.5 10172.5 46172.5 ;
      RECT  10487.5 46547.5 10552.5 46172.5 ;
      RECT  10657.5 46390.0 10722.5 46205.0 ;
      RECT  10657.5 47550.0 10722.5 47365.0 ;
      RECT  10107.5 46547.5 10172.5 46412.5 ;
      RECT  10297.5 46547.5 10362.5 46412.5 ;
      RECT  10297.5 46547.5 10362.5 46412.5 ;
      RECT  10107.5 46547.5 10172.5 46412.5 ;
      RECT  10297.5 46547.5 10362.5 46412.5 ;
      RECT  10487.5 46547.5 10552.5 46412.5 ;
      RECT  10487.5 46547.5 10552.5 46412.5 ;
      RECT  10297.5 46547.5 10362.5 46412.5 ;
      RECT  10107.5 47387.5 10172.5 47252.5 ;
      RECT  10297.5 47387.5 10362.5 47252.5 ;
      RECT  10297.5 47387.5 10362.5 47252.5 ;
      RECT  10107.5 47387.5 10172.5 47252.5 ;
      RECT  10297.5 47387.5 10362.5 47252.5 ;
      RECT  10487.5 47387.5 10552.5 47252.5 ;
      RECT  10487.5 47387.5 10552.5 47252.5 ;
      RECT  10297.5 47387.5 10362.5 47252.5 ;
      RECT  10657.5 46457.5 10722.5 46322.5 ;
      RECT  10657.5 47432.5 10722.5 47297.5 ;
      RECT  10492.5 47157.5 10357.5 47092.5 ;
      RECT  10235.0 46942.5 10100.0 46877.5 ;
      RECT  10297.5 46547.5 10362.5 46412.5 ;
      RECT  10487.5 47387.5 10552.5 47252.5 ;
      RECT  10587.5 46942.5 10452.5 46877.5 ;
      RECT  10100.0 46942.5 10235.0 46877.5 ;
      RECT  10357.5 47157.5 10492.5 47092.5 ;
      RECT  10452.5 46942.5 10587.5 46877.5 ;
      RECT  10040.0 46237.5 10960.0 46172.5 ;
      RECT  10040.0 47582.5 10960.0 47517.5 ;
      RECT  11387.5 46390.0 11452.5 46205.0 ;
      RECT  11387.5 47550.0 11452.5 47365.0 ;
      RECT  11027.5 47432.5 11092.5 47582.5 ;
      RECT  11027.5 46547.5 11092.5 46172.5 ;
      RECT  11217.5 47432.5 11282.5 46547.5 ;
      RECT  11027.5 46547.5 11092.5 46412.5 ;
      RECT  11217.5 46547.5 11282.5 46412.5 ;
      RECT  11217.5 46547.5 11282.5 46412.5 ;
      RECT  11027.5 46547.5 11092.5 46412.5 ;
      RECT  11027.5 47432.5 11092.5 47297.5 ;
      RECT  11217.5 47432.5 11282.5 47297.5 ;
      RECT  11217.5 47432.5 11282.5 47297.5 ;
      RECT  11027.5 47432.5 11092.5 47297.5 ;
      RECT  11387.5 46457.5 11452.5 46322.5 ;
      RECT  11387.5 47432.5 11452.5 47297.5 ;
      RECT  11085.0 46990.0 11150.0 46855.0 ;
      RECT  11085.0 46990.0 11150.0 46855.0 ;
      RECT  11250.0 46955.0 11315.0 46890.0 ;
      RECT  10960.0 46237.5 11520.0 46172.5 ;
      RECT  10960.0 47582.5 11520.0 47517.5 ;
      RECT  9222.5 46855.0 9287.5 46990.0 ;
      RECT  9362.5 47127.5 9427.5 47262.5 ;
      RECT  10357.5 47092.5 10222.5 47157.5 ;
      RECT  9907.5 48710.0 9972.5 48895.0 ;
      RECT  9907.5 47550.0 9972.5 47735.0 ;
      RECT  9547.5 47667.5 9612.5 47517.5 ;
      RECT  9547.5 48552.5 9612.5 48927.5 ;
      RECT  9737.5 47667.5 9802.5 48552.5 ;
      RECT  9547.5 48552.5 9612.5 48687.5 ;
      RECT  9737.5 48552.5 9802.5 48687.5 ;
      RECT  9737.5 48552.5 9802.5 48687.5 ;
      RECT  9547.5 48552.5 9612.5 48687.5 ;
      RECT  9547.5 47667.5 9612.5 47802.5 ;
      RECT  9737.5 47667.5 9802.5 47802.5 ;
      RECT  9737.5 47667.5 9802.5 47802.5 ;
      RECT  9547.5 47667.5 9612.5 47802.5 ;
      RECT  9907.5 48642.5 9972.5 48777.5 ;
      RECT  9907.5 47667.5 9972.5 47802.5 ;
      RECT  9605.0 48110.0 9670.0 48245.0 ;
      RECT  9605.0 48110.0 9670.0 48245.0 ;
      RECT  9770.0 48145.0 9835.0 48210.0 ;
      RECT  9480.0 48862.5 10040.0 48927.5 ;
      RECT  9480.0 47517.5 10040.0 47582.5 ;
      RECT  10107.5 47712.5 10172.5 47517.5 ;
      RECT  10107.5 48552.5 10172.5 48927.5 ;
      RECT  10487.5 48552.5 10552.5 48927.5 ;
      RECT  10657.5 48710.0 10722.5 48895.0 ;
      RECT  10657.5 47550.0 10722.5 47735.0 ;
      RECT  10107.5 48552.5 10172.5 48687.5 ;
      RECT  10297.5 48552.5 10362.5 48687.5 ;
      RECT  10297.5 48552.5 10362.5 48687.5 ;
      RECT  10107.5 48552.5 10172.5 48687.5 ;
      RECT  10297.5 48552.5 10362.5 48687.5 ;
      RECT  10487.5 48552.5 10552.5 48687.5 ;
      RECT  10487.5 48552.5 10552.5 48687.5 ;
      RECT  10297.5 48552.5 10362.5 48687.5 ;
      RECT  10107.5 47712.5 10172.5 47847.5 ;
      RECT  10297.5 47712.5 10362.5 47847.5 ;
      RECT  10297.5 47712.5 10362.5 47847.5 ;
      RECT  10107.5 47712.5 10172.5 47847.5 ;
      RECT  10297.5 47712.5 10362.5 47847.5 ;
      RECT  10487.5 47712.5 10552.5 47847.5 ;
      RECT  10487.5 47712.5 10552.5 47847.5 ;
      RECT  10297.5 47712.5 10362.5 47847.5 ;
      RECT  10657.5 48642.5 10722.5 48777.5 ;
      RECT  10657.5 47667.5 10722.5 47802.5 ;
      RECT  10492.5 47942.5 10357.5 48007.5 ;
      RECT  10235.0 48157.5 10100.0 48222.5 ;
      RECT  10297.5 48552.5 10362.5 48687.5 ;
      RECT  10487.5 47712.5 10552.5 47847.5 ;
      RECT  10587.5 48157.5 10452.5 48222.5 ;
      RECT  10100.0 48157.5 10235.0 48222.5 ;
      RECT  10357.5 47942.5 10492.5 48007.5 ;
      RECT  10452.5 48157.5 10587.5 48222.5 ;
      RECT  10040.0 48862.5 10960.0 48927.5 ;
      RECT  10040.0 47517.5 10960.0 47582.5 ;
      RECT  11387.5 48710.0 11452.5 48895.0 ;
      RECT  11387.5 47550.0 11452.5 47735.0 ;
      RECT  11027.5 47667.5 11092.5 47517.5 ;
      RECT  11027.5 48552.5 11092.5 48927.5 ;
      RECT  11217.5 47667.5 11282.5 48552.5 ;
      RECT  11027.5 48552.5 11092.5 48687.5 ;
      RECT  11217.5 48552.5 11282.5 48687.5 ;
      RECT  11217.5 48552.5 11282.5 48687.5 ;
      RECT  11027.5 48552.5 11092.5 48687.5 ;
      RECT  11027.5 47667.5 11092.5 47802.5 ;
      RECT  11217.5 47667.5 11282.5 47802.5 ;
      RECT  11217.5 47667.5 11282.5 47802.5 ;
      RECT  11027.5 47667.5 11092.5 47802.5 ;
      RECT  11387.5 48642.5 11452.5 48777.5 ;
      RECT  11387.5 47667.5 11452.5 47802.5 ;
      RECT  11085.0 48110.0 11150.0 48245.0 ;
      RECT  11085.0 48110.0 11150.0 48245.0 ;
      RECT  11250.0 48145.0 11315.0 48210.0 ;
      RECT  10960.0 48862.5 11520.0 48927.5 ;
      RECT  10960.0 47517.5 11520.0 47582.5 ;
      RECT  9222.5 48110.0 9287.5 48245.0 ;
      RECT  9362.5 47837.5 9427.5 47972.5 ;
      RECT  10357.5 47942.5 10222.5 48007.5 ;
      RECT  9907.5 49080.0 9972.5 48895.0 ;
      RECT  9907.5 50240.0 9972.5 50055.0 ;
      RECT  9547.5 50122.5 9612.5 50272.5 ;
      RECT  9547.5 49237.5 9612.5 48862.5 ;
      RECT  9737.5 50122.5 9802.5 49237.5 ;
      RECT  9547.5 49237.5 9612.5 49102.5 ;
      RECT  9737.5 49237.5 9802.5 49102.5 ;
      RECT  9737.5 49237.5 9802.5 49102.5 ;
      RECT  9547.5 49237.5 9612.5 49102.5 ;
      RECT  9547.5 50122.5 9612.5 49987.5 ;
      RECT  9737.5 50122.5 9802.5 49987.5 ;
      RECT  9737.5 50122.5 9802.5 49987.5 ;
      RECT  9547.5 50122.5 9612.5 49987.5 ;
      RECT  9907.5 49147.5 9972.5 49012.5 ;
      RECT  9907.5 50122.5 9972.5 49987.5 ;
      RECT  9605.0 49680.0 9670.0 49545.0 ;
      RECT  9605.0 49680.0 9670.0 49545.0 ;
      RECT  9770.0 49645.0 9835.0 49580.0 ;
      RECT  9480.0 48927.5 10040.0 48862.5 ;
      RECT  9480.0 50272.5 10040.0 50207.5 ;
      RECT  10107.5 50077.5 10172.5 50272.5 ;
      RECT  10107.5 49237.5 10172.5 48862.5 ;
      RECT  10487.5 49237.5 10552.5 48862.5 ;
      RECT  10657.5 49080.0 10722.5 48895.0 ;
      RECT  10657.5 50240.0 10722.5 50055.0 ;
      RECT  10107.5 49237.5 10172.5 49102.5 ;
      RECT  10297.5 49237.5 10362.5 49102.5 ;
      RECT  10297.5 49237.5 10362.5 49102.5 ;
      RECT  10107.5 49237.5 10172.5 49102.5 ;
      RECT  10297.5 49237.5 10362.5 49102.5 ;
      RECT  10487.5 49237.5 10552.5 49102.5 ;
      RECT  10487.5 49237.5 10552.5 49102.5 ;
      RECT  10297.5 49237.5 10362.5 49102.5 ;
      RECT  10107.5 50077.5 10172.5 49942.5 ;
      RECT  10297.5 50077.5 10362.5 49942.5 ;
      RECT  10297.5 50077.5 10362.5 49942.5 ;
      RECT  10107.5 50077.5 10172.5 49942.5 ;
      RECT  10297.5 50077.5 10362.5 49942.5 ;
      RECT  10487.5 50077.5 10552.5 49942.5 ;
      RECT  10487.5 50077.5 10552.5 49942.5 ;
      RECT  10297.5 50077.5 10362.5 49942.5 ;
      RECT  10657.5 49147.5 10722.5 49012.5 ;
      RECT  10657.5 50122.5 10722.5 49987.5 ;
      RECT  10492.5 49847.5 10357.5 49782.5 ;
      RECT  10235.0 49632.5 10100.0 49567.5 ;
      RECT  10297.5 49237.5 10362.5 49102.5 ;
      RECT  10487.5 50077.5 10552.5 49942.5 ;
      RECT  10587.5 49632.5 10452.5 49567.5 ;
      RECT  10100.0 49632.5 10235.0 49567.5 ;
      RECT  10357.5 49847.5 10492.5 49782.5 ;
      RECT  10452.5 49632.5 10587.5 49567.5 ;
      RECT  10040.0 48927.5 10960.0 48862.5 ;
      RECT  10040.0 50272.5 10960.0 50207.5 ;
      RECT  11387.5 49080.0 11452.5 48895.0 ;
      RECT  11387.5 50240.0 11452.5 50055.0 ;
      RECT  11027.5 50122.5 11092.5 50272.5 ;
      RECT  11027.5 49237.5 11092.5 48862.5 ;
      RECT  11217.5 50122.5 11282.5 49237.5 ;
      RECT  11027.5 49237.5 11092.5 49102.5 ;
      RECT  11217.5 49237.5 11282.5 49102.5 ;
      RECT  11217.5 49237.5 11282.5 49102.5 ;
      RECT  11027.5 49237.5 11092.5 49102.5 ;
      RECT  11027.5 50122.5 11092.5 49987.5 ;
      RECT  11217.5 50122.5 11282.5 49987.5 ;
      RECT  11217.5 50122.5 11282.5 49987.5 ;
      RECT  11027.5 50122.5 11092.5 49987.5 ;
      RECT  11387.5 49147.5 11452.5 49012.5 ;
      RECT  11387.5 50122.5 11452.5 49987.5 ;
      RECT  11085.0 49680.0 11150.0 49545.0 ;
      RECT  11085.0 49680.0 11150.0 49545.0 ;
      RECT  11250.0 49645.0 11315.0 49580.0 ;
      RECT  10960.0 48927.5 11520.0 48862.5 ;
      RECT  10960.0 50272.5 11520.0 50207.5 ;
      RECT  9222.5 49545.0 9287.5 49680.0 ;
      RECT  9362.5 49817.5 9427.5 49952.5 ;
      RECT  10357.5 49782.5 10222.5 49847.5 ;
      RECT  9907.5 51400.0 9972.5 51585.0 ;
      RECT  9907.5 50240.0 9972.5 50425.0 ;
      RECT  9547.5 50357.5 9612.5 50207.5 ;
      RECT  9547.5 51242.5 9612.5 51617.5 ;
      RECT  9737.5 50357.5 9802.5 51242.5 ;
      RECT  9547.5 51242.5 9612.5 51377.5 ;
      RECT  9737.5 51242.5 9802.5 51377.5 ;
      RECT  9737.5 51242.5 9802.5 51377.5 ;
      RECT  9547.5 51242.5 9612.5 51377.5 ;
      RECT  9547.5 50357.5 9612.5 50492.5 ;
      RECT  9737.5 50357.5 9802.5 50492.5 ;
      RECT  9737.5 50357.5 9802.5 50492.5 ;
      RECT  9547.5 50357.5 9612.5 50492.5 ;
      RECT  9907.5 51332.5 9972.5 51467.5 ;
      RECT  9907.5 50357.5 9972.5 50492.5 ;
      RECT  9605.0 50800.0 9670.0 50935.0 ;
      RECT  9605.0 50800.0 9670.0 50935.0 ;
      RECT  9770.0 50835.0 9835.0 50900.0 ;
      RECT  9480.0 51552.5 10040.0 51617.5 ;
      RECT  9480.0 50207.5 10040.0 50272.5 ;
      RECT  10107.5 50402.5 10172.5 50207.5 ;
      RECT  10107.5 51242.5 10172.5 51617.5 ;
      RECT  10487.5 51242.5 10552.5 51617.5 ;
      RECT  10657.5 51400.0 10722.5 51585.0 ;
      RECT  10657.5 50240.0 10722.5 50425.0 ;
      RECT  10107.5 51242.5 10172.5 51377.5 ;
      RECT  10297.5 51242.5 10362.5 51377.5 ;
      RECT  10297.5 51242.5 10362.5 51377.5 ;
      RECT  10107.5 51242.5 10172.5 51377.5 ;
      RECT  10297.5 51242.5 10362.5 51377.5 ;
      RECT  10487.5 51242.5 10552.5 51377.5 ;
      RECT  10487.5 51242.5 10552.5 51377.5 ;
      RECT  10297.5 51242.5 10362.5 51377.5 ;
      RECT  10107.5 50402.5 10172.5 50537.5 ;
      RECT  10297.5 50402.5 10362.5 50537.5 ;
      RECT  10297.5 50402.5 10362.5 50537.5 ;
      RECT  10107.5 50402.5 10172.5 50537.5 ;
      RECT  10297.5 50402.5 10362.5 50537.5 ;
      RECT  10487.5 50402.5 10552.5 50537.5 ;
      RECT  10487.5 50402.5 10552.5 50537.5 ;
      RECT  10297.5 50402.5 10362.5 50537.5 ;
      RECT  10657.5 51332.5 10722.5 51467.5 ;
      RECT  10657.5 50357.5 10722.5 50492.5 ;
      RECT  10492.5 50632.5 10357.5 50697.5 ;
      RECT  10235.0 50847.5 10100.0 50912.5 ;
      RECT  10297.5 51242.5 10362.5 51377.5 ;
      RECT  10487.5 50402.5 10552.5 50537.5 ;
      RECT  10587.5 50847.5 10452.5 50912.5 ;
      RECT  10100.0 50847.5 10235.0 50912.5 ;
      RECT  10357.5 50632.5 10492.5 50697.5 ;
      RECT  10452.5 50847.5 10587.5 50912.5 ;
      RECT  10040.0 51552.5 10960.0 51617.5 ;
      RECT  10040.0 50207.5 10960.0 50272.5 ;
      RECT  11387.5 51400.0 11452.5 51585.0 ;
      RECT  11387.5 50240.0 11452.5 50425.0 ;
      RECT  11027.5 50357.5 11092.5 50207.5 ;
      RECT  11027.5 51242.5 11092.5 51617.5 ;
      RECT  11217.5 50357.5 11282.5 51242.5 ;
      RECT  11027.5 51242.5 11092.5 51377.5 ;
      RECT  11217.5 51242.5 11282.5 51377.5 ;
      RECT  11217.5 51242.5 11282.5 51377.5 ;
      RECT  11027.5 51242.5 11092.5 51377.5 ;
      RECT  11027.5 50357.5 11092.5 50492.5 ;
      RECT  11217.5 50357.5 11282.5 50492.5 ;
      RECT  11217.5 50357.5 11282.5 50492.5 ;
      RECT  11027.5 50357.5 11092.5 50492.5 ;
      RECT  11387.5 51332.5 11452.5 51467.5 ;
      RECT  11387.5 50357.5 11452.5 50492.5 ;
      RECT  11085.0 50800.0 11150.0 50935.0 ;
      RECT  11085.0 50800.0 11150.0 50935.0 ;
      RECT  11250.0 50835.0 11315.0 50900.0 ;
      RECT  10960.0 51552.5 11520.0 51617.5 ;
      RECT  10960.0 50207.5 11520.0 50272.5 ;
      RECT  9222.5 50800.0 9287.5 50935.0 ;
      RECT  9362.5 50527.5 9427.5 50662.5 ;
      RECT  10357.5 50632.5 10222.5 50697.5 ;
      RECT  9907.5 51770.0 9972.5 51585.0 ;
      RECT  9907.5 52930.0 9972.5 52745.0 ;
      RECT  9547.5 52812.5 9612.5 52962.5 ;
      RECT  9547.5 51927.5 9612.5 51552.5 ;
      RECT  9737.5 52812.5 9802.5 51927.5 ;
      RECT  9547.5 51927.5 9612.5 51792.5 ;
      RECT  9737.5 51927.5 9802.5 51792.5 ;
      RECT  9737.5 51927.5 9802.5 51792.5 ;
      RECT  9547.5 51927.5 9612.5 51792.5 ;
      RECT  9547.5 52812.5 9612.5 52677.5 ;
      RECT  9737.5 52812.5 9802.5 52677.5 ;
      RECT  9737.5 52812.5 9802.5 52677.5 ;
      RECT  9547.5 52812.5 9612.5 52677.5 ;
      RECT  9907.5 51837.5 9972.5 51702.5 ;
      RECT  9907.5 52812.5 9972.5 52677.5 ;
      RECT  9605.0 52370.0 9670.0 52235.0 ;
      RECT  9605.0 52370.0 9670.0 52235.0 ;
      RECT  9770.0 52335.0 9835.0 52270.0 ;
      RECT  9480.0 51617.5 10040.0 51552.5 ;
      RECT  9480.0 52962.5 10040.0 52897.5 ;
      RECT  10107.5 52767.5 10172.5 52962.5 ;
      RECT  10107.5 51927.5 10172.5 51552.5 ;
      RECT  10487.5 51927.5 10552.5 51552.5 ;
      RECT  10657.5 51770.0 10722.5 51585.0 ;
      RECT  10657.5 52930.0 10722.5 52745.0 ;
      RECT  10107.5 51927.5 10172.5 51792.5 ;
      RECT  10297.5 51927.5 10362.5 51792.5 ;
      RECT  10297.5 51927.5 10362.5 51792.5 ;
      RECT  10107.5 51927.5 10172.5 51792.5 ;
      RECT  10297.5 51927.5 10362.5 51792.5 ;
      RECT  10487.5 51927.5 10552.5 51792.5 ;
      RECT  10487.5 51927.5 10552.5 51792.5 ;
      RECT  10297.5 51927.5 10362.5 51792.5 ;
      RECT  10107.5 52767.5 10172.5 52632.5 ;
      RECT  10297.5 52767.5 10362.5 52632.5 ;
      RECT  10297.5 52767.5 10362.5 52632.5 ;
      RECT  10107.5 52767.5 10172.5 52632.5 ;
      RECT  10297.5 52767.5 10362.5 52632.5 ;
      RECT  10487.5 52767.5 10552.5 52632.5 ;
      RECT  10487.5 52767.5 10552.5 52632.5 ;
      RECT  10297.5 52767.5 10362.5 52632.5 ;
      RECT  10657.5 51837.5 10722.5 51702.5 ;
      RECT  10657.5 52812.5 10722.5 52677.5 ;
      RECT  10492.5 52537.5 10357.5 52472.5 ;
      RECT  10235.0 52322.5 10100.0 52257.5 ;
      RECT  10297.5 51927.5 10362.5 51792.5 ;
      RECT  10487.5 52767.5 10552.5 52632.5 ;
      RECT  10587.5 52322.5 10452.5 52257.5 ;
      RECT  10100.0 52322.5 10235.0 52257.5 ;
      RECT  10357.5 52537.5 10492.5 52472.5 ;
      RECT  10452.5 52322.5 10587.5 52257.5 ;
      RECT  10040.0 51617.5 10960.0 51552.5 ;
      RECT  10040.0 52962.5 10960.0 52897.5 ;
      RECT  11387.5 51770.0 11452.5 51585.0 ;
      RECT  11387.5 52930.0 11452.5 52745.0 ;
      RECT  11027.5 52812.5 11092.5 52962.5 ;
      RECT  11027.5 51927.5 11092.5 51552.5 ;
      RECT  11217.5 52812.5 11282.5 51927.5 ;
      RECT  11027.5 51927.5 11092.5 51792.5 ;
      RECT  11217.5 51927.5 11282.5 51792.5 ;
      RECT  11217.5 51927.5 11282.5 51792.5 ;
      RECT  11027.5 51927.5 11092.5 51792.5 ;
      RECT  11027.5 52812.5 11092.5 52677.5 ;
      RECT  11217.5 52812.5 11282.5 52677.5 ;
      RECT  11217.5 52812.5 11282.5 52677.5 ;
      RECT  11027.5 52812.5 11092.5 52677.5 ;
      RECT  11387.5 51837.5 11452.5 51702.5 ;
      RECT  11387.5 52812.5 11452.5 52677.5 ;
      RECT  11085.0 52370.0 11150.0 52235.0 ;
      RECT  11085.0 52370.0 11150.0 52235.0 ;
      RECT  11250.0 52335.0 11315.0 52270.0 ;
      RECT  10960.0 51617.5 11520.0 51552.5 ;
      RECT  10960.0 52962.5 11520.0 52897.5 ;
      RECT  9222.5 52235.0 9287.5 52370.0 ;
      RECT  9362.5 52507.5 9427.5 52642.5 ;
      RECT  10357.5 52472.5 10222.5 52537.5 ;
      RECT  9907.5 54090.0 9972.5 54275.0 ;
      RECT  9907.5 52930.0 9972.5 53115.0 ;
      RECT  9547.5 53047.5 9612.5 52897.5 ;
      RECT  9547.5 53932.5 9612.5 54307.5 ;
      RECT  9737.5 53047.5 9802.5 53932.5 ;
      RECT  9547.5 53932.5 9612.5 54067.5 ;
      RECT  9737.5 53932.5 9802.5 54067.5 ;
      RECT  9737.5 53932.5 9802.5 54067.5 ;
      RECT  9547.5 53932.5 9612.5 54067.5 ;
      RECT  9547.5 53047.5 9612.5 53182.5 ;
      RECT  9737.5 53047.5 9802.5 53182.5 ;
      RECT  9737.5 53047.5 9802.5 53182.5 ;
      RECT  9547.5 53047.5 9612.5 53182.5 ;
      RECT  9907.5 54022.5 9972.5 54157.5 ;
      RECT  9907.5 53047.5 9972.5 53182.5 ;
      RECT  9605.0 53490.0 9670.0 53625.0 ;
      RECT  9605.0 53490.0 9670.0 53625.0 ;
      RECT  9770.0 53525.0 9835.0 53590.0 ;
      RECT  9480.0 54242.5 10040.0 54307.5 ;
      RECT  9480.0 52897.5 10040.0 52962.5 ;
      RECT  10107.5 53092.5 10172.5 52897.5 ;
      RECT  10107.5 53932.5 10172.5 54307.5 ;
      RECT  10487.5 53932.5 10552.5 54307.5 ;
      RECT  10657.5 54090.0 10722.5 54275.0 ;
      RECT  10657.5 52930.0 10722.5 53115.0 ;
      RECT  10107.5 53932.5 10172.5 54067.5 ;
      RECT  10297.5 53932.5 10362.5 54067.5 ;
      RECT  10297.5 53932.5 10362.5 54067.5 ;
      RECT  10107.5 53932.5 10172.5 54067.5 ;
      RECT  10297.5 53932.5 10362.5 54067.5 ;
      RECT  10487.5 53932.5 10552.5 54067.5 ;
      RECT  10487.5 53932.5 10552.5 54067.5 ;
      RECT  10297.5 53932.5 10362.5 54067.5 ;
      RECT  10107.5 53092.5 10172.5 53227.5 ;
      RECT  10297.5 53092.5 10362.5 53227.5 ;
      RECT  10297.5 53092.5 10362.5 53227.5 ;
      RECT  10107.5 53092.5 10172.5 53227.5 ;
      RECT  10297.5 53092.5 10362.5 53227.5 ;
      RECT  10487.5 53092.5 10552.5 53227.5 ;
      RECT  10487.5 53092.5 10552.5 53227.5 ;
      RECT  10297.5 53092.5 10362.5 53227.5 ;
      RECT  10657.5 54022.5 10722.5 54157.5 ;
      RECT  10657.5 53047.5 10722.5 53182.5 ;
      RECT  10492.5 53322.5 10357.5 53387.5 ;
      RECT  10235.0 53537.5 10100.0 53602.5 ;
      RECT  10297.5 53932.5 10362.5 54067.5 ;
      RECT  10487.5 53092.5 10552.5 53227.5 ;
      RECT  10587.5 53537.5 10452.5 53602.5 ;
      RECT  10100.0 53537.5 10235.0 53602.5 ;
      RECT  10357.5 53322.5 10492.5 53387.5 ;
      RECT  10452.5 53537.5 10587.5 53602.5 ;
      RECT  10040.0 54242.5 10960.0 54307.5 ;
      RECT  10040.0 52897.5 10960.0 52962.5 ;
      RECT  11387.5 54090.0 11452.5 54275.0 ;
      RECT  11387.5 52930.0 11452.5 53115.0 ;
      RECT  11027.5 53047.5 11092.5 52897.5 ;
      RECT  11027.5 53932.5 11092.5 54307.5 ;
      RECT  11217.5 53047.5 11282.5 53932.5 ;
      RECT  11027.5 53932.5 11092.5 54067.5 ;
      RECT  11217.5 53932.5 11282.5 54067.5 ;
      RECT  11217.5 53932.5 11282.5 54067.5 ;
      RECT  11027.5 53932.5 11092.5 54067.5 ;
      RECT  11027.5 53047.5 11092.5 53182.5 ;
      RECT  11217.5 53047.5 11282.5 53182.5 ;
      RECT  11217.5 53047.5 11282.5 53182.5 ;
      RECT  11027.5 53047.5 11092.5 53182.5 ;
      RECT  11387.5 54022.5 11452.5 54157.5 ;
      RECT  11387.5 53047.5 11452.5 53182.5 ;
      RECT  11085.0 53490.0 11150.0 53625.0 ;
      RECT  11085.0 53490.0 11150.0 53625.0 ;
      RECT  11250.0 53525.0 11315.0 53590.0 ;
      RECT  10960.0 54242.5 11520.0 54307.5 ;
      RECT  10960.0 52897.5 11520.0 52962.5 ;
      RECT  9222.5 53490.0 9287.5 53625.0 ;
      RECT  9362.5 53217.5 9427.5 53352.5 ;
      RECT  10357.5 53322.5 10222.5 53387.5 ;
      RECT  9907.5 54460.0 9972.5 54275.0 ;
      RECT  9907.5 55620.0 9972.5 55435.0 ;
      RECT  9547.5 55502.5 9612.5 55652.5 ;
      RECT  9547.5 54617.5 9612.5 54242.5 ;
      RECT  9737.5 55502.5 9802.5 54617.5 ;
      RECT  9547.5 54617.5 9612.5 54482.5 ;
      RECT  9737.5 54617.5 9802.5 54482.5 ;
      RECT  9737.5 54617.5 9802.5 54482.5 ;
      RECT  9547.5 54617.5 9612.5 54482.5 ;
      RECT  9547.5 55502.5 9612.5 55367.5 ;
      RECT  9737.5 55502.5 9802.5 55367.5 ;
      RECT  9737.5 55502.5 9802.5 55367.5 ;
      RECT  9547.5 55502.5 9612.5 55367.5 ;
      RECT  9907.5 54527.5 9972.5 54392.5 ;
      RECT  9907.5 55502.5 9972.5 55367.5 ;
      RECT  9605.0 55060.0 9670.0 54925.0 ;
      RECT  9605.0 55060.0 9670.0 54925.0 ;
      RECT  9770.0 55025.0 9835.0 54960.0 ;
      RECT  9480.0 54307.5 10040.0 54242.5 ;
      RECT  9480.0 55652.5 10040.0 55587.5 ;
      RECT  10107.5 55457.5 10172.5 55652.5 ;
      RECT  10107.5 54617.5 10172.5 54242.5 ;
      RECT  10487.5 54617.5 10552.5 54242.5 ;
      RECT  10657.5 54460.0 10722.5 54275.0 ;
      RECT  10657.5 55620.0 10722.5 55435.0 ;
      RECT  10107.5 54617.5 10172.5 54482.5 ;
      RECT  10297.5 54617.5 10362.5 54482.5 ;
      RECT  10297.5 54617.5 10362.5 54482.5 ;
      RECT  10107.5 54617.5 10172.5 54482.5 ;
      RECT  10297.5 54617.5 10362.5 54482.5 ;
      RECT  10487.5 54617.5 10552.5 54482.5 ;
      RECT  10487.5 54617.5 10552.5 54482.5 ;
      RECT  10297.5 54617.5 10362.5 54482.5 ;
      RECT  10107.5 55457.5 10172.5 55322.5 ;
      RECT  10297.5 55457.5 10362.5 55322.5 ;
      RECT  10297.5 55457.5 10362.5 55322.5 ;
      RECT  10107.5 55457.5 10172.5 55322.5 ;
      RECT  10297.5 55457.5 10362.5 55322.5 ;
      RECT  10487.5 55457.5 10552.5 55322.5 ;
      RECT  10487.5 55457.5 10552.5 55322.5 ;
      RECT  10297.5 55457.5 10362.5 55322.5 ;
      RECT  10657.5 54527.5 10722.5 54392.5 ;
      RECT  10657.5 55502.5 10722.5 55367.5 ;
      RECT  10492.5 55227.5 10357.5 55162.5 ;
      RECT  10235.0 55012.5 10100.0 54947.5 ;
      RECT  10297.5 54617.5 10362.5 54482.5 ;
      RECT  10487.5 55457.5 10552.5 55322.5 ;
      RECT  10587.5 55012.5 10452.5 54947.5 ;
      RECT  10100.0 55012.5 10235.0 54947.5 ;
      RECT  10357.5 55227.5 10492.5 55162.5 ;
      RECT  10452.5 55012.5 10587.5 54947.5 ;
      RECT  10040.0 54307.5 10960.0 54242.5 ;
      RECT  10040.0 55652.5 10960.0 55587.5 ;
      RECT  11387.5 54460.0 11452.5 54275.0 ;
      RECT  11387.5 55620.0 11452.5 55435.0 ;
      RECT  11027.5 55502.5 11092.5 55652.5 ;
      RECT  11027.5 54617.5 11092.5 54242.5 ;
      RECT  11217.5 55502.5 11282.5 54617.5 ;
      RECT  11027.5 54617.5 11092.5 54482.5 ;
      RECT  11217.5 54617.5 11282.5 54482.5 ;
      RECT  11217.5 54617.5 11282.5 54482.5 ;
      RECT  11027.5 54617.5 11092.5 54482.5 ;
      RECT  11027.5 55502.5 11092.5 55367.5 ;
      RECT  11217.5 55502.5 11282.5 55367.5 ;
      RECT  11217.5 55502.5 11282.5 55367.5 ;
      RECT  11027.5 55502.5 11092.5 55367.5 ;
      RECT  11387.5 54527.5 11452.5 54392.5 ;
      RECT  11387.5 55502.5 11452.5 55367.5 ;
      RECT  11085.0 55060.0 11150.0 54925.0 ;
      RECT  11085.0 55060.0 11150.0 54925.0 ;
      RECT  11250.0 55025.0 11315.0 54960.0 ;
      RECT  10960.0 54307.5 11520.0 54242.5 ;
      RECT  10960.0 55652.5 11520.0 55587.5 ;
      RECT  9222.5 54925.0 9287.5 55060.0 ;
      RECT  9362.5 55197.5 9427.5 55332.5 ;
      RECT  10357.5 55162.5 10222.5 55227.5 ;
      RECT  9907.5 56780.0 9972.5 56965.0 ;
      RECT  9907.5 55620.0 9972.5 55805.0 ;
      RECT  9547.5 55737.5 9612.5 55587.5 ;
      RECT  9547.5 56622.5 9612.5 56997.5 ;
      RECT  9737.5 55737.5 9802.5 56622.5 ;
      RECT  9547.5 56622.5 9612.5 56757.5 ;
      RECT  9737.5 56622.5 9802.5 56757.5 ;
      RECT  9737.5 56622.5 9802.5 56757.5 ;
      RECT  9547.5 56622.5 9612.5 56757.5 ;
      RECT  9547.5 55737.5 9612.5 55872.5 ;
      RECT  9737.5 55737.5 9802.5 55872.5 ;
      RECT  9737.5 55737.5 9802.5 55872.5 ;
      RECT  9547.5 55737.5 9612.5 55872.5 ;
      RECT  9907.5 56712.5 9972.5 56847.5 ;
      RECT  9907.5 55737.5 9972.5 55872.5 ;
      RECT  9605.0 56180.0 9670.0 56315.0 ;
      RECT  9605.0 56180.0 9670.0 56315.0 ;
      RECT  9770.0 56215.0 9835.0 56280.0 ;
      RECT  9480.0 56932.5 10040.0 56997.5 ;
      RECT  9480.0 55587.5 10040.0 55652.5 ;
      RECT  10107.5 55782.5 10172.5 55587.5 ;
      RECT  10107.5 56622.5 10172.5 56997.5 ;
      RECT  10487.5 56622.5 10552.5 56997.5 ;
      RECT  10657.5 56780.0 10722.5 56965.0 ;
      RECT  10657.5 55620.0 10722.5 55805.0 ;
      RECT  10107.5 56622.5 10172.5 56757.5 ;
      RECT  10297.5 56622.5 10362.5 56757.5 ;
      RECT  10297.5 56622.5 10362.5 56757.5 ;
      RECT  10107.5 56622.5 10172.5 56757.5 ;
      RECT  10297.5 56622.5 10362.5 56757.5 ;
      RECT  10487.5 56622.5 10552.5 56757.5 ;
      RECT  10487.5 56622.5 10552.5 56757.5 ;
      RECT  10297.5 56622.5 10362.5 56757.5 ;
      RECT  10107.5 55782.5 10172.5 55917.5 ;
      RECT  10297.5 55782.5 10362.5 55917.5 ;
      RECT  10297.5 55782.5 10362.5 55917.5 ;
      RECT  10107.5 55782.5 10172.5 55917.5 ;
      RECT  10297.5 55782.5 10362.5 55917.5 ;
      RECT  10487.5 55782.5 10552.5 55917.5 ;
      RECT  10487.5 55782.5 10552.5 55917.5 ;
      RECT  10297.5 55782.5 10362.5 55917.5 ;
      RECT  10657.5 56712.5 10722.5 56847.5 ;
      RECT  10657.5 55737.5 10722.5 55872.5 ;
      RECT  10492.5 56012.5 10357.5 56077.5 ;
      RECT  10235.0 56227.5 10100.0 56292.5 ;
      RECT  10297.5 56622.5 10362.5 56757.5 ;
      RECT  10487.5 55782.5 10552.5 55917.5 ;
      RECT  10587.5 56227.5 10452.5 56292.5 ;
      RECT  10100.0 56227.5 10235.0 56292.5 ;
      RECT  10357.5 56012.5 10492.5 56077.5 ;
      RECT  10452.5 56227.5 10587.5 56292.5 ;
      RECT  10040.0 56932.5 10960.0 56997.5 ;
      RECT  10040.0 55587.5 10960.0 55652.5 ;
      RECT  11387.5 56780.0 11452.5 56965.0 ;
      RECT  11387.5 55620.0 11452.5 55805.0 ;
      RECT  11027.5 55737.5 11092.5 55587.5 ;
      RECT  11027.5 56622.5 11092.5 56997.5 ;
      RECT  11217.5 55737.5 11282.5 56622.5 ;
      RECT  11027.5 56622.5 11092.5 56757.5 ;
      RECT  11217.5 56622.5 11282.5 56757.5 ;
      RECT  11217.5 56622.5 11282.5 56757.5 ;
      RECT  11027.5 56622.5 11092.5 56757.5 ;
      RECT  11027.5 55737.5 11092.5 55872.5 ;
      RECT  11217.5 55737.5 11282.5 55872.5 ;
      RECT  11217.5 55737.5 11282.5 55872.5 ;
      RECT  11027.5 55737.5 11092.5 55872.5 ;
      RECT  11387.5 56712.5 11452.5 56847.5 ;
      RECT  11387.5 55737.5 11452.5 55872.5 ;
      RECT  11085.0 56180.0 11150.0 56315.0 ;
      RECT  11085.0 56180.0 11150.0 56315.0 ;
      RECT  11250.0 56215.0 11315.0 56280.0 ;
      RECT  10960.0 56932.5 11520.0 56997.5 ;
      RECT  10960.0 55587.5 11520.0 55652.5 ;
      RECT  9222.5 56180.0 9287.5 56315.0 ;
      RECT  9362.5 55907.5 9427.5 56042.5 ;
      RECT  10357.5 56012.5 10222.5 56077.5 ;
      RECT  9907.5 57150.0 9972.5 56965.0 ;
      RECT  9907.5 58310.0 9972.5 58125.0 ;
      RECT  9547.5 58192.5 9612.5 58342.5 ;
      RECT  9547.5 57307.5 9612.5 56932.5 ;
      RECT  9737.5 58192.5 9802.5 57307.5 ;
      RECT  9547.5 57307.5 9612.5 57172.5 ;
      RECT  9737.5 57307.5 9802.5 57172.5 ;
      RECT  9737.5 57307.5 9802.5 57172.5 ;
      RECT  9547.5 57307.5 9612.5 57172.5 ;
      RECT  9547.5 58192.5 9612.5 58057.5 ;
      RECT  9737.5 58192.5 9802.5 58057.5 ;
      RECT  9737.5 58192.5 9802.5 58057.5 ;
      RECT  9547.5 58192.5 9612.5 58057.5 ;
      RECT  9907.5 57217.5 9972.5 57082.5 ;
      RECT  9907.5 58192.5 9972.5 58057.5 ;
      RECT  9605.0 57750.0 9670.0 57615.0 ;
      RECT  9605.0 57750.0 9670.0 57615.0 ;
      RECT  9770.0 57715.0 9835.0 57650.0 ;
      RECT  9480.0 56997.5 10040.0 56932.5 ;
      RECT  9480.0 58342.5 10040.0 58277.5 ;
      RECT  10107.5 58147.5 10172.5 58342.5 ;
      RECT  10107.5 57307.5 10172.5 56932.5 ;
      RECT  10487.5 57307.5 10552.5 56932.5 ;
      RECT  10657.5 57150.0 10722.5 56965.0 ;
      RECT  10657.5 58310.0 10722.5 58125.0 ;
      RECT  10107.5 57307.5 10172.5 57172.5 ;
      RECT  10297.5 57307.5 10362.5 57172.5 ;
      RECT  10297.5 57307.5 10362.5 57172.5 ;
      RECT  10107.5 57307.5 10172.5 57172.5 ;
      RECT  10297.5 57307.5 10362.5 57172.5 ;
      RECT  10487.5 57307.5 10552.5 57172.5 ;
      RECT  10487.5 57307.5 10552.5 57172.5 ;
      RECT  10297.5 57307.5 10362.5 57172.5 ;
      RECT  10107.5 58147.5 10172.5 58012.5 ;
      RECT  10297.5 58147.5 10362.5 58012.5 ;
      RECT  10297.5 58147.5 10362.5 58012.5 ;
      RECT  10107.5 58147.5 10172.5 58012.5 ;
      RECT  10297.5 58147.5 10362.5 58012.5 ;
      RECT  10487.5 58147.5 10552.5 58012.5 ;
      RECT  10487.5 58147.5 10552.5 58012.5 ;
      RECT  10297.5 58147.5 10362.5 58012.5 ;
      RECT  10657.5 57217.5 10722.5 57082.5 ;
      RECT  10657.5 58192.5 10722.5 58057.5 ;
      RECT  10492.5 57917.5 10357.5 57852.5 ;
      RECT  10235.0 57702.5 10100.0 57637.5 ;
      RECT  10297.5 57307.5 10362.5 57172.5 ;
      RECT  10487.5 58147.5 10552.5 58012.5 ;
      RECT  10587.5 57702.5 10452.5 57637.5 ;
      RECT  10100.0 57702.5 10235.0 57637.5 ;
      RECT  10357.5 57917.5 10492.5 57852.5 ;
      RECT  10452.5 57702.5 10587.5 57637.5 ;
      RECT  10040.0 56997.5 10960.0 56932.5 ;
      RECT  10040.0 58342.5 10960.0 58277.5 ;
      RECT  11387.5 57150.0 11452.5 56965.0 ;
      RECT  11387.5 58310.0 11452.5 58125.0 ;
      RECT  11027.5 58192.5 11092.5 58342.5 ;
      RECT  11027.5 57307.5 11092.5 56932.5 ;
      RECT  11217.5 58192.5 11282.5 57307.5 ;
      RECT  11027.5 57307.5 11092.5 57172.5 ;
      RECT  11217.5 57307.5 11282.5 57172.5 ;
      RECT  11217.5 57307.5 11282.5 57172.5 ;
      RECT  11027.5 57307.5 11092.5 57172.5 ;
      RECT  11027.5 58192.5 11092.5 58057.5 ;
      RECT  11217.5 58192.5 11282.5 58057.5 ;
      RECT  11217.5 58192.5 11282.5 58057.5 ;
      RECT  11027.5 58192.5 11092.5 58057.5 ;
      RECT  11387.5 57217.5 11452.5 57082.5 ;
      RECT  11387.5 58192.5 11452.5 58057.5 ;
      RECT  11085.0 57750.0 11150.0 57615.0 ;
      RECT  11085.0 57750.0 11150.0 57615.0 ;
      RECT  11250.0 57715.0 11315.0 57650.0 ;
      RECT  10960.0 56997.5 11520.0 56932.5 ;
      RECT  10960.0 58342.5 11520.0 58277.5 ;
      RECT  9222.5 57615.0 9287.5 57750.0 ;
      RECT  9362.5 57887.5 9427.5 58022.5 ;
      RECT  10357.5 57852.5 10222.5 57917.5 ;
      RECT  9907.5 59470.0 9972.5 59655.0 ;
      RECT  9907.5 58310.0 9972.5 58495.0 ;
      RECT  9547.5 58427.5 9612.5 58277.5 ;
      RECT  9547.5 59312.5 9612.5 59687.5 ;
      RECT  9737.5 58427.5 9802.5 59312.5 ;
      RECT  9547.5 59312.5 9612.5 59447.5 ;
      RECT  9737.5 59312.5 9802.5 59447.5 ;
      RECT  9737.5 59312.5 9802.5 59447.5 ;
      RECT  9547.5 59312.5 9612.5 59447.5 ;
      RECT  9547.5 58427.5 9612.5 58562.5 ;
      RECT  9737.5 58427.5 9802.5 58562.5 ;
      RECT  9737.5 58427.5 9802.5 58562.5 ;
      RECT  9547.5 58427.5 9612.5 58562.5 ;
      RECT  9907.5 59402.5 9972.5 59537.5 ;
      RECT  9907.5 58427.5 9972.5 58562.5 ;
      RECT  9605.0 58870.0 9670.0 59005.0 ;
      RECT  9605.0 58870.0 9670.0 59005.0 ;
      RECT  9770.0 58905.0 9835.0 58970.0 ;
      RECT  9480.0 59622.5 10040.0 59687.5 ;
      RECT  9480.0 58277.5 10040.0 58342.5 ;
      RECT  10107.5 58472.5 10172.5 58277.5 ;
      RECT  10107.5 59312.5 10172.5 59687.5 ;
      RECT  10487.5 59312.5 10552.5 59687.5 ;
      RECT  10657.5 59470.0 10722.5 59655.0 ;
      RECT  10657.5 58310.0 10722.5 58495.0 ;
      RECT  10107.5 59312.5 10172.5 59447.5 ;
      RECT  10297.5 59312.5 10362.5 59447.5 ;
      RECT  10297.5 59312.5 10362.5 59447.5 ;
      RECT  10107.5 59312.5 10172.5 59447.5 ;
      RECT  10297.5 59312.5 10362.5 59447.5 ;
      RECT  10487.5 59312.5 10552.5 59447.5 ;
      RECT  10487.5 59312.5 10552.5 59447.5 ;
      RECT  10297.5 59312.5 10362.5 59447.5 ;
      RECT  10107.5 58472.5 10172.5 58607.5 ;
      RECT  10297.5 58472.5 10362.5 58607.5 ;
      RECT  10297.5 58472.5 10362.5 58607.5 ;
      RECT  10107.5 58472.5 10172.5 58607.5 ;
      RECT  10297.5 58472.5 10362.5 58607.5 ;
      RECT  10487.5 58472.5 10552.5 58607.5 ;
      RECT  10487.5 58472.5 10552.5 58607.5 ;
      RECT  10297.5 58472.5 10362.5 58607.5 ;
      RECT  10657.5 59402.5 10722.5 59537.5 ;
      RECT  10657.5 58427.5 10722.5 58562.5 ;
      RECT  10492.5 58702.5 10357.5 58767.5 ;
      RECT  10235.0 58917.5 10100.0 58982.5 ;
      RECT  10297.5 59312.5 10362.5 59447.5 ;
      RECT  10487.5 58472.5 10552.5 58607.5 ;
      RECT  10587.5 58917.5 10452.5 58982.5 ;
      RECT  10100.0 58917.5 10235.0 58982.5 ;
      RECT  10357.5 58702.5 10492.5 58767.5 ;
      RECT  10452.5 58917.5 10587.5 58982.5 ;
      RECT  10040.0 59622.5 10960.0 59687.5 ;
      RECT  10040.0 58277.5 10960.0 58342.5 ;
      RECT  11387.5 59470.0 11452.5 59655.0 ;
      RECT  11387.5 58310.0 11452.5 58495.0 ;
      RECT  11027.5 58427.5 11092.5 58277.5 ;
      RECT  11027.5 59312.5 11092.5 59687.5 ;
      RECT  11217.5 58427.5 11282.5 59312.5 ;
      RECT  11027.5 59312.5 11092.5 59447.5 ;
      RECT  11217.5 59312.5 11282.5 59447.5 ;
      RECT  11217.5 59312.5 11282.5 59447.5 ;
      RECT  11027.5 59312.5 11092.5 59447.5 ;
      RECT  11027.5 58427.5 11092.5 58562.5 ;
      RECT  11217.5 58427.5 11282.5 58562.5 ;
      RECT  11217.5 58427.5 11282.5 58562.5 ;
      RECT  11027.5 58427.5 11092.5 58562.5 ;
      RECT  11387.5 59402.5 11452.5 59537.5 ;
      RECT  11387.5 58427.5 11452.5 58562.5 ;
      RECT  11085.0 58870.0 11150.0 59005.0 ;
      RECT  11085.0 58870.0 11150.0 59005.0 ;
      RECT  11250.0 58905.0 11315.0 58970.0 ;
      RECT  10960.0 59622.5 11520.0 59687.5 ;
      RECT  10960.0 58277.5 11520.0 58342.5 ;
      RECT  9222.5 58870.0 9287.5 59005.0 ;
      RECT  9362.5 58597.5 9427.5 58732.5 ;
      RECT  10357.5 58702.5 10222.5 58767.5 ;
      RECT  9907.5 59840.0 9972.5 59655.0 ;
      RECT  9907.5 61000.0 9972.5 60815.0 ;
      RECT  9547.5 60882.5 9612.5 61032.5 ;
      RECT  9547.5 59997.5 9612.5 59622.5 ;
      RECT  9737.5 60882.5 9802.5 59997.5 ;
      RECT  9547.5 59997.5 9612.5 59862.5 ;
      RECT  9737.5 59997.5 9802.5 59862.5 ;
      RECT  9737.5 59997.5 9802.5 59862.5 ;
      RECT  9547.5 59997.5 9612.5 59862.5 ;
      RECT  9547.5 60882.5 9612.5 60747.5 ;
      RECT  9737.5 60882.5 9802.5 60747.5 ;
      RECT  9737.5 60882.5 9802.5 60747.5 ;
      RECT  9547.5 60882.5 9612.5 60747.5 ;
      RECT  9907.5 59907.5 9972.5 59772.5 ;
      RECT  9907.5 60882.5 9972.5 60747.5 ;
      RECT  9605.0 60440.0 9670.0 60305.0 ;
      RECT  9605.0 60440.0 9670.0 60305.0 ;
      RECT  9770.0 60405.0 9835.0 60340.0 ;
      RECT  9480.0 59687.5 10040.0 59622.5 ;
      RECT  9480.0 61032.5 10040.0 60967.5 ;
      RECT  10107.5 60837.5 10172.5 61032.5 ;
      RECT  10107.5 59997.5 10172.5 59622.5 ;
      RECT  10487.5 59997.5 10552.5 59622.5 ;
      RECT  10657.5 59840.0 10722.5 59655.0 ;
      RECT  10657.5 61000.0 10722.5 60815.0 ;
      RECT  10107.5 59997.5 10172.5 59862.5 ;
      RECT  10297.5 59997.5 10362.5 59862.5 ;
      RECT  10297.5 59997.5 10362.5 59862.5 ;
      RECT  10107.5 59997.5 10172.5 59862.5 ;
      RECT  10297.5 59997.5 10362.5 59862.5 ;
      RECT  10487.5 59997.5 10552.5 59862.5 ;
      RECT  10487.5 59997.5 10552.5 59862.5 ;
      RECT  10297.5 59997.5 10362.5 59862.5 ;
      RECT  10107.5 60837.5 10172.5 60702.5 ;
      RECT  10297.5 60837.5 10362.5 60702.5 ;
      RECT  10297.5 60837.5 10362.5 60702.5 ;
      RECT  10107.5 60837.5 10172.5 60702.5 ;
      RECT  10297.5 60837.5 10362.5 60702.5 ;
      RECT  10487.5 60837.5 10552.5 60702.5 ;
      RECT  10487.5 60837.5 10552.5 60702.5 ;
      RECT  10297.5 60837.5 10362.5 60702.5 ;
      RECT  10657.5 59907.5 10722.5 59772.5 ;
      RECT  10657.5 60882.5 10722.5 60747.5 ;
      RECT  10492.5 60607.5 10357.5 60542.5 ;
      RECT  10235.0 60392.5 10100.0 60327.5 ;
      RECT  10297.5 59997.5 10362.5 59862.5 ;
      RECT  10487.5 60837.5 10552.5 60702.5 ;
      RECT  10587.5 60392.5 10452.5 60327.5 ;
      RECT  10100.0 60392.5 10235.0 60327.5 ;
      RECT  10357.5 60607.5 10492.5 60542.5 ;
      RECT  10452.5 60392.5 10587.5 60327.5 ;
      RECT  10040.0 59687.5 10960.0 59622.5 ;
      RECT  10040.0 61032.5 10960.0 60967.5 ;
      RECT  11387.5 59840.0 11452.5 59655.0 ;
      RECT  11387.5 61000.0 11452.5 60815.0 ;
      RECT  11027.5 60882.5 11092.5 61032.5 ;
      RECT  11027.5 59997.5 11092.5 59622.5 ;
      RECT  11217.5 60882.5 11282.5 59997.5 ;
      RECT  11027.5 59997.5 11092.5 59862.5 ;
      RECT  11217.5 59997.5 11282.5 59862.5 ;
      RECT  11217.5 59997.5 11282.5 59862.5 ;
      RECT  11027.5 59997.5 11092.5 59862.5 ;
      RECT  11027.5 60882.5 11092.5 60747.5 ;
      RECT  11217.5 60882.5 11282.5 60747.5 ;
      RECT  11217.5 60882.5 11282.5 60747.5 ;
      RECT  11027.5 60882.5 11092.5 60747.5 ;
      RECT  11387.5 59907.5 11452.5 59772.5 ;
      RECT  11387.5 60882.5 11452.5 60747.5 ;
      RECT  11085.0 60440.0 11150.0 60305.0 ;
      RECT  11085.0 60440.0 11150.0 60305.0 ;
      RECT  11250.0 60405.0 11315.0 60340.0 ;
      RECT  10960.0 59687.5 11520.0 59622.5 ;
      RECT  10960.0 61032.5 11520.0 60967.5 ;
      RECT  9222.5 60305.0 9287.5 60440.0 ;
      RECT  9362.5 60577.5 9427.5 60712.5 ;
      RECT  10357.5 60542.5 10222.5 60607.5 ;
      RECT  9907.5 62160.0 9972.5 62345.0 ;
      RECT  9907.5 61000.0 9972.5 61185.0 ;
      RECT  9547.5 61117.5 9612.5 60967.5 ;
      RECT  9547.5 62002.5 9612.5 62377.5 ;
      RECT  9737.5 61117.5 9802.5 62002.5 ;
      RECT  9547.5 62002.5 9612.5 62137.5 ;
      RECT  9737.5 62002.5 9802.5 62137.5 ;
      RECT  9737.5 62002.5 9802.5 62137.5 ;
      RECT  9547.5 62002.5 9612.5 62137.5 ;
      RECT  9547.5 61117.5 9612.5 61252.5 ;
      RECT  9737.5 61117.5 9802.5 61252.5 ;
      RECT  9737.5 61117.5 9802.5 61252.5 ;
      RECT  9547.5 61117.5 9612.5 61252.5 ;
      RECT  9907.5 62092.5 9972.5 62227.5 ;
      RECT  9907.5 61117.5 9972.5 61252.5 ;
      RECT  9605.0 61560.0 9670.0 61695.0 ;
      RECT  9605.0 61560.0 9670.0 61695.0 ;
      RECT  9770.0 61595.0 9835.0 61660.0 ;
      RECT  9480.0 62312.5 10040.0 62377.5 ;
      RECT  9480.0 60967.5 10040.0 61032.5 ;
      RECT  10107.5 61162.5 10172.5 60967.5 ;
      RECT  10107.5 62002.5 10172.5 62377.5 ;
      RECT  10487.5 62002.5 10552.5 62377.5 ;
      RECT  10657.5 62160.0 10722.5 62345.0 ;
      RECT  10657.5 61000.0 10722.5 61185.0 ;
      RECT  10107.5 62002.5 10172.5 62137.5 ;
      RECT  10297.5 62002.5 10362.5 62137.5 ;
      RECT  10297.5 62002.5 10362.5 62137.5 ;
      RECT  10107.5 62002.5 10172.5 62137.5 ;
      RECT  10297.5 62002.5 10362.5 62137.5 ;
      RECT  10487.5 62002.5 10552.5 62137.5 ;
      RECT  10487.5 62002.5 10552.5 62137.5 ;
      RECT  10297.5 62002.5 10362.5 62137.5 ;
      RECT  10107.5 61162.5 10172.5 61297.5 ;
      RECT  10297.5 61162.5 10362.5 61297.5 ;
      RECT  10297.5 61162.5 10362.5 61297.5 ;
      RECT  10107.5 61162.5 10172.5 61297.5 ;
      RECT  10297.5 61162.5 10362.5 61297.5 ;
      RECT  10487.5 61162.5 10552.5 61297.5 ;
      RECT  10487.5 61162.5 10552.5 61297.5 ;
      RECT  10297.5 61162.5 10362.5 61297.5 ;
      RECT  10657.5 62092.5 10722.5 62227.5 ;
      RECT  10657.5 61117.5 10722.5 61252.5 ;
      RECT  10492.5 61392.5 10357.5 61457.5 ;
      RECT  10235.0 61607.5 10100.0 61672.5 ;
      RECT  10297.5 62002.5 10362.5 62137.5 ;
      RECT  10487.5 61162.5 10552.5 61297.5 ;
      RECT  10587.5 61607.5 10452.5 61672.5 ;
      RECT  10100.0 61607.5 10235.0 61672.5 ;
      RECT  10357.5 61392.5 10492.5 61457.5 ;
      RECT  10452.5 61607.5 10587.5 61672.5 ;
      RECT  10040.0 62312.5 10960.0 62377.5 ;
      RECT  10040.0 60967.5 10960.0 61032.5 ;
      RECT  11387.5 62160.0 11452.5 62345.0 ;
      RECT  11387.5 61000.0 11452.5 61185.0 ;
      RECT  11027.5 61117.5 11092.5 60967.5 ;
      RECT  11027.5 62002.5 11092.5 62377.5 ;
      RECT  11217.5 61117.5 11282.5 62002.5 ;
      RECT  11027.5 62002.5 11092.5 62137.5 ;
      RECT  11217.5 62002.5 11282.5 62137.5 ;
      RECT  11217.5 62002.5 11282.5 62137.5 ;
      RECT  11027.5 62002.5 11092.5 62137.5 ;
      RECT  11027.5 61117.5 11092.5 61252.5 ;
      RECT  11217.5 61117.5 11282.5 61252.5 ;
      RECT  11217.5 61117.5 11282.5 61252.5 ;
      RECT  11027.5 61117.5 11092.5 61252.5 ;
      RECT  11387.5 62092.5 11452.5 62227.5 ;
      RECT  11387.5 61117.5 11452.5 61252.5 ;
      RECT  11085.0 61560.0 11150.0 61695.0 ;
      RECT  11085.0 61560.0 11150.0 61695.0 ;
      RECT  11250.0 61595.0 11315.0 61660.0 ;
      RECT  10960.0 62312.5 11520.0 62377.5 ;
      RECT  10960.0 60967.5 11520.0 61032.5 ;
      RECT  9222.5 61560.0 9287.5 61695.0 ;
      RECT  9362.5 61287.5 9427.5 61422.5 ;
      RECT  10357.5 61392.5 10222.5 61457.5 ;
      RECT  9907.5 62530.0 9972.5 62345.0 ;
      RECT  9907.5 63690.0 9972.5 63505.0 ;
      RECT  9547.5 63572.5 9612.5 63722.5 ;
      RECT  9547.5 62687.5 9612.5 62312.5 ;
      RECT  9737.5 63572.5 9802.5 62687.5 ;
      RECT  9547.5 62687.5 9612.5 62552.5 ;
      RECT  9737.5 62687.5 9802.5 62552.5 ;
      RECT  9737.5 62687.5 9802.5 62552.5 ;
      RECT  9547.5 62687.5 9612.5 62552.5 ;
      RECT  9547.5 63572.5 9612.5 63437.5 ;
      RECT  9737.5 63572.5 9802.5 63437.5 ;
      RECT  9737.5 63572.5 9802.5 63437.5 ;
      RECT  9547.5 63572.5 9612.5 63437.5 ;
      RECT  9907.5 62597.5 9972.5 62462.5 ;
      RECT  9907.5 63572.5 9972.5 63437.5 ;
      RECT  9605.0 63130.0 9670.0 62995.0 ;
      RECT  9605.0 63130.0 9670.0 62995.0 ;
      RECT  9770.0 63095.0 9835.0 63030.0 ;
      RECT  9480.0 62377.5 10040.0 62312.5 ;
      RECT  9480.0 63722.5 10040.0 63657.5 ;
      RECT  10107.5 63527.5 10172.5 63722.5 ;
      RECT  10107.5 62687.5 10172.5 62312.5 ;
      RECT  10487.5 62687.5 10552.5 62312.5 ;
      RECT  10657.5 62530.0 10722.5 62345.0 ;
      RECT  10657.5 63690.0 10722.5 63505.0 ;
      RECT  10107.5 62687.5 10172.5 62552.5 ;
      RECT  10297.5 62687.5 10362.5 62552.5 ;
      RECT  10297.5 62687.5 10362.5 62552.5 ;
      RECT  10107.5 62687.5 10172.5 62552.5 ;
      RECT  10297.5 62687.5 10362.5 62552.5 ;
      RECT  10487.5 62687.5 10552.5 62552.5 ;
      RECT  10487.5 62687.5 10552.5 62552.5 ;
      RECT  10297.5 62687.5 10362.5 62552.5 ;
      RECT  10107.5 63527.5 10172.5 63392.5 ;
      RECT  10297.5 63527.5 10362.5 63392.5 ;
      RECT  10297.5 63527.5 10362.5 63392.5 ;
      RECT  10107.5 63527.5 10172.5 63392.5 ;
      RECT  10297.5 63527.5 10362.5 63392.5 ;
      RECT  10487.5 63527.5 10552.5 63392.5 ;
      RECT  10487.5 63527.5 10552.5 63392.5 ;
      RECT  10297.5 63527.5 10362.5 63392.5 ;
      RECT  10657.5 62597.5 10722.5 62462.5 ;
      RECT  10657.5 63572.5 10722.5 63437.5 ;
      RECT  10492.5 63297.5 10357.5 63232.5 ;
      RECT  10235.0 63082.5 10100.0 63017.5 ;
      RECT  10297.5 62687.5 10362.5 62552.5 ;
      RECT  10487.5 63527.5 10552.5 63392.5 ;
      RECT  10587.5 63082.5 10452.5 63017.5 ;
      RECT  10100.0 63082.5 10235.0 63017.5 ;
      RECT  10357.5 63297.5 10492.5 63232.5 ;
      RECT  10452.5 63082.5 10587.5 63017.5 ;
      RECT  10040.0 62377.5 10960.0 62312.5 ;
      RECT  10040.0 63722.5 10960.0 63657.5 ;
      RECT  11387.5 62530.0 11452.5 62345.0 ;
      RECT  11387.5 63690.0 11452.5 63505.0 ;
      RECT  11027.5 63572.5 11092.5 63722.5 ;
      RECT  11027.5 62687.5 11092.5 62312.5 ;
      RECT  11217.5 63572.5 11282.5 62687.5 ;
      RECT  11027.5 62687.5 11092.5 62552.5 ;
      RECT  11217.5 62687.5 11282.5 62552.5 ;
      RECT  11217.5 62687.5 11282.5 62552.5 ;
      RECT  11027.5 62687.5 11092.5 62552.5 ;
      RECT  11027.5 63572.5 11092.5 63437.5 ;
      RECT  11217.5 63572.5 11282.5 63437.5 ;
      RECT  11217.5 63572.5 11282.5 63437.5 ;
      RECT  11027.5 63572.5 11092.5 63437.5 ;
      RECT  11387.5 62597.5 11452.5 62462.5 ;
      RECT  11387.5 63572.5 11452.5 63437.5 ;
      RECT  11085.0 63130.0 11150.0 62995.0 ;
      RECT  11085.0 63130.0 11150.0 62995.0 ;
      RECT  11250.0 63095.0 11315.0 63030.0 ;
      RECT  10960.0 62377.5 11520.0 62312.5 ;
      RECT  10960.0 63722.5 11520.0 63657.5 ;
      RECT  9222.5 62995.0 9287.5 63130.0 ;
      RECT  9362.5 63267.5 9427.5 63402.5 ;
      RECT  10357.5 63232.5 10222.5 63297.5 ;
      RECT  9907.5 64850.0 9972.5 65035.0 ;
      RECT  9907.5 63690.0 9972.5 63875.0 ;
      RECT  9547.5 63807.5 9612.5 63657.5 ;
      RECT  9547.5 64692.5 9612.5 65067.5 ;
      RECT  9737.5 63807.5 9802.5 64692.5 ;
      RECT  9547.5 64692.5 9612.5 64827.5 ;
      RECT  9737.5 64692.5 9802.5 64827.5 ;
      RECT  9737.5 64692.5 9802.5 64827.5 ;
      RECT  9547.5 64692.5 9612.5 64827.5 ;
      RECT  9547.5 63807.5 9612.5 63942.5 ;
      RECT  9737.5 63807.5 9802.5 63942.5 ;
      RECT  9737.5 63807.5 9802.5 63942.5 ;
      RECT  9547.5 63807.5 9612.5 63942.5 ;
      RECT  9907.5 64782.5 9972.5 64917.5 ;
      RECT  9907.5 63807.5 9972.5 63942.5 ;
      RECT  9605.0 64250.0 9670.0 64385.0 ;
      RECT  9605.0 64250.0 9670.0 64385.0 ;
      RECT  9770.0 64285.0 9835.0 64350.0 ;
      RECT  9480.0 65002.5 10040.0 65067.5 ;
      RECT  9480.0 63657.5 10040.0 63722.5 ;
      RECT  10107.5 63852.5 10172.5 63657.5 ;
      RECT  10107.5 64692.5 10172.5 65067.5 ;
      RECT  10487.5 64692.5 10552.5 65067.5 ;
      RECT  10657.5 64850.0 10722.5 65035.0 ;
      RECT  10657.5 63690.0 10722.5 63875.0 ;
      RECT  10107.5 64692.5 10172.5 64827.5 ;
      RECT  10297.5 64692.5 10362.5 64827.5 ;
      RECT  10297.5 64692.5 10362.5 64827.5 ;
      RECT  10107.5 64692.5 10172.5 64827.5 ;
      RECT  10297.5 64692.5 10362.5 64827.5 ;
      RECT  10487.5 64692.5 10552.5 64827.5 ;
      RECT  10487.5 64692.5 10552.5 64827.5 ;
      RECT  10297.5 64692.5 10362.5 64827.5 ;
      RECT  10107.5 63852.5 10172.5 63987.5 ;
      RECT  10297.5 63852.5 10362.5 63987.5 ;
      RECT  10297.5 63852.5 10362.5 63987.5 ;
      RECT  10107.5 63852.5 10172.5 63987.5 ;
      RECT  10297.5 63852.5 10362.5 63987.5 ;
      RECT  10487.5 63852.5 10552.5 63987.5 ;
      RECT  10487.5 63852.5 10552.5 63987.5 ;
      RECT  10297.5 63852.5 10362.5 63987.5 ;
      RECT  10657.5 64782.5 10722.5 64917.5 ;
      RECT  10657.5 63807.5 10722.5 63942.5 ;
      RECT  10492.5 64082.5 10357.5 64147.5 ;
      RECT  10235.0 64297.5 10100.0 64362.5 ;
      RECT  10297.5 64692.5 10362.5 64827.5 ;
      RECT  10487.5 63852.5 10552.5 63987.5 ;
      RECT  10587.5 64297.5 10452.5 64362.5 ;
      RECT  10100.0 64297.5 10235.0 64362.5 ;
      RECT  10357.5 64082.5 10492.5 64147.5 ;
      RECT  10452.5 64297.5 10587.5 64362.5 ;
      RECT  10040.0 65002.5 10960.0 65067.5 ;
      RECT  10040.0 63657.5 10960.0 63722.5 ;
      RECT  11387.5 64850.0 11452.5 65035.0 ;
      RECT  11387.5 63690.0 11452.5 63875.0 ;
      RECT  11027.5 63807.5 11092.5 63657.5 ;
      RECT  11027.5 64692.5 11092.5 65067.5 ;
      RECT  11217.5 63807.5 11282.5 64692.5 ;
      RECT  11027.5 64692.5 11092.5 64827.5 ;
      RECT  11217.5 64692.5 11282.5 64827.5 ;
      RECT  11217.5 64692.5 11282.5 64827.5 ;
      RECT  11027.5 64692.5 11092.5 64827.5 ;
      RECT  11027.5 63807.5 11092.5 63942.5 ;
      RECT  11217.5 63807.5 11282.5 63942.5 ;
      RECT  11217.5 63807.5 11282.5 63942.5 ;
      RECT  11027.5 63807.5 11092.5 63942.5 ;
      RECT  11387.5 64782.5 11452.5 64917.5 ;
      RECT  11387.5 63807.5 11452.5 63942.5 ;
      RECT  11085.0 64250.0 11150.0 64385.0 ;
      RECT  11085.0 64250.0 11150.0 64385.0 ;
      RECT  11250.0 64285.0 11315.0 64350.0 ;
      RECT  10960.0 65002.5 11520.0 65067.5 ;
      RECT  10960.0 63657.5 11520.0 63722.5 ;
      RECT  9222.5 64250.0 9287.5 64385.0 ;
      RECT  9362.5 63977.5 9427.5 64112.5 ;
      RECT  10357.5 64082.5 10222.5 64147.5 ;
      RECT  9907.5 65220.0 9972.5 65035.0 ;
      RECT  9907.5 66380.0 9972.5 66195.0 ;
      RECT  9547.5 66262.5 9612.5 66412.5 ;
      RECT  9547.5 65377.5 9612.5 65002.5 ;
      RECT  9737.5 66262.5 9802.5 65377.5 ;
      RECT  9547.5 65377.5 9612.5 65242.5 ;
      RECT  9737.5 65377.5 9802.5 65242.5 ;
      RECT  9737.5 65377.5 9802.5 65242.5 ;
      RECT  9547.5 65377.5 9612.5 65242.5 ;
      RECT  9547.5 66262.5 9612.5 66127.5 ;
      RECT  9737.5 66262.5 9802.5 66127.5 ;
      RECT  9737.5 66262.5 9802.5 66127.5 ;
      RECT  9547.5 66262.5 9612.5 66127.5 ;
      RECT  9907.5 65287.5 9972.5 65152.5 ;
      RECT  9907.5 66262.5 9972.5 66127.5 ;
      RECT  9605.0 65820.0 9670.0 65685.0 ;
      RECT  9605.0 65820.0 9670.0 65685.0 ;
      RECT  9770.0 65785.0 9835.0 65720.0 ;
      RECT  9480.0 65067.5 10040.0 65002.5 ;
      RECT  9480.0 66412.5 10040.0 66347.5 ;
      RECT  10107.5 66217.5 10172.5 66412.5 ;
      RECT  10107.5 65377.5 10172.5 65002.5 ;
      RECT  10487.5 65377.5 10552.5 65002.5 ;
      RECT  10657.5 65220.0 10722.5 65035.0 ;
      RECT  10657.5 66380.0 10722.5 66195.0 ;
      RECT  10107.5 65377.5 10172.5 65242.5 ;
      RECT  10297.5 65377.5 10362.5 65242.5 ;
      RECT  10297.5 65377.5 10362.5 65242.5 ;
      RECT  10107.5 65377.5 10172.5 65242.5 ;
      RECT  10297.5 65377.5 10362.5 65242.5 ;
      RECT  10487.5 65377.5 10552.5 65242.5 ;
      RECT  10487.5 65377.5 10552.5 65242.5 ;
      RECT  10297.5 65377.5 10362.5 65242.5 ;
      RECT  10107.5 66217.5 10172.5 66082.5 ;
      RECT  10297.5 66217.5 10362.5 66082.5 ;
      RECT  10297.5 66217.5 10362.5 66082.5 ;
      RECT  10107.5 66217.5 10172.5 66082.5 ;
      RECT  10297.5 66217.5 10362.5 66082.5 ;
      RECT  10487.5 66217.5 10552.5 66082.5 ;
      RECT  10487.5 66217.5 10552.5 66082.5 ;
      RECT  10297.5 66217.5 10362.5 66082.5 ;
      RECT  10657.5 65287.5 10722.5 65152.5 ;
      RECT  10657.5 66262.5 10722.5 66127.5 ;
      RECT  10492.5 65987.5 10357.5 65922.5 ;
      RECT  10235.0 65772.5 10100.0 65707.5 ;
      RECT  10297.5 65377.5 10362.5 65242.5 ;
      RECT  10487.5 66217.5 10552.5 66082.5 ;
      RECT  10587.5 65772.5 10452.5 65707.5 ;
      RECT  10100.0 65772.5 10235.0 65707.5 ;
      RECT  10357.5 65987.5 10492.5 65922.5 ;
      RECT  10452.5 65772.5 10587.5 65707.5 ;
      RECT  10040.0 65067.5 10960.0 65002.5 ;
      RECT  10040.0 66412.5 10960.0 66347.5 ;
      RECT  11387.5 65220.0 11452.5 65035.0 ;
      RECT  11387.5 66380.0 11452.5 66195.0 ;
      RECT  11027.5 66262.5 11092.5 66412.5 ;
      RECT  11027.5 65377.5 11092.5 65002.5 ;
      RECT  11217.5 66262.5 11282.5 65377.5 ;
      RECT  11027.5 65377.5 11092.5 65242.5 ;
      RECT  11217.5 65377.5 11282.5 65242.5 ;
      RECT  11217.5 65377.5 11282.5 65242.5 ;
      RECT  11027.5 65377.5 11092.5 65242.5 ;
      RECT  11027.5 66262.5 11092.5 66127.5 ;
      RECT  11217.5 66262.5 11282.5 66127.5 ;
      RECT  11217.5 66262.5 11282.5 66127.5 ;
      RECT  11027.5 66262.5 11092.5 66127.5 ;
      RECT  11387.5 65287.5 11452.5 65152.5 ;
      RECT  11387.5 66262.5 11452.5 66127.5 ;
      RECT  11085.0 65820.0 11150.0 65685.0 ;
      RECT  11085.0 65820.0 11150.0 65685.0 ;
      RECT  11250.0 65785.0 11315.0 65720.0 ;
      RECT  10960.0 65067.5 11520.0 65002.5 ;
      RECT  10960.0 66412.5 11520.0 66347.5 ;
      RECT  9222.5 65685.0 9287.5 65820.0 ;
      RECT  9362.5 65957.5 9427.5 66092.5 ;
      RECT  10357.5 65922.5 10222.5 65987.5 ;
      RECT  9907.5 67540.0 9972.5 67725.0 ;
      RECT  9907.5 66380.0 9972.5 66565.0 ;
      RECT  9547.5 66497.5 9612.5 66347.5 ;
      RECT  9547.5 67382.5 9612.5 67757.5 ;
      RECT  9737.5 66497.5 9802.5 67382.5 ;
      RECT  9547.5 67382.5 9612.5 67517.5 ;
      RECT  9737.5 67382.5 9802.5 67517.5 ;
      RECT  9737.5 67382.5 9802.5 67517.5 ;
      RECT  9547.5 67382.5 9612.5 67517.5 ;
      RECT  9547.5 66497.5 9612.5 66632.5 ;
      RECT  9737.5 66497.5 9802.5 66632.5 ;
      RECT  9737.5 66497.5 9802.5 66632.5 ;
      RECT  9547.5 66497.5 9612.5 66632.5 ;
      RECT  9907.5 67472.5 9972.5 67607.5 ;
      RECT  9907.5 66497.5 9972.5 66632.5 ;
      RECT  9605.0 66940.0 9670.0 67075.0 ;
      RECT  9605.0 66940.0 9670.0 67075.0 ;
      RECT  9770.0 66975.0 9835.0 67040.0 ;
      RECT  9480.0 67692.5 10040.0 67757.5 ;
      RECT  9480.0 66347.5 10040.0 66412.5 ;
      RECT  10107.5 66542.5 10172.5 66347.5 ;
      RECT  10107.5 67382.5 10172.5 67757.5 ;
      RECT  10487.5 67382.5 10552.5 67757.5 ;
      RECT  10657.5 67540.0 10722.5 67725.0 ;
      RECT  10657.5 66380.0 10722.5 66565.0 ;
      RECT  10107.5 67382.5 10172.5 67517.5 ;
      RECT  10297.5 67382.5 10362.5 67517.5 ;
      RECT  10297.5 67382.5 10362.5 67517.5 ;
      RECT  10107.5 67382.5 10172.5 67517.5 ;
      RECT  10297.5 67382.5 10362.5 67517.5 ;
      RECT  10487.5 67382.5 10552.5 67517.5 ;
      RECT  10487.5 67382.5 10552.5 67517.5 ;
      RECT  10297.5 67382.5 10362.5 67517.5 ;
      RECT  10107.5 66542.5 10172.5 66677.5 ;
      RECT  10297.5 66542.5 10362.5 66677.5 ;
      RECT  10297.5 66542.5 10362.5 66677.5 ;
      RECT  10107.5 66542.5 10172.5 66677.5 ;
      RECT  10297.5 66542.5 10362.5 66677.5 ;
      RECT  10487.5 66542.5 10552.5 66677.5 ;
      RECT  10487.5 66542.5 10552.5 66677.5 ;
      RECT  10297.5 66542.5 10362.5 66677.5 ;
      RECT  10657.5 67472.5 10722.5 67607.5 ;
      RECT  10657.5 66497.5 10722.5 66632.5 ;
      RECT  10492.5 66772.5 10357.5 66837.5 ;
      RECT  10235.0 66987.5 10100.0 67052.5 ;
      RECT  10297.5 67382.5 10362.5 67517.5 ;
      RECT  10487.5 66542.5 10552.5 66677.5 ;
      RECT  10587.5 66987.5 10452.5 67052.5 ;
      RECT  10100.0 66987.5 10235.0 67052.5 ;
      RECT  10357.5 66772.5 10492.5 66837.5 ;
      RECT  10452.5 66987.5 10587.5 67052.5 ;
      RECT  10040.0 67692.5 10960.0 67757.5 ;
      RECT  10040.0 66347.5 10960.0 66412.5 ;
      RECT  11387.5 67540.0 11452.5 67725.0 ;
      RECT  11387.5 66380.0 11452.5 66565.0 ;
      RECT  11027.5 66497.5 11092.5 66347.5 ;
      RECT  11027.5 67382.5 11092.5 67757.5 ;
      RECT  11217.5 66497.5 11282.5 67382.5 ;
      RECT  11027.5 67382.5 11092.5 67517.5 ;
      RECT  11217.5 67382.5 11282.5 67517.5 ;
      RECT  11217.5 67382.5 11282.5 67517.5 ;
      RECT  11027.5 67382.5 11092.5 67517.5 ;
      RECT  11027.5 66497.5 11092.5 66632.5 ;
      RECT  11217.5 66497.5 11282.5 66632.5 ;
      RECT  11217.5 66497.5 11282.5 66632.5 ;
      RECT  11027.5 66497.5 11092.5 66632.5 ;
      RECT  11387.5 67472.5 11452.5 67607.5 ;
      RECT  11387.5 66497.5 11452.5 66632.5 ;
      RECT  11085.0 66940.0 11150.0 67075.0 ;
      RECT  11085.0 66940.0 11150.0 67075.0 ;
      RECT  11250.0 66975.0 11315.0 67040.0 ;
      RECT  10960.0 67692.5 11520.0 67757.5 ;
      RECT  10960.0 66347.5 11520.0 66412.5 ;
      RECT  9222.5 66940.0 9287.5 67075.0 ;
      RECT  9362.5 66667.5 9427.5 66802.5 ;
      RECT  10357.5 66772.5 10222.5 66837.5 ;
      RECT  9907.5 67910.0 9972.5 67725.0 ;
      RECT  9907.5 69070.0 9972.5 68885.0 ;
      RECT  9547.5 68952.5 9612.5 69102.5 ;
      RECT  9547.5 68067.5 9612.5 67692.5 ;
      RECT  9737.5 68952.5 9802.5 68067.5 ;
      RECT  9547.5 68067.5 9612.5 67932.5 ;
      RECT  9737.5 68067.5 9802.5 67932.5 ;
      RECT  9737.5 68067.5 9802.5 67932.5 ;
      RECT  9547.5 68067.5 9612.5 67932.5 ;
      RECT  9547.5 68952.5 9612.5 68817.5 ;
      RECT  9737.5 68952.5 9802.5 68817.5 ;
      RECT  9737.5 68952.5 9802.5 68817.5 ;
      RECT  9547.5 68952.5 9612.5 68817.5 ;
      RECT  9907.5 67977.5 9972.5 67842.5 ;
      RECT  9907.5 68952.5 9972.5 68817.5 ;
      RECT  9605.0 68510.0 9670.0 68375.0 ;
      RECT  9605.0 68510.0 9670.0 68375.0 ;
      RECT  9770.0 68475.0 9835.0 68410.0 ;
      RECT  9480.0 67757.5 10040.0 67692.5 ;
      RECT  9480.0 69102.5 10040.0 69037.5 ;
      RECT  10107.5 68907.5 10172.5 69102.5 ;
      RECT  10107.5 68067.5 10172.5 67692.5 ;
      RECT  10487.5 68067.5 10552.5 67692.5 ;
      RECT  10657.5 67910.0 10722.5 67725.0 ;
      RECT  10657.5 69070.0 10722.5 68885.0 ;
      RECT  10107.5 68067.5 10172.5 67932.5 ;
      RECT  10297.5 68067.5 10362.5 67932.5 ;
      RECT  10297.5 68067.5 10362.5 67932.5 ;
      RECT  10107.5 68067.5 10172.5 67932.5 ;
      RECT  10297.5 68067.5 10362.5 67932.5 ;
      RECT  10487.5 68067.5 10552.5 67932.5 ;
      RECT  10487.5 68067.5 10552.5 67932.5 ;
      RECT  10297.5 68067.5 10362.5 67932.5 ;
      RECT  10107.5 68907.5 10172.5 68772.5 ;
      RECT  10297.5 68907.5 10362.5 68772.5 ;
      RECT  10297.5 68907.5 10362.5 68772.5 ;
      RECT  10107.5 68907.5 10172.5 68772.5 ;
      RECT  10297.5 68907.5 10362.5 68772.5 ;
      RECT  10487.5 68907.5 10552.5 68772.5 ;
      RECT  10487.5 68907.5 10552.5 68772.5 ;
      RECT  10297.5 68907.5 10362.5 68772.5 ;
      RECT  10657.5 67977.5 10722.5 67842.5 ;
      RECT  10657.5 68952.5 10722.5 68817.5 ;
      RECT  10492.5 68677.5 10357.5 68612.5 ;
      RECT  10235.0 68462.5 10100.0 68397.5 ;
      RECT  10297.5 68067.5 10362.5 67932.5 ;
      RECT  10487.5 68907.5 10552.5 68772.5 ;
      RECT  10587.5 68462.5 10452.5 68397.5 ;
      RECT  10100.0 68462.5 10235.0 68397.5 ;
      RECT  10357.5 68677.5 10492.5 68612.5 ;
      RECT  10452.5 68462.5 10587.5 68397.5 ;
      RECT  10040.0 67757.5 10960.0 67692.5 ;
      RECT  10040.0 69102.5 10960.0 69037.5 ;
      RECT  11387.5 67910.0 11452.5 67725.0 ;
      RECT  11387.5 69070.0 11452.5 68885.0 ;
      RECT  11027.5 68952.5 11092.5 69102.5 ;
      RECT  11027.5 68067.5 11092.5 67692.5 ;
      RECT  11217.5 68952.5 11282.5 68067.5 ;
      RECT  11027.5 68067.5 11092.5 67932.5 ;
      RECT  11217.5 68067.5 11282.5 67932.5 ;
      RECT  11217.5 68067.5 11282.5 67932.5 ;
      RECT  11027.5 68067.5 11092.5 67932.5 ;
      RECT  11027.5 68952.5 11092.5 68817.5 ;
      RECT  11217.5 68952.5 11282.5 68817.5 ;
      RECT  11217.5 68952.5 11282.5 68817.5 ;
      RECT  11027.5 68952.5 11092.5 68817.5 ;
      RECT  11387.5 67977.5 11452.5 67842.5 ;
      RECT  11387.5 68952.5 11452.5 68817.5 ;
      RECT  11085.0 68510.0 11150.0 68375.0 ;
      RECT  11085.0 68510.0 11150.0 68375.0 ;
      RECT  11250.0 68475.0 11315.0 68410.0 ;
      RECT  10960.0 67757.5 11520.0 67692.5 ;
      RECT  10960.0 69102.5 11520.0 69037.5 ;
      RECT  9222.5 68375.0 9287.5 68510.0 ;
      RECT  9362.5 68647.5 9427.5 68782.5 ;
      RECT  10357.5 68612.5 10222.5 68677.5 ;
      RECT  9907.5 70230.0 9972.5 70415.0 ;
      RECT  9907.5 69070.0 9972.5 69255.0 ;
      RECT  9547.5 69187.5 9612.5 69037.5 ;
      RECT  9547.5 70072.5 9612.5 70447.5 ;
      RECT  9737.5 69187.5 9802.5 70072.5 ;
      RECT  9547.5 70072.5 9612.5 70207.5 ;
      RECT  9737.5 70072.5 9802.5 70207.5 ;
      RECT  9737.5 70072.5 9802.5 70207.5 ;
      RECT  9547.5 70072.5 9612.5 70207.5 ;
      RECT  9547.5 69187.5 9612.5 69322.5 ;
      RECT  9737.5 69187.5 9802.5 69322.5 ;
      RECT  9737.5 69187.5 9802.5 69322.5 ;
      RECT  9547.5 69187.5 9612.5 69322.5 ;
      RECT  9907.5 70162.5 9972.5 70297.5 ;
      RECT  9907.5 69187.5 9972.5 69322.5 ;
      RECT  9605.0 69630.0 9670.0 69765.0 ;
      RECT  9605.0 69630.0 9670.0 69765.0 ;
      RECT  9770.0 69665.0 9835.0 69730.0 ;
      RECT  9480.0 70382.5 10040.0 70447.5 ;
      RECT  9480.0 69037.5 10040.0 69102.5 ;
      RECT  10107.5 69232.5 10172.5 69037.5 ;
      RECT  10107.5 70072.5 10172.5 70447.5 ;
      RECT  10487.5 70072.5 10552.5 70447.5 ;
      RECT  10657.5 70230.0 10722.5 70415.0 ;
      RECT  10657.5 69070.0 10722.5 69255.0 ;
      RECT  10107.5 70072.5 10172.5 70207.5 ;
      RECT  10297.5 70072.5 10362.5 70207.5 ;
      RECT  10297.5 70072.5 10362.5 70207.5 ;
      RECT  10107.5 70072.5 10172.5 70207.5 ;
      RECT  10297.5 70072.5 10362.5 70207.5 ;
      RECT  10487.5 70072.5 10552.5 70207.5 ;
      RECT  10487.5 70072.5 10552.5 70207.5 ;
      RECT  10297.5 70072.5 10362.5 70207.5 ;
      RECT  10107.5 69232.5 10172.5 69367.5 ;
      RECT  10297.5 69232.5 10362.5 69367.5 ;
      RECT  10297.5 69232.5 10362.5 69367.5 ;
      RECT  10107.5 69232.5 10172.5 69367.5 ;
      RECT  10297.5 69232.5 10362.5 69367.5 ;
      RECT  10487.5 69232.5 10552.5 69367.5 ;
      RECT  10487.5 69232.5 10552.5 69367.5 ;
      RECT  10297.5 69232.5 10362.5 69367.5 ;
      RECT  10657.5 70162.5 10722.5 70297.5 ;
      RECT  10657.5 69187.5 10722.5 69322.5 ;
      RECT  10492.5 69462.5 10357.5 69527.5 ;
      RECT  10235.0 69677.5 10100.0 69742.5 ;
      RECT  10297.5 70072.5 10362.5 70207.5 ;
      RECT  10487.5 69232.5 10552.5 69367.5 ;
      RECT  10587.5 69677.5 10452.5 69742.5 ;
      RECT  10100.0 69677.5 10235.0 69742.5 ;
      RECT  10357.5 69462.5 10492.5 69527.5 ;
      RECT  10452.5 69677.5 10587.5 69742.5 ;
      RECT  10040.0 70382.5 10960.0 70447.5 ;
      RECT  10040.0 69037.5 10960.0 69102.5 ;
      RECT  11387.5 70230.0 11452.5 70415.0 ;
      RECT  11387.5 69070.0 11452.5 69255.0 ;
      RECT  11027.5 69187.5 11092.5 69037.5 ;
      RECT  11027.5 70072.5 11092.5 70447.5 ;
      RECT  11217.5 69187.5 11282.5 70072.5 ;
      RECT  11027.5 70072.5 11092.5 70207.5 ;
      RECT  11217.5 70072.5 11282.5 70207.5 ;
      RECT  11217.5 70072.5 11282.5 70207.5 ;
      RECT  11027.5 70072.5 11092.5 70207.5 ;
      RECT  11027.5 69187.5 11092.5 69322.5 ;
      RECT  11217.5 69187.5 11282.5 69322.5 ;
      RECT  11217.5 69187.5 11282.5 69322.5 ;
      RECT  11027.5 69187.5 11092.5 69322.5 ;
      RECT  11387.5 70162.5 11452.5 70297.5 ;
      RECT  11387.5 69187.5 11452.5 69322.5 ;
      RECT  11085.0 69630.0 11150.0 69765.0 ;
      RECT  11085.0 69630.0 11150.0 69765.0 ;
      RECT  11250.0 69665.0 11315.0 69730.0 ;
      RECT  10960.0 70382.5 11520.0 70447.5 ;
      RECT  10960.0 69037.5 11520.0 69102.5 ;
      RECT  9222.5 69630.0 9287.5 69765.0 ;
      RECT  9362.5 69357.5 9427.5 69492.5 ;
      RECT  10357.5 69462.5 10222.5 69527.5 ;
      RECT  9907.5 70600.0 9972.5 70415.0 ;
      RECT  9907.5 71760.0 9972.5 71575.0 ;
      RECT  9547.5 71642.5 9612.5 71792.5 ;
      RECT  9547.5 70757.5 9612.5 70382.5 ;
      RECT  9737.5 71642.5 9802.5 70757.5 ;
      RECT  9547.5 70757.5 9612.5 70622.5 ;
      RECT  9737.5 70757.5 9802.5 70622.5 ;
      RECT  9737.5 70757.5 9802.5 70622.5 ;
      RECT  9547.5 70757.5 9612.5 70622.5 ;
      RECT  9547.5 71642.5 9612.5 71507.5 ;
      RECT  9737.5 71642.5 9802.5 71507.5 ;
      RECT  9737.5 71642.5 9802.5 71507.5 ;
      RECT  9547.5 71642.5 9612.5 71507.5 ;
      RECT  9907.5 70667.5 9972.5 70532.5 ;
      RECT  9907.5 71642.5 9972.5 71507.5 ;
      RECT  9605.0 71200.0 9670.0 71065.0 ;
      RECT  9605.0 71200.0 9670.0 71065.0 ;
      RECT  9770.0 71165.0 9835.0 71100.0 ;
      RECT  9480.0 70447.5 10040.0 70382.5 ;
      RECT  9480.0 71792.5 10040.0 71727.5 ;
      RECT  10107.5 71597.5 10172.5 71792.5 ;
      RECT  10107.5 70757.5 10172.5 70382.5 ;
      RECT  10487.5 70757.5 10552.5 70382.5 ;
      RECT  10657.5 70600.0 10722.5 70415.0 ;
      RECT  10657.5 71760.0 10722.5 71575.0 ;
      RECT  10107.5 70757.5 10172.5 70622.5 ;
      RECT  10297.5 70757.5 10362.5 70622.5 ;
      RECT  10297.5 70757.5 10362.5 70622.5 ;
      RECT  10107.5 70757.5 10172.5 70622.5 ;
      RECT  10297.5 70757.5 10362.5 70622.5 ;
      RECT  10487.5 70757.5 10552.5 70622.5 ;
      RECT  10487.5 70757.5 10552.5 70622.5 ;
      RECT  10297.5 70757.5 10362.5 70622.5 ;
      RECT  10107.5 71597.5 10172.5 71462.5 ;
      RECT  10297.5 71597.5 10362.5 71462.5 ;
      RECT  10297.5 71597.5 10362.5 71462.5 ;
      RECT  10107.5 71597.5 10172.5 71462.5 ;
      RECT  10297.5 71597.5 10362.5 71462.5 ;
      RECT  10487.5 71597.5 10552.5 71462.5 ;
      RECT  10487.5 71597.5 10552.5 71462.5 ;
      RECT  10297.5 71597.5 10362.5 71462.5 ;
      RECT  10657.5 70667.5 10722.5 70532.5 ;
      RECT  10657.5 71642.5 10722.5 71507.5 ;
      RECT  10492.5 71367.5 10357.5 71302.5 ;
      RECT  10235.0 71152.5 10100.0 71087.5 ;
      RECT  10297.5 70757.5 10362.5 70622.5 ;
      RECT  10487.5 71597.5 10552.5 71462.5 ;
      RECT  10587.5 71152.5 10452.5 71087.5 ;
      RECT  10100.0 71152.5 10235.0 71087.5 ;
      RECT  10357.5 71367.5 10492.5 71302.5 ;
      RECT  10452.5 71152.5 10587.5 71087.5 ;
      RECT  10040.0 70447.5 10960.0 70382.5 ;
      RECT  10040.0 71792.5 10960.0 71727.5 ;
      RECT  11387.5 70600.0 11452.5 70415.0 ;
      RECT  11387.5 71760.0 11452.5 71575.0 ;
      RECT  11027.5 71642.5 11092.5 71792.5 ;
      RECT  11027.5 70757.5 11092.5 70382.5 ;
      RECT  11217.5 71642.5 11282.5 70757.5 ;
      RECT  11027.5 70757.5 11092.5 70622.5 ;
      RECT  11217.5 70757.5 11282.5 70622.5 ;
      RECT  11217.5 70757.5 11282.5 70622.5 ;
      RECT  11027.5 70757.5 11092.5 70622.5 ;
      RECT  11027.5 71642.5 11092.5 71507.5 ;
      RECT  11217.5 71642.5 11282.5 71507.5 ;
      RECT  11217.5 71642.5 11282.5 71507.5 ;
      RECT  11027.5 71642.5 11092.5 71507.5 ;
      RECT  11387.5 70667.5 11452.5 70532.5 ;
      RECT  11387.5 71642.5 11452.5 71507.5 ;
      RECT  11085.0 71200.0 11150.0 71065.0 ;
      RECT  11085.0 71200.0 11150.0 71065.0 ;
      RECT  11250.0 71165.0 11315.0 71100.0 ;
      RECT  10960.0 70447.5 11520.0 70382.5 ;
      RECT  10960.0 71792.5 11520.0 71727.5 ;
      RECT  9222.5 71065.0 9287.5 71200.0 ;
      RECT  9362.5 71337.5 9427.5 71472.5 ;
      RECT  10357.5 71302.5 10222.5 71367.5 ;
      RECT  9907.5 72920.0 9972.5 73105.0 ;
      RECT  9907.5 71760.0 9972.5 71945.0 ;
      RECT  9547.5 71877.5 9612.5 71727.5 ;
      RECT  9547.5 72762.5 9612.5 73137.5 ;
      RECT  9737.5 71877.5 9802.5 72762.5 ;
      RECT  9547.5 72762.5 9612.5 72897.5 ;
      RECT  9737.5 72762.5 9802.5 72897.5 ;
      RECT  9737.5 72762.5 9802.5 72897.5 ;
      RECT  9547.5 72762.5 9612.5 72897.5 ;
      RECT  9547.5 71877.5 9612.5 72012.5 ;
      RECT  9737.5 71877.5 9802.5 72012.5 ;
      RECT  9737.5 71877.5 9802.5 72012.5 ;
      RECT  9547.5 71877.5 9612.5 72012.5 ;
      RECT  9907.5 72852.5 9972.5 72987.5 ;
      RECT  9907.5 71877.5 9972.5 72012.5 ;
      RECT  9605.0 72320.0 9670.0 72455.0 ;
      RECT  9605.0 72320.0 9670.0 72455.0 ;
      RECT  9770.0 72355.0 9835.0 72420.0 ;
      RECT  9480.0 73072.5 10040.0 73137.5 ;
      RECT  9480.0 71727.5 10040.0 71792.5 ;
      RECT  10107.5 71922.5 10172.5 71727.5 ;
      RECT  10107.5 72762.5 10172.5 73137.5 ;
      RECT  10487.5 72762.5 10552.5 73137.5 ;
      RECT  10657.5 72920.0 10722.5 73105.0 ;
      RECT  10657.5 71760.0 10722.5 71945.0 ;
      RECT  10107.5 72762.5 10172.5 72897.5 ;
      RECT  10297.5 72762.5 10362.5 72897.5 ;
      RECT  10297.5 72762.5 10362.5 72897.5 ;
      RECT  10107.5 72762.5 10172.5 72897.5 ;
      RECT  10297.5 72762.5 10362.5 72897.5 ;
      RECT  10487.5 72762.5 10552.5 72897.5 ;
      RECT  10487.5 72762.5 10552.5 72897.5 ;
      RECT  10297.5 72762.5 10362.5 72897.5 ;
      RECT  10107.5 71922.5 10172.5 72057.5 ;
      RECT  10297.5 71922.5 10362.5 72057.5 ;
      RECT  10297.5 71922.5 10362.5 72057.5 ;
      RECT  10107.5 71922.5 10172.5 72057.5 ;
      RECT  10297.5 71922.5 10362.5 72057.5 ;
      RECT  10487.5 71922.5 10552.5 72057.5 ;
      RECT  10487.5 71922.5 10552.5 72057.5 ;
      RECT  10297.5 71922.5 10362.5 72057.5 ;
      RECT  10657.5 72852.5 10722.5 72987.5 ;
      RECT  10657.5 71877.5 10722.5 72012.5 ;
      RECT  10492.5 72152.5 10357.5 72217.5 ;
      RECT  10235.0 72367.5 10100.0 72432.5 ;
      RECT  10297.5 72762.5 10362.5 72897.5 ;
      RECT  10487.5 71922.5 10552.5 72057.5 ;
      RECT  10587.5 72367.5 10452.5 72432.5 ;
      RECT  10100.0 72367.5 10235.0 72432.5 ;
      RECT  10357.5 72152.5 10492.5 72217.5 ;
      RECT  10452.5 72367.5 10587.5 72432.5 ;
      RECT  10040.0 73072.5 10960.0 73137.5 ;
      RECT  10040.0 71727.5 10960.0 71792.5 ;
      RECT  11387.5 72920.0 11452.5 73105.0 ;
      RECT  11387.5 71760.0 11452.5 71945.0 ;
      RECT  11027.5 71877.5 11092.5 71727.5 ;
      RECT  11027.5 72762.5 11092.5 73137.5 ;
      RECT  11217.5 71877.5 11282.5 72762.5 ;
      RECT  11027.5 72762.5 11092.5 72897.5 ;
      RECT  11217.5 72762.5 11282.5 72897.5 ;
      RECT  11217.5 72762.5 11282.5 72897.5 ;
      RECT  11027.5 72762.5 11092.5 72897.5 ;
      RECT  11027.5 71877.5 11092.5 72012.5 ;
      RECT  11217.5 71877.5 11282.5 72012.5 ;
      RECT  11217.5 71877.5 11282.5 72012.5 ;
      RECT  11027.5 71877.5 11092.5 72012.5 ;
      RECT  11387.5 72852.5 11452.5 72987.5 ;
      RECT  11387.5 71877.5 11452.5 72012.5 ;
      RECT  11085.0 72320.0 11150.0 72455.0 ;
      RECT  11085.0 72320.0 11150.0 72455.0 ;
      RECT  11250.0 72355.0 11315.0 72420.0 ;
      RECT  10960.0 73072.5 11520.0 73137.5 ;
      RECT  10960.0 71727.5 11520.0 71792.5 ;
      RECT  9222.5 72320.0 9287.5 72455.0 ;
      RECT  9362.5 72047.5 9427.5 72182.5 ;
      RECT  10357.5 72152.5 10222.5 72217.5 ;
      RECT  9907.5 73290.0 9972.5 73105.0 ;
      RECT  9907.5 74450.0 9972.5 74265.0 ;
      RECT  9547.5 74332.5 9612.5 74482.5 ;
      RECT  9547.5 73447.5 9612.5 73072.5 ;
      RECT  9737.5 74332.5 9802.5 73447.5 ;
      RECT  9547.5 73447.5 9612.5 73312.5 ;
      RECT  9737.5 73447.5 9802.5 73312.5 ;
      RECT  9737.5 73447.5 9802.5 73312.5 ;
      RECT  9547.5 73447.5 9612.5 73312.5 ;
      RECT  9547.5 74332.5 9612.5 74197.5 ;
      RECT  9737.5 74332.5 9802.5 74197.5 ;
      RECT  9737.5 74332.5 9802.5 74197.5 ;
      RECT  9547.5 74332.5 9612.5 74197.5 ;
      RECT  9907.5 73357.5 9972.5 73222.5 ;
      RECT  9907.5 74332.5 9972.5 74197.5 ;
      RECT  9605.0 73890.0 9670.0 73755.0 ;
      RECT  9605.0 73890.0 9670.0 73755.0 ;
      RECT  9770.0 73855.0 9835.0 73790.0 ;
      RECT  9480.0 73137.5 10040.0 73072.5 ;
      RECT  9480.0 74482.5 10040.0 74417.5 ;
      RECT  10107.5 74287.5 10172.5 74482.5 ;
      RECT  10107.5 73447.5 10172.5 73072.5 ;
      RECT  10487.5 73447.5 10552.5 73072.5 ;
      RECT  10657.5 73290.0 10722.5 73105.0 ;
      RECT  10657.5 74450.0 10722.5 74265.0 ;
      RECT  10107.5 73447.5 10172.5 73312.5 ;
      RECT  10297.5 73447.5 10362.5 73312.5 ;
      RECT  10297.5 73447.5 10362.5 73312.5 ;
      RECT  10107.5 73447.5 10172.5 73312.5 ;
      RECT  10297.5 73447.5 10362.5 73312.5 ;
      RECT  10487.5 73447.5 10552.5 73312.5 ;
      RECT  10487.5 73447.5 10552.5 73312.5 ;
      RECT  10297.5 73447.5 10362.5 73312.5 ;
      RECT  10107.5 74287.5 10172.5 74152.5 ;
      RECT  10297.5 74287.5 10362.5 74152.5 ;
      RECT  10297.5 74287.5 10362.5 74152.5 ;
      RECT  10107.5 74287.5 10172.5 74152.5 ;
      RECT  10297.5 74287.5 10362.5 74152.5 ;
      RECT  10487.5 74287.5 10552.5 74152.5 ;
      RECT  10487.5 74287.5 10552.5 74152.5 ;
      RECT  10297.5 74287.5 10362.5 74152.5 ;
      RECT  10657.5 73357.5 10722.5 73222.5 ;
      RECT  10657.5 74332.5 10722.5 74197.5 ;
      RECT  10492.5 74057.5 10357.5 73992.5 ;
      RECT  10235.0 73842.5 10100.0 73777.5 ;
      RECT  10297.5 73447.5 10362.5 73312.5 ;
      RECT  10487.5 74287.5 10552.5 74152.5 ;
      RECT  10587.5 73842.5 10452.5 73777.5 ;
      RECT  10100.0 73842.5 10235.0 73777.5 ;
      RECT  10357.5 74057.5 10492.5 73992.5 ;
      RECT  10452.5 73842.5 10587.5 73777.5 ;
      RECT  10040.0 73137.5 10960.0 73072.5 ;
      RECT  10040.0 74482.5 10960.0 74417.5 ;
      RECT  11387.5 73290.0 11452.5 73105.0 ;
      RECT  11387.5 74450.0 11452.5 74265.0 ;
      RECT  11027.5 74332.5 11092.5 74482.5 ;
      RECT  11027.5 73447.5 11092.5 73072.5 ;
      RECT  11217.5 74332.5 11282.5 73447.5 ;
      RECT  11027.5 73447.5 11092.5 73312.5 ;
      RECT  11217.5 73447.5 11282.5 73312.5 ;
      RECT  11217.5 73447.5 11282.5 73312.5 ;
      RECT  11027.5 73447.5 11092.5 73312.5 ;
      RECT  11027.5 74332.5 11092.5 74197.5 ;
      RECT  11217.5 74332.5 11282.5 74197.5 ;
      RECT  11217.5 74332.5 11282.5 74197.5 ;
      RECT  11027.5 74332.5 11092.5 74197.5 ;
      RECT  11387.5 73357.5 11452.5 73222.5 ;
      RECT  11387.5 74332.5 11452.5 74197.5 ;
      RECT  11085.0 73890.0 11150.0 73755.0 ;
      RECT  11085.0 73890.0 11150.0 73755.0 ;
      RECT  11250.0 73855.0 11315.0 73790.0 ;
      RECT  10960.0 73137.5 11520.0 73072.5 ;
      RECT  10960.0 74482.5 11520.0 74417.5 ;
      RECT  9222.5 73755.0 9287.5 73890.0 ;
      RECT  9362.5 74027.5 9427.5 74162.5 ;
      RECT  10357.5 73992.5 10222.5 74057.5 ;
      RECT  9907.5 75610.0 9972.5 75795.0 ;
      RECT  9907.5 74450.0 9972.5 74635.0 ;
      RECT  9547.5 74567.5 9612.5 74417.5 ;
      RECT  9547.5 75452.5 9612.5 75827.5 ;
      RECT  9737.5 74567.5 9802.5 75452.5 ;
      RECT  9547.5 75452.5 9612.5 75587.5 ;
      RECT  9737.5 75452.5 9802.5 75587.5 ;
      RECT  9737.5 75452.5 9802.5 75587.5 ;
      RECT  9547.5 75452.5 9612.5 75587.5 ;
      RECT  9547.5 74567.5 9612.5 74702.5 ;
      RECT  9737.5 74567.5 9802.5 74702.5 ;
      RECT  9737.5 74567.5 9802.5 74702.5 ;
      RECT  9547.5 74567.5 9612.5 74702.5 ;
      RECT  9907.5 75542.5 9972.5 75677.5 ;
      RECT  9907.5 74567.5 9972.5 74702.5 ;
      RECT  9605.0 75010.0 9670.0 75145.0 ;
      RECT  9605.0 75010.0 9670.0 75145.0 ;
      RECT  9770.0 75045.0 9835.0 75110.0 ;
      RECT  9480.0 75762.5 10040.0 75827.5 ;
      RECT  9480.0 74417.5 10040.0 74482.5 ;
      RECT  10107.5 74612.5 10172.5 74417.5 ;
      RECT  10107.5 75452.5 10172.5 75827.5 ;
      RECT  10487.5 75452.5 10552.5 75827.5 ;
      RECT  10657.5 75610.0 10722.5 75795.0 ;
      RECT  10657.5 74450.0 10722.5 74635.0 ;
      RECT  10107.5 75452.5 10172.5 75587.5 ;
      RECT  10297.5 75452.5 10362.5 75587.5 ;
      RECT  10297.5 75452.5 10362.5 75587.5 ;
      RECT  10107.5 75452.5 10172.5 75587.5 ;
      RECT  10297.5 75452.5 10362.5 75587.5 ;
      RECT  10487.5 75452.5 10552.5 75587.5 ;
      RECT  10487.5 75452.5 10552.5 75587.5 ;
      RECT  10297.5 75452.5 10362.5 75587.5 ;
      RECT  10107.5 74612.5 10172.5 74747.5 ;
      RECT  10297.5 74612.5 10362.5 74747.5 ;
      RECT  10297.5 74612.5 10362.5 74747.5 ;
      RECT  10107.5 74612.5 10172.5 74747.5 ;
      RECT  10297.5 74612.5 10362.5 74747.5 ;
      RECT  10487.5 74612.5 10552.5 74747.5 ;
      RECT  10487.5 74612.5 10552.5 74747.5 ;
      RECT  10297.5 74612.5 10362.5 74747.5 ;
      RECT  10657.5 75542.5 10722.5 75677.5 ;
      RECT  10657.5 74567.5 10722.5 74702.5 ;
      RECT  10492.5 74842.5 10357.5 74907.5 ;
      RECT  10235.0 75057.5 10100.0 75122.5 ;
      RECT  10297.5 75452.5 10362.5 75587.5 ;
      RECT  10487.5 74612.5 10552.5 74747.5 ;
      RECT  10587.5 75057.5 10452.5 75122.5 ;
      RECT  10100.0 75057.5 10235.0 75122.5 ;
      RECT  10357.5 74842.5 10492.5 74907.5 ;
      RECT  10452.5 75057.5 10587.5 75122.5 ;
      RECT  10040.0 75762.5 10960.0 75827.5 ;
      RECT  10040.0 74417.5 10960.0 74482.5 ;
      RECT  11387.5 75610.0 11452.5 75795.0 ;
      RECT  11387.5 74450.0 11452.5 74635.0 ;
      RECT  11027.5 74567.5 11092.5 74417.5 ;
      RECT  11027.5 75452.5 11092.5 75827.5 ;
      RECT  11217.5 74567.5 11282.5 75452.5 ;
      RECT  11027.5 75452.5 11092.5 75587.5 ;
      RECT  11217.5 75452.5 11282.5 75587.5 ;
      RECT  11217.5 75452.5 11282.5 75587.5 ;
      RECT  11027.5 75452.5 11092.5 75587.5 ;
      RECT  11027.5 74567.5 11092.5 74702.5 ;
      RECT  11217.5 74567.5 11282.5 74702.5 ;
      RECT  11217.5 74567.5 11282.5 74702.5 ;
      RECT  11027.5 74567.5 11092.5 74702.5 ;
      RECT  11387.5 75542.5 11452.5 75677.5 ;
      RECT  11387.5 74567.5 11452.5 74702.5 ;
      RECT  11085.0 75010.0 11150.0 75145.0 ;
      RECT  11085.0 75010.0 11150.0 75145.0 ;
      RECT  11250.0 75045.0 11315.0 75110.0 ;
      RECT  10960.0 75762.5 11520.0 75827.5 ;
      RECT  10960.0 74417.5 11520.0 74482.5 ;
      RECT  9222.5 75010.0 9287.5 75145.0 ;
      RECT  9362.5 74737.5 9427.5 74872.5 ;
      RECT  10357.5 74842.5 10222.5 74907.5 ;
      RECT  9907.5 75980.0 9972.5 75795.0 ;
      RECT  9907.5 77140.0 9972.5 76955.0 ;
      RECT  9547.5 77022.5 9612.5 77172.5 ;
      RECT  9547.5 76137.5 9612.5 75762.5 ;
      RECT  9737.5 77022.5 9802.5 76137.5 ;
      RECT  9547.5 76137.5 9612.5 76002.5 ;
      RECT  9737.5 76137.5 9802.5 76002.5 ;
      RECT  9737.5 76137.5 9802.5 76002.5 ;
      RECT  9547.5 76137.5 9612.5 76002.5 ;
      RECT  9547.5 77022.5 9612.5 76887.5 ;
      RECT  9737.5 77022.5 9802.5 76887.5 ;
      RECT  9737.5 77022.5 9802.5 76887.5 ;
      RECT  9547.5 77022.5 9612.5 76887.5 ;
      RECT  9907.5 76047.5 9972.5 75912.5 ;
      RECT  9907.5 77022.5 9972.5 76887.5 ;
      RECT  9605.0 76580.0 9670.0 76445.0 ;
      RECT  9605.0 76580.0 9670.0 76445.0 ;
      RECT  9770.0 76545.0 9835.0 76480.0 ;
      RECT  9480.0 75827.5 10040.0 75762.5 ;
      RECT  9480.0 77172.5 10040.0 77107.5 ;
      RECT  10107.5 76977.5 10172.5 77172.5 ;
      RECT  10107.5 76137.5 10172.5 75762.5 ;
      RECT  10487.5 76137.5 10552.5 75762.5 ;
      RECT  10657.5 75980.0 10722.5 75795.0 ;
      RECT  10657.5 77140.0 10722.5 76955.0 ;
      RECT  10107.5 76137.5 10172.5 76002.5 ;
      RECT  10297.5 76137.5 10362.5 76002.5 ;
      RECT  10297.5 76137.5 10362.5 76002.5 ;
      RECT  10107.5 76137.5 10172.5 76002.5 ;
      RECT  10297.5 76137.5 10362.5 76002.5 ;
      RECT  10487.5 76137.5 10552.5 76002.5 ;
      RECT  10487.5 76137.5 10552.5 76002.5 ;
      RECT  10297.5 76137.5 10362.5 76002.5 ;
      RECT  10107.5 76977.5 10172.5 76842.5 ;
      RECT  10297.5 76977.5 10362.5 76842.5 ;
      RECT  10297.5 76977.5 10362.5 76842.5 ;
      RECT  10107.5 76977.5 10172.5 76842.5 ;
      RECT  10297.5 76977.5 10362.5 76842.5 ;
      RECT  10487.5 76977.5 10552.5 76842.5 ;
      RECT  10487.5 76977.5 10552.5 76842.5 ;
      RECT  10297.5 76977.5 10362.5 76842.5 ;
      RECT  10657.5 76047.5 10722.5 75912.5 ;
      RECT  10657.5 77022.5 10722.5 76887.5 ;
      RECT  10492.5 76747.5 10357.5 76682.5 ;
      RECT  10235.0 76532.5 10100.0 76467.5 ;
      RECT  10297.5 76137.5 10362.5 76002.5 ;
      RECT  10487.5 76977.5 10552.5 76842.5 ;
      RECT  10587.5 76532.5 10452.5 76467.5 ;
      RECT  10100.0 76532.5 10235.0 76467.5 ;
      RECT  10357.5 76747.5 10492.5 76682.5 ;
      RECT  10452.5 76532.5 10587.5 76467.5 ;
      RECT  10040.0 75827.5 10960.0 75762.5 ;
      RECT  10040.0 77172.5 10960.0 77107.5 ;
      RECT  11387.5 75980.0 11452.5 75795.0 ;
      RECT  11387.5 77140.0 11452.5 76955.0 ;
      RECT  11027.5 77022.5 11092.5 77172.5 ;
      RECT  11027.5 76137.5 11092.5 75762.5 ;
      RECT  11217.5 77022.5 11282.5 76137.5 ;
      RECT  11027.5 76137.5 11092.5 76002.5 ;
      RECT  11217.5 76137.5 11282.5 76002.5 ;
      RECT  11217.5 76137.5 11282.5 76002.5 ;
      RECT  11027.5 76137.5 11092.5 76002.5 ;
      RECT  11027.5 77022.5 11092.5 76887.5 ;
      RECT  11217.5 77022.5 11282.5 76887.5 ;
      RECT  11217.5 77022.5 11282.5 76887.5 ;
      RECT  11027.5 77022.5 11092.5 76887.5 ;
      RECT  11387.5 76047.5 11452.5 75912.5 ;
      RECT  11387.5 77022.5 11452.5 76887.5 ;
      RECT  11085.0 76580.0 11150.0 76445.0 ;
      RECT  11085.0 76580.0 11150.0 76445.0 ;
      RECT  11250.0 76545.0 11315.0 76480.0 ;
      RECT  10960.0 75827.5 11520.0 75762.5 ;
      RECT  10960.0 77172.5 11520.0 77107.5 ;
      RECT  9222.5 76445.0 9287.5 76580.0 ;
      RECT  9362.5 76717.5 9427.5 76852.5 ;
      RECT  10357.5 76682.5 10222.5 76747.5 ;
      RECT  9907.5 78300.0 9972.5 78485.0 ;
      RECT  9907.5 77140.0 9972.5 77325.0 ;
      RECT  9547.5 77257.5 9612.5 77107.5 ;
      RECT  9547.5 78142.5 9612.5 78517.5 ;
      RECT  9737.5 77257.5 9802.5 78142.5 ;
      RECT  9547.5 78142.5 9612.5 78277.5 ;
      RECT  9737.5 78142.5 9802.5 78277.5 ;
      RECT  9737.5 78142.5 9802.5 78277.5 ;
      RECT  9547.5 78142.5 9612.5 78277.5 ;
      RECT  9547.5 77257.5 9612.5 77392.5 ;
      RECT  9737.5 77257.5 9802.5 77392.5 ;
      RECT  9737.5 77257.5 9802.5 77392.5 ;
      RECT  9547.5 77257.5 9612.5 77392.5 ;
      RECT  9907.5 78232.5 9972.5 78367.5 ;
      RECT  9907.5 77257.5 9972.5 77392.5 ;
      RECT  9605.0 77700.0 9670.0 77835.0 ;
      RECT  9605.0 77700.0 9670.0 77835.0 ;
      RECT  9770.0 77735.0 9835.0 77800.0 ;
      RECT  9480.0 78452.5 10040.0 78517.5 ;
      RECT  9480.0 77107.5 10040.0 77172.5 ;
      RECT  10107.5 77302.5 10172.5 77107.5 ;
      RECT  10107.5 78142.5 10172.5 78517.5 ;
      RECT  10487.5 78142.5 10552.5 78517.5 ;
      RECT  10657.5 78300.0 10722.5 78485.0 ;
      RECT  10657.5 77140.0 10722.5 77325.0 ;
      RECT  10107.5 78142.5 10172.5 78277.5 ;
      RECT  10297.5 78142.5 10362.5 78277.5 ;
      RECT  10297.5 78142.5 10362.5 78277.5 ;
      RECT  10107.5 78142.5 10172.5 78277.5 ;
      RECT  10297.5 78142.5 10362.5 78277.5 ;
      RECT  10487.5 78142.5 10552.5 78277.5 ;
      RECT  10487.5 78142.5 10552.5 78277.5 ;
      RECT  10297.5 78142.5 10362.5 78277.5 ;
      RECT  10107.5 77302.5 10172.5 77437.5 ;
      RECT  10297.5 77302.5 10362.5 77437.5 ;
      RECT  10297.5 77302.5 10362.5 77437.5 ;
      RECT  10107.5 77302.5 10172.5 77437.5 ;
      RECT  10297.5 77302.5 10362.5 77437.5 ;
      RECT  10487.5 77302.5 10552.5 77437.5 ;
      RECT  10487.5 77302.5 10552.5 77437.5 ;
      RECT  10297.5 77302.5 10362.5 77437.5 ;
      RECT  10657.5 78232.5 10722.5 78367.5 ;
      RECT  10657.5 77257.5 10722.5 77392.5 ;
      RECT  10492.5 77532.5 10357.5 77597.5 ;
      RECT  10235.0 77747.5 10100.0 77812.5 ;
      RECT  10297.5 78142.5 10362.5 78277.5 ;
      RECT  10487.5 77302.5 10552.5 77437.5 ;
      RECT  10587.5 77747.5 10452.5 77812.5 ;
      RECT  10100.0 77747.5 10235.0 77812.5 ;
      RECT  10357.5 77532.5 10492.5 77597.5 ;
      RECT  10452.5 77747.5 10587.5 77812.5 ;
      RECT  10040.0 78452.5 10960.0 78517.5 ;
      RECT  10040.0 77107.5 10960.0 77172.5 ;
      RECT  11387.5 78300.0 11452.5 78485.0 ;
      RECT  11387.5 77140.0 11452.5 77325.0 ;
      RECT  11027.5 77257.5 11092.5 77107.5 ;
      RECT  11027.5 78142.5 11092.5 78517.5 ;
      RECT  11217.5 77257.5 11282.5 78142.5 ;
      RECT  11027.5 78142.5 11092.5 78277.5 ;
      RECT  11217.5 78142.5 11282.5 78277.5 ;
      RECT  11217.5 78142.5 11282.5 78277.5 ;
      RECT  11027.5 78142.5 11092.5 78277.5 ;
      RECT  11027.5 77257.5 11092.5 77392.5 ;
      RECT  11217.5 77257.5 11282.5 77392.5 ;
      RECT  11217.5 77257.5 11282.5 77392.5 ;
      RECT  11027.5 77257.5 11092.5 77392.5 ;
      RECT  11387.5 78232.5 11452.5 78367.5 ;
      RECT  11387.5 77257.5 11452.5 77392.5 ;
      RECT  11085.0 77700.0 11150.0 77835.0 ;
      RECT  11085.0 77700.0 11150.0 77835.0 ;
      RECT  11250.0 77735.0 11315.0 77800.0 ;
      RECT  10960.0 78452.5 11520.0 78517.5 ;
      RECT  10960.0 77107.5 11520.0 77172.5 ;
      RECT  9222.5 77700.0 9287.5 77835.0 ;
      RECT  9362.5 77427.5 9427.5 77562.5 ;
      RECT  10357.5 77532.5 10222.5 77597.5 ;
      RECT  9907.5 78670.0 9972.5 78485.0 ;
      RECT  9907.5 79830.0 9972.5 79645.0 ;
      RECT  9547.5 79712.5 9612.5 79862.5 ;
      RECT  9547.5 78827.5 9612.5 78452.5 ;
      RECT  9737.5 79712.5 9802.5 78827.5 ;
      RECT  9547.5 78827.5 9612.5 78692.5 ;
      RECT  9737.5 78827.5 9802.5 78692.5 ;
      RECT  9737.5 78827.5 9802.5 78692.5 ;
      RECT  9547.5 78827.5 9612.5 78692.5 ;
      RECT  9547.5 79712.5 9612.5 79577.5 ;
      RECT  9737.5 79712.5 9802.5 79577.5 ;
      RECT  9737.5 79712.5 9802.5 79577.5 ;
      RECT  9547.5 79712.5 9612.5 79577.5 ;
      RECT  9907.5 78737.5 9972.5 78602.5 ;
      RECT  9907.5 79712.5 9972.5 79577.5 ;
      RECT  9605.0 79270.0 9670.0 79135.0 ;
      RECT  9605.0 79270.0 9670.0 79135.0 ;
      RECT  9770.0 79235.0 9835.0 79170.0 ;
      RECT  9480.0 78517.5 10040.0 78452.5 ;
      RECT  9480.0 79862.5 10040.0 79797.5 ;
      RECT  10107.5 79667.5 10172.5 79862.5 ;
      RECT  10107.5 78827.5 10172.5 78452.5 ;
      RECT  10487.5 78827.5 10552.5 78452.5 ;
      RECT  10657.5 78670.0 10722.5 78485.0 ;
      RECT  10657.5 79830.0 10722.5 79645.0 ;
      RECT  10107.5 78827.5 10172.5 78692.5 ;
      RECT  10297.5 78827.5 10362.5 78692.5 ;
      RECT  10297.5 78827.5 10362.5 78692.5 ;
      RECT  10107.5 78827.5 10172.5 78692.5 ;
      RECT  10297.5 78827.5 10362.5 78692.5 ;
      RECT  10487.5 78827.5 10552.5 78692.5 ;
      RECT  10487.5 78827.5 10552.5 78692.5 ;
      RECT  10297.5 78827.5 10362.5 78692.5 ;
      RECT  10107.5 79667.5 10172.5 79532.5 ;
      RECT  10297.5 79667.5 10362.5 79532.5 ;
      RECT  10297.5 79667.5 10362.5 79532.5 ;
      RECT  10107.5 79667.5 10172.5 79532.5 ;
      RECT  10297.5 79667.5 10362.5 79532.5 ;
      RECT  10487.5 79667.5 10552.5 79532.5 ;
      RECT  10487.5 79667.5 10552.5 79532.5 ;
      RECT  10297.5 79667.5 10362.5 79532.5 ;
      RECT  10657.5 78737.5 10722.5 78602.5 ;
      RECT  10657.5 79712.5 10722.5 79577.5 ;
      RECT  10492.5 79437.5 10357.5 79372.5 ;
      RECT  10235.0 79222.5 10100.0 79157.5 ;
      RECT  10297.5 78827.5 10362.5 78692.5 ;
      RECT  10487.5 79667.5 10552.5 79532.5 ;
      RECT  10587.5 79222.5 10452.5 79157.5 ;
      RECT  10100.0 79222.5 10235.0 79157.5 ;
      RECT  10357.5 79437.5 10492.5 79372.5 ;
      RECT  10452.5 79222.5 10587.5 79157.5 ;
      RECT  10040.0 78517.5 10960.0 78452.5 ;
      RECT  10040.0 79862.5 10960.0 79797.5 ;
      RECT  11387.5 78670.0 11452.5 78485.0 ;
      RECT  11387.5 79830.0 11452.5 79645.0 ;
      RECT  11027.5 79712.5 11092.5 79862.5 ;
      RECT  11027.5 78827.5 11092.5 78452.5 ;
      RECT  11217.5 79712.5 11282.5 78827.5 ;
      RECT  11027.5 78827.5 11092.5 78692.5 ;
      RECT  11217.5 78827.5 11282.5 78692.5 ;
      RECT  11217.5 78827.5 11282.5 78692.5 ;
      RECT  11027.5 78827.5 11092.5 78692.5 ;
      RECT  11027.5 79712.5 11092.5 79577.5 ;
      RECT  11217.5 79712.5 11282.5 79577.5 ;
      RECT  11217.5 79712.5 11282.5 79577.5 ;
      RECT  11027.5 79712.5 11092.5 79577.5 ;
      RECT  11387.5 78737.5 11452.5 78602.5 ;
      RECT  11387.5 79712.5 11452.5 79577.5 ;
      RECT  11085.0 79270.0 11150.0 79135.0 ;
      RECT  11085.0 79270.0 11150.0 79135.0 ;
      RECT  11250.0 79235.0 11315.0 79170.0 ;
      RECT  10960.0 78517.5 11520.0 78452.5 ;
      RECT  10960.0 79862.5 11520.0 79797.5 ;
      RECT  9222.5 79135.0 9287.5 79270.0 ;
      RECT  9362.5 79407.5 9427.5 79542.5 ;
      RECT  10357.5 79372.5 10222.5 79437.5 ;
      RECT  9907.5 80990.0 9972.5 81175.0 ;
      RECT  9907.5 79830.0 9972.5 80015.0 ;
      RECT  9547.5 79947.5 9612.5 79797.5 ;
      RECT  9547.5 80832.5 9612.5 81207.5 ;
      RECT  9737.5 79947.5 9802.5 80832.5 ;
      RECT  9547.5 80832.5 9612.5 80967.5 ;
      RECT  9737.5 80832.5 9802.5 80967.5 ;
      RECT  9737.5 80832.5 9802.5 80967.5 ;
      RECT  9547.5 80832.5 9612.5 80967.5 ;
      RECT  9547.5 79947.5 9612.5 80082.5 ;
      RECT  9737.5 79947.5 9802.5 80082.5 ;
      RECT  9737.5 79947.5 9802.5 80082.5 ;
      RECT  9547.5 79947.5 9612.5 80082.5 ;
      RECT  9907.5 80922.5 9972.5 81057.5 ;
      RECT  9907.5 79947.5 9972.5 80082.5 ;
      RECT  9605.0 80390.0 9670.0 80525.0 ;
      RECT  9605.0 80390.0 9670.0 80525.0 ;
      RECT  9770.0 80425.0 9835.0 80490.0 ;
      RECT  9480.0 81142.5 10040.0 81207.5 ;
      RECT  9480.0 79797.5 10040.0 79862.5 ;
      RECT  10107.5 79992.5 10172.5 79797.5 ;
      RECT  10107.5 80832.5 10172.5 81207.5 ;
      RECT  10487.5 80832.5 10552.5 81207.5 ;
      RECT  10657.5 80990.0 10722.5 81175.0 ;
      RECT  10657.5 79830.0 10722.5 80015.0 ;
      RECT  10107.5 80832.5 10172.5 80967.5 ;
      RECT  10297.5 80832.5 10362.5 80967.5 ;
      RECT  10297.5 80832.5 10362.5 80967.5 ;
      RECT  10107.5 80832.5 10172.5 80967.5 ;
      RECT  10297.5 80832.5 10362.5 80967.5 ;
      RECT  10487.5 80832.5 10552.5 80967.5 ;
      RECT  10487.5 80832.5 10552.5 80967.5 ;
      RECT  10297.5 80832.5 10362.5 80967.5 ;
      RECT  10107.5 79992.5 10172.5 80127.5 ;
      RECT  10297.5 79992.5 10362.5 80127.5 ;
      RECT  10297.5 79992.5 10362.5 80127.5 ;
      RECT  10107.5 79992.5 10172.5 80127.5 ;
      RECT  10297.5 79992.5 10362.5 80127.5 ;
      RECT  10487.5 79992.5 10552.5 80127.5 ;
      RECT  10487.5 79992.5 10552.5 80127.5 ;
      RECT  10297.5 79992.5 10362.5 80127.5 ;
      RECT  10657.5 80922.5 10722.5 81057.5 ;
      RECT  10657.5 79947.5 10722.5 80082.5 ;
      RECT  10492.5 80222.5 10357.5 80287.5 ;
      RECT  10235.0 80437.5 10100.0 80502.5 ;
      RECT  10297.5 80832.5 10362.5 80967.5 ;
      RECT  10487.5 79992.5 10552.5 80127.5 ;
      RECT  10587.5 80437.5 10452.5 80502.5 ;
      RECT  10100.0 80437.5 10235.0 80502.5 ;
      RECT  10357.5 80222.5 10492.5 80287.5 ;
      RECT  10452.5 80437.5 10587.5 80502.5 ;
      RECT  10040.0 81142.5 10960.0 81207.5 ;
      RECT  10040.0 79797.5 10960.0 79862.5 ;
      RECT  11387.5 80990.0 11452.5 81175.0 ;
      RECT  11387.5 79830.0 11452.5 80015.0 ;
      RECT  11027.5 79947.5 11092.5 79797.5 ;
      RECT  11027.5 80832.5 11092.5 81207.5 ;
      RECT  11217.5 79947.5 11282.5 80832.5 ;
      RECT  11027.5 80832.5 11092.5 80967.5 ;
      RECT  11217.5 80832.5 11282.5 80967.5 ;
      RECT  11217.5 80832.5 11282.5 80967.5 ;
      RECT  11027.5 80832.5 11092.5 80967.5 ;
      RECT  11027.5 79947.5 11092.5 80082.5 ;
      RECT  11217.5 79947.5 11282.5 80082.5 ;
      RECT  11217.5 79947.5 11282.5 80082.5 ;
      RECT  11027.5 79947.5 11092.5 80082.5 ;
      RECT  11387.5 80922.5 11452.5 81057.5 ;
      RECT  11387.5 79947.5 11452.5 80082.5 ;
      RECT  11085.0 80390.0 11150.0 80525.0 ;
      RECT  11085.0 80390.0 11150.0 80525.0 ;
      RECT  11250.0 80425.0 11315.0 80490.0 ;
      RECT  10960.0 81142.5 11520.0 81207.5 ;
      RECT  10960.0 79797.5 11520.0 79862.5 ;
      RECT  9222.5 80390.0 9287.5 80525.0 ;
      RECT  9362.5 80117.5 9427.5 80252.5 ;
      RECT  10357.5 80222.5 10222.5 80287.5 ;
      RECT  9907.5 81360.0 9972.5 81175.0 ;
      RECT  9907.5 82520.0 9972.5 82335.0 ;
      RECT  9547.5 82402.5 9612.5 82552.5 ;
      RECT  9547.5 81517.5 9612.5 81142.5 ;
      RECT  9737.5 82402.5 9802.5 81517.5 ;
      RECT  9547.5 81517.5 9612.5 81382.5 ;
      RECT  9737.5 81517.5 9802.5 81382.5 ;
      RECT  9737.5 81517.5 9802.5 81382.5 ;
      RECT  9547.5 81517.5 9612.5 81382.5 ;
      RECT  9547.5 82402.5 9612.5 82267.5 ;
      RECT  9737.5 82402.5 9802.5 82267.5 ;
      RECT  9737.5 82402.5 9802.5 82267.5 ;
      RECT  9547.5 82402.5 9612.5 82267.5 ;
      RECT  9907.5 81427.5 9972.5 81292.5 ;
      RECT  9907.5 82402.5 9972.5 82267.5 ;
      RECT  9605.0 81960.0 9670.0 81825.0 ;
      RECT  9605.0 81960.0 9670.0 81825.0 ;
      RECT  9770.0 81925.0 9835.0 81860.0 ;
      RECT  9480.0 81207.5 10040.0 81142.5 ;
      RECT  9480.0 82552.5 10040.0 82487.5 ;
      RECT  10107.5 82357.5 10172.5 82552.5 ;
      RECT  10107.5 81517.5 10172.5 81142.5 ;
      RECT  10487.5 81517.5 10552.5 81142.5 ;
      RECT  10657.5 81360.0 10722.5 81175.0 ;
      RECT  10657.5 82520.0 10722.5 82335.0 ;
      RECT  10107.5 81517.5 10172.5 81382.5 ;
      RECT  10297.5 81517.5 10362.5 81382.5 ;
      RECT  10297.5 81517.5 10362.5 81382.5 ;
      RECT  10107.5 81517.5 10172.5 81382.5 ;
      RECT  10297.5 81517.5 10362.5 81382.5 ;
      RECT  10487.5 81517.5 10552.5 81382.5 ;
      RECT  10487.5 81517.5 10552.5 81382.5 ;
      RECT  10297.5 81517.5 10362.5 81382.5 ;
      RECT  10107.5 82357.5 10172.5 82222.5 ;
      RECT  10297.5 82357.5 10362.5 82222.5 ;
      RECT  10297.5 82357.5 10362.5 82222.5 ;
      RECT  10107.5 82357.5 10172.5 82222.5 ;
      RECT  10297.5 82357.5 10362.5 82222.5 ;
      RECT  10487.5 82357.5 10552.5 82222.5 ;
      RECT  10487.5 82357.5 10552.5 82222.5 ;
      RECT  10297.5 82357.5 10362.5 82222.5 ;
      RECT  10657.5 81427.5 10722.5 81292.5 ;
      RECT  10657.5 82402.5 10722.5 82267.5 ;
      RECT  10492.5 82127.5 10357.5 82062.5 ;
      RECT  10235.0 81912.5 10100.0 81847.5 ;
      RECT  10297.5 81517.5 10362.5 81382.5 ;
      RECT  10487.5 82357.5 10552.5 82222.5 ;
      RECT  10587.5 81912.5 10452.5 81847.5 ;
      RECT  10100.0 81912.5 10235.0 81847.5 ;
      RECT  10357.5 82127.5 10492.5 82062.5 ;
      RECT  10452.5 81912.5 10587.5 81847.5 ;
      RECT  10040.0 81207.5 10960.0 81142.5 ;
      RECT  10040.0 82552.5 10960.0 82487.5 ;
      RECT  11387.5 81360.0 11452.5 81175.0 ;
      RECT  11387.5 82520.0 11452.5 82335.0 ;
      RECT  11027.5 82402.5 11092.5 82552.5 ;
      RECT  11027.5 81517.5 11092.5 81142.5 ;
      RECT  11217.5 82402.5 11282.5 81517.5 ;
      RECT  11027.5 81517.5 11092.5 81382.5 ;
      RECT  11217.5 81517.5 11282.5 81382.5 ;
      RECT  11217.5 81517.5 11282.5 81382.5 ;
      RECT  11027.5 81517.5 11092.5 81382.5 ;
      RECT  11027.5 82402.5 11092.5 82267.5 ;
      RECT  11217.5 82402.5 11282.5 82267.5 ;
      RECT  11217.5 82402.5 11282.5 82267.5 ;
      RECT  11027.5 82402.5 11092.5 82267.5 ;
      RECT  11387.5 81427.5 11452.5 81292.5 ;
      RECT  11387.5 82402.5 11452.5 82267.5 ;
      RECT  11085.0 81960.0 11150.0 81825.0 ;
      RECT  11085.0 81960.0 11150.0 81825.0 ;
      RECT  11250.0 81925.0 11315.0 81860.0 ;
      RECT  10960.0 81207.5 11520.0 81142.5 ;
      RECT  10960.0 82552.5 11520.0 82487.5 ;
      RECT  9222.5 81825.0 9287.5 81960.0 ;
      RECT  9362.5 82097.5 9427.5 82232.5 ;
      RECT  10357.5 82062.5 10222.5 82127.5 ;
      RECT  9907.5 83680.0 9972.5 83865.0 ;
      RECT  9907.5 82520.0 9972.5 82705.0 ;
      RECT  9547.5 82637.5 9612.5 82487.5 ;
      RECT  9547.5 83522.5 9612.5 83897.5 ;
      RECT  9737.5 82637.5 9802.5 83522.5 ;
      RECT  9547.5 83522.5 9612.5 83657.5 ;
      RECT  9737.5 83522.5 9802.5 83657.5 ;
      RECT  9737.5 83522.5 9802.5 83657.5 ;
      RECT  9547.5 83522.5 9612.5 83657.5 ;
      RECT  9547.5 82637.5 9612.5 82772.5 ;
      RECT  9737.5 82637.5 9802.5 82772.5 ;
      RECT  9737.5 82637.5 9802.5 82772.5 ;
      RECT  9547.5 82637.5 9612.5 82772.5 ;
      RECT  9907.5 83612.5 9972.5 83747.5 ;
      RECT  9907.5 82637.5 9972.5 82772.5 ;
      RECT  9605.0 83080.0 9670.0 83215.0 ;
      RECT  9605.0 83080.0 9670.0 83215.0 ;
      RECT  9770.0 83115.0 9835.0 83180.0 ;
      RECT  9480.0 83832.5 10040.0 83897.5 ;
      RECT  9480.0 82487.5 10040.0 82552.5 ;
      RECT  10107.5 82682.5 10172.5 82487.5 ;
      RECT  10107.5 83522.5 10172.5 83897.5 ;
      RECT  10487.5 83522.5 10552.5 83897.5 ;
      RECT  10657.5 83680.0 10722.5 83865.0 ;
      RECT  10657.5 82520.0 10722.5 82705.0 ;
      RECT  10107.5 83522.5 10172.5 83657.5 ;
      RECT  10297.5 83522.5 10362.5 83657.5 ;
      RECT  10297.5 83522.5 10362.5 83657.5 ;
      RECT  10107.5 83522.5 10172.5 83657.5 ;
      RECT  10297.5 83522.5 10362.5 83657.5 ;
      RECT  10487.5 83522.5 10552.5 83657.5 ;
      RECT  10487.5 83522.5 10552.5 83657.5 ;
      RECT  10297.5 83522.5 10362.5 83657.5 ;
      RECT  10107.5 82682.5 10172.5 82817.5 ;
      RECT  10297.5 82682.5 10362.5 82817.5 ;
      RECT  10297.5 82682.5 10362.5 82817.5 ;
      RECT  10107.5 82682.5 10172.5 82817.5 ;
      RECT  10297.5 82682.5 10362.5 82817.5 ;
      RECT  10487.5 82682.5 10552.5 82817.5 ;
      RECT  10487.5 82682.5 10552.5 82817.5 ;
      RECT  10297.5 82682.5 10362.5 82817.5 ;
      RECT  10657.5 83612.5 10722.5 83747.5 ;
      RECT  10657.5 82637.5 10722.5 82772.5 ;
      RECT  10492.5 82912.5 10357.5 82977.5 ;
      RECT  10235.0 83127.5 10100.0 83192.5 ;
      RECT  10297.5 83522.5 10362.5 83657.5 ;
      RECT  10487.5 82682.5 10552.5 82817.5 ;
      RECT  10587.5 83127.5 10452.5 83192.5 ;
      RECT  10100.0 83127.5 10235.0 83192.5 ;
      RECT  10357.5 82912.5 10492.5 82977.5 ;
      RECT  10452.5 83127.5 10587.5 83192.5 ;
      RECT  10040.0 83832.5 10960.0 83897.5 ;
      RECT  10040.0 82487.5 10960.0 82552.5 ;
      RECT  11387.5 83680.0 11452.5 83865.0 ;
      RECT  11387.5 82520.0 11452.5 82705.0 ;
      RECT  11027.5 82637.5 11092.5 82487.5 ;
      RECT  11027.5 83522.5 11092.5 83897.5 ;
      RECT  11217.5 82637.5 11282.5 83522.5 ;
      RECT  11027.5 83522.5 11092.5 83657.5 ;
      RECT  11217.5 83522.5 11282.5 83657.5 ;
      RECT  11217.5 83522.5 11282.5 83657.5 ;
      RECT  11027.5 83522.5 11092.5 83657.5 ;
      RECT  11027.5 82637.5 11092.5 82772.5 ;
      RECT  11217.5 82637.5 11282.5 82772.5 ;
      RECT  11217.5 82637.5 11282.5 82772.5 ;
      RECT  11027.5 82637.5 11092.5 82772.5 ;
      RECT  11387.5 83612.5 11452.5 83747.5 ;
      RECT  11387.5 82637.5 11452.5 82772.5 ;
      RECT  11085.0 83080.0 11150.0 83215.0 ;
      RECT  11085.0 83080.0 11150.0 83215.0 ;
      RECT  11250.0 83115.0 11315.0 83180.0 ;
      RECT  10960.0 83832.5 11520.0 83897.5 ;
      RECT  10960.0 82487.5 11520.0 82552.5 ;
      RECT  9222.5 83080.0 9287.5 83215.0 ;
      RECT  9362.5 82807.5 9427.5 82942.5 ;
      RECT  10357.5 82912.5 10222.5 82977.5 ;
      RECT  9907.5 84050.0 9972.5 83865.0 ;
      RECT  9907.5 85210.0 9972.5 85025.0 ;
      RECT  9547.5 85092.5 9612.5 85242.5 ;
      RECT  9547.5 84207.5 9612.5 83832.5 ;
      RECT  9737.5 85092.5 9802.5 84207.5 ;
      RECT  9547.5 84207.5 9612.5 84072.5 ;
      RECT  9737.5 84207.5 9802.5 84072.5 ;
      RECT  9737.5 84207.5 9802.5 84072.5 ;
      RECT  9547.5 84207.5 9612.5 84072.5 ;
      RECT  9547.5 85092.5 9612.5 84957.5 ;
      RECT  9737.5 85092.5 9802.5 84957.5 ;
      RECT  9737.5 85092.5 9802.5 84957.5 ;
      RECT  9547.5 85092.5 9612.5 84957.5 ;
      RECT  9907.5 84117.5 9972.5 83982.5 ;
      RECT  9907.5 85092.5 9972.5 84957.5 ;
      RECT  9605.0 84650.0 9670.0 84515.0 ;
      RECT  9605.0 84650.0 9670.0 84515.0 ;
      RECT  9770.0 84615.0 9835.0 84550.0 ;
      RECT  9480.0 83897.5 10040.0 83832.5 ;
      RECT  9480.0 85242.5 10040.0 85177.5 ;
      RECT  10107.5 85047.5 10172.5 85242.5 ;
      RECT  10107.5 84207.5 10172.5 83832.5 ;
      RECT  10487.5 84207.5 10552.5 83832.5 ;
      RECT  10657.5 84050.0 10722.5 83865.0 ;
      RECT  10657.5 85210.0 10722.5 85025.0 ;
      RECT  10107.5 84207.5 10172.5 84072.5 ;
      RECT  10297.5 84207.5 10362.5 84072.5 ;
      RECT  10297.5 84207.5 10362.5 84072.5 ;
      RECT  10107.5 84207.5 10172.5 84072.5 ;
      RECT  10297.5 84207.5 10362.5 84072.5 ;
      RECT  10487.5 84207.5 10552.5 84072.5 ;
      RECT  10487.5 84207.5 10552.5 84072.5 ;
      RECT  10297.5 84207.5 10362.5 84072.5 ;
      RECT  10107.5 85047.5 10172.5 84912.5 ;
      RECT  10297.5 85047.5 10362.5 84912.5 ;
      RECT  10297.5 85047.5 10362.5 84912.5 ;
      RECT  10107.5 85047.5 10172.5 84912.5 ;
      RECT  10297.5 85047.5 10362.5 84912.5 ;
      RECT  10487.5 85047.5 10552.5 84912.5 ;
      RECT  10487.5 85047.5 10552.5 84912.5 ;
      RECT  10297.5 85047.5 10362.5 84912.5 ;
      RECT  10657.5 84117.5 10722.5 83982.5 ;
      RECT  10657.5 85092.5 10722.5 84957.5 ;
      RECT  10492.5 84817.5 10357.5 84752.5 ;
      RECT  10235.0 84602.5 10100.0 84537.5 ;
      RECT  10297.5 84207.5 10362.5 84072.5 ;
      RECT  10487.5 85047.5 10552.5 84912.5 ;
      RECT  10587.5 84602.5 10452.5 84537.5 ;
      RECT  10100.0 84602.5 10235.0 84537.5 ;
      RECT  10357.5 84817.5 10492.5 84752.5 ;
      RECT  10452.5 84602.5 10587.5 84537.5 ;
      RECT  10040.0 83897.5 10960.0 83832.5 ;
      RECT  10040.0 85242.5 10960.0 85177.5 ;
      RECT  11387.5 84050.0 11452.5 83865.0 ;
      RECT  11387.5 85210.0 11452.5 85025.0 ;
      RECT  11027.5 85092.5 11092.5 85242.5 ;
      RECT  11027.5 84207.5 11092.5 83832.5 ;
      RECT  11217.5 85092.5 11282.5 84207.5 ;
      RECT  11027.5 84207.5 11092.5 84072.5 ;
      RECT  11217.5 84207.5 11282.5 84072.5 ;
      RECT  11217.5 84207.5 11282.5 84072.5 ;
      RECT  11027.5 84207.5 11092.5 84072.5 ;
      RECT  11027.5 85092.5 11092.5 84957.5 ;
      RECT  11217.5 85092.5 11282.5 84957.5 ;
      RECT  11217.5 85092.5 11282.5 84957.5 ;
      RECT  11027.5 85092.5 11092.5 84957.5 ;
      RECT  11387.5 84117.5 11452.5 83982.5 ;
      RECT  11387.5 85092.5 11452.5 84957.5 ;
      RECT  11085.0 84650.0 11150.0 84515.0 ;
      RECT  11085.0 84650.0 11150.0 84515.0 ;
      RECT  11250.0 84615.0 11315.0 84550.0 ;
      RECT  10960.0 83897.5 11520.0 83832.5 ;
      RECT  10960.0 85242.5 11520.0 85177.5 ;
      RECT  9222.5 84515.0 9287.5 84650.0 ;
      RECT  9362.5 84787.5 9427.5 84922.5 ;
      RECT  10357.5 84752.5 10222.5 84817.5 ;
      RECT  9907.5 86370.0 9972.5 86555.0 ;
      RECT  9907.5 85210.0 9972.5 85395.0 ;
      RECT  9547.5 85327.5 9612.5 85177.5 ;
      RECT  9547.5 86212.5 9612.5 86587.5 ;
      RECT  9737.5 85327.5 9802.5 86212.5 ;
      RECT  9547.5 86212.5 9612.5 86347.5 ;
      RECT  9737.5 86212.5 9802.5 86347.5 ;
      RECT  9737.5 86212.5 9802.5 86347.5 ;
      RECT  9547.5 86212.5 9612.5 86347.5 ;
      RECT  9547.5 85327.5 9612.5 85462.5 ;
      RECT  9737.5 85327.5 9802.5 85462.5 ;
      RECT  9737.5 85327.5 9802.5 85462.5 ;
      RECT  9547.5 85327.5 9612.5 85462.5 ;
      RECT  9907.5 86302.5 9972.5 86437.5 ;
      RECT  9907.5 85327.5 9972.5 85462.5 ;
      RECT  9605.0 85770.0 9670.0 85905.0 ;
      RECT  9605.0 85770.0 9670.0 85905.0 ;
      RECT  9770.0 85805.0 9835.0 85870.0 ;
      RECT  9480.0 86522.5 10040.0 86587.5 ;
      RECT  9480.0 85177.5 10040.0 85242.5 ;
      RECT  10107.5 85372.5 10172.5 85177.5 ;
      RECT  10107.5 86212.5 10172.5 86587.5 ;
      RECT  10487.5 86212.5 10552.5 86587.5 ;
      RECT  10657.5 86370.0 10722.5 86555.0 ;
      RECT  10657.5 85210.0 10722.5 85395.0 ;
      RECT  10107.5 86212.5 10172.5 86347.5 ;
      RECT  10297.5 86212.5 10362.5 86347.5 ;
      RECT  10297.5 86212.5 10362.5 86347.5 ;
      RECT  10107.5 86212.5 10172.5 86347.5 ;
      RECT  10297.5 86212.5 10362.5 86347.5 ;
      RECT  10487.5 86212.5 10552.5 86347.5 ;
      RECT  10487.5 86212.5 10552.5 86347.5 ;
      RECT  10297.5 86212.5 10362.5 86347.5 ;
      RECT  10107.5 85372.5 10172.5 85507.5 ;
      RECT  10297.5 85372.5 10362.5 85507.5 ;
      RECT  10297.5 85372.5 10362.5 85507.5 ;
      RECT  10107.5 85372.5 10172.5 85507.5 ;
      RECT  10297.5 85372.5 10362.5 85507.5 ;
      RECT  10487.5 85372.5 10552.5 85507.5 ;
      RECT  10487.5 85372.5 10552.5 85507.5 ;
      RECT  10297.5 85372.5 10362.5 85507.5 ;
      RECT  10657.5 86302.5 10722.5 86437.5 ;
      RECT  10657.5 85327.5 10722.5 85462.5 ;
      RECT  10492.5 85602.5 10357.5 85667.5 ;
      RECT  10235.0 85817.5 10100.0 85882.5 ;
      RECT  10297.5 86212.5 10362.5 86347.5 ;
      RECT  10487.5 85372.5 10552.5 85507.5 ;
      RECT  10587.5 85817.5 10452.5 85882.5 ;
      RECT  10100.0 85817.5 10235.0 85882.5 ;
      RECT  10357.5 85602.5 10492.5 85667.5 ;
      RECT  10452.5 85817.5 10587.5 85882.5 ;
      RECT  10040.0 86522.5 10960.0 86587.5 ;
      RECT  10040.0 85177.5 10960.0 85242.5 ;
      RECT  11387.5 86370.0 11452.5 86555.0 ;
      RECT  11387.5 85210.0 11452.5 85395.0 ;
      RECT  11027.5 85327.5 11092.5 85177.5 ;
      RECT  11027.5 86212.5 11092.5 86587.5 ;
      RECT  11217.5 85327.5 11282.5 86212.5 ;
      RECT  11027.5 86212.5 11092.5 86347.5 ;
      RECT  11217.5 86212.5 11282.5 86347.5 ;
      RECT  11217.5 86212.5 11282.5 86347.5 ;
      RECT  11027.5 86212.5 11092.5 86347.5 ;
      RECT  11027.5 85327.5 11092.5 85462.5 ;
      RECT  11217.5 85327.5 11282.5 85462.5 ;
      RECT  11217.5 85327.5 11282.5 85462.5 ;
      RECT  11027.5 85327.5 11092.5 85462.5 ;
      RECT  11387.5 86302.5 11452.5 86437.5 ;
      RECT  11387.5 85327.5 11452.5 85462.5 ;
      RECT  11085.0 85770.0 11150.0 85905.0 ;
      RECT  11085.0 85770.0 11150.0 85905.0 ;
      RECT  11250.0 85805.0 11315.0 85870.0 ;
      RECT  10960.0 86522.5 11520.0 86587.5 ;
      RECT  10960.0 85177.5 11520.0 85242.5 ;
      RECT  9222.5 85770.0 9287.5 85905.0 ;
      RECT  9362.5 85497.5 9427.5 85632.5 ;
      RECT  10357.5 85602.5 10222.5 85667.5 ;
      RECT  9907.5 86740.0 9972.5 86555.0 ;
      RECT  9907.5 87900.0 9972.5 87715.0 ;
      RECT  9547.5 87782.5 9612.5 87932.5 ;
      RECT  9547.5 86897.5 9612.5 86522.5 ;
      RECT  9737.5 87782.5 9802.5 86897.5 ;
      RECT  9547.5 86897.5 9612.5 86762.5 ;
      RECT  9737.5 86897.5 9802.5 86762.5 ;
      RECT  9737.5 86897.5 9802.5 86762.5 ;
      RECT  9547.5 86897.5 9612.5 86762.5 ;
      RECT  9547.5 87782.5 9612.5 87647.5 ;
      RECT  9737.5 87782.5 9802.5 87647.5 ;
      RECT  9737.5 87782.5 9802.5 87647.5 ;
      RECT  9547.5 87782.5 9612.5 87647.5 ;
      RECT  9907.5 86807.5 9972.5 86672.5 ;
      RECT  9907.5 87782.5 9972.5 87647.5 ;
      RECT  9605.0 87340.0 9670.0 87205.0 ;
      RECT  9605.0 87340.0 9670.0 87205.0 ;
      RECT  9770.0 87305.0 9835.0 87240.0 ;
      RECT  9480.0 86587.5 10040.0 86522.5 ;
      RECT  9480.0 87932.5 10040.0 87867.5 ;
      RECT  10107.5 87737.5 10172.5 87932.5 ;
      RECT  10107.5 86897.5 10172.5 86522.5 ;
      RECT  10487.5 86897.5 10552.5 86522.5 ;
      RECT  10657.5 86740.0 10722.5 86555.0 ;
      RECT  10657.5 87900.0 10722.5 87715.0 ;
      RECT  10107.5 86897.5 10172.5 86762.5 ;
      RECT  10297.5 86897.5 10362.5 86762.5 ;
      RECT  10297.5 86897.5 10362.5 86762.5 ;
      RECT  10107.5 86897.5 10172.5 86762.5 ;
      RECT  10297.5 86897.5 10362.5 86762.5 ;
      RECT  10487.5 86897.5 10552.5 86762.5 ;
      RECT  10487.5 86897.5 10552.5 86762.5 ;
      RECT  10297.5 86897.5 10362.5 86762.5 ;
      RECT  10107.5 87737.5 10172.5 87602.5 ;
      RECT  10297.5 87737.5 10362.5 87602.5 ;
      RECT  10297.5 87737.5 10362.5 87602.5 ;
      RECT  10107.5 87737.5 10172.5 87602.5 ;
      RECT  10297.5 87737.5 10362.5 87602.5 ;
      RECT  10487.5 87737.5 10552.5 87602.5 ;
      RECT  10487.5 87737.5 10552.5 87602.5 ;
      RECT  10297.5 87737.5 10362.5 87602.5 ;
      RECT  10657.5 86807.5 10722.5 86672.5 ;
      RECT  10657.5 87782.5 10722.5 87647.5 ;
      RECT  10492.5 87507.5 10357.5 87442.5 ;
      RECT  10235.0 87292.5 10100.0 87227.5 ;
      RECT  10297.5 86897.5 10362.5 86762.5 ;
      RECT  10487.5 87737.5 10552.5 87602.5 ;
      RECT  10587.5 87292.5 10452.5 87227.5 ;
      RECT  10100.0 87292.5 10235.0 87227.5 ;
      RECT  10357.5 87507.5 10492.5 87442.5 ;
      RECT  10452.5 87292.5 10587.5 87227.5 ;
      RECT  10040.0 86587.5 10960.0 86522.5 ;
      RECT  10040.0 87932.5 10960.0 87867.5 ;
      RECT  11387.5 86740.0 11452.5 86555.0 ;
      RECT  11387.5 87900.0 11452.5 87715.0 ;
      RECT  11027.5 87782.5 11092.5 87932.5 ;
      RECT  11027.5 86897.5 11092.5 86522.5 ;
      RECT  11217.5 87782.5 11282.5 86897.5 ;
      RECT  11027.5 86897.5 11092.5 86762.5 ;
      RECT  11217.5 86897.5 11282.5 86762.5 ;
      RECT  11217.5 86897.5 11282.5 86762.5 ;
      RECT  11027.5 86897.5 11092.5 86762.5 ;
      RECT  11027.5 87782.5 11092.5 87647.5 ;
      RECT  11217.5 87782.5 11282.5 87647.5 ;
      RECT  11217.5 87782.5 11282.5 87647.5 ;
      RECT  11027.5 87782.5 11092.5 87647.5 ;
      RECT  11387.5 86807.5 11452.5 86672.5 ;
      RECT  11387.5 87782.5 11452.5 87647.5 ;
      RECT  11085.0 87340.0 11150.0 87205.0 ;
      RECT  11085.0 87340.0 11150.0 87205.0 ;
      RECT  11250.0 87305.0 11315.0 87240.0 ;
      RECT  10960.0 86587.5 11520.0 86522.5 ;
      RECT  10960.0 87932.5 11520.0 87867.5 ;
      RECT  9222.5 87205.0 9287.5 87340.0 ;
      RECT  9362.5 87477.5 9427.5 87612.5 ;
      RECT  10357.5 87442.5 10222.5 87507.5 ;
      RECT  9907.5 89060.0 9972.5 89245.0 ;
      RECT  9907.5 87900.0 9972.5 88085.0 ;
      RECT  9547.5 88017.5 9612.5 87867.5 ;
      RECT  9547.5 88902.5 9612.5 89277.5 ;
      RECT  9737.5 88017.5 9802.5 88902.5 ;
      RECT  9547.5 88902.5 9612.5 89037.5 ;
      RECT  9737.5 88902.5 9802.5 89037.5 ;
      RECT  9737.5 88902.5 9802.5 89037.5 ;
      RECT  9547.5 88902.5 9612.5 89037.5 ;
      RECT  9547.5 88017.5 9612.5 88152.5 ;
      RECT  9737.5 88017.5 9802.5 88152.5 ;
      RECT  9737.5 88017.5 9802.5 88152.5 ;
      RECT  9547.5 88017.5 9612.5 88152.5 ;
      RECT  9907.5 88992.5 9972.5 89127.5 ;
      RECT  9907.5 88017.5 9972.5 88152.5 ;
      RECT  9605.0 88460.0 9670.0 88595.0 ;
      RECT  9605.0 88460.0 9670.0 88595.0 ;
      RECT  9770.0 88495.0 9835.0 88560.0 ;
      RECT  9480.0 89212.5 10040.0 89277.5 ;
      RECT  9480.0 87867.5 10040.0 87932.5 ;
      RECT  10107.5 88062.5 10172.5 87867.5 ;
      RECT  10107.5 88902.5 10172.5 89277.5 ;
      RECT  10487.5 88902.5 10552.5 89277.5 ;
      RECT  10657.5 89060.0 10722.5 89245.0 ;
      RECT  10657.5 87900.0 10722.5 88085.0 ;
      RECT  10107.5 88902.5 10172.5 89037.5 ;
      RECT  10297.5 88902.5 10362.5 89037.5 ;
      RECT  10297.5 88902.5 10362.5 89037.5 ;
      RECT  10107.5 88902.5 10172.5 89037.5 ;
      RECT  10297.5 88902.5 10362.5 89037.5 ;
      RECT  10487.5 88902.5 10552.5 89037.5 ;
      RECT  10487.5 88902.5 10552.5 89037.5 ;
      RECT  10297.5 88902.5 10362.5 89037.5 ;
      RECT  10107.5 88062.5 10172.5 88197.5 ;
      RECT  10297.5 88062.5 10362.5 88197.5 ;
      RECT  10297.5 88062.5 10362.5 88197.5 ;
      RECT  10107.5 88062.5 10172.5 88197.5 ;
      RECT  10297.5 88062.5 10362.5 88197.5 ;
      RECT  10487.5 88062.5 10552.5 88197.5 ;
      RECT  10487.5 88062.5 10552.5 88197.5 ;
      RECT  10297.5 88062.5 10362.5 88197.5 ;
      RECT  10657.5 88992.5 10722.5 89127.5 ;
      RECT  10657.5 88017.5 10722.5 88152.5 ;
      RECT  10492.5 88292.5 10357.5 88357.5 ;
      RECT  10235.0 88507.5 10100.0 88572.5 ;
      RECT  10297.5 88902.5 10362.5 89037.5 ;
      RECT  10487.5 88062.5 10552.5 88197.5 ;
      RECT  10587.5 88507.5 10452.5 88572.5 ;
      RECT  10100.0 88507.5 10235.0 88572.5 ;
      RECT  10357.5 88292.5 10492.5 88357.5 ;
      RECT  10452.5 88507.5 10587.5 88572.5 ;
      RECT  10040.0 89212.5 10960.0 89277.5 ;
      RECT  10040.0 87867.5 10960.0 87932.5 ;
      RECT  11387.5 89060.0 11452.5 89245.0 ;
      RECT  11387.5 87900.0 11452.5 88085.0 ;
      RECT  11027.5 88017.5 11092.5 87867.5 ;
      RECT  11027.5 88902.5 11092.5 89277.5 ;
      RECT  11217.5 88017.5 11282.5 88902.5 ;
      RECT  11027.5 88902.5 11092.5 89037.5 ;
      RECT  11217.5 88902.5 11282.5 89037.5 ;
      RECT  11217.5 88902.5 11282.5 89037.5 ;
      RECT  11027.5 88902.5 11092.5 89037.5 ;
      RECT  11027.5 88017.5 11092.5 88152.5 ;
      RECT  11217.5 88017.5 11282.5 88152.5 ;
      RECT  11217.5 88017.5 11282.5 88152.5 ;
      RECT  11027.5 88017.5 11092.5 88152.5 ;
      RECT  11387.5 88992.5 11452.5 89127.5 ;
      RECT  11387.5 88017.5 11452.5 88152.5 ;
      RECT  11085.0 88460.0 11150.0 88595.0 ;
      RECT  11085.0 88460.0 11150.0 88595.0 ;
      RECT  11250.0 88495.0 11315.0 88560.0 ;
      RECT  10960.0 89212.5 11520.0 89277.5 ;
      RECT  10960.0 87867.5 11520.0 87932.5 ;
      RECT  9222.5 88460.0 9287.5 88595.0 ;
      RECT  9362.5 88187.5 9427.5 88322.5 ;
      RECT  10357.5 88292.5 10222.5 88357.5 ;
      RECT  9907.5 89430.0 9972.5 89245.0 ;
      RECT  9907.5 90590.0 9972.5 90405.0 ;
      RECT  9547.5 90472.5 9612.5 90622.5 ;
      RECT  9547.5 89587.5 9612.5 89212.5 ;
      RECT  9737.5 90472.5 9802.5 89587.5 ;
      RECT  9547.5 89587.5 9612.5 89452.5 ;
      RECT  9737.5 89587.5 9802.5 89452.5 ;
      RECT  9737.5 89587.5 9802.5 89452.5 ;
      RECT  9547.5 89587.5 9612.5 89452.5 ;
      RECT  9547.5 90472.5 9612.5 90337.5 ;
      RECT  9737.5 90472.5 9802.5 90337.5 ;
      RECT  9737.5 90472.5 9802.5 90337.5 ;
      RECT  9547.5 90472.5 9612.5 90337.5 ;
      RECT  9907.5 89497.5 9972.5 89362.5 ;
      RECT  9907.5 90472.5 9972.5 90337.5 ;
      RECT  9605.0 90030.0 9670.0 89895.0 ;
      RECT  9605.0 90030.0 9670.0 89895.0 ;
      RECT  9770.0 89995.0 9835.0 89930.0 ;
      RECT  9480.0 89277.5 10040.0 89212.5 ;
      RECT  9480.0 90622.5 10040.0 90557.5 ;
      RECT  10107.5 90427.5 10172.5 90622.5 ;
      RECT  10107.5 89587.5 10172.5 89212.5 ;
      RECT  10487.5 89587.5 10552.5 89212.5 ;
      RECT  10657.5 89430.0 10722.5 89245.0 ;
      RECT  10657.5 90590.0 10722.5 90405.0 ;
      RECT  10107.5 89587.5 10172.5 89452.5 ;
      RECT  10297.5 89587.5 10362.5 89452.5 ;
      RECT  10297.5 89587.5 10362.5 89452.5 ;
      RECT  10107.5 89587.5 10172.5 89452.5 ;
      RECT  10297.5 89587.5 10362.5 89452.5 ;
      RECT  10487.5 89587.5 10552.5 89452.5 ;
      RECT  10487.5 89587.5 10552.5 89452.5 ;
      RECT  10297.5 89587.5 10362.5 89452.5 ;
      RECT  10107.5 90427.5 10172.5 90292.5 ;
      RECT  10297.5 90427.5 10362.5 90292.5 ;
      RECT  10297.5 90427.5 10362.5 90292.5 ;
      RECT  10107.5 90427.5 10172.5 90292.5 ;
      RECT  10297.5 90427.5 10362.5 90292.5 ;
      RECT  10487.5 90427.5 10552.5 90292.5 ;
      RECT  10487.5 90427.5 10552.5 90292.5 ;
      RECT  10297.5 90427.5 10362.5 90292.5 ;
      RECT  10657.5 89497.5 10722.5 89362.5 ;
      RECT  10657.5 90472.5 10722.5 90337.5 ;
      RECT  10492.5 90197.5 10357.5 90132.5 ;
      RECT  10235.0 89982.5 10100.0 89917.5 ;
      RECT  10297.5 89587.5 10362.5 89452.5 ;
      RECT  10487.5 90427.5 10552.5 90292.5 ;
      RECT  10587.5 89982.5 10452.5 89917.5 ;
      RECT  10100.0 89982.5 10235.0 89917.5 ;
      RECT  10357.5 90197.5 10492.5 90132.5 ;
      RECT  10452.5 89982.5 10587.5 89917.5 ;
      RECT  10040.0 89277.5 10960.0 89212.5 ;
      RECT  10040.0 90622.5 10960.0 90557.5 ;
      RECT  11387.5 89430.0 11452.5 89245.0 ;
      RECT  11387.5 90590.0 11452.5 90405.0 ;
      RECT  11027.5 90472.5 11092.5 90622.5 ;
      RECT  11027.5 89587.5 11092.5 89212.5 ;
      RECT  11217.5 90472.5 11282.5 89587.5 ;
      RECT  11027.5 89587.5 11092.5 89452.5 ;
      RECT  11217.5 89587.5 11282.5 89452.5 ;
      RECT  11217.5 89587.5 11282.5 89452.5 ;
      RECT  11027.5 89587.5 11092.5 89452.5 ;
      RECT  11027.5 90472.5 11092.5 90337.5 ;
      RECT  11217.5 90472.5 11282.5 90337.5 ;
      RECT  11217.5 90472.5 11282.5 90337.5 ;
      RECT  11027.5 90472.5 11092.5 90337.5 ;
      RECT  11387.5 89497.5 11452.5 89362.5 ;
      RECT  11387.5 90472.5 11452.5 90337.5 ;
      RECT  11085.0 90030.0 11150.0 89895.0 ;
      RECT  11085.0 90030.0 11150.0 89895.0 ;
      RECT  11250.0 89995.0 11315.0 89930.0 ;
      RECT  10960.0 89277.5 11520.0 89212.5 ;
      RECT  10960.0 90622.5 11520.0 90557.5 ;
      RECT  9222.5 89895.0 9287.5 90030.0 ;
      RECT  9362.5 90167.5 9427.5 90302.5 ;
      RECT  10357.5 90132.5 10222.5 90197.5 ;
      RECT  9907.5 91750.0 9972.5 91935.0 ;
      RECT  9907.5 90590.0 9972.5 90775.0 ;
      RECT  9547.5 90707.5 9612.5 90557.5 ;
      RECT  9547.5 91592.5 9612.5 91967.5 ;
      RECT  9737.5 90707.5 9802.5 91592.5 ;
      RECT  9547.5 91592.5 9612.5 91727.5 ;
      RECT  9737.5 91592.5 9802.5 91727.5 ;
      RECT  9737.5 91592.5 9802.5 91727.5 ;
      RECT  9547.5 91592.5 9612.5 91727.5 ;
      RECT  9547.5 90707.5 9612.5 90842.5 ;
      RECT  9737.5 90707.5 9802.5 90842.5 ;
      RECT  9737.5 90707.5 9802.5 90842.5 ;
      RECT  9547.5 90707.5 9612.5 90842.5 ;
      RECT  9907.5 91682.5 9972.5 91817.5 ;
      RECT  9907.5 90707.5 9972.5 90842.5 ;
      RECT  9605.0 91150.0 9670.0 91285.0 ;
      RECT  9605.0 91150.0 9670.0 91285.0 ;
      RECT  9770.0 91185.0 9835.0 91250.0 ;
      RECT  9480.0 91902.5 10040.0 91967.5 ;
      RECT  9480.0 90557.5 10040.0 90622.5 ;
      RECT  10107.5 90752.5 10172.5 90557.5 ;
      RECT  10107.5 91592.5 10172.5 91967.5 ;
      RECT  10487.5 91592.5 10552.5 91967.5 ;
      RECT  10657.5 91750.0 10722.5 91935.0 ;
      RECT  10657.5 90590.0 10722.5 90775.0 ;
      RECT  10107.5 91592.5 10172.5 91727.5 ;
      RECT  10297.5 91592.5 10362.5 91727.5 ;
      RECT  10297.5 91592.5 10362.5 91727.5 ;
      RECT  10107.5 91592.5 10172.5 91727.5 ;
      RECT  10297.5 91592.5 10362.5 91727.5 ;
      RECT  10487.5 91592.5 10552.5 91727.5 ;
      RECT  10487.5 91592.5 10552.5 91727.5 ;
      RECT  10297.5 91592.5 10362.5 91727.5 ;
      RECT  10107.5 90752.5 10172.5 90887.5 ;
      RECT  10297.5 90752.5 10362.5 90887.5 ;
      RECT  10297.5 90752.5 10362.5 90887.5 ;
      RECT  10107.5 90752.5 10172.5 90887.5 ;
      RECT  10297.5 90752.5 10362.5 90887.5 ;
      RECT  10487.5 90752.5 10552.5 90887.5 ;
      RECT  10487.5 90752.5 10552.5 90887.5 ;
      RECT  10297.5 90752.5 10362.5 90887.5 ;
      RECT  10657.5 91682.5 10722.5 91817.5 ;
      RECT  10657.5 90707.5 10722.5 90842.5 ;
      RECT  10492.5 90982.5 10357.5 91047.5 ;
      RECT  10235.0 91197.5 10100.0 91262.5 ;
      RECT  10297.5 91592.5 10362.5 91727.5 ;
      RECT  10487.5 90752.5 10552.5 90887.5 ;
      RECT  10587.5 91197.5 10452.5 91262.5 ;
      RECT  10100.0 91197.5 10235.0 91262.5 ;
      RECT  10357.5 90982.5 10492.5 91047.5 ;
      RECT  10452.5 91197.5 10587.5 91262.5 ;
      RECT  10040.0 91902.5 10960.0 91967.5 ;
      RECT  10040.0 90557.5 10960.0 90622.5 ;
      RECT  11387.5 91750.0 11452.5 91935.0 ;
      RECT  11387.5 90590.0 11452.5 90775.0 ;
      RECT  11027.5 90707.5 11092.5 90557.5 ;
      RECT  11027.5 91592.5 11092.5 91967.5 ;
      RECT  11217.5 90707.5 11282.5 91592.5 ;
      RECT  11027.5 91592.5 11092.5 91727.5 ;
      RECT  11217.5 91592.5 11282.5 91727.5 ;
      RECT  11217.5 91592.5 11282.5 91727.5 ;
      RECT  11027.5 91592.5 11092.5 91727.5 ;
      RECT  11027.5 90707.5 11092.5 90842.5 ;
      RECT  11217.5 90707.5 11282.5 90842.5 ;
      RECT  11217.5 90707.5 11282.5 90842.5 ;
      RECT  11027.5 90707.5 11092.5 90842.5 ;
      RECT  11387.5 91682.5 11452.5 91817.5 ;
      RECT  11387.5 90707.5 11452.5 90842.5 ;
      RECT  11085.0 91150.0 11150.0 91285.0 ;
      RECT  11085.0 91150.0 11150.0 91285.0 ;
      RECT  11250.0 91185.0 11315.0 91250.0 ;
      RECT  10960.0 91902.5 11520.0 91967.5 ;
      RECT  10960.0 90557.5 11520.0 90622.5 ;
      RECT  9222.5 91150.0 9287.5 91285.0 ;
      RECT  9362.5 90877.5 9427.5 91012.5 ;
      RECT  10357.5 90982.5 10222.5 91047.5 ;
      RECT  9907.5 92120.0 9972.5 91935.0 ;
      RECT  9907.5 93280.0 9972.5 93095.0 ;
      RECT  9547.5 93162.5 9612.5 93312.5 ;
      RECT  9547.5 92277.5 9612.5 91902.5 ;
      RECT  9737.5 93162.5 9802.5 92277.5 ;
      RECT  9547.5 92277.5 9612.5 92142.5 ;
      RECT  9737.5 92277.5 9802.5 92142.5 ;
      RECT  9737.5 92277.5 9802.5 92142.5 ;
      RECT  9547.5 92277.5 9612.5 92142.5 ;
      RECT  9547.5 93162.5 9612.5 93027.5 ;
      RECT  9737.5 93162.5 9802.5 93027.5 ;
      RECT  9737.5 93162.5 9802.5 93027.5 ;
      RECT  9547.5 93162.5 9612.5 93027.5 ;
      RECT  9907.5 92187.5 9972.5 92052.5 ;
      RECT  9907.5 93162.5 9972.5 93027.5 ;
      RECT  9605.0 92720.0 9670.0 92585.0 ;
      RECT  9605.0 92720.0 9670.0 92585.0 ;
      RECT  9770.0 92685.0 9835.0 92620.0 ;
      RECT  9480.0 91967.5 10040.0 91902.5 ;
      RECT  9480.0 93312.5 10040.0 93247.5 ;
      RECT  10107.5 93117.5 10172.5 93312.5 ;
      RECT  10107.5 92277.5 10172.5 91902.5 ;
      RECT  10487.5 92277.5 10552.5 91902.5 ;
      RECT  10657.5 92120.0 10722.5 91935.0 ;
      RECT  10657.5 93280.0 10722.5 93095.0 ;
      RECT  10107.5 92277.5 10172.5 92142.5 ;
      RECT  10297.5 92277.5 10362.5 92142.5 ;
      RECT  10297.5 92277.5 10362.5 92142.5 ;
      RECT  10107.5 92277.5 10172.5 92142.5 ;
      RECT  10297.5 92277.5 10362.5 92142.5 ;
      RECT  10487.5 92277.5 10552.5 92142.5 ;
      RECT  10487.5 92277.5 10552.5 92142.5 ;
      RECT  10297.5 92277.5 10362.5 92142.5 ;
      RECT  10107.5 93117.5 10172.5 92982.5 ;
      RECT  10297.5 93117.5 10362.5 92982.5 ;
      RECT  10297.5 93117.5 10362.5 92982.5 ;
      RECT  10107.5 93117.5 10172.5 92982.5 ;
      RECT  10297.5 93117.5 10362.5 92982.5 ;
      RECT  10487.5 93117.5 10552.5 92982.5 ;
      RECT  10487.5 93117.5 10552.5 92982.5 ;
      RECT  10297.5 93117.5 10362.5 92982.5 ;
      RECT  10657.5 92187.5 10722.5 92052.5 ;
      RECT  10657.5 93162.5 10722.5 93027.5 ;
      RECT  10492.5 92887.5 10357.5 92822.5 ;
      RECT  10235.0 92672.5 10100.0 92607.5 ;
      RECT  10297.5 92277.5 10362.5 92142.5 ;
      RECT  10487.5 93117.5 10552.5 92982.5 ;
      RECT  10587.5 92672.5 10452.5 92607.5 ;
      RECT  10100.0 92672.5 10235.0 92607.5 ;
      RECT  10357.5 92887.5 10492.5 92822.5 ;
      RECT  10452.5 92672.5 10587.5 92607.5 ;
      RECT  10040.0 91967.5 10960.0 91902.5 ;
      RECT  10040.0 93312.5 10960.0 93247.5 ;
      RECT  11387.5 92120.0 11452.5 91935.0 ;
      RECT  11387.5 93280.0 11452.5 93095.0 ;
      RECT  11027.5 93162.5 11092.5 93312.5 ;
      RECT  11027.5 92277.5 11092.5 91902.5 ;
      RECT  11217.5 93162.5 11282.5 92277.5 ;
      RECT  11027.5 92277.5 11092.5 92142.5 ;
      RECT  11217.5 92277.5 11282.5 92142.5 ;
      RECT  11217.5 92277.5 11282.5 92142.5 ;
      RECT  11027.5 92277.5 11092.5 92142.5 ;
      RECT  11027.5 93162.5 11092.5 93027.5 ;
      RECT  11217.5 93162.5 11282.5 93027.5 ;
      RECT  11217.5 93162.5 11282.5 93027.5 ;
      RECT  11027.5 93162.5 11092.5 93027.5 ;
      RECT  11387.5 92187.5 11452.5 92052.5 ;
      RECT  11387.5 93162.5 11452.5 93027.5 ;
      RECT  11085.0 92720.0 11150.0 92585.0 ;
      RECT  11085.0 92720.0 11150.0 92585.0 ;
      RECT  11250.0 92685.0 11315.0 92620.0 ;
      RECT  10960.0 91967.5 11520.0 91902.5 ;
      RECT  10960.0 93312.5 11520.0 93247.5 ;
      RECT  9222.5 92585.0 9287.5 92720.0 ;
      RECT  9362.5 92857.5 9427.5 92992.5 ;
      RECT  10357.5 92822.5 10222.5 92887.5 ;
      RECT  9907.5 94440.0 9972.5 94625.0 ;
      RECT  9907.5 93280.0 9972.5 93465.0 ;
      RECT  9547.5 93397.5 9612.5 93247.5 ;
      RECT  9547.5 94282.5 9612.5 94657.5 ;
      RECT  9737.5 93397.5 9802.5 94282.5 ;
      RECT  9547.5 94282.5 9612.5 94417.5 ;
      RECT  9737.5 94282.5 9802.5 94417.5 ;
      RECT  9737.5 94282.5 9802.5 94417.5 ;
      RECT  9547.5 94282.5 9612.5 94417.5 ;
      RECT  9547.5 93397.5 9612.5 93532.5 ;
      RECT  9737.5 93397.5 9802.5 93532.5 ;
      RECT  9737.5 93397.5 9802.5 93532.5 ;
      RECT  9547.5 93397.5 9612.5 93532.5 ;
      RECT  9907.5 94372.5 9972.5 94507.5 ;
      RECT  9907.5 93397.5 9972.5 93532.5 ;
      RECT  9605.0 93840.0 9670.0 93975.0 ;
      RECT  9605.0 93840.0 9670.0 93975.0 ;
      RECT  9770.0 93875.0 9835.0 93940.0 ;
      RECT  9480.0 94592.5 10040.0 94657.5 ;
      RECT  9480.0 93247.5 10040.0 93312.5 ;
      RECT  10107.5 93442.5 10172.5 93247.5 ;
      RECT  10107.5 94282.5 10172.5 94657.5 ;
      RECT  10487.5 94282.5 10552.5 94657.5 ;
      RECT  10657.5 94440.0 10722.5 94625.0 ;
      RECT  10657.5 93280.0 10722.5 93465.0 ;
      RECT  10107.5 94282.5 10172.5 94417.5 ;
      RECT  10297.5 94282.5 10362.5 94417.5 ;
      RECT  10297.5 94282.5 10362.5 94417.5 ;
      RECT  10107.5 94282.5 10172.5 94417.5 ;
      RECT  10297.5 94282.5 10362.5 94417.5 ;
      RECT  10487.5 94282.5 10552.5 94417.5 ;
      RECT  10487.5 94282.5 10552.5 94417.5 ;
      RECT  10297.5 94282.5 10362.5 94417.5 ;
      RECT  10107.5 93442.5 10172.5 93577.5 ;
      RECT  10297.5 93442.5 10362.5 93577.5 ;
      RECT  10297.5 93442.5 10362.5 93577.5 ;
      RECT  10107.5 93442.5 10172.5 93577.5 ;
      RECT  10297.5 93442.5 10362.5 93577.5 ;
      RECT  10487.5 93442.5 10552.5 93577.5 ;
      RECT  10487.5 93442.5 10552.5 93577.5 ;
      RECT  10297.5 93442.5 10362.5 93577.5 ;
      RECT  10657.5 94372.5 10722.5 94507.5 ;
      RECT  10657.5 93397.5 10722.5 93532.5 ;
      RECT  10492.5 93672.5 10357.5 93737.5 ;
      RECT  10235.0 93887.5 10100.0 93952.5 ;
      RECT  10297.5 94282.5 10362.5 94417.5 ;
      RECT  10487.5 93442.5 10552.5 93577.5 ;
      RECT  10587.5 93887.5 10452.5 93952.5 ;
      RECT  10100.0 93887.5 10235.0 93952.5 ;
      RECT  10357.5 93672.5 10492.5 93737.5 ;
      RECT  10452.5 93887.5 10587.5 93952.5 ;
      RECT  10040.0 94592.5 10960.0 94657.5 ;
      RECT  10040.0 93247.5 10960.0 93312.5 ;
      RECT  11387.5 94440.0 11452.5 94625.0 ;
      RECT  11387.5 93280.0 11452.5 93465.0 ;
      RECT  11027.5 93397.5 11092.5 93247.5 ;
      RECT  11027.5 94282.5 11092.5 94657.5 ;
      RECT  11217.5 93397.5 11282.5 94282.5 ;
      RECT  11027.5 94282.5 11092.5 94417.5 ;
      RECT  11217.5 94282.5 11282.5 94417.5 ;
      RECT  11217.5 94282.5 11282.5 94417.5 ;
      RECT  11027.5 94282.5 11092.5 94417.5 ;
      RECT  11027.5 93397.5 11092.5 93532.5 ;
      RECT  11217.5 93397.5 11282.5 93532.5 ;
      RECT  11217.5 93397.5 11282.5 93532.5 ;
      RECT  11027.5 93397.5 11092.5 93532.5 ;
      RECT  11387.5 94372.5 11452.5 94507.5 ;
      RECT  11387.5 93397.5 11452.5 93532.5 ;
      RECT  11085.0 93840.0 11150.0 93975.0 ;
      RECT  11085.0 93840.0 11150.0 93975.0 ;
      RECT  11250.0 93875.0 11315.0 93940.0 ;
      RECT  10960.0 94592.5 11520.0 94657.5 ;
      RECT  10960.0 93247.5 11520.0 93312.5 ;
      RECT  9222.5 93840.0 9287.5 93975.0 ;
      RECT  9362.5 93567.5 9427.5 93702.5 ;
      RECT  10357.5 93672.5 10222.5 93737.5 ;
      RECT  9907.5 94810.0 9972.5 94625.0 ;
      RECT  9907.5 95970.0 9972.5 95785.0 ;
      RECT  9547.5 95852.5 9612.5 96002.5 ;
      RECT  9547.5 94967.5 9612.5 94592.5 ;
      RECT  9737.5 95852.5 9802.5 94967.5 ;
      RECT  9547.5 94967.5 9612.5 94832.5 ;
      RECT  9737.5 94967.5 9802.5 94832.5 ;
      RECT  9737.5 94967.5 9802.5 94832.5 ;
      RECT  9547.5 94967.5 9612.5 94832.5 ;
      RECT  9547.5 95852.5 9612.5 95717.5 ;
      RECT  9737.5 95852.5 9802.5 95717.5 ;
      RECT  9737.5 95852.5 9802.5 95717.5 ;
      RECT  9547.5 95852.5 9612.5 95717.5 ;
      RECT  9907.5 94877.5 9972.5 94742.5 ;
      RECT  9907.5 95852.5 9972.5 95717.5 ;
      RECT  9605.0 95410.0 9670.0 95275.0 ;
      RECT  9605.0 95410.0 9670.0 95275.0 ;
      RECT  9770.0 95375.0 9835.0 95310.0 ;
      RECT  9480.0 94657.5 10040.0 94592.5 ;
      RECT  9480.0 96002.5 10040.0 95937.5 ;
      RECT  10107.5 95807.5 10172.5 96002.5 ;
      RECT  10107.5 94967.5 10172.5 94592.5 ;
      RECT  10487.5 94967.5 10552.5 94592.5 ;
      RECT  10657.5 94810.0 10722.5 94625.0 ;
      RECT  10657.5 95970.0 10722.5 95785.0 ;
      RECT  10107.5 94967.5 10172.5 94832.5 ;
      RECT  10297.5 94967.5 10362.5 94832.5 ;
      RECT  10297.5 94967.5 10362.5 94832.5 ;
      RECT  10107.5 94967.5 10172.5 94832.5 ;
      RECT  10297.5 94967.5 10362.5 94832.5 ;
      RECT  10487.5 94967.5 10552.5 94832.5 ;
      RECT  10487.5 94967.5 10552.5 94832.5 ;
      RECT  10297.5 94967.5 10362.5 94832.5 ;
      RECT  10107.5 95807.5 10172.5 95672.5 ;
      RECT  10297.5 95807.5 10362.5 95672.5 ;
      RECT  10297.5 95807.5 10362.5 95672.5 ;
      RECT  10107.5 95807.5 10172.5 95672.5 ;
      RECT  10297.5 95807.5 10362.5 95672.5 ;
      RECT  10487.5 95807.5 10552.5 95672.5 ;
      RECT  10487.5 95807.5 10552.5 95672.5 ;
      RECT  10297.5 95807.5 10362.5 95672.5 ;
      RECT  10657.5 94877.5 10722.5 94742.5 ;
      RECT  10657.5 95852.5 10722.5 95717.5 ;
      RECT  10492.5 95577.5 10357.5 95512.5 ;
      RECT  10235.0 95362.5 10100.0 95297.5 ;
      RECT  10297.5 94967.5 10362.5 94832.5 ;
      RECT  10487.5 95807.5 10552.5 95672.5 ;
      RECT  10587.5 95362.5 10452.5 95297.5 ;
      RECT  10100.0 95362.5 10235.0 95297.5 ;
      RECT  10357.5 95577.5 10492.5 95512.5 ;
      RECT  10452.5 95362.5 10587.5 95297.5 ;
      RECT  10040.0 94657.5 10960.0 94592.5 ;
      RECT  10040.0 96002.5 10960.0 95937.5 ;
      RECT  11387.5 94810.0 11452.5 94625.0 ;
      RECT  11387.5 95970.0 11452.5 95785.0 ;
      RECT  11027.5 95852.5 11092.5 96002.5 ;
      RECT  11027.5 94967.5 11092.5 94592.5 ;
      RECT  11217.5 95852.5 11282.5 94967.5 ;
      RECT  11027.5 94967.5 11092.5 94832.5 ;
      RECT  11217.5 94967.5 11282.5 94832.5 ;
      RECT  11217.5 94967.5 11282.5 94832.5 ;
      RECT  11027.5 94967.5 11092.5 94832.5 ;
      RECT  11027.5 95852.5 11092.5 95717.5 ;
      RECT  11217.5 95852.5 11282.5 95717.5 ;
      RECT  11217.5 95852.5 11282.5 95717.5 ;
      RECT  11027.5 95852.5 11092.5 95717.5 ;
      RECT  11387.5 94877.5 11452.5 94742.5 ;
      RECT  11387.5 95852.5 11452.5 95717.5 ;
      RECT  11085.0 95410.0 11150.0 95275.0 ;
      RECT  11085.0 95410.0 11150.0 95275.0 ;
      RECT  11250.0 95375.0 11315.0 95310.0 ;
      RECT  10960.0 94657.5 11520.0 94592.5 ;
      RECT  10960.0 96002.5 11520.0 95937.5 ;
      RECT  9222.5 95275.0 9287.5 95410.0 ;
      RECT  9362.5 95547.5 9427.5 95682.5 ;
      RECT  10357.5 95512.5 10222.5 95577.5 ;
      RECT  9907.5 97130.0 9972.5 97315.0 ;
      RECT  9907.5 95970.0 9972.5 96155.0 ;
      RECT  9547.5 96087.5 9612.5 95937.5 ;
      RECT  9547.5 96972.5 9612.5 97347.5 ;
      RECT  9737.5 96087.5 9802.5 96972.5 ;
      RECT  9547.5 96972.5 9612.5 97107.5 ;
      RECT  9737.5 96972.5 9802.5 97107.5 ;
      RECT  9737.5 96972.5 9802.5 97107.5 ;
      RECT  9547.5 96972.5 9612.5 97107.5 ;
      RECT  9547.5 96087.5 9612.5 96222.5 ;
      RECT  9737.5 96087.5 9802.5 96222.5 ;
      RECT  9737.5 96087.5 9802.5 96222.5 ;
      RECT  9547.5 96087.5 9612.5 96222.5 ;
      RECT  9907.5 97062.5 9972.5 97197.5 ;
      RECT  9907.5 96087.5 9972.5 96222.5 ;
      RECT  9605.0 96530.0 9670.0 96665.0 ;
      RECT  9605.0 96530.0 9670.0 96665.0 ;
      RECT  9770.0 96565.0 9835.0 96630.0 ;
      RECT  9480.0 97282.5 10040.0 97347.5 ;
      RECT  9480.0 95937.5 10040.0 96002.5 ;
      RECT  10107.5 96132.5 10172.5 95937.5 ;
      RECT  10107.5 96972.5 10172.5 97347.5 ;
      RECT  10487.5 96972.5 10552.5 97347.5 ;
      RECT  10657.5 97130.0 10722.5 97315.0 ;
      RECT  10657.5 95970.0 10722.5 96155.0 ;
      RECT  10107.5 96972.5 10172.5 97107.5 ;
      RECT  10297.5 96972.5 10362.5 97107.5 ;
      RECT  10297.5 96972.5 10362.5 97107.5 ;
      RECT  10107.5 96972.5 10172.5 97107.5 ;
      RECT  10297.5 96972.5 10362.5 97107.5 ;
      RECT  10487.5 96972.5 10552.5 97107.5 ;
      RECT  10487.5 96972.5 10552.5 97107.5 ;
      RECT  10297.5 96972.5 10362.5 97107.5 ;
      RECT  10107.5 96132.5 10172.5 96267.5 ;
      RECT  10297.5 96132.5 10362.5 96267.5 ;
      RECT  10297.5 96132.5 10362.5 96267.5 ;
      RECT  10107.5 96132.5 10172.5 96267.5 ;
      RECT  10297.5 96132.5 10362.5 96267.5 ;
      RECT  10487.5 96132.5 10552.5 96267.5 ;
      RECT  10487.5 96132.5 10552.5 96267.5 ;
      RECT  10297.5 96132.5 10362.5 96267.5 ;
      RECT  10657.5 97062.5 10722.5 97197.5 ;
      RECT  10657.5 96087.5 10722.5 96222.5 ;
      RECT  10492.5 96362.5 10357.5 96427.5 ;
      RECT  10235.0 96577.5 10100.0 96642.5 ;
      RECT  10297.5 96972.5 10362.5 97107.5 ;
      RECT  10487.5 96132.5 10552.5 96267.5 ;
      RECT  10587.5 96577.5 10452.5 96642.5 ;
      RECT  10100.0 96577.5 10235.0 96642.5 ;
      RECT  10357.5 96362.5 10492.5 96427.5 ;
      RECT  10452.5 96577.5 10587.5 96642.5 ;
      RECT  10040.0 97282.5 10960.0 97347.5 ;
      RECT  10040.0 95937.5 10960.0 96002.5 ;
      RECT  11387.5 97130.0 11452.5 97315.0 ;
      RECT  11387.5 95970.0 11452.5 96155.0 ;
      RECT  11027.5 96087.5 11092.5 95937.5 ;
      RECT  11027.5 96972.5 11092.5 97347.5 ;
      RECT  11217.5 96087.5 11282.5 96972.5 ;
      RECT  11027.5 96972.5 11092.5 97107.5 ;
      RECT  11217.5 96972.5 11282.5 97107.5 ;
      RECT  11217.5 96972.5 11282.5 97107.5 ;
      RECT  11027.5 96972.5 11092.5 97107.5 ;
      RECT  11027.5 96087.5 11092.5 96222.5 ;
      RECT  11217.5 96087.5 11282.5 96222.5 ;
      RECT  11217.5 96087.5 11282.5 96222.5 ;
      RECT  11027.5 96087.5 11092.5 96222.5 ;
      RECT  11387.5 97062.5 11452.5 97197.5 ;
      RECT  11387.5 96087.5 11452.5 96222.5 ;
      RECT  11085.0 96530.0 11150.0 96665.0 ;
      RECT  11085.0 96530.0 11150.0 96665.0 ;
      RECT  11250.0 96565.0 11315.0 96630.0 ;
      RECT  10960.0 97282.5 11520.0 97347.5 ;
      RECT  10960.0 95937.5 11520.0 96002.5 ;
      RECT  9222.5 96530.0 9287.5 96665.0 ;
      RECT  9362.5 96257.5 9427.5 96392.5 ;
      RECT  10357.5 96362.5 10222.5 96427.5 ;
      RECT  9907.5 97500.0 9972.5 97315.0 ;
      RECT  9907.5 98660.0 9972.5 98475.0 ;
      RECT  9547.5 98542.5 9612.5 98692.5 ;
      RECT  9547.5 97657.5 9612.5 97282.5 ;
      RECT  9737.5 98542.5 9802.5 97657.5 ;
      RECT  9547.5 97657.5 9612.5 97522.5 ;
      RECT  9737.5 97657.5 9802.5 97522.5 ;
      RECT  9737.5 97657.5 9802.5 97522.5 ;
      RECT  9547.5 97657.5 9612.5 97522.5 ;
      RECT  9547.5 98542.5 9612.5 98407.5 ;
      RECT  9737.5 98542.5 9802.5 98407.5 ;
      RECT  9737.5 98542.5 9802.5 98407.5 ;
      RECT  9547.5 98542.5 9612.5 98407.5 ;
      RECT  9907.5 97567.5 9972.5 97432.5 ;
      RECT  9907.5 98542.5 9972.5 98407.5 ;
      RECT  9605.0 98100.0 9670.0 97965.0 ;
      RECT  9605.0 98100.0 9670.0 97965.0 ;
      RECT  9770.0 98065.0 9835.0 98000.0 ;
      RECT  9480.0 97347.5 10040.0 97282.5 ;
      RECT  9480.0 98692.5 10040.0 98627.5 ;
      RECT  10107.5 98497.5 10172.5 98692.5 ;
      RECT  10107.5 97657.5 10172.5 97282.5 ;
      RECT  10487.5 97657.5 10552.5 97282.5 ;
      RECT  10657.5 97500.0 10722.5 97315.0 ;
      RECT  10657.5 98660.0 10722.5 98475.0 ;
      RECT  10107.5 97657.5 10172.5 97522.5 ;
      RECT  10297.5 97657.5 10362.5 97522.5 ;
      RECT  10297.5 97657.5 10362.5 97522.5 ;
      RECT  10107.5 97657.5 10172.5 97522.5 ;
      RECT  10297.5 97657.5 10362.5 97522.5 ;
      RECT  10487.5 97657.5 10552.5 97522.5 ;
      RECT  10487.5 97657.5 10552.5 97522.5 ;
      RECT  10297.5 97657.5 10362.5 97522.5 ;
      RECT  10107.5 98497.5 10172.5 98362.5 ;
      RECT  10297.5 98497.5 10362.5 98362.5 ;
      RECT  10297.5 98497.5 10362.5 98362.5 ;
      RECT  10107.5 98497.5 10172.5 98362.5 ;
      RECT  10297.5 98497.5 10362.5 98362.5 ;
      RECT  10487.5 98497.5 10552.5 98362.5 ;
      RECT  10487.5 98497.5 10552.5 98362.5 ;
      RECT  10297.5 98497.5 10362.5 98362.5 ;
      RECT  10657.5 97567.5 10722.5 97432.5 ;
      RECT  10657.5 98542.5 10722.5 98407.5 ;
      RECT  10492.5 98267.5 10357.5 98202.5 ;
      RECT  10235.0 98052.5 10100.0 97987.5 ;
      RECT  10297.5 97657.5 10362.5 97522.5 ;
      RECT  10487.5 98497.5 10552.5 98362.5 ;
      RECT  10587.5 98052.5 10452.5 97987.5 ;
      RECT  10100.0 98052.5 10235.0 97987.5 ;
      RECT  10357.5 98267.5 10492.5 98202.5 ;
      RECT  10452.5 98052.5 10587.5 97987.5 ;
      RECT  10040.0 97347.5 10960.0 97282.5 ;
      RECT  10040.0 98692.5 10960.0 98627.5 ;
      RECT  11387.5 97500.0 11452.5 97315.0 ;
      RECT  11387.5 98660.0 11452.5 98475.0 ;
      RECT  11027.5 98542.5 11092.5 98692.5 ;
      RECT  11027.5 97657.5 11092.5 97282.5 ;
      RECT  11217.5 98542.5 11282.5 97657.5 ;
      RECT  11027.5 97657.5 11092.5 97522.5 ;
      RECT  11217.5 97657.5 11282.5 97522.5 ;
      RECT  11217.5 97657.5 11282.5 97522.5 ;
      RECT  11027.5 97657.5 11092.5 97522.5 ;
      RECT  11027.5 98542.5 11092.5 98407.5 ;
      RECT  11217.5 98542.5 11282.5 98407.5 ;
      RECT  11217.5 98542.5 11282.5 98407.5 ;
      RECT  11027.5 98542.5 11092.5 98407.5 ;
      RECT  11387.5 97567.5 11452.5 97432.5 ;
      RECT  11387.5 98542.5 11452.5 98407.5 ;
      RECT  11085.0 98100.0 11150.0 97965.0 ;
      RECT  11085.0 98100.0 11150.0 97965.0 ;
      RECT  11250.0 98065.0 11315.0 98000.0 ;
      RECT  10960.0 97347.5 11520.0 97282.5 ;
      RECT  10960.0 98692.5 11520.0 98627.5 ;
      RECT  9222.5 97965.0 9287.5 98100.0 ;
      RECT  9362.5 98237.5 9427.5 98372.5 ;
      RECT  10357.5 98202.5 10222.5 98267.5 ;
      RECT  9907.5 99820.0 9972.5 100005.0 ;
      RECT  9907.5 98660.0 9972.5 98845.0 ;
      RECT  9547.5 98777.5 9612.5 98627.5 ;
      RECT  9547.5 99662.5 9612.5 100037.5 ;
      RECT  9737.5 98777.5 9802.5 99662.5 ;
      RECT  9547.5 99662.5 9612.5 99797.5 ;
      RECT  9737.5 99662.5 9802.5 99797.5 ;
      RECT  9737.5 99662.5 9802.5 99797.5 ;
      RECT  9547.5 99662.5 9612.5 99797.5 ;
      RECT  9547.5 98777.5 9612.5 98912.5 ;
      RECT  9737.5 98777.5 9802.5 98912.5 ;
      RECT  9737.5 98777.5 9802.5 98912.5 ;
      RECT  9547.5 98777.5 9612.5 98912.5 ;
      RECT  9907.5 99752.5 9972.5 99887.5 ;
      RECT  9907.5 98777.5 9972.5 98912.5 ;
      RECT  9605.0 99220.0 9670.0 99355.0 ;
      RECT  9605.0 99220.0 9670.0 99355.0 ;
      RECT  9770.0 99255.0 9835.0 99320.0 ;
      RECT  9480.0 99972.5 10040.0 100037.5 ;
      RECT  9480.0 98627.5 10040.0 98692.5 ;
      RECT  10107.5 98822.5 10172.5 98627.5 ;
      RECT  10107.5 99662.5 10172.5 100037.5 ;
      RECT  10487.5 99662.5 10552.5 100037.5 ;
      RECT  10657.5 99820.0 10722.5 100005.0 ;
      RECT  10657.5 98660.0 10722.5 98845.0 ;
      RECT  10107.5 99662.5 10172.5 99797.5 ;
      RECT  10297.5 99662.5 10362.5 99797.5 ;
      RECT  10297.5 99662.5 10362.5 99797.5 ;
      RECT  10107.5 99662.5 10172.5 99797.5 ;
      RECT  10297.5 99662.5 10362.5 99797.5 ;
      RECT  10487.5 99662.5 10552.5 99797.5 ;
      RECT  10487.5 99662.5 10552.5 99797.5 ;
      RECT  10297.5 99662.5 10362.5 99797.5 ;
      RECT  10107.5 98822.5 10172.5 98957.5 ;
      RECT  10297.5 98822.5 10362.5 98957.5 ;
      RECT  10297.5 98822.5 10362.5 98957.5 ;
      RECT  10107.5 98822.5 10172.5 98957.5 ;
      RECT  10297.5 98822.5 10362.5 98957.5 ;
      RECT  10487.5 98822.5 10552.5 98957.5 ;
      RECT  10487.5 98822.5 10552.5 98957.5 ;
      RECT  10297.5 98822.5 10362.5 98957.5 ;
      RECT  10657.5 99752.5 10722.5 99887.5 ;
      RECT  10657.5 98777.5 10722.5 98912.5 ;
      RECT  10492.5 99052.5 10357.5 99117.5 ;
      RECT  10235.0 99267.5 10100.0 99332.5 ;
      RECT  10297.5 99662.5 10362.5 99797.5 ;
      RECT  10487.5 98822.5 10552.5 98957.5 ;
      RECT  10587.5 99267.5 10452.5 99332.5 ;
      RECT  10100.0 99267.5 10235.0 99332.5 ;
      RECT  10357.5 99052.5 10492.5 99117.5 ;
      RECT  10452.5 99267.5 10587.5 99332.5 ;
      RECT  10040.0 99972.5 10960.0 100037.5 ;
      RECT  10040.0 98627.5 10960.0 98692.5 ;
      RECT  11387.5 99820.0 11452.5 100005.0 ;
      RECT  11387.5 98660.0 11452.5 98845.0 ;
      RECT  11027.5 98777.5 11092.5 98627.5 ;
      RECT  11027.5 99662.5 11092.5 100037.5 ;
      RECT  11217.5 98777.5 11282.5 99662.5 ;
      RECT  11027.5 99662.5 11092.5 99797.5 ;
      RECT  11217.5 99662.5 11282.5 99797.5 ;
      RECT  11217.5 99662.5 11282.5 99797.5 ;
      RECT  11027.5 99662.5 11092.5 99797.5 ;
      RECT  11027.5 98777.5 11092.5 98912.5 ;
      RECT  11217.5 98777.5 11282.5 98912.5 ;
      RECT  11217.5 98777.5 11282.5 98912.5 ;
      RECT  11027.5 98777.5 11092.5 98912.5 ;
      RECT  11387.5 99752.5 11452.5 99887.5 ;
      RECT  11387.5 98777.5 11452.5 98912.5 ;
      RECT  11085.0 99220.0 11150.0 99355.0 ;
      RECT  11085.0 99220.0 11150.0 99355.0 ;
      RECT  11250.0 99255.0 11315.0 99320.0 ;
      RECT  10960.0 99972.5 11520.0 100037.5 ;
      RECT  10960.0 98627.5 11520.0 98692.5 ;
      RECT  9222.5 99220.0 9287.5 99355.0 ;
      RECT  9362.5 98947.5 9427.5 99082.5 ;
      RECT  10357.5 99052.5 10222.5 99117.5 ;
      RECT  9907.5 100190.0 9972.5 100005.0 ;
      RECT  9907.5 101350.0 9972.5 101165.0 ;
      RECT  9547.5 101232.5 9612.5 101382.5 ;
      RECT  9547.5 100347.5 9612.5 99972.5 ;
      RECT  9737.5 101232.5 9802.5 100347.5 ;
      RECT  9547.5 100347.5 9612.5 100212.5 ;
      RECT  9737.5 100347.5 9802.5 100212.5 ;
      RECT  9737.5 100347.5 9802.5 100212.5 ;
      RECT  9547.5 100347.5 9612.5 100212.5 ;
      RECT  9547.5 101232.5 9612.5 101097.5 ;
      RECT  9737.5 101232.5 9802.5 101097.5 ;
      RECT  9737.5 101232.5 9802.5 101097.5 ;
      RECT  9547.5 101232.5 9612.5 101097.5 ;
      RECT  9907.5 100257.5 9972.5 100122.5 ;
      RECT  9907.5 101232.5 9972.5 101097.5 ;
      RECT  9605.0 100790.0 9670.0 100655.0 ;
      RECT  9605.0 100790.0 9670.0 100655.0 ;
      RECT  9770.0 100755.0 9835.0 100690.0 ;
      RECT  9480.0 100037.5 10040.0 99972.5 ;
      RECT  9480.0 101382.5 10040.0 101317.5 ;
      RECT  10107.5 101187.5 10172.5 101382.5 ;
      RECT  10107.5 100347.5 10172.5 99972.5 ;
      RECT  10487.5 100347.5 10552.5 99972.5 ;
      RECT  10657.5 100190.0 10722.5 100005.0 ;
      RECT  10657.5 101350.0 10722.5 101165.0 ;
      RECT  10107.5 100347.5 10172.5 100212.5 ;
      RECT  10297.5 100347.5 10362.5 100212.5 ;
      RECT  10297.5 100347.5 10362.5 100212.5 ;
      RECT  10107.5 100347.5 10172.5 100212.5 ;
      RECT  10297.5 100347.5 10362.5 100212.5 ;
      RECT  10487.5 100347.5 10552.5 100212.5 ;
      RECT  10487.5 100347.5 10552.5 100212.5 ;
      RECT  10297.5 100347.5 10362.5 100212.5 ;
      RECT  10107.5 101187.5 10172.5 101052.5 ;
      RECT  10297.5 101187.5 10362.5 101052.5 ;
      RECT  10297.5 101187.5 10362.5 101052.5 ;
      RECT  10107.5 101187.5 10172.5 101052.5 ;
      RECT  10297.5 101187.5 10362.5 101052.5 ;
      RECT  10487.5 101187.5 10552.5 101052.5 ;
      RECT  10487.5 101187.5 10552.5 101052.5 ;
      RECT  10297.5 101187.5 10362.5 101052.5 ;
      RECT  10657.5 100257.5 10722.5 100122.5 ;
      RECT  10657.5 101232.5 10722.5 101097.5 ;
      RECT  10492.5 100957.5 10357.5 100892.5 ;
      RECT  10235.0 100742.5 10100.0 100677.5 ;
      RECT  10297.5 100347.5 10362.5 100212.5 ;
      RECT  10487.5 101187.5 10552.5 101052.5 ;
      RECT  10587.5 100742.5 10452.5 100677.5 ;
      RECT  10100.0 100742.5 10235.0 100677.5 ;
      RECT  10357.5 100957.5 10492.5 100892.5 ;
      RECT  10452.5 100742.5 10587.5 100677.5 ;
      RECT  10040.0 100037.5 10960.0 99972.5 ;
      RECT  10040.0 101382.5 10960.0 101317.5 ;
      RECT  11387.5 100190.0 11452.5 100005.0 ;
      RECT  11387.5 101350.0 11452.5 101165.0 ;
      RECT  11027.5 101232.5 11092.5 101382.5 ;
      RECT  11027.5 100347.5 11092.5 99972.5 ;
      RECT  11217.5 101232.5 11282.5 100347.5 ;
      RECT  11027.5 100347.5 11092.5 100212.5 ;
      RECT  11217.5 100347.5 11282.5 100212.5 ;
      RECT  11217.5 100347.5 11282.5 100212.5 ;
      RECT  11027.5 100347.5 11092.5 100212.5 ;
      RECT  11027.5 101232.5 11092.5 101097.5 ;
      RECT  11217.5 101232.5 11282.5 101097.5 ;
      RECT  11217.5 101232.5 11282.5 101097.5 ;
      RECT  11027.5 101232.5 11092.5 101097.5 ;
      RECT  11387.5 100257.5 11452.5 100122.5 ;
      RECT  11387.5 101232.5 11452.5 101097.5 ;
      RECT  11085.0 100790.0 11150.0 100655.0 ;
      RECT  11085.0 100790.0 11150.0 100655.0 ;
      RECT  11250.0 100755.0 11315.0 100690.0 ;
      RECT  10960.0 100037.5 11520.0 99972.5 ;
      RECT  10960.0 101382.5 11520.0 101317.5 ;
      RECT  9222.5 100655.0 9287.5 100790.0 ;
      RECT  9362.5 100927.5 9427.5 101062.5 ;
      RECT  10357.5 100892.5 10222.5 100957.5 ;
      RECT  9907.5 102510.0 9972.5 102695.0 ;
      RECT  9907.5 101350.0 9972.5 101535.0 ;
      RECT  9547.5 101467.5 9612.5 101317.5 ;
      RECT  9547.5 102352.5 9612.5 102727.5 ;
      RECT  9737.5 101467.5 9802.5 102352.5 ;
      RECT  9547.5 102352.5 9612.5 102487.5 ;
      RECT  9737.5 102352.5 9802.5 102487.5 ;
      RECT  9737.5 102352.5 9802.5 102487.5 ;
      RECT  9547.5 102352.5 9612.5 102487.5 ;
      RECT  9547.5 101467.5 9612.5 101602.5 ;
      RECT  9737.5 101467.5 9802.5 101602.5 ;
      RECT  9737.5 101467.5 9802.5 101602.5 ;
      RECT  9547.5 101467.5 9612.5 101602.5 ;
      RECT  9907.5 102442.5 9972.5 102577.5 ;
      RECT  9907.5 101467.5 9972.5 101602.5 ;
      RECT  9605.0 101910.0 9670.0 102045.0 ;
      RECT  9605.0 101910.0 9670.0 102045.0 ;
      RECT  9770.0 101945.0 9835.0 102010.0 ;
      RECT  9480.0 102662.5 10040.0 102727.5 ;
      RECT  9480.0 101317.5 10040.0 101382.5 ;
      RECT  10107.5 101512.5 10172.5 101317.5 ;
      RECT  10107.5 102352.5 10172.5 102727.5 ;
      RECT  10487.5 102352.5 10552.5 102727.5 ;
      RECT  10657.5 102510.0 10722.5 102695.0 ;
      RECT  10657.5 101350.0 10722.5 101535.0 ;
      RECT  10107.5 102352.5 10172.5 102487.5 ;
      RECT  10297.5 102352.5 10362.5 102487.5 ;
      RECT  10297.5 102352.5 10362.5 102487.5 ;
      RECT  10107.5 102352.5 10172.5 102487.5 ;
      RECT  10297.5 102352.5 10362.5 102487.5 ;
      RECT  10487.5 102352.5 10552.5 102487.5 ;
      RECT  10487.5 102352.5 10552.5 102487.5 ;
      RECT  10297.5 102352.5 10362.5 102487.5 ;
      RECT  10107.5 101512.5 10172.5 101647.5 ;
      RECT  10297.5 101512.5 10362.5 101647.5 ;
      RECT  10297.5 101512.5 10362.5 101647.5 ;
      RECT  10107.5 101512.5 10172.5 101647.5 ;
      RECT  10297.5 101512.5 10362.5 101647.5 ;
      RECT  10487.5 101512.5 10552.5 101647.5 ;
      RECT  10487.5 101512.5 10552.5 101647.5 ;
      RECT  10297.5 101512.5 10362.5 101647.5 ;
      RECT  10657.5 102442.5 10722.5 102577.5 ;
      RECT  10657.5 101467.5 10722.5 101602.5 ;
      RECT  10492.5 101742.5 10357.5 101807.5 ;
      RECT  10235.0 101957.5 10100.0 102022.5 ;
      RECT  10297.5 102352.5 10362.5 102487.5 ;
      RECT  10487.5 101512.5 10552.5 101647.5 ;
      RECT  10587.5 101957.5 10452.5 102022.5 ;
      RECT  10100.0 101957.5 10235.0 102022.5 ;
      RECT  10357.5 101742.5 10492.5 101807.5 ;
      RECT  10452.5 101957.5 10587.5 102022.5 ;
      RECT  10040.0 102662.5 10960.0 102727.5 ;
      RECT  10040.0 101317.5 10960.0 101382.5 ;
      RECT  11387.5 102510.0 11452.5 102695.0 ;
      RECT  11387.5 101350.0 11452.5 101535.0 ;
      RECT  11027.5 101467.5 11092.5 101317.5 ;
      RECT  11027.5 102352.5 11092.5 102727.5 ;
      RECT  11217.5 101467.5 11282.5 102352.5 ;
      RECT  11027.5 102352.5 11092.5 102487.5 ;
      RECT  11217.5 102352.5 11282.5 102487.5 ;
      RECT  11217.5 102352.5 11282.5 102487.5 ;
      RECT  11027.5 102352.5 11092.5 102487.5 ;
      RECT  11027.5 101467.5 11092.5 101602.5 ;
      RECT  11217.5 101467.5 11282.5 101602.5 ;
      RECT  11217.5 101467.5 11282.5 101602.5 ;
      RECT  11027.5 101467.5 11092.5 101602.5 ;
      RECT  11387.5 102442.5 11452.5 102577.5 ;
      RECT  11387.5 101467.5 11452.5 101602.5 ;
      RECT  11085.0 101910.0 11150.0 102045.0 ;
      RECT  11085.0 101910.0 11150.0 102045.0 ;
      RECT  11250.0 101945.0 11315.0 102010.0 ;
      RECT  10960.0 102662.5 11520.0 102727.5 ;
      RECT  10960.0 101317.5 11520.0 101382.5 ;
      RECT  9222.5 101910.0 9287.5 102045.0 ;
      RECT  9362.5 101637.5 9427.5 101772.5 ;
      RECT  10357.5 101742.5 10222.5 101807.5 ;
      RECT  9907.5 102880.0 9972.5 102695.0 ;
      RECT  9907.5 104040.0 9972.5 103855.0 ;
      RECT  9547.5 103922.5 9612.5 104072.5 ;
      RECT  9547.5 103037.5 9612.5 102662.5 ;
      RECT  9737.5 103922.5 9802.5 103037.5 ;
      RECT  9547.5 103037.5 9612.5 102902.5 ;
      RECT  9737.5 103037.5 9802.5 102902.5 ;
      RECT  9737.5 103037.5 9802.5 102902.5 ;
      RECT  9547.5 103037.5 9612.5 102902.5 ;
      RECT  9547.5 103922.5 9612.5 103787.5 ;
      RECT  9737.5 103922.5 9802.5 103787.5 ;
      RECT  9737.5 103922.5 9802.5 103787.5 ;
      RECT  9547.5 103922.5 9612.5 103787.5 ;
      RECT  9907.5 102947.5 9972.5 102812.5 ;
      RECT  9907.5 103922.5 9972.5 103787.5 ;
      RECT  9605.0 103480.0 9670.0 103345.0 ;
      RECT  9605.0 103480.0 9670.0 103345.0 ;
      RECT  9770.0 103445.0 9835.0 103380.0 ;
      RECT  9480.0 102727.5 10040.0 102662.5 ;
      RECT  9480.0 104072.5 10040.0 104007.5 ;
      RECT  10107.5 103877.5 10172.5 104072.5 ;
      RECT  10107.5 103037.5 10172.5 102662.5 ;
      RECT  10487.5 103037.5 10552.5 102662.5 ;
      RECT  10657.5 102880.0 10722.5 102695.0 ;
      RECT  10657.5 104040.0 10722.5 103855.0 ;
      RECT  10107.5 103037.5 10172.5 102902.5 ;
      RECT  10297.5 103037.5 10362.5 102902.5 ;
      RECT  10297.5 103037.5 10362.5 102902.5 ;
      RECT  10107.5 103037.5 10172.5 102902.5 ;
      RECT  10297.5 103037.5 10362.5 102902.5 ;
      RECT  10487.5 103037.5 10552.5 102902.5 ;
      RECT  10487.5 103037.5 10552.5 102902.5 ;
      RECT  10297.5 103037.5 10362.5 102902.5 ;
      RECT  10107.5 103877.5 10172.5 103742.5 ;
      RECT  10297.5 103877.5 10362.5 103742.5 ;
      RECT  10297.5 103877.5 10362.5 103742.5 ;
      RECT  10107.5 103877.5 10172.5 103742.5 ;
      RECT  10297.5 103877.5 10362.5 103742.5 ;
      RECT  10487.5 103877.5 10552.5 103742.5 ;
      RECT  10487.5 103877.5 10552.5 103742.5 ;
      RECT  10297.5 103877.5 10362.5 103742.5 ;
      RECT  10657.5 102947.5 10722.5 102812.5 ;
      RECT  10657.5 103922.5 10722.5 103787.5 ;
      RECT  10492.5 103647.5 10357.5 103582.5 ;
      RECT  10235.0 103432.5 10100.0 103367.5 ;
      RECT  10297.5 103037.5 10362.5 102902.5 ;
      RECT  10487.5 103877.5 10552.5 103742.5 ;
      RECT  10587.5 103432.5 10452.5 103367.5 ;
      RECT  10100.0 103432.5 10235.0 103367.5 ;
      RECT  10357.5 103647.5 10492.5 103582.5 ;
      RECT  10452.5 103432.5 10587.5 103367.5 ;
      RECT  10040.0 102727.5 10960.0 102662.5 ;
      RECT  10040.0 104072.5 10960.0 104007.5 ;
      RECT  11387.5 102880.0 11452.5 102695.0 ;
      RECT  11387.5 104040.0 11452.5 103855.0 ;
      RECT  11027.5 103922.5 11092.5 104072.5 ;
      RECT  11027.5 103037.5 11092.5 102662.5 ;
      RECT  11217.5 103922.5 11282.5 103037.5 ;
      RECT  11027.5 103037.5 11092.5 102902.5 ;
      RECT  11217.5 103037.5 11282.5 102902.5 ;
      RECT  11217.5 103037.5 11282.5 102902.5 ;
      RECT  11027.5 103037.5 11092.5 102902.5 ;
      RECT  11027.5 103922.5 11092.5 103787.5 ;
      RECT  11217.5 103922.5 11282.5 103787.5 ;
      RECT  11217.5 103922.5 11282.5 103787.5 ;
      RECT  11027.5 103922.5 11092.5 103787.5 ;
      RECT  11387.5 102947.5 11452.5 102812.5 ;
      RECT  11387.5 103922.5 11452.5 103787.5 ;
      RECT  11085.0 103480.0 11150.0 103345.0 ;
      RECT  11085.0 103480.0 11150.0 103345.0 ;
      RECT  11250.0 103445.0 11315.0 103380.0 ;
      RECT  10960.0 102727.5 11520.0 102662.5 ;
      RECT  10960.0 104072.5 11520.0 104007.5 ;
      RECT  9222.5 103345.0 9287.5 103480.0 ;
      RECT  9362.5 103617.5 9427.5 103752.5 ;
      RECT  10357.5 103582.5 10222.5 103647.5 ;
      RECT  9907.5 105200.0 9972.5 105385.0 ;
      RECT  9907.5 104040.0 9972.5 104225.0 ;
      RECT  9547.5 104157.5 9612.5 104007.5 ;
      RECT  9547.5 105042.5 9612.5 105417.5 ;
      RECT  9737.5 104157.5 9802.5 105042.5 ;
      RECT  9547.5 105042.5 9612.5 105177.5 ;
      RECT  9737.5 105042.5 9802.5 105177.5 ;
      RECT  9737.5 105042.5 9802.5 105177.5 ;
      RECT  9547.5 105042.5 9612.5 105177.5 ;
      RECT  9547.5 104157.5 9612.5 104292.5 ;
      RECT  9737.5 104157.5 9802.5 104292.5 ;
      RECT  9737.5 104157.5 9802.5 104292.5 ;
      RECT  9547.5 104157.5 9612.5 104292.5 ;
      RECT  9907.5 105132.5 9972.5 105267.5 ;
      RECT  9907.5 104157.5 9972.5 104292.5 ;
      RECT  9605.0 104600.0 9670.0 104735.0 ;
      RECT  9605.0 104600.0 9670.0 104735.0 ;
      RECT  9770.0 104635.0 9835.0 104700.0 ;
      RECT  9480.0 105352.5 10040.0 105417.5 ;
      RECT  9480.0 104007.5 10040.0 104072.5 ;
      RECT  10107.5 104202.5 10172.5 104007.5 ;
      RECT  10107.5 105042.5 10172.5 105417.5 ;
      RECT  10487.5 105042.5 10552.5 105417.5 ;
      RECT  10657.5 105200.0 10722.5 105385.0 ;
      RECT  10657.5 104040.0 10722.5 104225.0 ;
      RECT  10107.5 105042.5 10172.5 105177.5 ;
      RECT  10297.5 105042.5 10362.5 105177.5 ;
      RECT  10297.5 105042.5 10362.5 105177.5 ;
      RECT  10107.5 105042.5 10172.5 105177.5 ;
      RECT  10297.5 105042.5 10362.5 105177.5 ;
      RECT  10487.5 105042.5 10552.5 105177.5 ;
      RECT  10487.5 105042.5 10552.5 105177.5 ;
      RECT  10297.5 105042.5 10362.5 105177.5 ;
      RECT  10107.5 104202.5 10172.5 104337.5 ;
      RECT  10297.5 104202.5 10362.5 104337.5 ;
      RECT  10297.5 104202.5 10362.5 104337.5 ;
      RECT  10107.5 104202.5 10172.5 104337.5 ;
      RECT  10297.5 104202.5 10362.5 104337.5 ;
      RECT  10487.5 104202.5 10552.5 104337.5 ;
      RECT  10487.5 104202.5 10552.5 104337.5 ;
      RECT  10297.5 104202.5 10362.5 104337.5 ;
      RECT  10657.5 105132.5 10722.5 105267.5 ;
      RECT  10657.5 104157.5 10722.5 104292.5 ;
      RECT  10492.5 104432.5 10357.5 104497.5 ;
      RECT  10235.0 104647.5 10100.0 104712.5 ;
      RECT  10297.5 105042.5 10362.5 105177.5 ;
      RECT  10487.5 104202.5 10552.5 104337.5 ;
      RECT  10587.5 104647.5 10452.5 104712.5 ;
      RECT  10100.0 104647.5 10235.0 104712.5 ;
      RECT  10357.5 104432.5 10492.5 104497.5 ;
      RECT  10452.5 104647.5 10587.5 104712.5 ;
      RECT  10040.0 105352.5 10960.0 105417.5 ;
      RECT  10040.0 104007.5 10960.0 104072.5 ;
      RECT  11387.5 105200.0 11452.5 105385.0 ;
      RECT  11387.5 104040.0 11452.5 104225.0 ;
      RECT  11027.5 104157.5 11092.5 104007.5 ;
      RECT  11027.5 105042.5 11092.5 105417.5 ;
      RECT  11217.5 104157.5 11282.5 105042.5 ;
      RECT  11027.5 105042.5 11092.5 105177.5 ;
      RECT  11217.5 105042.5 11282.5 105177.5 ;
      RECT  11217.5 105042.5 11282.5 105177.5 ;
      RECT  11027.5 105042.5 11092.5 105177.5 ;
      RECT  11027.5 104157.5 11092.5 104292.5 ;
      RECT  11217.5 104157.5 11282.5 104292.5 ;
      RECT  11217.5 104157.5 11282.5 104292.5 ;
      RECT  11027.5 104157.5 11092.5 104292.5 ;
      RECT  11387.5 105132.5 11452.5 105267.5 ;
      RECT  11387.5 104157.5 11452.5 104292.5 ;
      RECT  11085.0 104600.0 11150.0 104735.0 ;
      RECT  11085.0 104600.0 11150.0 104735.0 ;
      RECT  11250.0 104635.0 11315.0 104700.0 ;
      RECT  10960.0 105352.5 11520.0 105417.5 ;
      RECT  10960.0 104007.5 11520.0 104072.5 ;
      RECT  9222.5 104600.0 9287.5 104735.0 ;
      RECT  9362.5 104327.5 9427.5 104462.5 ;
      RECT  10357.5 104432.5 10222.5 104497.5 ;
      RECT  9907.5 105570.0 9972.5 105385.0 ;
      RECT  9907.5 106730.0 9972.5 106545.0 ;
      RECT  9547.5 106612.5 9612.5 106762.5 ;
      RECT  9547.5 105727.5 9612.5 105352.5 ;
      RECT  9737.5 106612.5 9802.5 105727.5 ;
      RECT  9547.5 105727.5 9612.5 105592.5 ;
      RECT  9737.5 105727.5 9802.5 105592.5 ;
      RECT  9737.5 105727.5 9802.5 105592.5 ;
      RECT  9547.5 105727.5 9612.5 105592.5 ;
      RECT  9547.5 106612.5 9612.5 106477.5 ;
      RECT  9737.5 106612.5 9802.5 106477.5 ;
      RECT  9737.5 106612.5 9802.5 106477.5 ;
      RECT  9547.5 106612.5 9612.5 106477.5 ;
      RECT  9907.5 105637.5 9972.5 105502.5 ;
      RECT  9907.5 106612.5 9972.5 106477.5 ;
      RECT  9605.0 106170.0 9670.0 106035.0 ;
      RECT  9605.0 106170.0 9670.0 106035.0 ;
      RECT  9770.0 106135.0 9835.0 106070.0 ;
      RECT  9480.0 105417.5 10040.0 105352.5 ;
      RECT  9480.0 106762.5 10040.0 106697.5 ;
      RECT  10107.5 106567.5 10172.5 106762.5 ;
      RECT  10107.5 105727.5 10172.5 105352.5 ;
      RECT  10487.5 105727.5 10552.5 105352.5 ;
      RECT  10657.5 105570.0 10722.5 105385.0 ;
      RECT  10657.5 106730.0 10722.5 106545.0 ;
      RECT  10107.5 105727.5 10172.5 105592.5 ;
      RECT  10297.5 105727.5 10362.5 105592.5 ;
      RECT  10297.5 105727.5 10362.5 105592.5 ;
      RECT  10107.5 105727.5 10172.5 105592.5 ;
      RECT  10297.5 105727.5 10362.5 105592.5 ;
      RECT  10487.5 105727.5 10552.5 105592.5 ;
      RECT  10487.5 105727.5 10552.5 105592.5 ;
      RECT  10297.5 105727.5 10362.5 105592.5 ;
      RECT  10107.5 106567.5 10172.5 106432.5 ;
      RECT  10297.5 106567.5 10362.5 106432.5 ;
      RECT  10297.5 106567.5 10362.5 106432.5 ;
      RECT  10107.5 106567.5 10172.5 106432.5 ;
      RECT  10297.5 106567.5 10362.5 106432.5 ;
      RECT  10487.5 106567.5 10552.5 106432.5 ;
      RECT  10487.5 106567.5 10552.5 106432.5 ;
      RECT  10297.5 106567.5 10362.5 106432.5 ;
      RECT  10657.5 105637.5 10722.5 105502.5 ;
      RECT  10657.5 106612.5 10722.5 106477.5 ;
      RECT  10492.5 106337.5 10357.5 106272.5 ;
      RECT  10235.0 106122.5 10100.0 106057.5 ;
      RECT  10297.5 105727.5 10362.5 105592.5 ;
      RECT  10487.5 106567.5 10552.5 106432.5 ;
      RECT  10587.5 106122.5 10452.5 106057.5 ;
      RECT  10100.0 106122.5 10235.0 106057.5 ;
      RECT  10357.5 106337.5 10492.5 106272.5 ;
      RECT  10452.5 106122.5 10587.5 106057.5 ;
      RECT  10040.0 105417.5 10960.0 105352.5 ;
      RECT  10040.0 106762.5 10960.0 106697.5 ;
      RECT  11387.5 105570.0 11452.5 105385.0 ;
      RECT  11387.5 106730.0 11452.5 106545.0 ;
      RECT  11027.5 106612.5 11092.5 106762.5 ;
      RECT  11027.5 105727.5 11092.5 105352.5 ;
      RECT  11217.5 106612.5 11282.5 105727.5 ;
      RECT  11027.5 105727.5 11092.5 105592.5 ;
      RECT  11217.5 105727.5 11282.5 105592.5 ;
      RECT  11217.5 105727.5 11282.5 105592.5 ;
      RECT  11027.5 105727.5 11092.5 105592.5 ;
      RECT  11027.5 106612.5 11092.5 106477.5 ;
      RECT  11217.5 106612.5 11282.5 106477.5 ;
      RECT  11217.5 106612.5 11282.5 106477.5 ;
      RECT  11027.5 106612.5 11092.5 106477.5 ;
      RECT  11387.5 105637.5 11452.5 105502.5 ;
      RECT  11387.5 106612.5 11452.5 106477.5 ;
      RECT  11085.0 106170.0 11150.0 106035.0 ;
      RECT  11085.0 106170.0 11150.0 106035.0 ;
      RECT  11250.0 106135.0 11315.0 106070.0 ;
      RECT  10960.0 105417.5 11520.0 105352.5 ;
      RECT  10960.0 106762.5 11520.0 106697.5 ;
      RECT  9222.5 106035.0 9287.5 106170.0 ;
      RECT  9362.5 106307.5 9427.5 106442.5 ;
      RECT  10357.5 106272.5 10222.5 106337.5 ;
      RECT  9907.5 107890.0 9972.5 108075.0 ;
      RECT  9907.5 106730.0 9972.5 106915.0 ;
      RECT  9547.5 106847.5 9612.5 106697.5 ;
      RECT  9547.5 107732.5 9612.5 108107.5 ;
      RECT  9737.5 106847.5 9802.5 107732.5 ;
      RECT  9547.5 107732.5 9612.5 107867.5 ;
      RECT  9737.5 107732.5 9802.5 107867.5 ;
      RECT  9737.5 107732.5 9802.5 107867.5 ;
      RECT  9547.5 107732.5 9612.5 107867.5 ;
      RECT  9547.5 106847.5 9612.5 106982.5 ;
      RECT  9737.5 106847.5 9802.5 106982.5 ;
      RECT  9737.5 106847.5 9802.5 106982.5 ;
      RECT  9547.5 106847.5 9612.5 106982.5 ;
      RECT  9907.5 107822.5 9972.5 107957.5 ;
      RECT  9907.5 106847.5 9972.5 106982.5 ;
      RECT  9605.0 107290.0 9670.0 107425.0 ;
      RECT  9605.0 107290.0 9670.0 107425.0 ;
      RECT  9770.0 107325.0 9835.0 107390.0 ;
      RECT  9480.0 108042.5 10040.0 108107.5 ;
      RECT  9480.0 106697.5 10040.0 106762.5 ;
      RECT  10107.5 106892.5 10172.5 106697.5 ;
      RECT  10107.5 107732.5 10172.5 108107.5 ;
      RECT  10487.5 107732.5 10552.5 108107.5 ;
      RECT  10657.5 107890.0 10722.5 108075.0 ;
      RECT  10657.5 106730.0 10722.5 106915.0 ;
      RECT  10107.5 107732.5 10172.5 107867.5 ;
      RECT  10297.5 107732.5 10362.5 107867.5 ;
      RECT  10297.5 107732.5 10362.5 107867.5 ;
      RECT  10107.5 107732.5 10172.5 107867.5 ;
      RECT  10297.5 107732.5 10362.5 107867.5 ;
      RECT  10487.5 107732.5 10552.5 107867.5 ;
      RECT  10487.5 107732.5 10552.5 107867.5 ;
      RECT  10297.5 107732.5 10362.5 107867.5 ;
      RECT  10107.5 106892.5 10172.5 107027.5 ;
      RECT  10297.5 106892.5 10362.5 107027.5 ;
      RECT  10297.5 106892.5 10362.5 107027.5 ;
      RECT  10107.5 106892.5 10172.5 107027.5 ;
      RECT  10297.5 106892.5 10362.5 107027.5 ;
      RECT  10487.5 106892.5 10552.5 107027.5 ;
      RECT  10487.5 106892.5 10552.5 107027.5 ;
      RECT  10297.5 106892.5 10362.5 107027.5 ;
      RECT  10657.5 107822.5 10722.5 107957.5 ;
      RECT  10657.5 106847.5 10722.5 106982.5 ;
      RECT  10492.5 107122.5 10357.5 107187.5 ;
      RECT  10235.0 107337.5 10100.0 107402.5 ;
      RECT  10297.5 107732.5 10362.5 107867.5 ;
      RECT  10487.5 106892.5 10552.5 107027.5 ;
      RECT  10587.5 107337.5 10452.5 107402.5 ;
      RECT  10100.0 107337.5 10235.0 107402.5 ;
      RECT  10357.5 107122.5 10492.5 107187.5 ;
      RECT  10452.5 107337.5 10587.5 107402.5 ;
      RECT  10040.0 108042.5 10960.0 108107.5 ;
      RECT  10040.0 106697.5 10960.0 106762.5 ;
      RECT  11387.5 107890.0 11452.5 108075.0 ;
      RECT  11387.5 106730.0 11452.5 106915.0 ;
      RECT  11027.5 106847.5 11092.5 106697.5 ;
      RECT  11027.5 107732.5 11092.5 108107.5 ;
      RECT  11217.5 106847.5 11282.5 107732.5 ;
      RECT  11027.5 107732.5 11092.5 107867.5 ;
      RECT  11217.5 107732.5 11282.5 107867.5 ;
      RECT  11217.5 107732.5 11282.5 107867.5 ;
      RECT  11027.5 107732.5 11092.5 107867.5 ;
      RECT  11027.5 106847.5 11092.5 106982.5 ;
      RECT  11217.5 106847.5 11282.5 106982.5 ;
      RECT  11217.5 106847.5 11282.5 106982.5 ;
      RECT  11027.5 106847.5 11092.5 106982.5 ;
      RECT  11387.5 107822.5 11452.5 107957.5 ;
      RECT  11387.5 106847.5 11452.5 106982.5 ;
      RECT  11085.0 107290.0 11150.0 107425.0 ;
      RECT  11085.0 107290.0 11150.0 107425.0 ;
      RECT  11250.0 107325.0 11315.0 107390.0 ;
      RECT  10960.0 108042.5 11520.0 108107.5 ;
      RECT  10960.0 106697.5 11520.0 106762.5 ;
      RECT  9222.5 107290.0 9287.5 107425.0 ;
      RECT  9362.5 107017.5 9427.5 107152.5 ;
      RECT  10357.5 107122.5 10222.5 107187.5 ;
      RECT  9907.5 108260.0 9972.5 108075.0 ;
      RECT  9907.5 109420.0 9972.5 109235.0 ;
      RECT  9547.5 109302.5 9612.5 109452.5 ;
      RECT  9547.5 108417.5 9612.5 108042.5 ;
      RECT  9737.5 109302.5 9802.5 108417.5 ;
      RECT  9547.5 108417.5 9612.5 108282.5 ;
      RECT  9737.5 108417.5 9802.5 108282.5 ;
      RECT  9737.5 108417.5 9802.5 108282.5 ;
      RECT  9547.5 108417.5 9612.5 108282.5 ;
      RECT  9547.5 109302.5 9612.5 109167.5 ;
      RECT  9737.5 109302.5 9802.5 109167.5 ;
      RECT  9737.5 109302.5 9802.5 109167.5 ;
      RECT  9547.5 109302.5 9612.5 109167.5 ;
      RECT  9907.5 108327.5 9972.5 108192.5 ;
      RECT  9907.5 109302.5 9972.5 109167.5 ;
      RECT  9605.0 108860.0 9670.0 108725.0 ;
      RECT  9605.0 108860.0 9670.0 108725.0 ;
      RECT  9770.0 108825.0 9835.0 108760.0 ;
      RECT  9480.0 108107.5 10040.0 108042.5 ;
      RECT  9480.0 109452.5 10040.0 109387.5 ;
      RECT  10107.5 109257.5 10172.5 109452.5 ;
      RECT  10107.5 108417.5 10172.5 108042.5 ;
      RECT  10487.5 108417.5 10552.5 108042.5 ;
      RECT  10657.5 108260.0 10722.5 108075.0 ;
      RECT  10657.5 109420.0 10722.5 109235.0 ;
      RECT  10107.5 108417.5 10172.5 108282.5 ;
      RECT  10297.5 108417.5 10362.5 108282.5 ;
      RECT  10297.5 108417.5 10362.5 108282.5 ;
      RECT  10107.5 108417.5 10172.5 108282.5 ;
      RECT  10297.5 108417.5 10362.5 108282.5 ;
      RECT  10487.5 108417.5 10552.5 108282.5 ;
      RECT  10487.5 108417.5 10552.5 108282.5 ;
      RECT  10297.5 108417.5 10362.5 108282.5 ;
      RECT  10107.5 109257.5 10172.5 109122.5 ;
      RECT  10297.5 109257.5 10362.5 109122.5 ;
      RECT  10297.5 109257.5 10362.5 109122.5 ;
      RECT  10107.5 109257.5 10172.5 109122.5 ;
      RECT  10297.5 109257.5 10362.5 109122.5 ;
      RECT  10487.5 109257.5 10552.5 109122.5 ;
      RECT  10487.5 109257.5 10552.5 109122.5 ;
      RECT  10297.5 109257.5 10362.5 109122.5 ;
      RECT  10657.5 108327.5 10722.5 108192.5 ;
      RECT  10657.5 109302.5 10722.5 109167.5 ;
      RECT  10492.5 109027.5 10357.5 108962.5 ;
      RECT  10235.0 108812.5 10100.0 108747.5 ;
      RECT  10297.5 108417.5 10362.5 108282.5 ;
      RECT  10487.5 109257.5 10552.5 109122.5 ;
      RECT  10587.5 108812.5 10452.5 108747.5 ;
      RECT  10100.0 108812.5 10235.0 108747.5 ;
      RECT  10357.5 109027.5 10492.5 108962.5 ;
      RECT  10452.5 108812.5 10587.5 108747.5 ;
      RECT  10040.0 108107.5 10960.0 108042.5 ;
      RECT  10040.0 109452.5 10960.0 109387.5 ;
      RECT  11387.5 108260.0 11452.5 108075.0 ;
      RECT  11387.5 109420.0 11452.5 109235.0 ;
      RECT  11027.5 109302.5 11092.5 109452.5 ;
      RECT  11027.5 108417.5 11092.5 108042.5 ;
      RECT  11217.5 109302.5 11282.5 108417.5 ;
      RECT  11027.5 108417.5 11092.5 108282.5 ;
      RECT  11217.5 108417.5 11282.5 108282.5 ;
      RECT  11217.5 108417.5 11282.5 108282.5 ;
      RECT  11027.5 108417.5 11092.5 108282.5 ;
      RECT  11027.5 109302.5 11092.5 109167.5 ;
      RECT  11217.5 109302.5 11282.5 109167.5 ;
      RECT  11217.5 109302.5 11282.5 109167.5 ;
      RECT  11027.5 109302.5 11092.5 109167.5 ;
      RECT  11387.5 108327.5 11452.5 108192.5 ;
      RECT  11387.5 109302.5 11452.5 109167.5 ;
      RECT  11085.0 108860.0 11150.0 108725.0 ;
      RECT  11085.0 108860.0 11150.0 108725.0 ;
      RECT  11250.0 108825.0 11315.0 108760.0 ;
      RECT  10960.0 108107.5 11520.0 108042.5 ;
      RECT  10960.0 109452.5 11520.0 109387.5 ;
      RECT  9222.5 108725.0 9287.5 108860.0 ;
      RECT  9362.5 108997.5 9427.5 109132.5 ;
      RECT  10357.5 108962.5 10222.5 109027.5 ;
      RECT  9907.5 110580.0 9972.5 110765.0 ;
      RECT  9907.5 109420.0 9972.5 109605.0 ;
      RECT  9547.5 109537.5 9612.5 109387.5 ;
      RECT  9547.5 110422.5 9612.5 110797.5 ;
      RECT  9737.5 109537.5 9802.5 110422.5 ;
      RECT  9547.5 110422.5 9612.5 110557.5 ;
      RECT  9737.5 110422.5 9802.5 110557.5 ;
      RECT  9737.5 110422.5 9802.5 110557.5 ;
      RECT  9547.5 110422.5 9612.5 110557.5 ;
      RECT  9547.5 109537.5 9612.5 109672.5 ;
      RECT  9737.5 109537.5 9802.5 109672.5 ;
      RECT  9737.5 109537.5 9802.5 109672.5 ;
      RECT  9547.5 109537.5 9612.5 109672.5 ;
      RECT  9907.5 110512.5 9972.5 110647.5 ;
      RECT  9907.5 109537.5 9972.5 109672.5 ;
      RECT  9605.0 109980.0 9670.0 110115.0 ;
      RECT  9605.0 109980.0 9670.0 110115.0 ;
      RECT  9770.0 110015.0 9835.0 110080.0 ;
      RECT  9480.0 110732.5 10040.0 110797.5 ;
      RECT  9480.0 109387.5 10040.0 109452.5 ;
      RECT  10107.5 109582.5 10172.5 109387.5 ;
      RECT  10107.5 110422.5 10172.5 110797.5 ;
      RECT  10487.5 110422.5 10552.5 110797.5 ;
      RECT  10657.5 110580.0 10722.5 110765.0 ;
      RECT  10657.5 109420.0 10722.5 109605.0 ;
      RECT  10107.5 110422.5 10172.5 110557.5 ;
      RECT  10297.5 110422.5 10362.5 110557.5 ;
      RECT  10297.5 110422.5 10362.5 110557.5 ;
      RECT  10107.5 110422.5 10172.5 110557.5 ;
      RECT  10297.5 110422.5 10362.5 110557.5 ;
      RECT  10487.5 110422.5 10552.5 110557.5 ;
      RECT  10487.5 110422.5 10552.5 110557.5 ;
      RECT  10297.5 110422.5 10362.5 110557.5 ;
      RECT  10107.5 109582.5 10172.5 109717.5 ;
      RECT  10297.5 109582.5 10362.5 109717.5 ;
      RECT  10297.5 109582.5 10362.5 109717.5 ;
      RECT  10107.5 109582.5 10172.5 109717.5 ;
      RECT  10297.5 109582.5 10362.5 109717.5 ;
      RECT  10487.5 109582.5 10552.5 109717.5 ;
      RECT  10487.5 109582.5 10552.5 109717.5 ;
      RECT  10297.5 109582.5 10362.5 109717.5 ;
      RECT  10657.5 110512.5 10722.5 110647.5 ;
      RECT  10657.5 109537.5 10722.5 109672.5 ;
      RECT  10492.5 109812.5 10357.5 109877.5 ;
      RECT  10235.0 110027.5 10100.0 110092.5 ;
      RECT  10297.5 110422.5 10362.5 110557.5 ;
      RECT  10487.5 109582.5 10552.5 109717.5 ;
      RECT  10587.5 110027.5 10452.5 110092.5 ;
      RECT  10100.0 110027.5 10235.0 110092.5 ;
      RECT  10357.5 109812.5 10492.5 109877.5 ;
      RECT  10452.5 110027.5 10587.5 110092.5 ;
      RECT  10040.0 110732.5 10960.0 110797.5 ;
      RECT  10040.0 109387.5 10960.0 109452.5 ;
      RECT  11387.5 110580.0 11452.5 110765.0 ;
      RECT  11387.5 109420.0 11452.5 109605.0 ;
      RECT  11027.5 109537.5 11092.5 109387.5 ;
      RECT  11027.5 110422.5 11092.5 110797.5 ;
      RECT  11217.5 109537.5 11282.5 110422.5 ;
      RECT  11027.5 110422.5 11092.5 110557.5 ;
      RECT  11217.5 110422.5 11282.5 110557.5 ;
      RECT  11217.5 110422.5 11282.5 110557.5 ;
      RECT  11027.5 110422.5 11092.5 110557.5 ;
      RECT  11027.5 109537.5 11092.5 109672.5 ;
      RECT  11217.5 109537.5 11282.5 109672.5 ;
      RECT  11217.5 109537.5 11282.5 109672.5 ;
      RECT  11027.5 109537.5 11092.5 109672.5 ;
      RECT  11387.5 110512.5 11452.5 110647.5 ;
      RECT  11387.5 109537.5 11452.5 109672.5 ;
      RECT  11085.0 109980.0 11150.0 110115.0 ;
      RECT  11085.0 109980.0 11150.0 110115.0 ;
      RECT  11250.0 110015.0 11315.0 110080.0 ;
      RECT  10960.0 110732.5 11520.0 110797.5 ;
      RECT  10960.0 109387.5 11520.0 109452.5 ;
      RECT  9222.5 109980.0 9287.5 110115.0 ;
      RECT  9362.5 109707.5 9427.5 109842.5 ;
      RECT  10357.5 109812.5 10222.5 109877.5 ;
      RECT  9907.5 110950.0 9972.5 110765.0 ;
      RECT  9907.5 112110.0 9972.5 111925.0 ;
      RECT  9547.5 111992.5 9612.5 112142.5 ;
      RECT  9547.5 111107.5 9612.5 110732.5 ;
      RECT  9737.5 111992.5 9802.5 111107.5 ;
      RECT  9547.5 111107.5 9612.5 110972.5 ;
      RECT  9737.5 111107.5 9802.5 110972.5 ;
      RECT  9737.5 111107.5 9802.5 110972.5 ;
      RECT  9547.5 111107.5 9612.5 110972.5 ;
      RECT  9547.5 111992.5 9612.5 111857.5 ;
      RECT  9737.5 111992.5 9802.5 111857.5 ;
      RECT  9737.5 111992.5 9802.5 111857.5 ;
      RECT  9547.5 111992.5 9612.5 111857.5 ;
      RECT  9907.5 111017.5 9972.5 110882.5 ;
      RECT  9907.5 111992.5 9972.5 111857.5 ;
      RECT  9605.0 111550.0 9670.0 111415.0 ;
      RECT  9605.0 111550.0 9670.0 111415.0 ;
      RECT  9770.0 111515.0 9835.0 111450.0 ;
      RECT  9480.0 110797.5 10040.0 110732.5 ;
      RECT  9480.0 112142.5 10040.0 112077.5 ;
      RECT  10107.5 111947.5 10172.5 112142.5 ;
      RECT  10107.5 111107.5 10172.5 110732.5 ;
      RECT  10487.5 111107.5 10552.5 110732.5 ;
      RECT  10657.5 110950.0 10722.5 110765.0 ;
      RECT  10657.5 112110.0 10722.5 111925.0 ;
      RECT  10107.5 111107.5 10172.5 110972.5 ;
      RECT  10297.5 111107.5 10362.5 110972.5 ;
      RECT  10297.5 111107.5 10362.5 110972.5 ;
      RECT  10107.5 111107.5 10172.5 110972.5 ;
      RECT  10297.5 111107.5 10362.5 110972.5 ;
      RECT  10487.5 111107.5 10552.5 110972.5 ;
      RECT  10487.5 111107.5 10552.5 110972.5 ;
      RECT  10297.5 111107.5 10362.5 110972.5 ;
      RECT  10107.5 111947.5 10172.5 111812.5 ;
      RECT  10297.5 111947.5 10362.5 111812.5 ;
      RECT  10297.5 111947.5 10362.5 111812.5 ;
      RECT  10107.5 111947.5 10172.5 111812.5 ;
      RECT  10297.5 111947.5 10362.5 111812.5 ;
      RECT  10487.5 111947.5 10552.5 111812.5 ;
      RECT  10487.5 111947.5 10552.5 111812.5 ;
      RECT  10297.5 111947.5 10362.5 111812.5 ;
      RECT  10657.5 111017.5 10722.5 110882.5 ;
      RECT  10657.5 111992.5 10722.5 111857.5 ;
      RECT  10492.5 111717.5 10357.5 111652.5 ;
      RECT  10235.0 111502.5 10100.0 111437.5 ;
      RECT  10297.5 111107.5 10362.5 110972.5 ;
      RECT  10487.5 111947.5 10552.5 111812.5 ;
      RECT  10587.5 111502.5 10452.5 111437.5 ;
      RECT  10100.0 111502.5 10235.0 111437.5 ;
      RECT  10357.5 111717.5 10492.5 111652.5 ;
      RECT  10452.5 111502.5 10587.5 111437.5 ;
      RECT  10040.0 110797.5 10960.0 110732.5 ;
      RECT  10040.0 112142.5 10960.0 112077.5 ;
      RECT  11387.5 110950.0 11452.5 110765.0 ;
      RECT  11387.5 112110.0 11452.5 111925.0 ;
      RECT  11027.5 111992.5 11092.5 112142.5 ;
      RECT  11027.5 111107.5 11092.5 110732.5 ;
      RECT  11217.5 111992.5 11282.5 111107.5 ;
      RECT  11027.5 111107.5 11092.5 110972.5 ;
      RECT  11217.5 111107.5 11282.5 110972.5 ;
      RECT  11217.5 111107.5 11282.5 110972.5 ;
      RECT  11027.5 111107.5 11092.5 110972.5 ;
      RECT  11027.5 111992.5 11092.5 111857.5 ;
      RECT  11217.5 111992.5 11282.5 111857.5 ;
      RECT  11217.5 111992.5 11282.5 111857.5 ;
      RECT  11027.5 111992.5 11092.5 111857.5 ;
      RECT  11387.5 111017.5 11452.5 110882.5 ;
      RECT  11387.5 111992.5 11452.5 111857.5 ;
      RECT  11085.0 111550.0 11150.0 111415.0 ;
      RECT  11085.0 111550.0 11150.0 111415.0 ;
      RECT  11250.0 111515.0 11315.0 111450.0 ;
      RECT  10960.0 110797.5 11520.0 110732.5 ;
      RECT  10960.0 112142.5 11520.0 112077.5 ;
      RECT  9222.5 111415.0 9287.5 111550.0 ;
      RECT  9362.5 111687.5 9427.5 111822.5 ;
      RECT  10357.5 111652.5 10222.5 111717.5 ;
      RECT  9907.5 113270.0 9972.5 113455.0 ;
      RECT  9907.5 112110.0 9972.5 112295.0 ;
      RECT  9547.5 112227.5 9612.5 112077.5 ;
      RECT  9547.5 113112.5 9612.5 113487.5 ;
      RECT  9737.5 112227.5 9802.5 113112.5 ;
      RECT  9547.5 113112.5 9612.5 113247.5 ;
      RECT  9737.5 113112.5 9802.5 113247.5 ;
      RECT  9737.5 113112.5 9802.5 113247.5 ;
      RECT  9547.5 113112.5 9612.5 113247.5 ;
      RECT  9547.5 112227.5 9612.5 112362.5 ;
      RECT  9737.5 112227.5 9802.5 112362.5 ;
      RECT  9737.5 112227.5 9802.5 112362.5 ;
      RECT  9547.5 112227.5 9612.5 112362.5 ;
      RECT  9907.5 113202.5 9972.5 113337.5 ;
      RECT  9907.5 112227.5 9972.5 112362.5 ;
      RECT  9605.0 112670.0 9670.0 112805.0 ;
      RECT  9605.0 112670.0 9670.0 112805.0 ;
      RECT  9770.0 112705.0 9835.0 112770.0 ;
      RECT  9480.0 113422.5 10040.0 113487.5 ;
      RECT  9480.0 112077.5 10040.0 112142.5 ;
      RECT  10107.5 112272.5 10172.5 112077.5 ;
      RECT  10107.5 113112.5 10172.5 113487.5 ;
      RECT  10487.5 113112.5 10552.5 113487.5 ;
      RECT  10657.5 113270.0 10722.5 113455.0 ;
      RECT  10657.5 112110.0 10722.5 112295.0 ;
      RECT  10107.5 113112.5 10172.5 113247.5 ;
      RECT  10297.5 113112.5 10362.5 113247.5 ;
      RECT  10297.5 113112.5 10362.5 113247.5 ;
      RECT  10107.5 113112.5 10172.5 113247.5 ;
      RECT  10297.5 113112.5 10362.5 113247.5 ;
      RECT  10487.5 113112.5 10552.5 113247.5 ;
      RECT  10487.5 113112.5 10552.5 113247.5 ;
      RECT  10297.5 113112.5 10362.5 113247.5 ;
      RECT  10107.5 112272.5 10172.5 112407.5 ;
      RECT  10297.5 112272.5 10362.5 112407.5 ;
      RECT  10297.5 112272.5 10362.5 112407.5 ;
      RECT  10107.5 112272.5 10172.5 112407.5 ;
      RECT  10297.5 112272.5 10362.5 112407.5 ;
      RECT  10487.5 112272.5 10552.5 112407.5 ;
      RECT  10487.5 112272.5 10552.5 112407.5 ;
      RECT  10297.5 112272.5 10362.5 112407.5 ;
      RECT  10657.5 113202.5 10722.5 113337.5 ;
      RECT  10657.5 112227.5 10722.5 112362.5 ;
      RECT  10492.5 112502.5 10357.5 112567.5 ;
      RECT  10235.0 112717.5 10100.0 112782.5 ;
      RECT  10297.5 113112.5 10362.5 113247.5 ;
      RECT  10487.5 112272.5 10552.5 112407.5 ;
      RECT  10587.5 112717.5 10452.5 112782.5 ;
      RECT  10100.0 112717.5 10235.0 112782.5 ;
      RECT  10357.5 112502.5 10492.5 112567.5 ;
      RECT  10452.5 112717.5 10587.5 112782.5 ;
      RECT  10040.0 113422.5 10960.0 113487.5 ;
      RECT  10040.0 112077.5 10960.0 112142.5 ;
      RECT  11387.5 113270.0 11452.5 113455.0 ;
      RECT  11387.5 112110.0 11452.5 112295.0 ;
      RECT  11027.5 112227.5 11092.5 112077.5 ;
      RECT  11027.5 113112.5 11092.5 113487.5 ;
      RECT  11217.5 112227.5 11282.5 113112.5 ;
      RECT  11027.5 113112.5 11092.5 113247.5 ;
      RECT  11217.5 113112.5 11282.5 113247.5 ;
      RECT  11217.5 113112.5 11282.5 113247.5 ;
      RECT  11027.5 113112.5 11092.5 113247.5 ;
      RECT  11027.5 112227.5 11092.5 112362.5 ;
      RECT  11217.5 112227.5 11282.5 112362.5 ;
      RECT  11217.5 112227.5 11282.5 112362.5 ;
      RECT  11027.5 112227.5 11092.5 112362.5 ;
      RECT  11387.5 113202.5 11452.5 113337.5 ;
      RECT  11387.5 112227.5 11452.5 112362.5 ;
      RECT  11085.0 112670.0 11150.0 112805.0 ;
      RECT  11085.0 112670.0 11150.0 112805.0 ;
      RECT  11250.0 112705.0 11315.0 112770.0 ;
      RECT  10960.0 113422.5 11520.0 113487.5 ;
      RECT  10960.0 112077.5 11520.0 112142.5 ;
      RECT  9222.5 112670.0 9287.5 112805.0 ;
      RECT  9362.5 112397.5 9427.5 112532.5 ;
      RECT  10357.5 112502.5 10222.5 112567.5 ;
      RECT  9907.5 113640.0 9972.5 113455.0 ;
      RECT  9907.5 114800.0 9972.5 114615.0 ;
      RECT  9547.5 114682.5 9612.5 114832.5 ;
      RECT  9547.5 113797.5 9612.5 113422.5 ;
      RECT  9737.5 114682.5 9802.5 113797.5 ;
      RECT  9547.5 113797.5 9612.5 113662.5 ;
      RECT  9737.5 113797.5 9802.5 113662.5 ;
      RECT  9737.5 113797.5 9802.5 113662.5 ;
      RECT  9547.5 113797.5 9612.5 113662.5 ;
      RECT  9547.5 114682.5 9612.5 114547.5 ;
      RECT  9737.5 114682.5 9802.5 114547.5 ;
      RECT  9737.5 114682.5 9802.5 114547.5 ;
      RECT  9547.5 114682.5 9612.5 114547.5 ;
      RECT  9907.5 113707.5 9972.5 113572.5 ;
      RECT  9907.5 114682.5 9972.5 114547.5 ;
      RECT  9605.0 114240.0 9670.0 114105.0 ;
      RECT  9605.0 114240.0 9670.0 114105.0 ;
      RECT  9770.0 114205.0 9835.0 114140.0 ;
      RECT  9480.0 113487.5 10040.0 113422.5 ;
      RECT  9480.0 114832.5 10040.0 114767.5 ;
      RECT  10107.5 114637.5 10172.5 114832.5 ;
      RECT  10107.5 113797.5 10172.5 113422.5 ;
      RECT  10487.5 113797.5 10552.5 113422.5 ;
      RECT  10657.5 113640.0 10722.5 113455.0 ;
      RECT  10657.5 114800.0 10722.5 114615.0 ;
      RECT  10107.5 113797.5 10172.5 113662.5 ;
      RECT  10297.5 113797.5 10362.5 113662.5 ;
      RECT  10297.5 113797.5 10362.5 113662.5 ;
      RECT  10107.5 113797.5 10172.5 113662.5 ;
      RECT  10297.5 113797.5 10362.5 113662.5 ;
      RECT  10487.5 113797.5 10552.5 113662.5 ;
      RECT  10487.5 113797.5 10552.5 113662.5 ;
      RECT  10297.5 113797.5 10362.5 113662.5 ;
      RECT  10107.5 114637.5 10172.5 114502.5 ;
      RECT  10297.5 114637.5 10362.5 114502.5 ;
      RECT  10297.5 114637.5 10362.5 114502.5 ;
      RECT  10107.5 114637.5 10172.5 114502.5 ;
      RECT  10297.5 114637.5 10362.5 114502.5 ;
      RECT  10487.5 114637.5 10552.5 114502.5 ;
      RECT  10487.5 114637.5 10552.5 114502.5 ;
      RECT  10297.5 114637.5 10362.5 114502.5 ;
      RECT  10657.5 113707.5 10722.5 113572.5 ;
      RECT  10657.5 114682.5 10722.5 114547.5 ;
      RECT  10492.5 114407.5 10357.5 114342.5 ;
      RECT  10235.0 114192.5 10100.0 114127.5 ;
      RECT  10297.5 113797.5 10362.5 113662.5 ;
      RECT  10487.5 114637.5 10552.5 114502.5 ;
      RECT  10587.5 114192.5 10452.5 114127.5 ;
      RECT  10100.0 114192.5 10235.0 114127.5 ;
      RECT  10357.5 114407.5 10492.5 114342.5 ;
      RECT  10452.5 114192.5 10587.5 114127.5 ;
      RECT  10040.0 113487.5 10960.0 113422.5 ;
      RECT  10040.0 114832.5 10960.0 114767.5 ;
      RECT  11387.5 113640.0 11452.5 113455.0 ;
      RECT  11387.5 114800.0 11452.5 114615.0 ;
      RECT  11027.5 114682.5 11092.5 114832.5 ;
      RECT  11027.5 113797.5 11092.5 113422.5 ;
      RECT  11217.5 114682.5 11282.5 113797.5 ;
      RECT  11027.5 113797.5 11092.5 113662.5 ;
      RECT  11217.5 113797.5 11282.5 113662.5 ;
      RECT  11217.5 113797.5 11282.5 113662.5 ;
      RECT  11027.5 113797.5 11092.5 113662.5 ;
      RECT  11027.5 114682.5 11092.5 114547.5 ;
      RECT  11217.5 114682.5 11282.5 114547.5 ;
      RECT  11217.5 114682.5 11282.5 114547.5 ;
      RECT  11027.5 114682.5 11092.5 114547.5 ;
      RECT  11387.5 113707.5 11452.5 113572.5 ;
      RECT  11387.5 114682.5 11452.5 114547.5 ;
      RECT  11085.0 114240.0 11150.0 114105.0 ;
      RECT  11085.0 114240.0 11150.0 114105.0 ;
      RECT  11250.0 114205.0 11315.0 114140.0 ;
      RECT  10960.0 113487.5 11520.0 113422.5 ;
      RECT  10960.0 114832.5 11520.0 114767.5 ;
      RECT  9222.5 114105.0 9287.5 114240.0 ;
      RECT  9362.5 114377.5 9427.5 114512.5 ;
      RECT  10357.5 114342.5 10222.5 114407.5 ;
      RECT  9907.5 115960.0 9972.5 116145.0 ;
      RECT  9907.5 114800.0 9972.5 114985.0 ;
      RECT  9547.5 114917.5 9612.5 114767.5 ;
      RECT  9547.5 115802.5 9612.5 116177.5 ;
      RECT  9737.5 114917.5 9802.5 115802.5 ;
      RECT  9547.5 115802.5 9612.5 115937.5 ;
      RECT  9737.5 115802.5 9802.5 115937.5 ;
      RECT  9737.5 115802.5 9802.5 115937.5 ;
      RECT  9547.5 115802.5 9612.5 115937.5 ;
      RECT  9547.5 114917.5 9612.5 115052.5 ;
      RECT  9737.5 114917.5 9802.5 115052.5 ;
      RECT  9737.5 114917.5 9802.5 115052.5 ;
      RECT  9547.5 114917.5 9612.5 115052.5 ;
      RECT  9907.5 115892.5 9972.5 116027.5 ;
      RECT  9907.5 114917.5 9972.5 115052.5 ;
      RECT  9605.0 115360.0 9670.0 115495.0 ;
      RECT  9605.0 115360.0 9670.0 115495.0 ;
      RECT  9770.0 115395.0 9835.0 115460.0 ;
      RECT  9480.0 116112.5 10040.0 116177.5 ;
      RECT  9480.0 114767.5 10040.0 114832.5 ;
      RECT  10107.5 114962.5 10172.5 114767.5 ;
      RECT  10107.5 115802.5 10172.5 116177.5 ;
      RECT  10487.5 115802.5 10552.5 116177.5 ;
      RECT  10657.5 115960.0 10722.5 116145.0 ;
      RECT  10657.5 114800.0 10722.5 114985.0 ;
      RECT  10107.5 115802.5 10172.5 115937.5 ;
      RECT  10297.5 115802.5 10362.5 115937.5 ;
      RECT  10297.5 115802.5 10362.5 115937.5 ;
      RECT  10107.5 115802.5 10172.5 115937.5 ;
      RECT  10297.5 115802.5 10362.5 115937.5 ;
      RECT  10487.5 115802.5 10552.5 115937.5 ;
      RECT  10487.5 115802.5 10552.5 115937.5 ;
      RECT  10297.5 115802.5 10362.5 115937.5 ;
      RECT  10107.5 114962.5 10172.5 115097.5 ;
      RECT  10297.5 114962.5 10362.5 115097.5 ;
      RECT  10297.5 114962.5 10362.5 115097.5 ;
      RECT  10107.5 114962.5 10172.5 115097.5 ;
      RECT  10297.5 114962.5 10362.5 115097.5 ;
      RECT  10487.5 114962.5 10552.5 115097.5 ;
      RECT  10487.5 114962.5 10552.5 115097.5 ;
      RECT  10297.5 114962.5 10362.5 115097.5 ;
      RECT  10657.5 115892.5 10722.5 116027.5 ;
      RECT  10657.5 114917.5 10722.5 115052.5 ;
      RECT  10492.5 115192.5 10357.5 115257.5 ;
      RECT  10235.0 115407.5 10100.0 115472.5 ;
      RECT  10297.5 115802.5 10362.5 115937.5 ;
      RECT  10487.5 114962.5 10552.5 115097.5 ;
      RECT  10587.5 115407.5 10452.5 115472.5 ;
      RECT  10100.0 115407.5 10235.0 115472.5 ;
      RECT  10357.5 115192.5 10492.5 115257.5 ;
      RECT  10452.5 115407.5 10587.5 115472.5 ;
      RECT  10040.0 116112.5 10960.0 116177.5 ;
      RECT  10040.0 114767.5 10960.0 114832.5 ;
      RECT  11387.5 115960.0 11452.5 116145.0 ;
      RECT  11387.5 114800.0 11452.5 114985.0 ;
      RECT  11027.5 114917.5 11092.5 114767.5 ;
      RECT  11027.5 115802.5 11092.5 116177.5 ;
      RECT  11217.5 114917.5 11282.5 115802.5 ;
      RECT  11027.5 115802.5 11092.5 115937.5 ;
      RECT  11217.5 115802.5 11282.5 115937.5 ;
      RECT  11217.5 115802.5 11282.5 115937.5 ;
      RECT  11027.5 115802.5 11092.5 115937.5 ;
      RECT  11027.5 114917.5 11092.5 115052.5 ;
      RECT  11217.5 114917.5 11282.5 115052.5 ;
      RECT  11217.5 114917.5 11282.5 115052.5 ;
      RECT  11027.5 114917.5 11092.5 115052.5 ;
      RECT  11387.5 115892.5 11452.5 116027.5 ;
      RECT  11387.5 114917.5 11452.5 115052.5 ;
      RECT  11085.0 115360.0 11150.0 115495.0 ;
      RECT  11085.0 115360.0 11150.0 115495.0 ;
      RECT  11250.0 115395.0 11315.0 115460.0 ;
      RECT  10960.0 116112.5 11520.0 116177.5 ;
      RECT  10960.0 114767.5 11520.0 114832.5 ;
      RECT  9222.5 115360.0 9287.5 115495.0 ;
      RECT  9362.5 115087.5 9427.5 115222.5 ;
      RECT  10357.5 115192.5 10222.5 115257.5 ;
      RECT  9907.5 116330.0 9972.5 116145.0 ;
      RECT  9907.5 117490.0 9972.5 117305.0 ;
      RECT  9547.5 117372.5 9612.5 117522.5 ;
      RECT  9547.5 116487.5 9612.5 116112.5 ;
      RECT  9737.5 117372.5 9802.5 116487.5 ;
      RECT  9547.5 116487.5 9612.5 116352.5 ;
      RECT  9737.5 116487.5 9802.5 116352.5 ;
      RECT  9737.5 116487.5 9802.5 116352.5 ;
      RECT  9547.5 116487.5 9612.5 116352.5 ;
      RECT  9547.5 117372.5 9612.5 117237.5 ;
      RECT  9737.5 117372.5 9802.5 117237.5 ;
      RECT  9737.5 117372.5 9802.5 117237.5 ;
      RECT  9547.5 117372.5 9612.5 117237.5 ;
      RECT  9907.5 116397.5 9972.5 116262.5 ;
      RECT  9907.5 117372.5 9972.5 117237.5 ;
      RECT  9605.0 116930.0 9670.0 116795.0 ;
      RECT  9605.0 116930.0 9670.0 116795.0 ;
      RECT  9770.0 116895.0 9835.0 116830.0 ;
      RECT  9480.0 116177.5 10040.0 116112.5 ;
      RECT  9480.0 117522.5 10040.0 117457.5 ;
      RECT  10107.5 117327.5 10172.5 117522.5 ;
      RECT  10107.5 116487.5 10172.5 116112.5 ;
      RECT  10487.5 116487.5 10552.5 116112.5 ;
      RECT  10657.5 116330.0 10722.5 116145.0 ;
      RECT  10657.5 117490.0 10722.5 117305.0 ;
      RECT  10107.5 116487.5 10172.5 116352.5 ;
      RECT  10297.5 116487.5 10362.5 116352.5 ;
      RECT  10297.5 116487.5 10362.5 116352.5 ;
      RECT  10107.5 116487.5 10172.5 116352.5 ;
      RECT  10297.5 116487.5 10362.5 116352.5 ;
      RECT  10487.5 116487.5 10552.5 116352.5 ;
      RECT  10487.5 116487.5 10552.5 116352.5 ;
      RECT  10297.5 116487.5 10362.5 116352.5 ;
      RECT  10107.5 117327.5 10172.5 117192.5 ;
      RECT  10297.5 117327.5 10362.5 117192.5 ;
      RECT  10297.5 117327.5 10362.5 117192.5 ;
      RECT  10107.5 117327.5 10172.5 117192.5 ;
      RECT  10297.5 117327.5 10362.5 117192.5 ;
      RECT  10487.5 117327.5 10552.5 117192.5 ;
      RECT  10487.5 117327.5 10552.5 117192.5 ;
      RECT  10297.5 117327.5 10362.5 117192.5 ;
      RECT  10657.5 116397.5 10722.5 116262.5 ;
      RECT  10657.5 117372.5 10722.5 117237.5 ;
      RECT  10492.5 117097.5 10357.5 117032.5 ;
      RECT  10235.0 116882.5 10100.0 116817.5 ;
      RECT  10297.5 116487.5 10362.5 116352.5 ;
      RECT  10487.5 117327.5 10552.5 117192.5 ;
      RECT  10587.5 116882.5 10452.5 116817.5 ;
      RECT  10100.0 116882.5 10235.0 116817.5 ;
      RECT  10357.5 117097.5 10492.5 117032.5 ;
      RECT  10452.5 116882.5 10587.5 116817.5 ;
      RECT  10040.0 116177.5 10960.0 116112.5 ;
      RECT  10040.0 117522.5 10960.0 117457.5 ;
      RECT  11387.5 116330.0 11452.5 116145.0 ;
      RECT  11387.5 117490.0 11452.5 117305.0 ;
      RECT  11027.5 117372.5 11092.5 117522.5 ;
      RECT  11027.5 116487.5 11092.5 116112.5 ;
      RECT  11217.5 117372.5 11282.5 116487.5 ;
      RECT  11027.5 116487.5 11092.5 116352.5 ;
      RECT  11217.5 116487.5 11282.5 116352.5 ;
      RECT  11217.5 116487.5 11282.5 116352.5 ;
      RECT  11027.5 116487.5 11092.5 116352.5 ;
      RECT  11027.5 117372.5 11092.5 117237.5 ;
      RECT  11217.5 117372.5 11282.5 117237.5 ;
      RECT  11217.5 117372.5 11282.5 117237.5 ;
      RECT  11027.5 117372.5 11092.5 117237.5 ;
      RECT  11387.5 116397.5 11452.5 116262.5 ;
      RECT  11387.5 117372.5 11452.5 117237.5 ;
      RECT  11085.0 116930.0 11150.0 116795.0 ;
      RECT  11085.0 116930.0 11150.0 116795.0 ;
      RECT  11250.0 116895.0 11315.0 116830.0 ;
      RECT  10960.0 116177.5 11520.0 116112.5 ;
      RECT  10960.0 117522.5 11520.0 117457.5 ;
      RECT  9222.5 116795.0 9287.5 116930.0 ;
      RECT  9362.5 117067.5 9427.5 117202.5 ;
      RECT  10357.5 117032.5 10222.5 117097.5 ;
      RECT  9907.5 118650.0 9972.5 118835.0 ;
      RECT  9907.5 117490.0 9972.5 117675.0 ;
      RECT  9547.5 117607.5 9612.5 117457.5 ;
      RECT  9547.5 118492.5 9612.5 118867.5 ;
      RECT  9737.5 117607.5 9802.5 118492.5 ;
      RECT  9547.5 118492.5 9612.5 118627.5 ;
      RECT  9737.5 118492.5 9802.5 118627.5 ;
      RECT  9737.5 118492.5 9802.5 118627.5 ;
      RECT  9547.5 118492.5 9612.5 118627.5 ;
      RECT  9547.5 117607.5 9612.5 117742.5 ;
      RECT  9737.5 117607.5 9802.5 117742.5 ;
      RECT  9737.5 117607.5 9802.5 117742.5 ;
      RECT  9547.5 117607.5 9612.5 117742.5 ;
      RECT  9907.5 118582.5 9972.5 118717.5 ;
      RECT  9907.5 117607.5 9972.5 117742.5 ;
      RECT  9605.0 118050.0 9670.0 118185.0 ;
      RECT  9605.0 118050.0 9670.0 118185.0 ;
      RECT  9770.0 118085.0 9835.0 118150.0 ;
      RECT  9480.0 118802.5 10040.0 118867.5 ;
      RECT  9480.0 117457.5 10040.0 117522.5 ;
      RECT  10107.5 117652.5 10172.5 117457.5 ;
      RECT  10107.5 118492.5 10172.5 118867.5 ;
      RECT  10487.5 118492.5 10552.5 118867.5 ;
      RECT  10657.5 118650.0 10722.5 118835.0 ;
      RECT  10657.5 117490.0 10722.5 117675.0 ;
      RECT  10107.5 118492.5 10172.5 118627.5 ;
      RECT  10297.5 118492.5 10362.5 118627.5 ;
      RECT  10297.5 118492.5 10362.5 118627.5 ;
      RECT  10107.5 118492.5 10172.5 118627.5 ;
      RECT  10297.5 118492.5 10362.5 118627.5 ;
      RECT  10487.5 118492.5 10552.5 118627.5 ;
      RECT  10487.5 118492.5 10552.5 118627.5 ;
      RECT  10297.5 118492.5 10362.5 118627.5 ;
      RECT  10107.5 117652.5 10172.5 117787.5 ;
      RECT  10297.5 117652.5 10362.5 117787.5 ;
      RECT  10297.5 117652.5 10362.5 117787.5 ;
      RECT  10107.5 117652.5 10172.5 117787.5 ;
      RECT  10297.5 117652.5 10362.5 117787.5 ;
      RECT  10487.5 117652.5 10552.5 117787.5 ;
      RECT  10487.5 117652.5 10552.5 117787.5 ;
      RECT  10297.5 117652.5 10362.5 117787.5 ;
      RECT  10657.5 118582.5 10722.5 118717.5 ;
      RECT  10657.5 117607.5 10722.5 117742.5 ;
      RECT  10492.5 117882.5 10357.5 117947.5 ;
      RECT  10235.0 118097.5 10100.0 118162.5 ;
      RECT  10297.5 118492.5 10362.5 118627.5 ;
      RECT  10487.5 117652.5 10552.5 117787.5 ;
      RECT  10587.5 118097.5 10452.5 118162.5 ;
      RECT  10100.0 118097.5 10235.0 118162.5 ;
      RECT  10357.5 117882.5 10492.5 117947.5 ;
      RECT  10452.5 118097.5 10587.5 118162.5 ;
      RECT  10040.0 118802.5 10960.0 118867.5 ;
      RECT  10040.0 117457.5 10960.0 117522.5 ;
      RECT  11387.5 118650.0 11452.5 118835.0 ;
      RECT  11387.5 117490.0 11452.5 117675.0 ;
      RECT  11027.5 117607.5 11092.5 117457.5 ;
      RECT  11027.5 118492.5 11092.5 118867.5 ;
      RECT  11217.5 117607.5 11282.5 118492.5 ;
      RECT  11027.5 118492.5 11092.5 118627.5 ;
      RECT  11217.5 118492.5 11282.5 118627.5 ;
      RECT  11217.5 118492.5 11282.5 118627.5 ;
      RECT  11027.5 118492.5 11092.5 118627.5 ;
      RECT  11027.5 117607.5 11092.5 117742.5 ;
      RECT  11217.5 117607.5 11282.5 117742.5 ;
      RECT  11217.5 117607.5 11282.5 117742.5 ;
      RECT  11027.5 117607.5 11092.5 117742.5 ;
      RECT  11387.5 118582.5 11452.5 118717.5 ;
      RECT  11387.5 117607.5 11452.5 117742.5 ;
      RECT  11085.0 118050.0 11150.0 118185.0 ;
      RECT  11085.0 118050.0 11150.0 118185.0 ;
      RECT  11250.0 118085.0 11315.0 118150.0 ;
      RECT  10960.0 118802.5 11520.0 118867.5 ;
      RECT  10960.0 117457.5 11520.0 117522.5 ;
      RECT  9222.5 118050.0 9287.5 118185.0 ;
      RECT  9362.5 117777.5 9427.5 117912.5 ;
      RECT  10357.5 117882.5 10222.5 117947.5 ;
      RECT  9907.5 119020.0 9972.5 118835.0 ;
      RECT  9907.5 120180.0 9972.5 119995.0 ;
      RECT  9547.5 120062.5 9612.5 120212.5 ;
      RECT  9547.5 119177.5 9612.5 118802.5 ;
      RECT  9737.5 120062.5 9802.5 119177.5 ;
      RECT  9547.5 119177.5 9612.5 119042.5 ;
      RECT  9737.5 119177.5 9802.5 119042.5 ;
      RECT  9737.5 119177.5 9802.5 119042.5 ;
      RECT  9547.5 119177.5 9612.5 119042.5 ;
      RECT  9547.5 120062.5 9612.5 119927.5 ;
      RECT  9737.5 120062.5 9802.5 119927.5 ;
      RECT  9737.5 120062.5 9802.5 119927.5 ;
      RECT  9547.5 120062.5 9612.5 119927.5 ;
      RECT  9907.5 119087.5 9972.5 118952.5 ;
      RECT  9907.5 120062.5 9972.5 119927.5 ;
      RECT  9605.0 119620.0 9670.0 119485.0 ;
      RECT  9605.0 119620.0 9670.0 119485.0 ;
      RECT  9770.0 119585.0 9835.0 119520.0 ;
      RECT  9480.0 118867.5 10040.0 118802.5 ;
      RECT  9480.0 120212.5 10040.0 120147.5 ;
      RECT  10107.5 120017.5 10172.5 120212.5 ;
      RECT  10107.5 119177.5 10172.5 118802.5 ;
      RECT  10487.5 119177.5 10552.5 118802.5 ;
      RECT  10657.5 119020.0 10722.5 118835.0 ;
      RECT  10657.5 120180.0 10722.5 119995.0 ;
      RECT  10107.5 119177.5 10172.5 119042.5 ;
      RECT  10297.5 119177.5 10362.5 119042.5 ;
      RECT  10297.5 119177.5 10362.5 119042.5 ;
      RECT  10107.5 119177.5 10172.5 119042.5 ;
      RECT  10297.5 119177.5 10362.5 119042.5 ;
      RECT  10487.5 119177.5 10552.5 119042.5 ;
      RECT  10487.5 119177.5 10552.5 119042.5 ;
      RECT  10297.5 119177.5 10362.5 119042.5 ;
      RECT  10107.5 120017.5 10172.5 119882.5 ;
      RECT  10297.5 120017.5 10362.5 119882.5 ;
      RECT  10297.5 120017.5 10362.5 119882.5 ;
      RECT  10107.5 120017.5 10172.5 119882.5 ;
      RECT  10297.5 120017.5 10362.5 119882.5 ;
      RECT  10487.5 120017.5 10552.5 119882.5 ;
      RECT  10487.5 120017.5 10552.5 119882.5 ;
      RECT  10297.5 120017.5 10362.5 119882.5 ;
      RECT  10657.5 119087.5 10722.5 118952.5 ;
      RECT  10657.5 120062.5 10722.5 119927.5 ;
      RECT  10492.5 119787.5 10357.5 119722.5 ;
      RECT  10235.0 119572.5 10100.0 119507.5 ;
      RECT  10297.5 119177.5 10362.5 119042.5 ;
      RECT  10487.5 120017.5 10552.5 119882.5 ;
      RECT  10587.5 119572.5 10452.5 119507.5 ;
      RECT  10100.0 119572.5 10235.0 119507.5 ;
      RECT  10357.5 119787.5 10492.5 119722.5 ;
      RECT  10452.5 119572.5 10587.5 119507.5 ;
      RECT  10040.0 118867.5 10960.0 118802.5 ;
      RECT  10040.0 120212.5 10960.0 120147.5 ;
      RECT  11387.5 119020.0 11452.5 118835.0 ;
      RECT  11387.5 120180.0 11452.5 119995.0 ;
      RECT  11027.5 120062.5 11092.5 120212.5 ;
      RECT  11027.5 119177.5 11092.5 118802.5 ;
      RECT  11217.5 120062.5 11282.5 119177.5 ;
      RECT  11027.5 119177.5 11092.5 119042.5 ;
      RECT  11217.5 119177.5 11282.5 119042.5 ;
      RECT  11217.5 119177.5 11282.5 119042.5 ;
      RECT  11027.5 119177.5 11092.5 119042.5 ;
      RECT  11027.5 120062.5 11092.5 119927.5 ;
      RECT  11217.5 120062.5 11282.5 119927.5 ;
      RECT  11217.5 120062.5 11282.5 119927.5 ;
      RECT  11027.5 120062.5 11092.5 119927.5 ;
      RECT  11387.5 119087.5 11452.5 118952.5 ;
      RECT  11387.5 120062.5 11452.5 119927.5 ;
      RECT  11085.0 119620.0 11150.0 119485.0 ;
      RECT  11085.0 119620.0 11150.0 119485.0 ;
      RECT  11250.0 119585.0 11315.0 119520.0 ;
      RECT  10960.0 118867.5 11520.0 118802.5 ;
      RECT  10960.0 120212.5 11520.0 120147.5 ;
      RECT  9222.5 119485.0 9287.5 119620.0 ;
      RECT  9362.5 119757.5 9427.5 119892.5 ;
      RECT  10357.5 119722.5 10222.5 119787.5 ;
      RECT  9907.5 121340.0 9972.5 121525.0 ;
      RECT  9907.5 120180.0 9972.5 120365.0 ;
      RECT  9547.5 120297.5 9612.5 120147.5 ;
      RECT  9547.5 121182.5 9612.5 121557.5 ;
      RECT  9737.5 120297.5 9802.5 121182.5 ;
      RECT  9547.5 121182.5 9612.5 121317.5 ;
      RECT  9737.5 121182.5 9802.5 121317.5 ;
      RECT  9737.5 121182.5 9802.5 121317.5 ;
      RECT  9547.5 121182.5 9612.5 121317.5 ;
      RECT  9547.5 120297.5 9612.5 120432.5 ;
      RECT  9737.5 120297.5 9802.5 120432.5 ;
      RECT  9737.5 120297.5 9802.5 120432.5 ;
      RECT  9547.5 120297.5 9612.5 120432.5 ;
      RECT  9907.5 121272.5 9972.5 121407.5 ;
      RECT  9907.5 120297.5 9972.5 120432.5 ;
      RECT  9605.0 120740.0 9670.0 120875.0 ;
      RECT  9605.0 120740.0 9670.0 120875.0 ;
      RECT  9770.0 120775.0 9835.0 120840.0 ;
      RECT  9480.0 121492.5 10040.0 121557.5 ;
      RECT  9480.0 120147.5 10040.0 120212.5 ;
      RECT  10107.5 120342.5 10172.5 120147.5 ;
      RECT  10107.5 121182.5 10172.5 121557.5 ;
      RECT  10487.5 121182.5 10552.5 121557.5 ;
      RECT  10657.5 121340.0 10722.5 121525.0 ;
      RECT  10657.5 120180.0 10722.5 120365.0 ;
      RECT  10107.5 121182.5 10172.5 121317.5 ;
      RECT  10297.5 121182.5 10362.5 121317.5 ;
      RECT  10297.5 121182.5 10362.5 121317.5 ;
      RECT  10107.5 121182.5 10172.5 121317.5 ;
      RECT  10297.5 121182.5 10362.5 121317.5 ;
      RECT  10487.5 121182.5 10552.5 121317.5 ;
      RECT  10487.5 121182.5 10552.5 121317.5 ;
      RECT  10297.5 121182.5 10362.5 121317.5 ;
      RECT  10107.5 120342.5 10172.5 120477.5 ;
      RECT  10297.5 120342.5 10362.5 120477.5 ;
      RECT  10297.5 120342.5 10362.5 120477.5 ;
      RECT  10107.5 120342.5 10172.5 120477.5 ;
      RECT  10297.5 120342.5 10362.5 120477.5 ;
      RECT  10487.5 120342.5 10552.5 120477.5 ;
      RECT  10487.5 120342.5 10552.5 120477.5 ;
      RECT  10297.5 120342.5 10362.5 120477.5 ;
      RECT  10657.5 121272.5 10722.5 121407.5 ;
      RECT  10657.5 120297.5 10722.5 120432.5 ;
      RECT  10492.5 120572.5 10357.5 120637.5 ;
      RECT  10235.0 120787.5 10100.0 120852.5 ;
      RECT  10297.5 121182.5 10362.5 121317.5 ;
      RECT  10487.5 120342.5 10552.5 120477.5 ;
      RECT  10587.5 120787.5 10452.5 120852.5 ;
      RECT  10100.0 120787.5 10235.0 120852.5 ;
      RECT  10357.5 120572.5 10492.5 120637.5 ;
      RECT  10452.5 120787.5 10587.5 120852.5 ;
      RECT  10040.0 121492.5 10960.0 121557.5 ;
      RECT  10040.0 120147.5 10960.0 120212.5 ;
      RECT  11387.5 121340.0 11452.5 121525.0 ;
      RECT  11387.5 120180.0 11452.5 120365.0 ;
      RECT  11027.5 120297.5 11092.5 120147.5 ;
      RECT  11027.5 121182.5 11092.5 121557.5 ;
      RECT  11217.5 120297.5 11282.5 121182.5 ;
      RECT  11027.5 121182.5 11092.5 121317.5 ;
      RECT  11217.5 121182.5 11282.5 121317.5 ;
      RECT  11217.5 121182.5 11282.5 121317.5 ;
      RECT  11027.5 121182.5 11092.5 121317.5 ;
      RECT  11027.5 120297.5 11092.5 120432.5 ;
      RECT  11217.5 120297.5 11282.5 120432.5 ;
      RECT  11217.5 120297.5 11282.5 120432.5 ;
      RECT  11027.5 120297.5 11092.5 120432.5 ;
      RECT  11387.5 121272.5 11452.5 121407.5 ;
      RECT  11387.5 120297.5 11452.5 120432.5 ;
      RECT  11085.0 120740.0 11150.0 120875.0 ;
      RECT  11085.0 120740.0 11150.0 120875.0 ;
      RECT  11250.0 120775.0 11315.0 120840.0 ;
      RECT  10960.0 121492.5 11520.0 121557.5 ;
      RECT  10960.0 120147.5 11520.0 120212.5 ;
      RECT  9222.5 120740.0 9287.5 120875.0 ;
      RECT  9362.5 120467.5 9427.5 120602.5 ;
      RECT  10357.5 120572.5 10222.5 120637.5 ;
      RECT  9907.5 121710.0 9972.5 121525.0 ;
      RECT  9907.5 122870.0 9972.5 122685.0 ;
      RECT  9547.5 122752.5 9612.5 122902.5 ;
      RECT  9547.5 121867.5 9612.5 121492.5 ;
      RECT  9737.5 122752.5 9802.5 121867.5 ;
      RECT  9547.5 121867.5 9612.5 121732.5 ;
      RECT  9737.5 121867.5 9802.5 121732.5 ;
      RECT  9737.5 121867.5 9802.5 121732.5 ;
      RECT  9547.5 121867.5 9612.5 121732.5 ;
      RECT  9547.5 122752.5 9612.5 122617.5 ;
      RECT  9737.5 122752.5 9802.5 122617.5 ;
      RECT  9737.5 122752.5 9802.5 122617.5 ;
      RECT  9547.5 122752.5 9612.5 122617.5 ;
      RECT  9907.5 121777.5 9972.5 121642.5 ;
      RECT  9907.5 122752.5 9972.5 122617.5 ;
      RECT  9605.0 122310.0 9670.0 122175.0 ;
      RECT  9605.0 122310.0 9670.0 122175.0 ;
      RECT  9770.0 122275.0 9835.0 122210.0 ;
      RECT  9480.0 121557.5 10040.0 121492.5 ;
      RECT  9480.0 122902.5 10040.0 122837.5 ;
      RECT  10107.5 122707.5 10172.5 122902.5 ;
      RECT  10107.5 121867.5 10172.5 121492.5 ;
      RECT  10487.5 121867.5 10552.5 121492.5 ;
      RECT  10657.5 121710.0 10722.5 121525.0 ;
      RECT  10657.5 122870.0 10722.5 122685.0 ;
      RECT  10107.5 121867.5 10172.5 121732.5 ;
      RECT  10297.5 121867.5 10362.5 121732.5 ;
      RECT  10297.5 121867.5 10362.5 121732.5 ;
      RECT  10107.5 121867.5 10172.5 121732.5 ;
      RECT  10297.5 121867.5 10362.5 121732.5 ;
      RECT  10487.5 121867.5 10552.5 121732.5 ;
      RECT  10487.5 121867.5 10552.5 121732.5 ;
      RECT  10297.5 121867.5 10362.5 121732.5 ;
      RECT  10107.5 122707.5 10172.5 122572.5 ;
      RECT  10297.5 122707.5 10362.5 122572.5 ;
      RECT  10297.5 122707.5 10362.5 122572.5 ;
      RECT  10107.5 122707.5 10172.5 122572.5 ;
      RECT  10297.5 122707.5 10362.5 122572.5 ;
      RECT  10487.5 122707.5 10552.5 122572.5 ;
      RECT  10487.5 122707.5 10552.5 122572.5 ;
      RECT  10297.5 122707.5 10362.5 122572.5 ;
      RECT  10657.5 121777.5 10722.5 121642.5 ;
      RECT  10657.5 122752.5 10722.5 122617.5 ;
      RECT  10492.5 122477.5 10357.5 122412.5 ;
      RECT  10235.0 122262.5 10100.0 122197.5 ;
      RECT  10297.5 121867.5 10362.5 121732.5 ;
      RECT  10487.5 122707.5 10552.5 122572.5 ;
      RECT  10587.5 122262.5 10452.5 122197.5 ;
      RECT  10100.0 122262.5 10235.0 122197.5 ;
      RECT  10357.5 122477.5 10492.5 122412.5 ;
      RECT  10452.5 122262.5 10587.5 122197.5 ;
      RECT  10040.0 121557.5 10960.0 121492.5 ;
      RECT  10040.0 122902.5 10960.0 122837.5 ;
      RECT  11387.5 121710.0 11452.5 121525.0 ;
      RECT  11387.5 122870.0 11452.5 122685.0 ;
      RECT  11027.5 122752.5 11092.5 122902.5 ;
      RECT  11027.5 121867.5 11092.5 121492.5 ;
      RECT  11217.5 122752.5 11282.5 121867.5 ;
      RECT  11027.5 121867.5 11092.5 121732.5 ;
      RECT  11217.5 121867.5 11282.5 121732.5 ;
      RECT  11217.5 121867.5 11282.5 121732.5 ;
      RECT  11027.5 121867.5 11092.5 121732.5 ;
      RECT  11027.5 122752.5 11092.5 122617.5 ;
      RECT  11217.5 122752.5 11282.5 122617.5 ;
      RECT  11217.5 122752.5 11282.5 122617.5 ;
      RECT  11027.5 122752.5 11092.5 122617.5 ;
      RECT  11387.5 121777.5 11452.5 121642.5 ;
      RECT  11387.5 122752.5 11452.5 122617.5 ;
      RECT  11085.0 122310.0 11150.0 122175.0 ;
      RECT  11085.0 122310.0 11150.0 122175.0 ;
      RECT  11250.0 122275.0 11315.0 122210.0 ;
      RECT  10960.0 121557.5 11520.0 121492.5 ;
      RECT  10960.0 122902.5 11520.0 122837.5 ;
      RECT  9222.5 122175.0 9287.5 122310.0 ;
      RECT  9362.5 122447.5 9427.5 122582.5 ;
      RECT  10357.5 122412.5 10222.5 122477.5 ;
      RECT  9907.5 124030.0 9972.5 124215.0 ;
      RECT  9907.5 122870.0 9972.5 123055.0 ;
      RECT  9547.5 122987.5 9612.5 122837.5 ;
      RECT  9547.5 123872.5 9612.5 124247.5 ;
      RECT  9737.5 122987.5 9802.5 123872.5 ;
      RECT  9547.5 123872.5 9612.5 124007.5 ;
      RECT  9737.5 123872.5 9802.5 124007.5 ;
      RECT  9737.5 123872.5 9802.5 124007.5 ;
      RECT  9547.5 123872.5 9612.5 124007.5 ;
      RECT  9547.5 122987.5 9612.5 123122.5 ;
      RECT  9737.5 122987.5 9802.5 123122.5 ;
      RECT  9737.5 122987.5 9802.5 123122.5 ;
      RECT  9547.5 122987.5 9612.5 123122.5 ;
      RECT  9907.5 123962.5 9972.5 124097.5 ;
      RECT  9907.5 122987.5 9972.5 123122.5 ;
      RECT  9605.0 123430.0 9670.0 123565.0 ;
      RECT  9605.0 123430.0 9670.0 123565.0 ;
      RECT  9770.0 123465.0 9835.0 123530.0 ;
      RECT  9480.0 124182.5 10040.0 124247.5 ;
      RECT  9480.0 122837.5 10040.0 122902.5 ;
      RECT  10107.5 123032.5 10172.5 122837.5 ;
      RECT  10107.5 123872.5 10172.5 124247.5 ;
      RECT  10487.5 123872.5 10552.5 124247.5 ;
      RECT  10657.5 124030.0 10722.5 124215.0 ;
      RECT  10657.5 122870.0 10722.5 123055.0 ;
      RECT  10107.5 123872.5 10172.5 124007.5 ;
      RECT  10297.5 123872.5 10362.5 124007.5 ;
      RECT  10297.5 123872.5 10362.5 124007.5 ;
      RECT  10107.5 123872.5 10172.5 124007.5 ;
      RECT  10297.5 123872.5 10362.5 124007.5 ;
      RECT  10487.5 123872.5 10552.5 124007.5 ;
      RECT  10487.5 123872.5 10552.5 124007.5 ;
      RECT  10297.5 123872.5 10362.5 124007.5 ;
      RECT  10107.5 123032.5 10172.5 123167.5 ;
      RECT  10297.5 123032.5 10362.5 123167.5 ;
      RECT  10297.5 123032.5 10362.5 123167.5 ;
      RECT  10107.5 123032.5 10172.5 123167.5 ;
      RECT  10297.5 123032.5 10362.5 123167.5 ;
      RECT  10487.5 123032.5 10552.5 123167.5 ;
      RECT  10487.5 123032.5 10552.5 123167.5 ;
      RECT  10297.5 123032.5 10362.5 123167.5 ;
      RECT  10657.5 123962.5 10722.5 124097.5 ;
      RECT  10657.5 122987.5 10722.5 123122.5 ;
      RECT  10492.5 123262.5 10357.5 123327.5 ;
      RECT  10235.0 123477.5 10100.0 123542.5 ;
      RECT  10297.5 123872.5 10362.5 124007.5 ;
      RECT  10487.5 123032.5 10552.5 123167.5 ;
      RECT  10587.5 123477.5 10452.5 123542.5 ;
      RECT  10100.0 123477.5 10235.0 123542.5 ;
      RECT  10357.5 123262.5 10492.5 123327.5 ;
      RECT  10452.5 123477.5 10587.5 123542.5 ;
      RECT  10040.0 124182.5 10960.0 124247.5 ;
      RECT  10040.0 122837.5 10960.0 122902.5 ;
      RECT  11387.5 124030.0 11452.5 124215.0 ;
      RECT  11387.5 122870.0 11452.5 123055.0 ;
      RECT  11027.5 122987.5 11092.5 122837.5 ;
      RECT  11027.5 123872.5 11092.5 124247.5 ;
      RECT  11217.5 122987.5 11282.5 123872.5 ;
      RECT  11027.5 123872.5 11092.5 124007.5 ;
      RECT  11217.5 123872.5 11282.5 124007.5 ;
      RECT  11217.5 123872.5 11282.5 124007.5 ;
      RECT  11027.5 123872.5 11092.5 124007.5 ;
      RECT  11027.5 122987.5 11092.5 123122.5 ;
      RECT  11217.5 122987.5 11282.5 123122.5 ;
      RECT  11217.5 122987.5 11282.5 123122.5 ;
      RECT  11027.5 122987.5 11092.5 123122.5 ;
      RECT  11387.5 123962.5 11452.5 124097.5 ;
      RECT  11387.5 122987.5 11452.5 123122.5 ;
      RECT  11085.0 123430.0 11150.0 123565.0 ;
      RECT  11085.0 123430.0 11150.0 123565.0 ;
      RECT  11250.0 123465.0 11315.0 123530.0 ;
      RECT  10960.0 124182.5 11520.0 124247.5 ;
      RECT  10960.0 122837.5 11520.0 122902.5 ;
      RECT  9222.5 123430.0 9287.5 123565.0 ;
      RECT  9362.5 123157.5 9427.5 123292.5 ;
      RECT  10357.5 123262.5 10222.5 123327.5 ;
      RECT  9907.5 124400.0 9972.5 124215.0 ;
      RECT  9907.5 125560.0 9972.5 125375.0 ;
      RECT  9547.5 125442.5 9612.5 125592.5 ;
      RECT  9547.5 124557.5 9612.5 124182.5 ;
      RECT  9737.5 125442.5 9802.5 124557.5 ;
      RECT  9547.5 124557.5 9612.5 124422.5 ;
      RECT  9737.5 124557.5 9802.5 124422.5 ;
      RECT  9737.5 124557.5 9802.5 124422.5 ;
      RECT  9547.5 124557.5 9612.5 124422.5 ;
      RECT  9547.5 125442.5 9612.5 125307.5 ;
      RECT  9737.5 125442.5 9802.5 125307.5 ;
      RECT  9737.5 125442.5 9802.5 125307.5 ;
      RECT  9547.5 125442.5 9612.5 125307.5 ;
      RECT  9907.5 124467.5 9972.5 124332.5 ;
      RECT  9907.5 125442.5 9972.5 125307.5 ;
      RECT  9605.0 125000.0 9670.0 124865.0 ;
      RECT  9605.0 125000.0 9670.0 124865.0 ;
      RECT  9770.0 124965.0 9835.0 124900.0 ;
      RECT  9480.0 124247.5 10040.0 124182.5 ;
      RECT  9480.0 125592.5 10040.0 125527.5 ;
      RECT  10107.5 125397.5 10172.5 125592.5 ;
      RECT  10107.5 124557.5 10172.5 124182.5 ;
      RECT  10487.5 124557.5 10552.5 124182.5 ;
      RECT  10657.5 124400.0 10722.5 124215.0 ;
      RECT  10657.5 125560.0 10722.5 125375.0 ;
      RECT  10107.5 124557.5 10172.5 124422.5 ;
      RECT  10297.5 124557.5 10362.5 124422.5 ;
      RECT  10297.5 124557.5 10362.5 124422.5 ;
      RECT  10107.5 124557.5 10172.5 124422.5 ;
      RECT  10297.5 124557.5 10362.5 124422.5 ;
      RECT  10487.5 124557.5 10552.5 124422.5 ;
      RECT  10487.5 124557.5 10552.5 124422.5 ;
      RECT  10297.5 124557.5 10362.5 124422.5 ;
      RECT  10107.5 125397.5 10172.5 125262.5 ;
      RECT  10297.5 125397.5 10362.5 125262.5 ;
      RECT  10297.5 125397.5 10362.5 125262.5 ;
      RECT  10107.5 125397.5 10172.5 125262.5 ;
      RECT  10297.5 125397.5 10362.5 125262.5 ;
      RECT  10487.5 125397.5 10552.5 125262.5 ;
      RECT  10487.5 125397.5 10552.5 125262.5 ;
      RECT  10297.5 125397.5 10362.5 125262.5 ;
      RECT  10657.5 124467.5 10722.5 124332.5 ;
      RECT  10657.5 125442.5 10722.5 125307.5 ;
      RECT  10492.5 125167.5 10357.5 125102.5 ;
      RECT  10235.0 124952.5 10100.0 124887.5 ;
      RECT  10297.5 124557.5 10362.5 124422.5 ;
      RECT  10487.5 125397.5 10552.5 125262.5 ;
      RECT  10587.5 124952.5 10452.5 124887.5 ;
      RECT  10100.0 124952.5 10235.0 124887.5 ;
      RECT  10357.5 125167.5 10492.5 125102.5 ;
      RECT  10452.5 124952.5 10587.5 124887.5 ;
      RECT  10040.0 124247.5 10960.0 124182.5 ;
      RECT  10040.0 125592.5 10960.0 125527.5 ;
      RECT  11387.5 124400.0 11452.5 124215.0 ;
      RECT  11387.5 125560.0 11452.5 125375.0 ;
      RECT  11027.5 125442.5 11092.5 125592.5 ;
      RECT  11027.5 124557.5 11092.5 124182.5 ;
      RECT  11217.5 125442.5 11282.5 124557.5 ;
      RECT  11027.5 124557.5 11092.5 124422.5 ;
      RECT  11217.5 124557.5 11282.5 124422.5 ;
      RECT  11217.5 124557.5 11282.5 124422.5 ;
      RECT  11027.5 124557.5 11092.5 124422.5 ;
      RECT  11027.5 125442.5 11092.5 125307.5 ;
      RECT  11217.5 125442.5 11282.5 125307.5 ;
      RECT  11217.5 125442.5 11282.5 125307.5 ;
      RECT  11027.5 125442.5 11092.5 125307.5 ;
      RECT  11387.5 124467.5 11452.5 124332.5 ;
      RECT  11387.5 125442.5 11452.5 125307.5 ;
      RECT  11085.0 125000.0 11150.0 124865.0 ;
      RECT  11085.0 125000.0 11150.0 124865.0 ;
      RECT  11250.0 124965.0 11315.0 124900.0 ;
      RECT  10960.0 124247.5 11520.0 124182.5 ;
      RECT  10960.0 125592.5 11520.0 125527.5 ;
      RECT  9222.5 124865.0 9287.5 125000.0 ;
      RECT  9362.5 125137.5 9427.5 125272.5 ;
      RECT  10357.5 125102.5 10222.5 125167.5 ;
      RECT  9907.5 126720.0 9972.5 126905.0 ;
      RECT  9907.5 125560.0 9972.5 125745.0 ;
      RECT  9547.5 125677.5 9612.5 125527.5 ;
      RECT  9547.5 126562.5 9612.5 126937.5 ;
      RECT  9737.5 125677.5 9802.5 126562.5 ;
      RECT  9547.5 126562.5 9612.5 126697.5 ;
      RECT  9737.5 126562.5 9802.5 126697.5 ;
      RECT  9737.5 126562.5 9802.5 126697.5 ;
      RECT  9547.5 126562.5 9612.5 126697.5 ;
      RECT  9547.5 125677.5 9612.5 125812.5 ;
      RECT  9737.5 125677.5 9802.5 125812.5 ;
      RECT  9737.5 125677.5 9802.5 125812.5 ;
      RECT  9547.5 125677.5 9612.5 125812.5 ;
      RECT  9907.5 126652.5 9972.5 126787.5 ;
      RECT  9907.5 125677.5 9972.5 125812.5 ;
      RECT  9605.0 126120.0 9670.0 126255.0 ;
      RECT  9605.0 126120.0 9670.0 126255.0 ;
      RECT  9770.0 126155.0 9835.0 126220.0 ;
      RECT  9480.0 126872.5 10040.0 126937.5 ;
      RECT  9480.0 125527.5 10040.0 125592.5 ;
      RECT  10107.5 125722.5 10172.5 125527.5 ;
      RECT  10107.5 126562.5 10172.5 126937.5 ;
      RECT  10487.5 126562.5 10552.5 126937.5 ;
      RECT  10657.5 126720.0 10722.5 126905.0 ;
      RECT  10657.5 125560.0 10722.5 125745.0 ;
      RECT  10107.5 126562.5 10172.5 126697.5 ;
      RECT  10297.5 126562.5 10362.5 126697.5 ;
      RECT  10297.5 126562.5 10362.5 126697.5 ;
      RECT  10107.5 126562.5 10172.5 126697.5 ;
      RECT  10297.5 126562.5 10362.5 126697.5 ;
      RECT  10487.5 126562.5 10552.5 126697.5 ;
      RECT  10487.5 126562.5 10552.5 126697.5 ;
      RECT  10297.5 126562.5 10362.5 126697.5 ;
      RECT  10107.5 125722.5 10172.5 125857.5 ;
      RECT  10297.5 125722.5 10362.5 125857.5 ;
      RECT  10297.5 125722.5 10362.5 125857.5 ;
      RECT  10107.5 125722.5 10172.5 125857.5 ;
      RECT  10297.5 125722.5 10362.5 125857.5 ;
      RECT  10487.5 125722.5 10552.5 125857.5 ;
      RECT  10487.5 125722.5 10552.5 125857.5 ;
      RECT  10297.5 125722.5 10362.5 125857.5 ;
      RECT  10657.5 126652.5 10722.5 126787.5 ;
      RECT  10657.5 125677.5 10722.5 125812.5 ;
      RECT  10492.5 125952.5 10357.5 126017.5 ;
      RECT  10235.0 126167.5 10100.0 126232.5 ;
      RECT  10297.5 126562.5 10362.5 126697.5 ;
      RECT  10487.5 125722.5 10552.5 125857.5 ;
      RECT  10587.5 126167.5 10452.5 126232.5 ;
      RECT  10100.0 126167.5 10235.0 126232.5 ;
      RECT  10357.5 125952.5 10492.5 126017.5 ;
      RECT  10452.5 126167.5 10587.5 126232.5 ;
      RECT  10040.0 126872.5 10960.0 126937.5 ;
      RECT  10040.0 125527.5 10960.0 125592.5 ;
      RECT  11387.5 126720.0 11452.5 126905.0 ;
      RECT  11387.5 125560.0 11452.5 125745.0 ;
      RECT  11027.5 125677.5 11092.5 125527.5 ;
      RECT  11027.5 126562.5 11092.5 126937.5 ;
      RECT  11217.5 125677.5 11282.5 126562.5 ;
      RECT  11027.5 126562.5 11092.5 126697.5 ;
      RECT  11217.5 126562.5 11282.5 126697.5 ;
      RECT  11217.5 126562.5 11282.5 126697.5 ;
      RECT  11027.5 126562.5 11092.5 126697.5 ;
      RECT  11027.5 125677.5 11092.5 125812.5 ;
      RECT  11217.5 125677.5 11282.5 125812.5 ;
      RECT  11217.5 125677.5 11282.5 125812.5 ;
      RECT  11027.5 125677.5 11092.5 125812.5 ;
      RECT  11387.5 126652.5 11452.5 126787.5 ;
      RECT  11387.5 125677.5 11452.5 125812.5 ;
      RECT  11085.0 126120.0 11150.0 126255.0 ;
      RECT  11085.0 126120.0 11150.0 126255.0 ;
      RECT  11250.0 126155.0 11315.0 126220.0 ;
      RECT  10960.0 126872.5 11520.0 126937.5 ;
      RECT  10960.0 125527.5 11520.0 125592.5 ;
      RECT  9222.5 126120.0 9287.5 126255.0 ;
      RECT  9362.5 125847.5 9427.5 125982.5 ;
      RECT  10357.5 125952.5 10222.5 126017.5 ;
      RECT  9907.5 127090.0 9972.5 126905.0 ;
      RECT  9907.5 128250.0 9972.5 128065.0 ;
      RECT  9547.5 128132.5 9612.5 128282.5 ;
      RECT  9547.5 127247.5 9612.5 126872.5 ;
      RECT  9737.5 128132.5 9802.5 127247.5 ;
      RECT  9547.5 127247.5 9612.5 127112.5 ;
      RECT  9737.5 127247.5 9802.5 127112.5 ;
      RECT  9737.5 127247.5 9802.5 127112.5 ;
      RECT  9547.5 127247.5 9612.5 127112.5 ;
      RECT  9547.5 128132.5 9612.5 127997.5 ;
      RECT  9737.5 128132.5 9802.5 127997.5 ;
      RECT  9737.5 128132.5 9802.5 127997.5 ;
      RECT  9547.5 128132.5 9612.5 127997.5 ;
      RECT  9907.5 127157.5 9972.5 127022.5 ;
      RECT  9907.5 128132.5 9972.5 127997.5 ;
      RECT  9605.0 127690.0 9670.0 127555.0 ;
      RECT  9605.0 127690.0 9670.0 127555.0 ;
      RECT  9770.0 127655.0 9835.0 127590.0 ;
      RECT  9480.0 126937.5 10040.0 126872.5 ;
      RECT  9480.0 128282.5 10040.0 128217.5 ;
      RECT  10107.5 128087.5 10172.5 128282.5 ;
      RECT  10107.5 127247.5 10172.5 126872.5 ;
      RECT  10487.5 127247.5 10552.5 126872.5 ;
      RECT  10657.5 127090.0 10722.5 126905.0 ;
      RECT  10657.5 128250.0 10722.5 128065.0 ;
      RECT  10107.5 127247.5 10172.5 127112.5 ;
      RECT  10297.5 127247.5 10362.5 127112.5 ;
      RECT  10297.5 127247.5 10362.5 127112.5 ;
      RECT  10107.5 127247.5 10172.5 127112.5 ;
      RECT  10297.5 127247.5 10362.5 127112.5 ;
      RECT  10487.5 127247.5 10552.5 127112.5 ;
      RECT  10487.5 127247.5 10552.5 127112.5 ;
      RECT  10297.5 127247.5 10362.5 127112.5 ;
      RECT  10107.5 128087.5 10172.5 127952.5 ;
      RECT  10297.5 128087.5 10362.5 127952.5 ;
      RECT  10297.5 128087.5 10362.5 127952.5 ;
      RECT  10107.5 128087.5 10172.5 127952.5 ;
      RECT  10297.5 128087.5 10362.5 127952.5 ;
      RECT  10487.5 128087.5 10552.5 127952.5 ;
      RECT  10487.5 128087.5 10552.5 127952.5 ;
      RECT  10297.5 128087.5 10362.5 127952.5 ;
      RECT  10657.5 127157.5 10722.5 127022.5 ;
      RECT  10657.5 128132.5 10722.5 127997.5 ;
      RECT  10492.5 127857.5 10357.5 127792.5 ;
      RECT  10235.0 127642.5 10100.0 127577.5 ;
      RECT  10297.5 127247.5 10362.5 127112.5 ;
      RECT  10487.5 128087.5 10552.5 127952.5 ;
      RECT  10587.5 127642.5 10452.5 127577.5 ;
      RECT  10100.0 127642.5 10235.0 127577.5 ;
      RECT  10357.5 127857.5 10492.5 127792.5 ;
      RECT  10452.5 127642.5 10587.5 127577.5 ;
      RECT  10040.0 126937.5 10960.0 126872.5 ;
      RECT  10040.0 128282.5 10960.0 128217.5 ;
      RECT  11387.5 127090.0 11452.5 126905.0 ;
      RECT  11387.5 128250.0 11452.5 128065.0 ;
      RECT  11027.5 128132.5 11092.5 128282.5 ;
      RECT  11027.5 127247.5 11092.5 126872.5 ;
      RECT  11217.5 128132.5 11282.5 127247.5 ;
      RECT  11027.5 127247.5 11092.5 127112.5 ;
      RECT  11217.5 127247.5 11282.5 127112.5 ;
      RECT  11217.5 127247.5 11282.5 127112.5 ;
      RECT  11027.5 127247.5 11092.5 127112.5 ;
      RECT  11027.5 128132.5 11092.5 127997.5 ;
      RECT  11217.5 128132.5 11282.5 127997.5 ;
      RECT  11217.5 128132.5 11282.5 127997.5 ;
      RECT  11027.5 128132.5 11092.5 127997.5 ;
      RECT  11387.5 127157.5 11452.5 127022.5 ;
      RECT  11387.5 128132.5 11452.5 127997.5 ;
      RECT  11085.0 127690.0 11150.0 127555.0 ;
      RECT  11085.0 127690.0 11150.0 127555.0 ;
      RECT  11250.0 127655.0 11315.0 127590.0 ;
      RECT  10960.0 126937.5 11520.0 126872.5 ;
      RECT  10960.0 128282.5 11520.0 128217.5 ;
      RECT  9222.5 127555.0 9287.5 127690.0 ;
      RECT  9362.5 127827.5 9427.5 127962.5 ;
      RECT  10357.5 127792.5 10222.5 127857.5 ;
      RECT  9907.5 129410.0 9972.5 129595.0 ;
      RECT  9907.5 128250.0 9972.5 128435.0 ;
      RECT  9547.5 128367.5 9612.5 128217.5 ;
      RECT  9547.5 129252.5 9612.5 129627.5 ;
      RECT  9737.5 128367.5 9802.5 129252.5 ;
      RECT  9547.5 129252.5 9612.5 129387.5 ;
      RECT  9737.5 129252.5 9802.5 129387.5 ;
      RECT  9737.5 129252.5 9802.5 129387.5 ;
      RECT  9547.5 129252.5 9612.5 129387.5 ;
      RECT  9547.5 128367.5 9612.5 128502.5 ;
      RECT  9737.5 128367.5 9802.5 128502.5 ;
      RECT  9737.5 128367.5 9802.5 128502.5 ;
      RECT  9547.5 128367.5 9612.5 128502.5 ;
      RECT  9907.5 129342.5 9972.5 129477.5 ;
      RECT  9907.5 128367.5 9972.5 128502.5 ;
      RECT  9605.0 128810.0 9670.0 128945.0 ;
      RECT  9605.0 128810.0 9670.0 128945.0 ;
      RECT  9770.0 128845.0 9835.0 128910.0 ;
      RECT  9480.0 129562.5 10040.0 129627.5 ;
      RECT  9480.0 128217.5 10040.0 128282.5 ;
      RECT  10107.5 128412.5 10172.5 128217.5 ;
      RECT  10107.5 129252.5 10172.5 129627.5 ;
      RECT  10487.5 129252.5 10552.5 129627.5 ;
      RECT  10657.5 129410.0 10722.5 129595.0 ;
      RECT  10657.5 128250.0 10722.5 128435.0 ;
      RECT  10107.5 129252.5 10172.5 129387.5 ;
      RECT  10297.5 129252.5 10362.5 129387.5 ;
      RECT  10297.5 129252.5 10362.5 129387.5 ;
      RECT  10107.5 129252.5 10172.5 129387.5 ;
      RECT  10297.5 129252.5 10362.5 129387.5 ;
      RECT  10487.5 129252.5 10552.5 129387.5 ;
      RECT  10487.5 129252.5 10552.5 129387.5 ;
      RECT  10297.5 129252.5 10362.5 129387.5 ;
      RECT  10107.5 128412.5 10172.5 128547.5 ;
      RECT  10297.5 128412.5 10362.5 128547.5 ;
      RECT  10297.5 128412.5 10362.5 128547.5 ;
      RECT  10107.5 128412.5 10172.5 128547.5 ;
      RECT  10297.5 128412.5 10362.5 128547.5 ;
      RECT  10487.5 128412.5 10552.5 128547.5 ;
      RECT  10487.5 128412.5 10552.5 128547.5 ;
      RECT  10297.5 128412.5 10362.5 128547.5 ;
      RECT  10657.5 129342.5 10722.5 129477.5 ;
      RECT  10657.5 128367.5 10722.5 128502.5 ;
      RECT  10492.5 128642.5 10357.5 128707.5 ;
      RECT  10235.0 128857.5 10100.0 128922.5 ;
      RECT  10297.5 129252.5 10362.5 129387.5 ;
      RECT  10487.5 128412.5 10552.5 128547.5 ;
      RECT  10587.5 128857.5 10452.5 128922.5 ;
      RECT  10100.0 128857.5 10235.0 128922.5 ;
      RECT  10357.5 128642.5 10492.5 128707.5 ;
      RECT  10452.5 128857.5 10587.5 128922.5 ;
      RECT  10040.0 129562.5 10960.0 129627.5 ;
      RECT  10040.0 128217.5 10960.0 128282.5 ;
      RECT  11387.5 129410.0 11452.5 129595.0 ;
      RECT  11387.5 128250.0 11452.5 128435.0 ;
      RECT  11027.5 128367.5 11092.5 128217.5 ;
      RECT  11027.5 129252.5 11092.5 129627.5 ;
      RECT  11217.5 128367.5 11282.5 129252.5 ;
      RECT  11027.5 129252.5 11092.5 129387.5 ;
      RECT  11217.5 129252.5 11282.5 129387.5 ;
      RECT  11217.5 129252.5 11282.5 129387.5 ;
      RECT  11027.5 129252.5 11092.5 129387.5 ;
      RECT  11027.5 128367.5 11092.5 128502.5 ;
      RECT  11217.5 128367.5 11282.5 128502.5 ;
      RECT  11217.5 128367.5 11282.5 128502.5 ;
      RECT  11027.5 128367.5 11092.5 128502.5 ;
      RECT  11387.5 129342.5 11452.5 129477.5 ;
      RECT  11387.5 128367.5 11452.5 128502.5 ;
      RECT  11085.0 128810.0 11150.0 128945.0 ;
      RECT  11085.0 128810.0 11150.0 128945.0 ;
      RECT  11250.0 128845.0 11315.0 128910.0 ;
      RECT  10960.0 129562.5 11520.0 129627.5 ;
      RECT  10960.0 128217.5 11520.0 128282.5 ;
      RECT  9222.5 128810.0 9287.5 128945.0 ;
      RECT  9362.5 128537.5 9427.5 128672.5 ;
      RECT  10357.5 128642.5 10222.5 128707.5 ;
      RECT  9907.5 129780.0 9972.5 129595.0 ;
      RECT  9907.5 130940.0 9972.5 130755.0 ;
      RECT  9547.5 130822.5 9612.5 130972.5 ;
      RECT  9547.5 129937.5 9612.5 129562.5 ;
      RECT  9737.5 130822.5 9802.5 129937.5 ;
      RECT  9547.5 129937.5 9612.5 129802.5 ;
      RECT  9737.5 129937.5 9802.5 129802.5 ;
      RECT  9737.5 129937.5 9802.5 129802.5 ;
      RECT  9547.5 129937.5 9612.5 129802.5 ;
      RECT  9547.5 130822.5 9612.5 130687.5 ;
      RECT  9737.5 130822.5 9802.5 130687.5 ;
      RECT  9737.5 130822.5 9802.5 130687.5 ;
      RECT  9547.5 130822.5 9612.5 130687.5 ;
      RECT  9907.5 129847.5 9972.5 129712.5 ;
      RECT  9907.5 130822.5 9972.5 130687.5 ;
      RECT  9605.0 130380.0 9670.0 130245.0 ;
      RECT  9605.0 130380.0 9670.0 130245.0 ;
      RECT  9770.0 130345.0 9835.0 130280.0 ;
      RECT  9480.0 129627.5 10040.0 129562.5 ;
      RECT  9480.0 130972.5 10040.0 130907.5 ;
      RECT  10107.5 130777.5 10172.5 130972.5 ;
      RECT  10107.5 129937.5 10172.5 129562.5 ;
      RECT  10487.5 129937.5 10552.5 129562.5 ;
      RECT  10657.5 129780.0 10722.5 129595.0 ;
      RECT  10657.5 130940.0 10722.5 130755.0 ;
      RECT  10107.5 129937.5 10172.5 129802.5 ;
      RECT  10297.5 129937.5 10362.5 129802.5 ;
      RECT  10297.5 129937.5 10362.5 129802.5 ;
      RECT  10107.5 129937.5 10172.5 129802.5 ;
      RECT  10297.5 129937.5 10362.5 129802.5 ;
      RECT  10487.5 129937.5 10552.5 129802.5 ;
      RECT  10487.5 129937.5 10552.5 129802.5 ;
      RECT  10297.5 129937.5 10362.5 129802.5 ;
      RECT  10107.5 130777.5 10172.5 130642.5 ;
      RECT  10297.5 130777.5 10362.5 130642.5 ;
      RECT  10297.5 130777.5 10362.5 130642.5 ;
      RECT  10107.5 130777.5 10172.5 130642.5 ;
      RECT  10297.5 130777.5 10362.5 130642.5 ;
      RECT  10487.5 130777.5 10552.5 130642.5 ;
      RECT  10487.5 130777.5 10552.5 130642.5 ;
      RECT  10297.5 130777.5 10362.5 130642.5 ;
      RECT  10657.5 129847.5 10722.5 129712.5 ;
      RECT  10657.5 130822.5 10722.5 130687.5 ;
      RECT  10492.5 130547.5 10357.5 130482.5 ;
      RECT  10235.0 130332.5 10100.0 130267.5 ;
      RECT  10297.5 129937.5 10362.5 129802.5 ;
      RECT  10487.5 130777.5 10552.5 130642.5 ;
      RECT  10587.5 130332.5 10452.5 130267.5 ;
      RECT  10100.0 130332.5 10235.0 130267.5 ;
      RECT  10357.5 130547.5 10492.5 130482.5 ;
      RECT  10452.5 130332.5 10587.5 130267.5 ;
      RECT  10040.0 129627.5 10960.0 129562.5 ;
      RECT  10040.0 130972.5 10960.0 130907.5 ;
      RECT  11387.5 129780.0 11452.5 129595.0 ;
      RECT  11387.5 130940.0 11452.5 130755.0 ;
      RECT  11027.5 130822.5 11092.5 130972.5 ;
      RECT  11027.5 129937.5 11092.5 129562.5 ;
      RECT  11217.5 130822.5 11282.5 129937.5 ;
      RECT  11027.5 129937.5 11092.5 129802.5 ;
      RECT  11217.5 129937.5 11282.5 129802.5 ;
      RECT  11217.5 129937.5 11282.5 129802.5 ;
      RECT  11027.5 129937.5 11092.5 129802.5 ;
      RECT  11027.5 130822.5 11092.5 130687.5 ;
      RECT  11217.5 130822.5 11282.5 130687.5 ;
      RECT  11217.5 130822.5 11282.5 130687.5 ;
      RECT  11027.5 130822.5 11092.5 130687.5 ;
      RECT  11387.5 129847.5 11452.5 129712.5 ;
      RECT  11387.5 130822.5 11452.5 130687.5 ;
      RECT  11085.0 130380.0 11150.0 130245.0 ;
      RECT  11085.0 130380.0 11150.0 130245.0 ;
      RECT  11250.0 130345.0 11315.0 130280.0 ;
      RECT  10960.0 129627.5 11520.0 129562.5 ;
      RECT  10960.0 130972.5 11520.0 130907.5 ;
      RECT  9222.5 130245.0 9287.5 130380.0 ;
      RECT  9362.5 130517.5 9427.5 130652.5 ;
      RECT  10357.5 130482.5 10222.5 130547.5 ;
      RECT  9907.5 132100.0 9972.5 132285.0 ;
      RECT  9907.5 130940.0 9972.5 131125.0 ;
      RECT  9547.5 131057.5 9612.5 130907.5 ;
      RECT  9547.5 131942.5 9612.5 132317.5 ;
      RECT  9737.5 131057.5 9802.5 131942.5 ;
      RECT  9547.5 131942.5 9612.5 132077.5 ;
      RECT  9737.5 131942.5 9802.5 132077.5 ;
      RECT  9737.5 131942.5 9802.5 132077.5 ;
      RECT  9547.5 131942.5 9612.5 132077.5 ;
      RECT  9547.5 131057.5 9612.5 131192.5 ;
      RECT  9737.5 131057.5 9802.5 131192.5 ;
      RECT  9737.5 131057.5 9802.5 131192.5 ;
      RECT  9547.5 131057.5 9612.5 131192.5 ;
      RECT  9907.5 132032.5 9972.5 132167.5 ;
      RECT  9907.5 131057.5 9972.5 131192.5 ;
      RECT  9605.0 131500.0 9670.0 131635.0 ;
      RECT  9605.0 131500.0 9670.0 131635.0 ;
      RECT  9770.0 131535.0 9835.0 131600.0 ;
      RECT  9480.0 132252.5 10040.0 132317.5 ;
      RECT  9480.0 130907.5 10040.0 130972.5 ;
      RECT  10107.5 131102.5 10172.5 130907.5 ;
      RECT  10107.5 131942.5 10172.5 132317.5 ;
      RECT  10487.5 131942.5 10552.5 132317.5 ;
      RECT  10657.5 132100.0 10722.5 132285.0 ;
      RECT  10657.5 130940.0 10722.5 131125.0 ;
      RECT  10107.5 131942.5 10172.5 132077.5 ;
      RECT  10297.5 131942.5 10362.5 132077.5 ;
      RECT  10297.5 131942.5 10362.5 132077.5 ;
      RECT  10107.5 131942.5 10172.5 132077.5 ;
      RECT  10297.5 131942.5 10362.5 132077.5 ;
      RECT  10487.5 131942.5 10552.5 132077.5 ;
      RECT  10487.5 131942.5 10552.5 132077.5 ;
      RECT  10297.5 131942.5 10362.5 132077.5 ;
      RECT  10107.5 131102.5 10172.5 131237.5 ;
      RECT  10297.5 131102.5 10362.5 131237.5 ;
      RECT  10297.5 131102.5 10362.5 131237.5 ;
      RECT  10107.5 131102.5 10172.5 131237.5 ;
      RECT  10297.5 131102.5 10362.5 131237.5 ;
      RECT  10487.5 131102.5 10552.5 131237.5 ;
      RECT  10487.5 131102.5 10552.5 131237.5 ;
      RECT  10297.5 131102.5 10362.5 131237.5 ;
      RECT  10657.5 132032.5 10722.5 132167.5 ;
      RECT  10657.5 131057.5 10722.5 131192.5 ;
      RECT  10492.5 131332.5 10357.5 131397.5 ;
      RECT  10235.0 131547.5 10100.0 131612.5 ;
      RECT  10297.5 131942.5 10362.5 132077.5 ;
      RECT  10487.5 131102.5 10552.5 131237.5 ;
      RECT  10587.5 131547.5 10452.5 131612.5 ;
      RECT  10100.0 131547.5 10235.0 131612.5 ;
      RECT  10357.5 131332.5 10492.5 131397.5 ;
      RECT  10452.5 131547.5 10587.5 131612.5 ;
      RECT  10040.0 132252.5 10960.0 132317.5 ;
      RECT  10040.0 130907.5 10960.0 130972.5 ;
      RECT  11387.5 132100.0 11452.5 132285.0 ;
      RECT  11387.5 130940.0 11452.5 131125.0 ;
      RECT  11027.5 131057.5 11092.5 130907.5 ;
      RECT  11027.5 131942.5 11092.5 132317.5 ;
      RECT  11217.5 131057.5 11282.5 131942.5 ;
      RECT  11027.5 131942.5 11092.5 132077.5 ;
      RECT  11217.5 131942.5 11282.5 132077.5 ;
      RECT  11217.5 131942.5 11282.5 132077.5 ;
      RECT  11027.5 131942.5 11092.5 132077.5 ;
      RECT  11027.5 131057.5 11092.5 131192.5 ;
      RECT  11217.5 131057.5 11282.5 131192.5 ;
      RECT  11217.5 131057.5 11282.5 131192.5 ;
      RECT  11027.5 131057.5 11092.5 131192.5 ;
      RECT  11387.5 132032.5 11452.5 132167.5 ;
      RECT  11387.5 131057.5 11452.5 131192.5 ;
      RECT  11085.0 131500.0 11150.0 131635.0 ;
      RECT  11085.0 131500.0 11150.0 131635.0 ;
      RECT  11250.0 131535.0 11315.0 131600.0 ;
      RECT  10960.0 132252.5 11520.0 132317.5 ;
      RECT  10960.0 130907.5 11520.0 130972.5 ;
      RECT  9222.5 131500.0 9287.5 131635.0 ;
      RECT  9362.5 131227.5 9427.5 131362.5 ;
      RECT  10357.5 131332.5 10222.5 131397.5 ;
      RECT  9907.5 132470.0 9972.5 132285.0 ;
      RECT  9907.5 133630.0 9972.5 133445.0 ;
      RECT  9547.5 133512.5 9612.5 133662.5 ;
      RECT  9547.5 132627.5 9612.5 132252.5 ;
      RECT  9737.5 133512.5 9802.5 132627.5 ;
      RECT  9547.5 132627.5 9612.5 132492.5 ;
      RECT  9737.5 132627.5 9802.5 132492.5 ;
      RECT  9737.5 132627.5 9802.5 132492.5 ;
      RECT  9547.5 132627.5 9612.5 132492.5 ;
      RECT  9547.5 133512.5 9612.5 133377.5 ;
      RECT  9737.5 133512.5 9802.5 133377.5 ;
      RECT  9737.5 133512.5 9802.5 133377.5 ;
      RECT  9547.5 133512.5 9612.5 133377.5 ;
      RECT  9907.5 132537.5 9972.5 132402.5 ;
      RECT  9907.5 133512.5 9972.5 133377.5 ;
      RECT  9605.0 133070.0 9670.0 132935.0 ;
      RECT  9605.0 133070.0 9670.0 132935.0 ;
      RECT  9770.0 133035.0 9835.0 132970.0 ;
      RECT  9480.0 132317.5 10040.0 132252.5 ;
      RECT  9480.0 133662.5 10040.0 133597.5 ;
      RECT  10107.5 133467.5 10172.5 133662.5 ;
      RECT  10107.5 132627.5 10172.5 132252.5 ;
      RECT  10487.5 132627.5 10552.5 132252.5 ;
      RECT  10657.5 132470.0 10722.5 132285.0 ;
      RECT  10657.5 133630.0 10722.5 133445.0 ;
      RECT  10107.5 132627.5 10172.5 132492.5 ;
      RECT  10297.5 132627.5 10362.5 132492.5 ;
      RECT  10297.5 132627.5 10362.5 132492.5 ;
      RECT  10107.5 132627.5 10172.5 132492.5 ;
      RECT  10297.5 132627.5 10362.5 132492.5 ;
      RECT  10487.5 132627.5 10552.5 132492.5 ;
      RECT  10487.5 132627.5 10552.5 132492.5 ;
      RECT  10297.5 132627.5 10362.5 132492.5 ;
      RECT  10107.5 133467.5 10172.5 133332.5 ;
      RECT  10297.5 133467.5 10362.5 133332.5 ;
      RECT  10297.5 133467.5 10362.5 133332.5 ;
      RECT  10107.5 133467.5 10172.5 133332.5 ;
      RECT  10297.5 133467.5 10362.5 133332.5 ;
      RECT  10487.5 133467.5 10552.5 133332.5 ;
      RECT  10487.5 133467.5 10552.5 133332.5 ;
      RECT  10297.5 133467.5 10362.5 133332.5 ;
      RECT  10657.5 132537.5 10722.5 132402.5 ;
      RECT  10657.5 133512.5 10722.5 133377.5 ;
      RECT  10492.5 133237.5 10357.5 133172.5 ;
      RECT  10235.0 133022.5 10100.0 132957.5 ;
      RECT  10297.5 132627.5 10362.5 132492.5 ;
      RECT  10487.5 133467.5 10552.5 133332.5 ;
      RECT  10587.5 133022.5 10452.5 132957.5 ;
      RECT  10100.0 133022.5 10235.0 132957.5 ;
      RECT  10357.5 133237.5 10492.5 133172.5 ;
      RECT  10452.5 133022.5 10587.5 132957.5 ;
      RECT  10040.0 132317.5 10960.0 132252.5 ;
      RECT  10040.0 133662.5 10960.0 133597.5 ;
      RECT  11387.5 132470.0 11452.5 132285.0 ;
      RECT  11387.5 133630.0 11452.5 133445.0 ;
      RECT  11027.5 133512.5 11092.5 133662.5 ;
      RECT  11027.5 132627.5 11092.5 132252.5 ;
      RECT  11217.5 133512.5 11282.5 132627.5 ;
      RECT  11027.5 132627.5 11092.5 132492.5 ;
      RECT  11217.5 132627.5 11282.5 132492.5 ;
      RECT  11217.5 132627.5 11282.5 132492.5 ;
      RECT  11027.5 132627.5 11092.5 132492.5 ;
      RECT  11027.5 133512.5 11092.5 133377.5 ;
      RECT  11217.5 133512.5 11282.5 133377.5 ;
      RECT  11217.5 133512.5 11282.5 133377.5 ;
      RECT  11027.5 133512.5 11092.5 133377.5 ;
      RECT  11387.5 132537.5 11452.5 132402.5 ;
      RECT  11387.5 133512.5 11452.5 133377.5 ;
      RECT  11085.0 133070.0 11150.0 132935.0 ;
      RECT  11085.0 133070.0 11150.0 132935.0 ;
      RECT  11250.0 133035.0 11315.0 132970.0 ;
      RECT  10960.0 132317.5 11520.0 132252.5 ;
      RECT  10960.0 133662.5 11520.0 133597.5 ;
      RECT  9222.5 132935.0 9287.5 133070.0 ;
      RECT  9362.5 133207.5 9427.5 133342.5 ;
      RECT  10357.5 133172.5 10222.5 133237.5 ;
      RECT  9907.5 134790.0 9972.5 134975.0 ;
      RECT  9907.5 133630.0 9972.5 133815.0 ;
      RECT  9547.5 133747.5 9612.5 133597.5 ;
      RECT  9547.5 134632.5 9612.5 135007.5 ;
      RECT  9737.5 133747.5 9802.5 134632.5 ;
      RECT  9547.5 134632.5 9612.5 134767.5 ;
      RECT  9737.5 134632.5 9802.5 134767.5 ;
      RECT  9737.5 134632.5 9802.5 134767.5 ;
      RECT  9547.5 134632.5 9612.5 134767.5 ;
      RECT  9547.5 133747.5 9612.5 133882.5 ;
      RECT  9737.5 133747.5 9802.5 133882.5 ;
      RECT  9737.5 133747.5 9802.5 133882.5 ;
      RECT  9547.5 133747.5 9612.5 133882.5 ;
      RECT  9907.5 134722.5 9972.5 134857.5 ;
      RECT  9907.5 133747.5 9972.5 133882.5 ;
      RECT  9605.0 134190.0 9670.0 134325.0 ;
      RECT  9605.0 134190.0 9670.0 134325.0 ;
      RECT  9770.0 134225.0 9835.0 134290.0 ;
      RECT  9480.0 134942.5 10040.0 135007.5 ;
      RECT  9480.0 133597.5 10040.0 133662.5 ;
      RECT  10107.5 133792.5 10172.5 133597.5 ;
      RECT  10107.5 134632.5 10172.5 135007.5 ;
      RECT  10487.5 134632.5 10552.5 135007.5 ;
      RECT  10657.5 134790.0 10722.5 134975.0 ;
      RECT  10657.5 133630.0 10722.5 133815.0 ;
      RECT  10107.5 134632.5 10172.5 134767.5 ;
      RECT  10297.5 134632.5 10362.5 134767.5 ;
      RECT  10297.5 134632.5 10362.5 134767.5 ;
      RECT  10107.5 134632.5 10172.5 134767.5 ;
      RECT  10297.5 134632.5 10362.5 134767.5 ;
      RECT  10487.5 134632.5 10552.5 134767.5 ;
      RECT  10487.5 134632.5 10552.5 134767.5 ;
      RECT  10297.5 134632.5 10362.5 134767.5 ;
      RECT  10107.5 133792.5 10172.5 133927.5 ;
      RECT  10297.5 133792.5 10362.5 133927.5 ;
      RECT  10297.5 133792.5 10362.5 133927.5 ;
      RECT  10107.5 133792.5 10172.5 133927.5 ;
      RECT  10297.5 133792.5 10362.5 133927.5 ;
      RECT  10487.5 133792.5 10552.5 133927.5 ;
      RECT  10487.5 133792.5 10552.5 133927.5 ;
      RECT  10297.5 133792.5 10362.5 133927.5 ;
      RECT  10657.5 134722.5 10722.5 134857.5 ;
      RECT  10657.5 133747.5 10722.5 133882.5 ;
      RECT  10492.5 134022.5 10357.5 134087.5 ;
      RECT  10235.0 134237.5 10100.0 134302.5 ;
      RECT  10297.5 134632.5 10362.5 134767.5 ;
      RECT  10487.5 133792.5 10552.5 133927.5 ;
      RECT  10587.5 134237.5 10452.5 134302.5 ;
      RECT  10100.0 134237.5 10235.0 134302.5 ;
      RECT  10357.5 134022.5 10492.5 134087.5 ;
      RECT  10452.5 134237.5 10587.5 134302.5 ;
      RECT  10040.0 134942.5 10960.0 135007.5 ;
      RECT  10040.0 133597.5 10960.0 133662.5 ;
      RECT  11387.5 134790.0 11452.5 134975.0 ;
      RECT  11387.5 133630.0 11452.5 133815.0 ;
      RECT  11027.5 133747.5 11092.5 133597.5 ;
      RECT  11027.5 134632.5 11092.5 135007.5 ;
      RECT  11217.5 133747.5 11282.5 134632.5 ;
      RECT  11027.5 134632.5 11092.5 134767.5 ;
      RECT  11217.5 134632.5 11282.5 134767.5 ;
      RECT  11217.5 134632.5 11282.5 134767.5 ;
      RECT  11027.5 134632.5 11092.5 134767.5 ;
      RECT  11027.5 133747.5 11092.5 133882.5 ;
      RECT  11217.5 133747.5 11282.5 133882.5 ;
      RECT  11217.5 133747.5 11282.5 133882.5 ;
      RECT  11027.5 133747.5 11092.5 133882.5 ;
      RECT  11387.5 134722.5 11452.5 134857.5 ;
      RECT  11387.5 133747.5 11452.5 133882.5 ;
      RECT  11085.0 134190.0 11150.0 134325.0 ;
      RECT  11085.0 134190.0 11150.0 134325.0 ;
      RECT  11250.0 134225.0 11315.0 134290.0 ;
      RECT  10960.0 134942.5 11520.0 135007.5 ;
      RECT  10960.0 133597.5 11520.0 133662.5 ;
      RECT  9222.5 134190.0 9287.5 134325.0 ;
      RECT  9362.5 133917.5 9427.5 134052.5 ;
      RECT  10357.5 134022.5 10222.5 134087.5 ;
      RECT  9907.5 135160.0 9972.5 134975.0 ;
      RECT  9907.5 136320.0 9972.5 136135.0 ;
      RECT  9547.5 136202.5 9612.5 136352.5 ;
      RECT  9547.5 135317.5 9612.5 134942.5 ;
      RECT  9737.5 136202.5 9802.5 135317.5 ;
      RECT  9547.5 135317.5 9612.5 135182.5 ;
      RECT  9737.5 135317.5 9802.5 135182.5 ;
      RECT  9737.5 135317.5 9802.5 135182.5 ;
      RECT  9547.5 135317.5 9612.5 135182.5 ;
      RECT  9547.5 136202.5 9612.5 136067.5 ;
      RECT  9737.5 136202.5 9802.5 136067.5 ;
      RECT  9737.5 136202.5 9802.5 136067.5 ;
      RECT  9547.5 136202.5 9612.5 136067.5 ;
      RECT  9907.5 135227.5 9972.5 135092.5 ;
      RECT  9907.5 136202.5 9972.5 136067.5 ;
      RECT  9605.0 135760.0 9670.0 135625.0 ;
      RECT  9605.0 135760.0 9670.0 135625.0 ;
      RECT  9770.0 135725.0 9835.0 135660.0 ;
      RECT  9480.0 135007.5 10040.0 134942.5 ;
      RECT  9480.0 136352.5 10040.0 136287.5 ;
      RECT  10107.5 136157.5 10172.5 136352.5 ;
      RECT  10107.5 135317.5 10172.5 134942.5 ;
      RECT  10487.5 135317.5 10552.5 134942.5 ;
      RECT  10657.5 135160.0 10722.5 134975.0 ;
      RECT  10657.5 136320.0 10722.5 136135.0 ;
      RECT  10107.5 135317.5 10172.5 135182.5 ;
      RECT  10297.5 135317.5 10362.5 135182.5 ;
      RECT  10297.5 135317.5 10362.5 135182.5 ;
      RECT  10107.5 135317.5 10172.5 135182.5 ;
      RECT  10297.5 135317.5 10362.5 135182.5 ;
      RECT  10487.5 135317.5 10552.5 135182.5 ;
      RECT  10487.5 135317.5 10552.5 135182.5 ;
      RECT  10297.5 135317.5 10362.5 135182.5 ;
      RECT  10107.5 136157.5 10172.5 136022.5 ;
      RECT  10297.5 136157.5 10362.5 136022.5 ;
      RECT  10297.5 136157.5 10362.5 136022.5 ;
      RECT  10107.5 136157.5 10172.5 136022.5 ;
      RECT  10297.5 136157.5 10362.5 136022.5 ;
      RECT  10487.5 136157.5 10552.5 136022.5 ;
      RECT  10487.5 136157.5 10552.5 136022.5 ;
      RECT  10297.5 136157.5 10362.5 136022.5 ;
      RECT  10657.5 135227.5 10722.5 135092.5 ;
      RECT  10657.5 136202.5 10722.5 136067.5 ;
      RECT  10492.5 135927.5 10357.5 135862.5 ;
      RECT  10235.0 135712.5 10100.0 135647.5 ;
      RECT  10297.5 135317.5 10362.5 135182.5 ;
      RECT  10487.5 136157.5 10552.5 136022.5 ;
      RECT  10587.5 135712.5 10452.5 135647.5 ;
      RECT  10100.0 135712.5 10235.0 135647.5 ;
      RECT  10357.5 135927.5 10492.5 135862.5 ;
      RECT  10452.5 135712.5 10587.5 135647.5 ;
      RECT  10040.0 135007.5 10960.0 134942.5 ;
      RECT  10040.0 136352.5 10960.0 136287.5 ;
      RECT  11387.5 135160.0 11452.5 134975.0 ;
      RECT  11387.5 136320.0 11452.5 136135.0 ;
      RECT  11027.5 136202.5 11092.5 136352.5 ;
      RECT  11027.5 135317.5 11092.5 134942.5 ;
      RECT  11217.5 136202.5 11282.5 135317.5 ;
      RECT  11027.5 135317.5 11092.5 135182.5 ;
      RECT  11217.5 135317.5 11282.5 135182.5 ;
      RECT  11217.5 135317.5 11282.5 135182.5 ;
      RECT  11027.5 135317.5 11092.5 135182.5 ;
      RECT  11027.5 136202.5 11092.5 136067.5 ;
      RECT  11217.5 136202.5 11282.5 136067.5 ;
      RECT  11217.5 136202.5 11282.5 136067.5 ;
      RECT  11027.5 136202.5 11092.5 136067.5 ;
      RECT  11387.5 135227.5 11452.5 135092.5 ;
      RECT  11387.5 136202.5 11452.5 136067.5 ;
      RECT  11085.0 135760.0 11150.0 135625.0 ;
      RECT  11085.0 135760.0 11150.0 135625.0 ;
      RECT  11250.0 135725.0 11315.0 135660.0 ;
      RECT  10960.0 135007.5 11520.0 134942.5 ;
      RECT  10960.0 136352.5 11520.0 136287.5 ;
      RECT  9222.5 135625.0 9287.5 135760.0 ;
      RECT  9362.5 135897.5 9427.5 136032.5 ;
      RECT  10357.5 135862.5 10222.5 135927.5 ;
      RECT  9907.5 137480.0 9972.5 137665.0 ;
      RECT  9907.5 136320.0 9972.5 136505.0 ;
      RECT  9547.5 136437.5 9612.5 136287.5 ;
      RECT  9547.5 137322.5 9612.5 137697.5 ;
      RECT  9737.5 136437.5 9802.5 137322.5 ;
      RECT  9547.5 137322.5 9612.5 137457.5 ;
      RECT  9737.5 137322.5 9802.5 137457.5 ;
      RECT  9737.5 137322.5 9802.5 137457.5 ;
      RECT  9547.5 137322.5 9612.5 137457.5 ;
      RECT  9547.5 136437.5 9612.5 136572.5 ;
      RECT  9737.5 136437.5 9802.5 136572.5 ;
      RECT  9737.5 136437.5 9802.5 136572.5 ;
      RECT  9547.5 136437.5 9612.5 136572.5 ;
      RECT  9907.5 137412.5 9972.5 137547.5 ;
      RECT  9907.5 136437.5 9972.5 136572.5 ;
      RECT  9605.0 136880.0 9670.0 137015.0 ;
      RECT  9605.0 136880.0 9670.0 137015.0 ;
      RECT  9770.0 136915.0 9835.0 136980.0 ;
      RECT  9480.0 137632.5 10040.0 137697.5 ;
      RECT  9480.0 136287.5 10040.0 136352.5 ;
      RECT  10107.5 136482.5 10172.5 136287.5 ;
      RECT  10107.5 137322.5 10172.5 137697.5 ;
      RECT  10487.5 137322.5 10552.5 137697.5 ;
      RECT  10657.5 137480.0 10722.5 137665.0 ;
      RECT  10657.5 136320.0 10722.5 136505.0 ;
      RECT  10107.5 137322.5 10172.5 137457.5 ;
      RECT  10297.5 137322.5 10362.5 137457.5 ;
      RECT  10297.5 137322.5 10362.5 137457.5 ;
      RECT  10107.5 137322.5 10172.5 137457.5 ;
      RECT  10297.5 137322.5 10362.5 137457.5 ;
      RECT  10487.5 137322.5 10552.5 137457.5 ;
      RECT  10487.5 137322.5 10552.5 137457.5 ;
      RECT  10297.5 137322.5 10362.5 137457.5 ;
      RECT  10107.5 136482.5 10172.5 136617.5 ;
      RECT  10297.5 136482.5 10362.5 136617.5 ;
      RECT  10297.5 136482.5 10362.5 136617.5 ;
      RECT  10107.5 136482.5 10172.5 136617.5 ;
      RECT  10297.5 136482.5 10362.5 136617.5 ;
      RECT  10487.5 136482.5 10552.5 136617.5 ;
      RECT  10487.5 136482.5 10552.5 136617.5 ;
      RECT  10297.5 136482.5 10362.5 136617.5 ;
      RECT  10657.5 137412.5 10722.5 137547.5 ;
      RECT  10657.5 136437.5 10722.5 136572.5 ;
      RECT  10492.5 136712.5 10357.5 136777.5 ;
      RECT  10235.0 136927.5 10100.0 136992.5 ;
      RECT  10297.5 137322.5 10362.5 137457.5 ;
      RECT  10487.5 136482.5 10552.5 136617.5 ;
      RECT  10587.5 136927.5 10452.5 136992.5 ;
      RECT  10100.0 136927.5 10235.0 136992.5 ;
      RECT  10357.5 136712.5 10492.5 136777.5 ;
      RECT  10452.5 136927.5 10587.5 136992.5 ;
      RECT  10040.0 137632.5 10960.0 137697.5 ;
      RECT  10040.0 136287.5 10960.0 136352.5 ;
      RECT  11387.5 137480.0 11452.5 137665.0 ;
      RECT  11387.5 136320.0 11452.5 136505.0 ;
      RECT  11027.5 136437.5 11092.5 136287.5 ;
      RECT  11027.5 137322.5 11092.5 137697.5 ;
      RECT  11217.5 136437.5 11282.5 137322.5 ;
      RECT  11027.5 137322.5 11092.5 137457.5 ;
      RECT  11217.5 137322.5 11282.5 137457.5 ;
      RECT  11217.5 137322.5 11282.5 137457.5 ;
      RECT  11027.5 137322.5 11092.5 137457.5 ;
      RECT  11027.5 136437.5 11092.5 136572.5 ;
      RECT  11217.5 136437.5 11282.5 136572.5 ;
      RECT  11217.5 136437.5 11282.5 136572.5 ;
      RECT  11027.5 136437.5 11092.5 136572.5 ;
      RECT  11387.5 137412.5 11452.5 137547.5 ;
      RECT  11387.5 136437.5 11452.5 136572.5 ;
      RECT  11085.0 136880.0 11150.0 137015.0 ;
      RECT  11085.0 136880.0 11150.0 137015.0 ;
      RECT  11250.0 136915.0 11315.0 136980.0 ;
      RECT  10960.0 137632.5 11520.0 137697.5 ;
      RECT  10960.0 136287.5 11520.0 136352.5 ;
      RECT  9222.5 136880.0 9287.5 137015.0 ;
      RECT  9362.5 136607.5 9427.5 136742.5 ;
      RECT  10357.5 136712.5 10222.5 136777.5 ;
      RECT  9907.5 137850.0 9972.5 137665.0 ;
      RECT  9907.5 139010.0 9972.5 138825.0 ;
      RECT  9547.5 138892.5 9612.5 139042.5 ;
      RECT  9547.5 138007.5 9612.5 137632.5 ;
      RECT  9737.5 138892.5 9802.5 138007.5 ;
      RECT  9547.5 138007.5 9612.5 137872.5 ;
      RECT  9737.5 138007.5 9802.5 137872.5 ;
      RECT  9737.5 138007.5 9802.5 137872.5 ;
      RECT  9547.5 138007.5 9612.5 137872.5 ;
      RECT  9547.5 138892.5 9612.5 138757.5 ;
      RECT  9737.5 138892.5 9802.5 138757.5 ;
      RECT  9737.5 138892.5 9802.5 138757.5 ;
      RECT  9547.5 138892.5 9612.5 138757.5 ;
      RECT  9907.5 137917.5 9972.5 137782.5 ;
      RECT  9907.5 138892.5 9972.5 138757.5 ;
      RECT  9605.0 138450.0 9670.0 138315.0 ;
      RECT  9605.0 138450.0 9670.0 138315.0 ;
      RECT  9770.0 138415.0 9835.0 138350.0 ;
      RECT  9480.0 137697.5 10040.0 137632.5 ;
      RECT  9480.0 139042.5 10040.0 138977.5 ;
      RECT  10107.5 138847.5 10172.5 139042.5 ;
      RECT  10107.5 138007.5 10172.5 137632.5 ;
      RECT  10487.5 138007.5 10552.5 137632.5 ;
      RECT  10657.5 137850.0 10722.5 137665.0 ;
      RECT  10657.5 139010.0 10722.5 138825.0 ;
      RECT  10107.5 138007.5 10172.5 137872.5 ;
      RECT  10297.5 138007.5 10362.5 137872.5 ;
      RECT  10297.5 138007.5 10362.5 137872.5 ;
      RECT  10107.5 138007.5 10172.5 137872.5 ;
      RECT  10297.5 138007.5 10362.5 137872.5 ;
      RECT  10487.5 138007.5 10552.5 137872.5 ;
      RECT  10487.5 138007.5 10552.5 137872.5 ;
      RECT  10297.5 138007.5 10362.5 137872.5 ;
      RECT  10107.5 138847.5 10172.5 138712.5 ;
      RECT  10297.5 138847.5 10362.5 138712.5 ;
      RECT  10297.5 138847.5 10362.5 138712.5 ;
      RECT  10107.5 138847.5 10172.5 138712.5 ;
      RECT  10297.5 138847.5 10362.5 138712.5 ;
      RECT  10487.5 138847.5 10552.5 138712.5 ;
      RECT  10487.5 138847.5 10552.5 138712.5 ;
      RECT  10297.5 138847.5 10362.5 138712.5 ;
      RECT  10657.5 137917.5 10722.5 137782.5 ;
      RECT  10657.5 138892.5 10722.5 138757.5 ;
      RECT  10492.5 138617.5 10357.5 138552.5 ;
      RECT  10235.0 138402.5 10100.0 138337.5 ;
      RECT  10297.5 138007.5 10362.5 137872.5 ;
      RECT  10487.5 138847.5 10552.5 138712.5 ;
      RECT  10587.5 138402.5 10452.5 138337.5 ;
      RECT  10100.0 138402.5 10235.0 138337.5 ;
      RECT  10357.5 138617.5 10492.5 138552.5 ;
      RECT  10452.5 138402.5 10587.5 138337.5 ;
      RECT  10040.0 137697.5 10960.0 137632.5 ;
      RECT  10040.0 139042.5 10960.0 138977.5 ;
      RECT  11387.5 137850.0 11452.5 137665.0 ;
      RECT  11387.5 139010.0 11452.5 138825.0 ;
      RECT  11027.5 138892.5 11092.5 139042.5 ;
      RECT  11027.5 138007.5 11092.5 137632.5 ;
      RECT  11217.5 138892.5 11282.5 138007.5 ;
      RECT  11027.5 138007.5 11092.5 137872.5 ;
      RECT  11217.5 138007.5 11282.5 137872.5 ;
      RECT  11217.5 138007.5 11282.5 137872.5 ;
      RECT  11027.5 138007.5 11092.5 137872.5 ;
      RECT  11027.5 138892.5 11092.5 138757.5 ;
      RECT  11217.5 138892.5 11282.5 138757.5 ;
      RECT  11217.5 138892.5 11282.5 138757.5 ;
      RECT  11027.5 138892.5 11092.5 138757.5 ;
      RECT  11387.5 137917.5 11452.5 137782.5 ;
      RECT  11387.5 138892.5 11452.5 138757.5 ;
      RECT  11085.0 138450.0 11150.0 138315.0 ;
      RECT  11085.0 138450.0 11150.0 138315.0 ;
      RECT  11250.0 138415.0 11315.0 138350.0 ;
      RECT  10960.0 137697.5 11520.0 137632.5 ;
      RECT  10960.0 139042.5 11520.0 138977.5 ;
      RECT  9222.5 138315.0 9287.5 138450.0 ;
      RECT  9362.5 138587.5 9427.5 138722.5 ;
      RECT  10357.5 138552.5 10222.5 138617.5 ;
      RECT  9907.5 140170.0 9972.5 140355.0 ;
      RECT  9907.5 139010.0 9972.5 139195.0 ;
      RECT  9547.5 139127.5 9612.5 138977.5 ;
      RECT  9547.5 140012.5 9612.5 140387.5 ;
      RECT  9737.5 139127.5 9802.5 140012.5 ;
      RECT  9547.5 140012.5 9612.5 140147.5 ;
      RECT  9737.5 140012.5 9802.5 140147.5 ;
      RECT  9737.5 140012.5 9802.5 140147.5 ;
      RECT  9547.5 140012.5 9612.5 140147.5 ;
      RECT  9547.5 139127.5 9612.5 139262.5 ;
      RECT  9737.5 139127.5 9802.5 139262.5 ;
      RECT  9737.5 139127.5 9802.5 139262.5 ;
      RECT  9547.5 139127.5 9612.5 139262.5 ;
      RECT  9907.5 140102.5 9972.5 140237.5 ;
      RECT  9907.5 139127.5 9972.5 139262.5 ;
      RECT  9605.0 139570.0 9670.0 139705.0 ;
      RECT  9605.0 139570.0 9670.0 139705.0 ;
      RECT  9770.0 139605.0 9835.0 139670.0 ;
      RECT  9480.0 140322.5 10040.0 140387.5 ;
      RECT  9480.0 138977.5 10040.0 139042.5 ;
      RECT  10107.5 139172.5 10172.5 138977.5 ;
      RECT  10107.5 140012.5 10172.5 140387.5 ;
      RECT  10487.5 140012.5 10552.5 140387.5 ;
      RECT  10657.5 140170.0 10722.5 140355.0 ;
      RECT  10657.5 139010.0 10722.5 139195.0 ;
      RECT  10107.5 140012.5 10172.5 140147.5 ;
      RECT  10297.5 140012.5 10362.5 140147.5 ;
      RECT  10297.5 140012.5 10362.5 140147.5 ;
      RECT  10107.5 140012.5 10172.5 140147.5 ;
      RECT  10297.5 140012.5 10362.5 140147.5 ;
      RECT  10487.5 140012.5 10552.5 140147.5 ;
      RECT  10487.5 140012.5 10552.5 140147.5 ;
      RECT  10297.5 140012.5 10362.5 140147.5 ;
      RECT  10107.5 139172.5 10172.5 139307.5 ;
      RECT  10297.5 139172.5 10362.5 139307.5 ;
      RECT  10297.5 139172.5 10362.5 139307.5 ;
      RECT  10107.5 139172.5 10172.5 139307.5 ;
      RECT  10297.5 139172.5 10362.5 139307.5 ;
      RECT  10487.5 139172.5 10552.5 139307.5 ;
      RECT  10487.5 139172.5 10552.5 139307.5 ;
      RECT  10297.5 139172.5 10362.5 139307.5 ;
      RECT  10657.5 140102.5 10722.5 140237.5 ;
      RECT  10657.5 139127.5 10722.5 139262.5 ;
      RECT  10492.5 139402.5 10357.5 139467.5 ;
      RECT  10235.0 139617.5 10100.0 139682.5 ;
      RECT  10297.5 140012.5 10362.5 140147.5 ;
      RECT  10487.5 139172.5 10552.5 139307.5 ;
      RECT  10587.5 139617.5 10452.5 139682.5 ;
      RECT  10100.0 139617.5 10235.0 139682.5 ;
      RECT  10357.5 139402.5 10492.5 139467.5 ;
      RECT  10452.5 139617.5 10587.5 139682.5 ;
      RECT  10040.0 140322.5 10960.0 140387.5 ;
      RECT  10040.0 138977.5 10960.0 139042.5 ;
      RECT  11387.5 140170.0 11452.5 140355.0 ;
      RECT  11387.5 139010.0 11452.5 139195.0 ;
      RECT  11027.5 139127.5 11092.5 138977.5 ;
      RECT  11027.5 140012.5 11092.5 140387.5 ;
      RECT  11217.5 139127.5 11282.5 140012.5 ;
      RECT  11027.5 140012.5 11092.5 140147.5 ;
      RECT  11217.5 140012.5 11282.5 140147.5 ;
      RECT  11217.5 140012.5 11282.5 140147.5 ;
      RECT  11027.5 140012.5 11092.5 140147.5 ;
      RECT  11027.5 139127.5 11092.5 139262.5 ;
      RECT  11217.5 139127.5 11282.5 139262.5 ;
      RECT  11217.5 139127.5 11282.5 139262.5 ;
      RECT  11027.5 139127.5 11092.5 139262.5 ;
      RECT  11387.5 140102.5 11452.5 140237.5 ;
      RECT  11387.5 139127.5 11452.5 139262.5 ;
      RECT  11085.0 139570.0 11150.0 139705.0 ;
      RECT  11085.0 139570.0 11150.0 139705.0 ;
      RECT  11250.0 139605.0 11315.0 139670.0 ;
      RECT  10960.0 140322.5 11520.0 140387.5 ;
      RECT  10960.0 138977.5 11520.0 139042.5 ;
      RECT  9222.5 139570.0 9287.5 139705.0 ;
      RECT  9362.5 139297.5 9427.5 139432.5 ;
      RECT  10357.5 139402.5 10222.5 139467.5 ;
      RECT  9907.5 140540.0 9972.5 140355.0 ;
      RECT  9907.5 141700.0 9972.5 141515.0 ;
      RECT  9547.5 141582.5 9612.5 141732.5 ;
      RECT  9547.5 140697.5 9612.5 140322.5 ;
      RECT  9737.5 141582.5 9802.5 140697.5 ;
      RECT  9547.5 140697.5 9612.5 140562.5 ;
      RECT  9737.5 140697.5 9802.5 140562.5 ;
      RECT  9737.5 140697.5 9802.5 140562.5 ;
      RECT  9547.5 140697.5 9612.5 140562.5 ;
      RECT  9547.5 141582.5 9612.5 141447.5 ;
      RECT  9737.5 141582.5 9802.5 141447.5 ;
      RECT  9737.5 141582.5 9802.5 141447.5 ;
      RECT  9547.5 141582.5 9612.5 141447.5 ;
      RECT  9907.5 140607.5 9972.5 140472.5 ;
      RECT  9907.5 141582.5 9972.5 141447.5 ;
      RECT  9605.0 141140.0 9670.0 141005.0 ;
      RECT  9605.0 141140.0 9670.0 141005.0 ;
      RECT  9770.0 141105.0 9835.0 141040.0 ;
      RECT  9480.0 140387.5 10040.0 140322.5 ;
      RECT  9480.0 141732.5 10040.0 141667.5 ;
      RECT  10107.5 141537.5 10172.5 141732.5 ;
      RECT  10107.5 140697.5 10172.5 140322.5 ;
      RECT  10487.5 140697.5 10552.5 140322.5 ;
      RECT  10657.5 140540.0 10722.5 140355.0 ;
      RECT  10657.5 141700.0 10722.5 141515.0 ;
      RECT  10107.5 140697.5 10172.5 140562.5 ;
      RECT  10297.5 140697.5 10362.5 140562.5 ;
      RECT  10297.5 140697.5 10362.5 140562.5 ;
      RECT  10107.5 140697.5 10172.5 140562.5 ;
      RECT  10297.5 140697.5 10362.5 140562.5 ;
      RECT  10487.5 140697.5 10552.5 140562.5 ;
      RECT  10487.5 140697.5 10552.5 140562.5 ;
      RECT  10297.5 140697.5 10362.5 140562.5 ;
      RECT  10107.5 141537.5 10172.5 141402.5 ;
      RECT  10297.5 141537.5 10362.5 141402.5 ;
      RECT  10297.5 141537.5 10362.5 141402.5 ;
      RECT  10107.5 141537.5 10172.5 141402.5 ;
      RECT  10297.5 141537.5 10362.5 141402.5 ;
      RECT  10487.5 141537.5 10552.5 141402.5 ;
      RECT  10487.5 141537.5 10552.5 141402.5 ;
      RECT  10297.5 141537.5 10362.5 141402.5 ;
      RECT  10657.5 140607.5 10722.5 140472.5 ;
      RECT  10657.5 141582.5 10722.5 141447.5 ;
      RECT  10492.5 141307.5 10357.5 141242.5 ;
      RECT  10235.0 141092.5 10100.0 141027.5 ;
      RECT  10297.5 140697.5 10362.5 140562.5 ;
      RECT  10487.5 141537.5 10552.5 141402.5 ;
      RECT  10587.5 141092.5 10452.5 141027.5 ;
      RECT  10100.0 141092.5 10235.0 141027.5 ;
      RECT  10357.5 141307.5 10492.5 141242.5 ;
      RECT  10452.5 141092.5 10587.5 141027.5 ;
      RECT  10040.0 140387.5 10960.0 140322.5 ;
      RECT  10040.0 141732.5 10960.0 141667.5 ;
      RECT  11387.5 140540.0 11452.5 140355.0 ;
      RECT  11387.5 141700.0 11452.5 141515.0 ;
      RECT  11027.5 141582.5 11092.5 141732.5 ;
      RECT  11027.5 140697.5 11092.5 140322.5 ;
      RECT  11217.5 141582.5 11282.5 140697.5 ;
      RECT  11027.5 140697.5 11092.5 140562.5 ;
      RECT  11217.5 140697.5 11282.5 140562.5 ;
      RECT  11217.5 140697.5 11282.5 140562.5 ;
      RECT  11027.5 140697.5 11092.5 140562.5 ;
      RECT  11027.5 141582.5 11092.5 141447.5 ;
      RECT  11217.5 141582.5 11282.5 141447.5 ;
      RECT  11217.5 141582.5 11282.5 141447.5 ;
      RECT  11027.5 141582.5 11092.5 141447.5 ;
      RECT  11387.5 140607.5 11452.5 140472.5 ;
      RECT  11387.5 141582.5 11452.5 141447.5 ;
      RECT  11085.0 141140.0 11150.0 141005.0 ;
      RECT  11085.0 141140.0 11150.0 141005.0 ;
      RECT  11250.0 141105.0 11315.0 141040.0 ;
      RECT  10960.0 140387.5 11520.0 140322.5 ;
      RECT  10960.0 141732.5 11520.0 141667.5 ;
      RECT  9222.5 141005.0 9287.5 141140.0 ;
      RECT  9362.5 141277.5 9427.5 141412.5 ;
      RECT  10357.5 141242.5 10222.5 141307.5 ;
      RECT  9907.5 142860.0 9972.5 143045.0 ;
      RECT  9907.5 141700.0 9972.5 141885.0 ;
      RECT  9547.5 141817.5 9612.5 141667.5 ;
      RECT  9547.5 142702.5 9612.5 143077.5 ;
      RECT  9737.5 141817.5 9802.5 142702.5 ;
      RECT  9547.5 142702.5 9612.5 142837.5 ;
      RECT  9737.5 142702.5 9802.5 142837.5 ;
      RECT  9737.5 142702.5 9802.5 142837.5 ;
      RECT  9547.5 142702.5 9612.5 142837.5 ;
      RECT  9547.5 141817.5 9612.5 141952.5 ;
      RECT  9737.5 141817.5 9802.5 141952.5 ;
      RECT  9737.5 141817.5 9802.5 141952.5 ;
      RECT  9547.5 141817.5 9612.5 141952.5 ;
      RECT  9907.5 142792.5 9972.5 142927.5 ;
      RECT  9907.5 141817.5 9972.5 141952.5 ;
      RECT  9605.0 142260.0 9670.0 142395.0 ;
      RECT  9605.0 142260.0 9670.0 142395.0 ;
      RECT  9770.0 142295.0 9835.0 142360.0 ;
      RECT  9480.0 143012.5 10040.0 143077.5 ;
      RECT  9480.0 141667.5 10040.0 141732.5 ;
      RECT  10107.5 141862.5 10172.5 141667.5 ;
      RECT  10107.5 142702.5 10172.5 143077.5 ;
      RECT  10487.5 142702.5 10552.5 143077.5 ;
      RECT  10657.5 142860.0 10722.5 143045.0 ;
      RECT  10657.5 141700.0 10722.5 141885.0 ;
      RECT  10107.5 142702.5 10172.5 142837.5 ;
      RECT  10297.5 142702.5 10362.5 142837.5 ;
      RECT  10297.5 142702.5 10362.5 142837.5 ;
      RECT  10107.5 142702.5 10172.5 142837.5 ;
      RECT  10297.5 142702.5 10362.5 142837.5 ;
      RECT  10487.5 142702.5 10552.5 142837.5 ;
      RECT  10487.5 142702.5 10552.5 142837.5 ;
      RECT  10297.5 142702.5 10362.5 142837.5 ;
      RECT  10107.5 141862.5 10172.5 141997.5 ;
      RECT  10297.5 141862.5 10362.5 141997.5 ;
      RECT  10297.5 141862.5 10362.5 141997.5 ;
      RECT  10107.5 141862.5 10172.5 141997.5 ;
      RECT  10297.5 141862.5 10362.5 141997.5 ;
      RECT  10487.5 141862.5 10552.5 141997.5 ;
      RECT  10487.5 141862.5 10552.5 141997.5 ;
      RECT  10297.5 141862.5 10362.5 141997.5 ;
      RECT  10657.5 142792.5 10722.5 142927.5 ;
      RECT  10657.5 141817.5 10722.5 141952.5 ;
      RECT  10492.5 142092.5 10357.5 142157.5 ;
      RECT  10235.0 142307.5 10100.0 142372.5 ;
      RECT  10297.5 142702.5 10362.5 142837.5 ;
      RECT  10487.5 141862.5 10552.5 141997.5 ;
      RECT  10587.5 142307.5 10452.5 142372.5 ;
      RECT  10100.0 142307.5 10235.0 142372.5 ;
      RECT  10357.5 142092.5 10492.5 142157.5 ;
      RECT  10452.5 142307.5 10587.5 142372.5 ;
      RECT  10040.0 143012.5 10960.0 143077.5 ;
      RECT  10040.0 141667.5 10960.0 141732.5 ;
      RECT  11387.5 142860.0 11452.5 143045.0 ;
      RECT  11387.5 141700.0 11452.5 141885.0 ;
      RECT  11027.5 141817.5 11092.5 141667.5 ;
      RECT  11027.5 142702.5 11092.5 143077.5 ;
      RECT  11217.5 141817.5 11282.5 142702.5 ;
      RECT  11027.5 142702.5 11092.5 142837.5 ;
      RECT  11217.5 142702.5 11282.5 142837.5 ;
      RECT  11217.5 142702.5 11282.5 142837.5 ;
      RECT  11027.5 142702.5 11092.5 142837.5 ;
      RECT  11027.5 141817.5 11092.5 141952.5 ;
      RECT  11217.5 141817.5 11282.5 141952.5 ;
      RECT  11217.5 141817.5 11282.5 141952.5 ;
      RECT  11027.5 141817.5 11092.5 141952.5 ;
      RECT  11387.5 142792.5 11452.5 142927.5 ;
      RECT  11387.5 141817.5 11452.5 141952.5 ;
      RECT  11085.0 142260.0 11150.0 142395.0 ;
      RECT  11085.0 142260.0 11150.0 142395.0 ;
      RECT  11250.0 142295.0 11315.0 142360.0 ;
      RECT  10960.0 143012.5 11520.0 143077.5 ;
      RECT  10960.0 141667.5 11520.0 141732.5 ;
      RECT  9222.5 142260.0 9287.5 142395.0 ;
      RECT  9362.5 141987.5 9427.5 142122.5 ;
      RECT  10357.5 142092.5 10222.5 142157.5 ;
      RECT  9907.5 143230.0 9972.5 143045.0 ;
      RECT  9907.5 144390.0 9972.5 144205.0 ;
      RECT  9547.5 144272.5 9612.5 144422.5 ;
      RECT  9547.5 143387.5 9612.5 143012.5 ;
      RECT  9737.5 144272.5 9802.5 143387.5 ;
      RECT  9547.5 143387.5 9612.5 143252.5 ;
      RECT  9737.5 143387.5 9802.5 143252.5 ;
      RECT  9737.5 143387.5 9802.5 143252.5 ;
      RECT  9547.5 143387.5 9612.5 143252.5 ;
      RECT  9547.5 144272.5 9612.5 144137.5 ;
      RECT  9737.5 144272.5 9802.5 144137.5 ;
      RECT  9737.5 144272.5 9802.5 144137.5 ;
      RECT  9547.5 144272.5 9612.5 144137.5 ;
      RECT  9907.5 143297.5 9972.5 143162.5 ;
      RECT  9907.5 144272.5 9972.5 144137.5 ;
      RECT  9605.0 143830.0 9670.0 143695.0 ;
      RECT  9605.0 143830.0 9670.0 143695.0 ;
      RECT  9770.0 143795.0 9835.0 143730.0 ;
      RECT  9480.0 143077.5 10040.0 143012.5 ;
      RECT  9480.0 144422.5 10040.0 144357.5 ;
      RECT  10107.5 144227.5 10172.5 144422.5 ;
      RECT  10107.5 143387.5 10172.5 143012.5 ;
      RECT  10487.5 143387.5 10552.5 143012.5 ;
      RECT  10657.5 143230.0 10722.5 143045.0 ;
      RECT  10657.5 144390.0 10722.5 144205.0 ;
      RECT  10107.5 143387.5 10172.5 143252.5 ;
      RECT  10297.5 143387.5 10362.5 143252.5 ;
      RECT  10297.5 143387.5 10362.5 143252.5 ;
      RECT  10107.5 143387.5 10172.5 143252.5 ;
      RECT  10297.5 143387.5 10362.5 143252.5 ;
      RECT  10487.5 143387.5 10552.5 143252.5 ;
      RECT  10487.5 143387.5 10552.5 143252.5 ;
      RECT  10297.5 143387.5 10362.5 143252.5 ;
      RECT  10107.5 144227.5 10172.5 144092.5 ;
      RECT  10297.5 144227.5 10362.5 144092.5 ;
      RECT  10297.5 144227.5 10362.5 144092.5 ;
      RECT  10107.5 144227.5 10172.5 144092.5 ;
      RECT  10297.5 144227.5 10362.5 144092.5 ;
      RECT  10487.5 144227.5 10552.5 144092.5 ;
      RECT  10487.5 144227.5 10552.5 144092.5 ;
      RECT  10297.5 144227.5 10362.5 144092.5 ;
      RECT  10657.5 143297.5 10722.5 143162.5 ;
      RECT  10657.5 144272.5 10722.5 144137.5 ;
      RECT  10492.5 143997.5 10357.5 143932.5 ;
      RECT  10235.0 143782.5 10100.0 143717.5 ;
      RECT  10297.5 143387.5 10362.5 143252.5 ;
      RECT  10487.5 144227.5 10552.5 144092.5 ;
      RECT  10587.5 143782.5 10452.5 143717.5 ;
      RECT  10100.0 143782.5 10235.0 143717.5 ;
      RECT  10357.5 143997.5 10492.5 143932.5 ;
      RECT  10452.5 143782.5 10587.5 143717.5 ;
      RECT  10040.0 143077.5 10960.0 143012.5 ;
      RECT  10040.0 144422.5 10960.0 144357.5 ;
      RECT  11387.5 143230.0 11452.5 143045.0 ;
      RECT  11387.5 144390.0 11452.5 144205.0 ;
      RECT  11027.5 144272.5 11092.5 144422.5 ;
      RECT  11027.5 143387.5 11092.5 143012.5 ;
      RECT  11217.5 144272.5 11282.5 143387.5 ;
      RECT  11027.5 143387.5 11092.5 143252.5 ;
      RECT  11217.5 143387.5 11282.5 143252.5 ;
      RECT  11217.5 143387.5 11282.5 143252.5 ;
      RECT  11027.5 143387.5 11092.5 143252.5 ;
      RECT  11027.5 144272.5 11092.5 144137.5 ;
      RECT  11217.5 144272.5 11282.5 144137.5 ;
      RECT  11217.5 144272.5 11282.5 144137.5 ;
      RECT  11027.5 144272.5 11092.5 144137.5 ;
      RECT  11387.5 143297.5 11452.5 143162.5 ;
      RECT  11387.5 144272.5 11452.5 144137.5 ;
      RECT  11085.0 143830.0 11150.0 143695.0 ;
      RECT  11085.0 143830.0 11150.0 143695.0 ;
      RECT  11250.0 143795.0 11315.0 143730.0 ;
      RECT  10960.0 143077.5 11520.0 143012.5 ;
      RECT  10960.0 144422.5 11520.0 144357.5 ;
      RECT  9222.5 143695.0 9287.5 143830.0 ;
      RECT  9362.5 143967.5 9427.5 144102.5 ;
      RECT  10357.5 143932.5 10222.5 143997.5 ;
      RECT  9907.5 145550.0 9972.5 145735.0 ;
      RECT  9907.5 144390.0 9972.5 144575.0 ;
      RECT  9547.5 144507.5 9612.5 144357.5 ;
      RECT  9547.5 145392.5 9612.5 145767.5 ;
      RECT  9737.5 144507.5 9802.5 145392.5 ;
      RECT  9547.5 145392.5 9612.5 145527.5 ;
      RECT  9737.5 145392.5 9802.5 145527.5 ;
      RECT  9737.5 145392.5 9802.5 145527.5 ;
      RECT  9547.5 145392.5 9612.5 145527.5 ;
      RECT  9547.5 144507.5 9612.5 144642.5 ;
      RECT  9737.5 144507.5 9802.5 144642.5 ;
      RECT  9737.5 144507.5 9802.5 144642.5 ;
      RECT  9547.5 144507.5 9612.5 144642.5 ;
      RECT  9907.5 145482.5 9972.5 145617.5 ;
      RECT  9907.5 144507.5 9972.5 144642.5 ;
      RECT  9605.0 144950.0 9670.0 145085.0 ;
      RECT  9605.0 144950.0 9670.0 145085.0 ;
      RECT  9770.0 144985.0 9835.0 145050.0 ;
      RECT  9480.0 145702.5 10040.0 145767.5 ;
      RECT  9480.0 144357.5 10040.0 144422.5 ;
      RECT  10107.5 144552.5 10172.5 144357.5 ;
      RECT  10107.5 145392.5 10172.5 145767.5 ;
      RECT  10487.5 145392.5 10552.5 145767.5 ;
      RECT  10657.5 145550.0 10722.5 145735.0 ;
      RECT  10657.5 144390.0 10722.5 144575.0 ;
      RECT  10107.5 145392.5 10172.5 145527.5 ;
      RECT  10297.5 145392.5 10362.5 145527.5 ;
      RECT  10297.5 145392.5 10362.5 145527.5 ;
      RECT  10107.5 145392.5 10172.5 145527.5 ;
      RECT  10297.5 145392.5 10362.5 145527.5 ;
      RECT  10487.5 145392.5 10552.5 145527.5 ;
      RECT  10487.5 145392.5 10552.5 145527.5 ;
      RECT  10297.5 145392.5 10362.5 145527.5 ;
      RECT  10107.5 144552.5 10172.5 144687.5 ;
      RECT  10297.5 144552.5 10362.5 144687.5 ;
      RECT  10297.5 144552.5 10362.5 144687.5 ;
      RECT  10107.5 144552.5 10172.5 144687.5 ;
      RECT  10297.5 144552.5 10362.5 144687.5 ;
      RECT  10487.5 144552.5 10552.5 144687.5 ;
      RECT  10487.5 144552.5 10552.5 144687.5 ;
      RECT  10297.5 144552.5 10362.5 144687.5 ;
      RECT  10657.5 145482.5 10722.5 145617.5 ;
      RECT  10657.5 144507.5 10722.5 144642.5 ;
      RECT  10492.5 144782.5 10357.5 144847.5 ;
      RECT  10235.0 144997.5 10100.0 145062.5 ;
      RECT  10297.5 145392.5 10362.5 145527.5 ;
      RECT  10487.5 144552.5 10552.5 144687.5 ;
      RECT  10587.5 144997.5 10452.5 145062.5 ;
      RECT  10100.0 144997.5 10235.0 145062.5 ;
      RECT  10357.5 144782.5 10492.5 144847.5 ;
      RECT  10452.5 144997.5 10587.5 145062.5 ;
      RECT  10040.0 145702.5 10960.0 145767.5 ;
      RECT  10040.0 144357.5 10960.0 144422.5 ;
      RECT  11387.5 145550.0 11452.5 145735.0 ;
      RECT  11387.5 144390.0 11452.5 144575.0 ;
      RECT  11027.5 144507.5 11092.5 144357.5 ;
      RECT  11027.5 145392.5 11092.5 145767.5 ;
      RECT  11217.5 144507.5 11282.5 145392.5 ;
      RECT  11027.5 145392.5 11092.5 145527.5 ;
      RECT  11217.5 145392.5 11282.5 145527.5 ;
      RECT  11217.5 145392.5 11282.5 145527.5 ;
      RECT  11027.5 145392.5 11092.5 145527.5 ;
      RECT  11027.5 144507.5 11092.5 144642.5 ;
      RECT  11217.5 144507.5 11282.5 144642.5 ;
      RECT  11217.5 144507.5 11282.5 144642.5 ;
      RECT  11027.5 144507.5 11092.5 144642.5 ;
      RECT  11387.5 145482.5 11452.5 145617.5 ;
      RECT  11387.5 144507.5 11452.5 144642.5 ;
      RECT  11085.0 144950.0 11150.0 145085.0 ;
      RECT  11085.0 144950.0 11150.0 145085.0 ;
      RECT  11250.0 144985.0 11315.0 145050.0 ;
      RECT  10960.0 145702.5 11520.0 145767.5 ;
      RECT  10960.0 144357.5 11520.0 144422.5 ;
      RECT  9222.5 144950.0 9287.5 145085.0 ;
      RECT  9362.5 144677.5 9427.5 144812.5 ;
      RECT  10357.5 144782.5 10222.5 144847.5 ;
      RECT  9907.5 145920.0 9972.5 145735.0 ;
      RECT  9907.5 147080.0 9972.5 146895.0 ;
      RECT  9547.5 146962.5 9612.5 147112.5 ;
      RECT  9547.5 146077.5 9612.5 145702.5 ;
      RECT  9737.5 146962.5 9802.5 146077.5 ;
      RECT  9547.5 146077.5 9612.5 145942.5 ;
      RECT  9737.5 146077.5 9802.5 145942.5 ;
      RECT  9737.5 146077.5 9802.5 145942.5 ;
      RECT  9547.5 146077.5 9612.5 145942.5 ;
      RECT  9547.5 146962.5 9612.5 146827.5 ;
      RECT  9737.5 146962.5 9802.5 146827.5 ;
      RECT  9737.5 146962.5 9802.5 146827.5 ;
      RECT  9547.5 146962.5 9612.5 146827.5 ;
      RECT  9907.5 145987.5 9972.5 145852.5 ;
      RECT  9907.5 146962.5 9972.5 146827.5 ;
      RECT  9605.0 146520.0 9670.0 146385.0 ;
      RECT  9605.0 146520.0 9670.0 146385.0 ;
      RECT  9770.0 146485.0 9835.0 146420.0 ;
      RECT  9480.0 145767.5 10040.0 145702.5 ;
      RECT  9480.0 147112.5 10040.0 147047.5 ;
      RECT  10107.5 146917.5 10172.5 147112.5 ;
      RECT  10107.5 146077.5 10172.5 145702.5 ;
      RECT  10487.5 146077.5 10552.5 145702.5 ;
      RECT  10657.5 145920.0 10722.5 145735.0 ;
      RECT  10657.5 147080.0 10722.5 146895.0 ;
      RECT  10107.5 146077.5 10172.5 145942.5 ;
      RECT  10297.5 146077.5 10362.5 145942.5 ;
      RECT  10297.5 146077.5 10362.5 145942.5 ;
      RECT  10107.5 146077.5 10172.5 145942.5 ;
      RECT  10297.5 146077.5 10362.5 145942.5 ;
      RECT  10487.5 146077.5 10552.5 145942.5 ;
      RECT  10487.5 146077.5 10552.5 145942.5 ;
      RECT  10297.5 146077.5 10362.5 145942.5 ;
      RECT  10107.5 146917.5 10172.5 146782.5 ;
      RECT  10297.5 146917.5 10362.5 146782.5 ;
      RECT  10297.5 146917.5 10362.5 146782.5 ;
      RECT  10107.5 146917.5 10172.5 146782.5 ;
      RECT  10297.5 146917.5 10362.5 146782.5 ;
      RECT  10487.5 146917.5 10552.5 146782.5 ;
      RECT  10487.5 146917.5 10552.5 146782.5 ;
      RECT  10297.5 146917.5 10362.5 146782.5 ;
      RECT  10657.5 145987.5 10722.5 145852.5 ;
      RECT  10657.5 146962.5 10722.5 146827.5 ;
      RECT  10492.5 146687.5 10357.5 146622.5 ;
      RECT  10235.0 146472.5 10100.0 146407.5 ;
      RECT  10297.5 146077.5 10362.5 145942.5 ;
      RECT  10487.5 146917.5 10552.5 146782.5 ;
      RECT  10587.5 146472.5 10452.5 146407.5 ;
      RECT  10100.0 146472.5 10235.0 146407.5 ;
      RECT  10357.5 146687.5 10492.5 146622.5 ;
      RECT  10452.5 146472.5 10587.5 146407.5 ;
      RECT  10040.0 145767.5 10960.0 145702.5 ;
      RECT  10040.0 147112.5 10960.0 147047.5 ;
      RECT  11387.5 145920.0 11452.5 145735.0 ;
      RECT  11387.5 147080.0 11452.5 146895.0 ;
      RECT  11027.5 146962.5 11092.5 147112.5 ;
      RECT  11027.5 146077.5 11092.5 145702.5 ;
      RECT  11217.5 146962.5 11282.5 146077.5 ;
      RECT  11027.5 146077.5 11092.5 145942.5 ;
      RECT  11217.5 146077.5 11282.5 145942.5 ;
      RECT  11217.5 146077.5 11282.5 145942.5 ;
      RECT  11027.5 146077.5 11092.5 145942.5 ;
      RECT  11027.5 146962.5 11092.5 146827.5 ;
      RECT  11217.5 146962.5 11282.5 146827.5 ;
      RECT  11217.5 146962.5 11282.5 146827.5 ;
      RECT  11027.5 146962.5 11092.5 146827.5 ;
      RECT  11387.5 145987.5 11452.5 145852.5 ;
      RECT  11387.5 146962.5 11452.5 146827.5 ;
      RECT  11085.0 146520.0 11150.0 146385.0 ;
      RECT  11085.0 146520.0 11150.0 146385.0 ;
      RECT  11250.0 146485.0 11315.0 146420.0 ;
      RECT  10960.0 145767.5 11520.0 145702.5 ;
      RECT  10960.0 147112.5 11520.0 147047.5 ;
      RECT  9222.5 146385.0 9287.5 146520.0 ;
      RECT  9362.5 146657.5 9427.5 146792.5 ;
      RECT  10357.5 146622.5 10222.5 146687.5 ;
      RECT  9907.5 148240.0 9972.5 148425.0 ;
      RECT  9907.5 147080.0 9972.5 147265.0 ;
      RECT  9547.5 147197.5 9612.5 147047.5 ;
      RECT  9547.5 148082.5 9612.5 148457.5 ;
      RECT  9737.5 147197.5 9802.5 148082.5 ;
      RECT  9547.5 148082.5 9612.5 148217.5 ;
      RECT  9737.5 148082.5 9802.5 148217.5 ;
      RECT  9737.5 148082.5 9802.5 148217.5 ;
      RECT  9547.5 148082.5 9612.5 148217.5 ;
      RECT  9547.5 147197.5 9612.5 147332.5 ;
      RECT  9737.5 147197.5 9802.5 147332.5 ;
      RECT  9737.5 147197.5 9802.5 147332.5 ;
      RECT  9547.5 147197.5 9612.5 147332.5 ;
      RECT  9907.5 148172.5 9972.5 148307.5 ;
      RECT  9907.5 147197.5 9972.5 147332.5 ;
      RECT  9605.0 147640.0 9670.0 147775.0 ;
      RECT  9605.0 147640.0 9670.0 147775.0 ;
      RECT  9770.0 147675.0 9835.0 147740.0 ;
      RECT  9480.0 148392.5 10040.0 148457.5 ;
      RECT  9480.0 147047.5 10040.0 147112.5 ;
      RECT  10107.5 147242.5 10172.5 147047.5 ;
      RECT  10107.5 148082.5 10172.5 148457.5 ;
      RECT  10487.5 148082.5 10552.5 148457.5 ;
      RECT  10657.5 148240.0 10722.5 148425.0 ;
      RECT  10657.5 147080.0 10722.5 147265.0 ;
      RECT  10107.5 148082.5 10172.5 148217.5 ;
      RECT  10297.5 148082.5 10362.5 148217.5 ;
      RECT  10297.5 148082.5 10362.5 148217.5 ;
      RECT  10107.5 148082.5 10172.5 148217.5 ;
      RECT  10297.5 148082.5 10362.5 148217.5 ;
      RECT  10487.5 148082.5 10552.5 148217.5 ;
      RECT  10487.5 148082.5 10552.5 148217.5 ;
      RECT  10297.5 148082.5 10362.5 148217.5 ;
      RECT  10107.5 147242.5 10172.5 147377.5 ;
      RECT  10297.5 147242.5 10362.5 147377.5 ;
      RECT  10297.5 147242.5 10362.5 147377.5 ;
      RECT  10107.5 147242.5 10172.5 147377.5 ;
      RECT  10297.5 147242.5 10362.5 147377.5 ;
      RECT  10487.5 147242.5 10552.5 147377.5 ;
      RECT  10487.5 147242.5 10552.5 147377.5 ;
      RECT  10297.5 147242.5 10362.5 147377.5 ;
      RECT  10657.5 148172.5 10722.5 148307.5 ;
      RECT  10657.5 147197.5 10722.5 147332.5 ;
      RECT  10492.5 147472.5 10357.5 147537.5 ;
      RECT  10235.0 147687.5 10100.0 147752.5 ;
      RECT  10297.5 148082.5 10362.5 148217.5 ;
      RECT  10487.5 147242.5 10552.5 147377.5 ;
      RECT  10587.5 147687.5 10452.5 147752.5 ;
      RECT  10100.0 147687.5 10235.0 147752.5 ;
      RECT  10357.5 147472.5 10492.5 147537.5 ;
      RECT  10452.5 147687.5 10587.5 147752.5 ;
      RECT  10040.0 148392.5 10960.0 148457.5 ;
      RECT  10040.0 147047.5 10960.0 147112.5 ;
      RECT  11387.5 148240.0 11452.5 148425.0 ;
      RECT  11387.5 147080.0 11452.5 147265.0 ;
      RECT  11027.5 147197.5 11092.5 147047.5 ;
      RECT  11027.5 148082.5 11092.5 148457.5 ;
      RECT  11217.5 147197.5 11282.5 148082.5 ;
      RECT  11027.5 148082.5 11092.5 148217.5 ;
      RECT  11217.5 148082.5 11282.5 148217.5 ;
      RECT  11217.5 148082.5 11282.5 148217.5 ;
      RECT  11027.5 148082.5 11092.5 148217.5 ;
      RECT  11027.5 147197.5 11092.5 147332.5 ;
      RECT  11217.5 147197.5 11282.5 147332.5 ;
      RECT  11217.5 147197.5 11282.5 147332.5 ;
      RECT  11027.5 147197.5 11092.5 147332.5 ;
      RECT  11387.5 148172.5 11452.5 148307.5 ;
      RECT  11387.5 147197.5 11452.5 147332.5 ;
      RECT  11085.0 147640.0 11150.0 147775.0 ;
      RECT  11085.0 147640.0 11150.0 147775.0 ;
      RECT  11250.0 147675.0 11315.0 147740.0 ;
      RECT  10960.0 148392.5 11520.0 148457.5 ;
      RECT  10960.0 147047.5 11520.0 147112.5 ;
      RECT  9222.5 147640.0 9287.5 147775.0 ;
      RECT  9362.5 147367.5 9427.5 147502.5 ;
      RECT  10357.5 147472.5 10222.5 147537.5 ;
      RECT  9907.5 148610.0 9972.5 148425.0 ;
      RECT  9907.5 149770.0 9972.5 149585.0 ;
      RECT  9547.5 149652.5 9612.5 149802.5 ;
      RECT  9547.5 148767.5 9612.5 148392.5 ;
      RECT  9737.5 149652.5 9802.5 148767.5 ;
      RECT  9547.5 148767.5 9612.5 148632.5 ;
      RECT  9737.5 148767.5 9802.5 148632.5 ;
      RECT  9737.5 148767.5 9802.5 148632.5 ;
      RECT  9547.5 148767.5 9612.5 148632.5 ;
      RECT  9547.5 149652.5 9612.5 149517.5 ;
      RECT  9737.5 149652.5 9802.5 149517.5 ;
      RECT  9737.5 149652.5 9802.5 149517.5 ;
      RECT  9547.5 149652.5 9612.5 149517.5 ;
      RECT  9907.5 148677.5 9972.5 148542.5 ;
      RECT  9907.5 149652.5 9972.5 149517.5 ;
      RECT  9605.0 149210.0 9670.0 149075.0 ;
      RECT  9605.0 149210.0 9670.0 149075.0 ;
      RECT  9770.0 149175.0 9835.0 149110.0 ;
      RECT  9480.0 148457.5 10040.0 148392.5 ;
      RECT  9480.0 149802.5 10040.0 149737.5 ;
      RECT  10107.5 149607.5 10172.5 149802.5 ;
      RECT  10107.5 148767.5 10172.5 148392.5 ;
      RECT  10487.5 148767.5 10552.5 148392.5 ;
      RECT  10657.5 148610.0 10722.5 148425.0 ;
      RECT  10657.5 149770.0 10722.5 149585.0 ;
      RECT  10107.5 148767.5 10172.5 148632.5 ;
      RECT  10297.5 148767.5 10362.5 148632.5 ;
      RECT  10297.5 148767.5 10362.5 148632.5 ;
      RECT  10107.5 148767.5 10172.5 148632.5 ;
      RECT  10297.5 148767.5 10362.5 148632.5 ;
      RECT  10487.5 148767.5 10552.5 148632.5 ;
      RECT  10487.5 148767.5 10552.5 148632.5 ;
      RECT  10297.5 148767.5 10362.5 148632.5 ;
      RECT  10107.5 149607.5 10172.5 149472.5 ;
      RECT  10297.5 149607.5 10362.5 149472.5 ;
      RECT  10297.5 149607.5 10362.5 149472.5 ;
      RECT  10107.5 149607.5 10172.5 149472.5 ;
      RECT  10297.5 149607.5 10362.5 149472.5 ;
      RECT  10487.5 149607.5 10552.5 149472.5 ;
      RECT  10487.5 149607.5 10552.5 149472.5 ;
      RECT  10297.5 149607.5 10362.5 149472.5 ;
      RECT  10657.5 148677.5 10722.5 148542.5 ;
      RECT  10657.5 149652.5 10722.5 149517.5 ;
      RECT  10492.5 149377.5 10357.5 149312.5 ;
      RECT  10235.0 149162.5 10100.0 149097.5 ;
      RECT  10297.5 148767.5 10362.5 148632.5 ;
      RECT  10487.5 149607.5 10552.5 149472.5 ;
      RECT  10587.5 149162.5 10452.5 149097.5 ;
      RECT  10100.0 149162.5 10235.0 149097.5 ;
      RECT  10357.5 149377.5 10492.5 149312.5 ;
      RECT  10452.5 149162.5 10587.5 149097.5 ;
      RECT  10040.0 148457.5 10960.0 148392.5 ;
      RECT  10040.0 149802.5 10960.0 149737.5 ;
      RECT  11387.5 148610.0 11452.5 148425.0 ;
      RECT  11387.5 149770.0 11452.5 149585.0 ;
      RECT  11027.5 149652.5 11092.5 149802.5 ;
      RECT  11027.5 148767.5 11092.5 148392.5 ;
      RECT  11217.5 149652.5 11282.5 148767.5 ;
      RECT  11027.5 148767.5 11092.5 148632.5 ;
      RECT  11217.5 148767.5 11282.5 148632.5 ;
      RECT  11217.5 148767.5 11282.5 148632.5 ;
      RECT  11027.5 148767.5 11092.5 148632.5 ;
      RECT  11027.5 149652.5 11092.5 149517.5 ;
      RECT  11217.5 149652.5 11282.5 149517.5 ;
      RECT  11217.5 149652.5 11282.5 149517.5 ;
      RECT  11027.5 149652.5 11092.5 149517.5 ;
      RECT  11387.5 148677.5 11452.5 148542.5 ;
      RECT  11387.5 149652.5 11452.5 149517.5 ;
      RECT  11085.0 149210.0 11150.0 149075.0 ;
      RECT  11085.0 149210.0 11150.0 149075.0 ;
      RECT  11250.0 149175.0 11315.0 149110.0 ;
      RECT  10960.0 148457.5 11520.0 148392.5 ;
      RECT  10960.0 149802.5 11520.0 149737.5 ;
      RECT  9222.5 149075.0 9287.5 149210.0 ;
      RECT  9362.5 149347.5 9427.5 149482.5 ;
      RECT  10357.5 149312.5 10222.5 149377.5 ;
      RECT  9907.5 150930.0 9972.5 151115.0 ;
      RECT  9907.5 149770.0 9972.5 149955.0 ;
      RECT  9547.5 149887.5 9612.5 149737.5 ;
      RECT  9547.5 150772.5 9612.5 151147.5 ;
      RECT  9737.5 149887.5 9802.5 150772.5 ;
      RECT  9547.5 150772.5 9612.5 150907.5 ;
      RECT  9737.5 150772.5 9802.5 150907.5 ;
      RECT  9737.5 150772.5 9802.5 150907.5 ;
      RECT  9547.5 150772.5 9612.5 150907.5 ;
      RECT  9547.5 149887.5 9612.5 150022.5 ;
      RECT  9737.5 149887.5 9802.5 150022.5 ;
      RECT  9737.5 149887.5 9802.5 150022.5 ;
      RECT  9547.5 149887.5 9612.5 150022.5 ;
      RECT  9907.5 150862.5 9972.5 150997.5 ;
      RECT  9907.5 149887.5 9972.5 150022.5 ;
      RECT  9605.0 150330.0 9670.0 150465.0 ;
      RECT  9605.0 150330.0 9670.0 150465.0 ;
      RECT  9770.0 150365.0 9835.0 150430.0 ;
      RECT  9480.0 151082.5 10040.0 151147.5 ;
      RECT  9480.0 149737.5 10040.0 149802.5 ;
      RECT  10107.5 149932.5 10172.5 149737.5 ;
      RECT  10107.5 150772.5 10172.5 151147.5 ;
      RECT  10487.5 150772.5 10552.5 151147.5 ;
      RECT  10657.5 150930.0 10722.5 151115.0 ;
      RECT  10657.5 149770.0 10722.5 149955.0 ;
      RECT  10107.5 150772.5 10172.5 150907.5 ;
      RECT  10297.5 150772.5 10362.5 150907.5 ;
      RECT  10297.5 150772.5 10362.5 150907.5 ;
      RECT  10107.5 150772.5 10172.5 150907.5 ;
      RECT  10297.5 150772.5 10362.5 150907.5 ;
      RECT  10487.5 150772.5 10552.5 150907.5 ;
      RECT  10487.5 150772.5 10552.5 150907.5 ;
      RECT  10297.5 150772.5 10362.5 150907.5 ;
      RECT  10107.5 149932.5 10172.5 150067.5 ;
      RECT  10297.5 149932.5 10362.5 150067.5 ;
      RECT  10297.5 149932.5 10362.5 150067.5 ;
      RECT  10107.5 149932.5 10172.5 150067.5 ;
      RECT  10297.5 149932.5 10362.5 150067.5 ;
      RECT  10487.5 149932.5 10552.5 150067.5 ;
      RECT  10487.5 149932.5 10552.5 150067.5 ;
      RECT  10297.5 149932.5 10362.5 150067.5 ;
      RECT  10657.5 150862.5 10722.5 150997.5 ;
      RECT  10657.5 149887.5 10722.5 150022.5 ;
      RECT  10492.5 150162.5 10357.5 150227.5 ;
      RECT  10235.0 150377.5 10100.0 150442.5 ;
      RECT  10297.5 150772.5 10362.5 150907.5 ;
      RECT  10487.5 149932.5 10552.5 150067.5 ;
      RECT  10587.5 150377.5 10452.5 150442.5 ;
      RECT  10100.0 150377.5 10235.0 150442.5 ;
      RECT  10357.5 150162.5 10492.5 150227.5 ;
      RECT  10452.5 150377.5 10587.5 150442.5 ;
      RECT  10040.0 151082.5 10960.0 151147.5 ;
      RECT  10040.0 149737.5 10960.0 149802.5 ;
      RECT  11387.5 150930.0 11452.5 151115.0 ;
      RECT  11387.5 149770.0 11452.5 149955.0 ;
      RECT  11027.5 149887.5 11092.5 149737.5 ;
      RECT  11027.5 150772.5 11092.5 151147.5 ;
      RECT  11217.5 149887.5 11282.5 150772.5 ;
      RECT  11027.5 150772.5 11092.5 150907.5 ;
      RECT  11217.5 150772.5 11282.5 150907.5 ;
      RECT  11217.5 150772.5 11282.5 150907.5 ;
      RECT  11027.5 150772.5 11092.5 150907.5 ;
      RECT  11027.5 149887.5 11092.5 150022.5 ;
      RECT  11217.5 149887.5 11282.5 150022.5 ;
      RECT  11217.5 149887.5 11282.5 150022.5 ;
      RECT  11027.5 149887.5 11092.5 150022.5 ;
      RECT  11387.5 150862.5 11452.5 150997.5 ;
      RECT  11387.5 149887.5 11452.5 150022.5 ;
      RECT  11085.0 150330.0 11150.0 150465.0 ;
      RECT  11085.0 150330.0 11150.0 150465.0 ;
      RECT  11250.0 150365.0 11315.0 150430.0 ;
      RECT  10960.0 151082.5 11520.0 151147.5 ;
      RECT  10960.0 149737.5 11520.0 149802.5 ;
      RECT  9222.5 150330.0 9287.5 150465.0 ;
      RECT  9362.5 150057.5 9427.5 150192.5 ;
      RECT  10357.5 150162.5 10222.5 150227.5 ;
      RECT  9907.5 151300.0 9972.5 151115.0 ;
      RECT  9907.5 152460.0 9972.5 152275.0 ;
      RECT  9547.5 152342.5 9612.5 152492.5 ;
      RECT  9547.5 151457.5 9612.5 151082.5 ;
      RECT  9737.5 152342.5 9802.5 151457.5 ;
      RECT  9547.5 151457.5 9612.5 151322.5 ;
      RECT  9737.5 151457.5 9802.5 151322.5 ;
      RECT  9737.5 151457.5 9802.5 151322.5 ;
      RECT  9547.5 151457.5 9612.5 151322.5 ;
      RECT  9547.5 152342.5 9612.5 152207.5 ;
      RECT  9737.5 152342.5 9802.5 152207.5 ;
      RECT  9737.5 152342.5 9802.5 152207.5 ;
      RECT  9547.5 152342.5 9612.5 152207.5 ;
      RECT  9907.5 151367.5 9972.5 151232.5 ;
      RECT  9907.5 152342.5 9972.5 152207.5 ;
      RECT  9605.0 151900.0 9670.0 151765.0 ;
      RECT  9605.0 151900.0 9670.0 151765.0 ;
      RECT  9770.0 151865.0 9835.0 151800.0 ;
      RECT  9480.0 151147.5 10040.0 151082.5 ;
      RECT  9480.0 152492.5 10040.0 152427.5 ;
      RECT  10107.5 152297.5 10172.5 152492.5 ;
      RECT  10107.5 151457.5 10172.5 151082.5 ;
      RECT  10487.5 151457.5 10552.5 151082.5 ;
      RECT  10657.5 151300.0 10722.5 151115.0 ;
      RECT  10657.5 152460.0 10722.5 152275.0 ;
      RECT  10107.5 151457.5 10172.5 151322.5 ;
      RECT  10297.5 151457.5 10362.5 151322.5 ;
      RECT  10297.5 151457.5 10362.5 151322.5 ;
      RECT  10107.5 151457.5 10172.5 151322.5 ;
      RECT  10297.5 151457.5 10362.5 151322.5 ;
      RECT  10487.5 151457.5 10552.5 151322.5 ;
      RECT  10487.5 151457.5 10552.5 151322.5 ;
      RECT  10297.5 151457.5 10362.5 151322.5 ;
      RECT  10107.5 152297.5 10172.5 152162.5 ;
      RECT  10297.5 152297.5 10362.5 152162.5 ;
      RECT  10297.5 152297.5 10362.5 152162.5 ;
      RECT  10107.5 152297.5 10172.5 152162.5 ;
      RECT  10297.5 152297.5 10362.5 152162.5 ;
      RECT  10487.5 152297.5 10552.5 152162.5 ;
      RECT  10487.5 152297.5 10552.5 152162.5 ;
      RECT  10297.5 152297.5 10362.5 152162.5 ;
      RECT  10657.5 151367.5 10722.5 151232.5 ;
      RECT  10657.5 152342.5 10722.5 152207.5 ;
      RECT  10492.5 152067.5 10357.5 152002.5 ;
      RECT  10235.0 151852.5 10100.0 151787.5 ;
      RECT  10297.5 151457.5 10362.5 151322.5 ;
      RECT  10487.5 152297.5 10552.5 152162.5 ;
      RECT  10587.5 151852.5 10452.5 151787.5 ;
      RECT  10100.0 151852.5 10235.0 151787.5 ;
      RECT  10357.5 152067.5 10492.5 152002.5 ;
      RECT  10452.5 151852.5 10587.5 151787.5 ;
      RECT  10040.0 151147.5 10960.0 151082.5 ;
      RECT  10040.0 152492.5 10960.0 152427.5 ;
      RECT  11387.5 151300.0 11452.5 151115.0 ;
      RECT  11387.5 152460.0 11452.5 152275.0 ;
      RECT  11027.5 152342.5 11092.5 152492.5 ;
      RECT  11027.5 151457.5 11092.5 151082.5 ;
      RECT  11217.5 152342.5 11282.5 151457.5 ;
      RECT  11027.5 151457.5 11092.5 151322.5 ;
      RECT  11217.5 151457.5 11282.5 151322.5 ;
      RECT  11217.5 151457.5 11282.5 151322.5 ;
      RECT  11027.5 151457.5 11092.5 151322.5 ;
      RECT  11027.5 152342.5 11092.5 152207.5 ;
      RECT  11217.5 152342.5 11282.5 152207.5 ;
      RECT  11217.5 152342.5 11282.5 152207.5 ;
      RECT  11027.5 152342.5 11092.5 152207.5 ;
      RECT  11387.5 151367.5 11452.5 151232.5 ;
      RECT  11387.5 152342.5 11452.5 152207.5 ;
      RECT  11085.0 151900.0 11150.0 151765.0 ;
      RECT  11085.0 151900.0 11150.0 151765.0 ;
      RECT  11250.0 151865.0 11315.0 151800.0 ;
      RECT  10960.0 151147.5 11520.0 151082.5 ;
      RECT  10960.0 152492.5 11520.0 152427.5 ;
      RECT  9222.5 151765.0 9287.5 151900.0 ;
      RECT  9362.5 152037.5 9427.5 152172.5 ;
      RECT  10357.5 152002.5 10222.5 152067.5 ;
      RECT  9907.5 153620.0 9972.5 153805.0 ;
      RECT  9907.5 152460.0 9972.5 152645.0 ;
      RECT  9547.5 152577.5 9612.5 152427.5 ;
      RECT  9547.5 153462.5 9612.5 153837.5 ;
      RECT  9737.5 152577.5 9802.5 153462.5 ;
      RECT  9547.5 153462.5 9612.5 153597.5 ;
      RECT  9737.5 153462.5 9802.5 153597.5 ;
      RECT  9737.5 153462.5 9802.5 153597.5 ;
      RECT  9547.5 153462.5 9612.5 153597.5 ;
      RECT  9547.5 152577.5 9612.5 152712.5 ;
      RECT  9737.5 152577.5 9802.5 152712.5 ;
      RECT  9737.5 152577.5 9802.5 152712.5 ;
      RECT  9547.5 152577.5 9612.5 152712.5 ;
      RECT  9907.5 153552.5 9972.5 153687.5 ;
      RECT  9907.5 152577.5 9972.5 152712.5 ;
      RECT  9605.0 153020.0 9670.0 153155.0 ;
      RECT  9605.0 153020.0 9670.0 153155.0 ;
      RECT  9770.0 153055.0 9835.0 153120.0 ;
      RECT  9480.0 153772.5 10040.0 153837.5 ;
      RECT  9480.0 152427.5 10040.0 152492.5 ;
      RECT  10107.5 152622.5 10172.5 152427.5 ;
      RECT  10107.5 153462.5 10172.5 153837.5 ;
      RECT  10487.5 153462.5 10552.5 153837.5 ;
      RECT  10657.5 153620.0 10722.5 153805.0 ;
      RECT  10657.5 152460.0 10722.5 152645.0 ;
      RECT  10107.5 153462.5 10172.5 153597.5 ;
      RECT  10297.5 153462.5 10362.5 153597.5 ;
      RECT  10297.5 153462.5 10362.5 153597.5 ;
      RECT  10107.5 153462.5 10172.5 153597.5 ;
      RECT  10297.5 153462.5 10362.5 153597.5 ;
      RECT  10487.5 153462.5 10552.5 153597.5 ;
      RECT  10487.5 153462.5 10552.5 153597.5 ;
      RECT  10297.5 153462.5 10362.5 153597.5 ;
      RECT  10107.5 152622.5 10172.5 152757.5 ;
      RECT  10297.5 152622.5 10362.5 152757.5 ;
      RECT  10297.5 152622.5 10362.5 152757.5 ;
      RECT  10107.5 152622.5 10172.5 152757.5 ;
      RECT  10297.5 152622.5 10362.5 152757.5 ;
      RECT  10487.5 152622.5 10552.5 152757.5 ;
      RECT  10487.5 152622.5 10552.5 152757.5 ;
      RECT  10297.5 152622.5 10362.5 152757.5 ;
      RECT  10657.5 153552.5 10722.5 153687.5 ;
      RECT  10657.5 152577.5 10722.5 152712.5 ;
      RECT  10492.5 152852.5 10357.5 152917.5 ;
      RECT  10235.0 153067.5 10100.0 153132.5 ;
      RECT  10297.5 153462.5 10362.5 153597.5 ;
      RECT  10487.5 152622.5 10552.5 152757.5 ;
      RECT  10587.5 153067.5 10452.5 153132.5 ;
      RECT  10100.0 153067.5 10235.0 153132.5 ;
      RECT  10357.5 152852.5 10492.5 152917.5 ;
      RECT  10452.5 153067.5 10587.5 153132.5 ;
      RECT  10040.0 153772.5 10960.0 153837.5 ;
      RECT  10040.0 152427.5 10960.0 152492.5 ;
      RECT  11387.5 153620.0 11452.5 153805.0 ;
      RECT  11387.5 152460.0 11452.5 152645.0 ;
      RECT  11027.5 152577.5 11092.5 152427.5 ;
      RECT  11027.5 153462.5 11092.5 153837.5 ;
      RECT  11217.5 152577.5 11282.5 153462.5 ;
      RECT  11027.5 153462.5 11092.5 153597.5 ;
      RECT  11217.5 153462.5 11282.5 153597.5 ;
      RECT  11217.5 153462.5 11282.5 153597.5 ;
      RECT  11027.5 153462.5 11092.5 153597.5 ;
      RECT  11027.5 152577.5 11092.5 152712.5 ;
      RECT  11217.5 152577.5 11282.5 152712.5 ;
      RECT  11217.5 152577.5 11282.5 152712.5 ;
      RECT  11027.5 152577.5 11092.5 152712.5 ;
      RECT  11387.5 153552.5 11452.5 153687.5 ;
      RECT  11387.5 152577.5 11452.5 152712.5 ;
      RECT  11085.0 153020.0 11150.0 153155.0 ;
      RECT  11085.0 153020.0 11150.0 153155.0 ;
      RECT  11250.0 153055.0 11315.0 153120.0 ;
      RECT  10960.0 153772.5 11520.0 153837.5 ;
      RECT  10960.0 152427.5 11520.0 152492.5 ;
      RECT  9222.5 153020.0 9287.5 153155.0 ;
      RECT  9362.5 152747.5 9427.5 152882.5 ;
      RECT  10357.5 152852.5 10222.5 152917.5 ;
      RECT  9907.5 153990.0 9972.5 153805.0 ;
      RECT  9907.5 155150.0 9972.5 154965.0 ;
      RECT  9547.5 155032.5 9612.5 155182.5 ;
      RECT  9547.5 154147.5 9612.5 153772.5 ;
      RECT  9737.5 155032.5 9802.5 154147.5 ;
      RECT  9547.5 154147.5 9612.5 154012.5 ;
      RECT  9737.5 154147.5 9802.5 154012.5 ;
      RECT  9737.5 154147.5 9802.5 154012.5 ;
      RECT  9547.5 154147.5 9612.5 154012.5 ;
      RECT  9547.5 155032.5 9612.5 154897.5 ;
      RECT  9737.5 155032.5 9802.5 154897.5 ;
      RECT  9737.5 155032.5 9802.5 154897.5 ;
      RECT  9547.5 155032.5 9612.5 154897.5 ;
      RECT  9907.5 154057.5 9972.5 153922.5 ;
      RECT  9907.5 155032.5 9972.5 154897.5 ;
      RECT  9605.0 154590.0 9670.0 154455.0 ;
      RECT  9605.0 154590.0 9670.0 154455.0 ;
      RECT  9770.0 154555.0 9835.0 154490.0 ;
      RECT  9480.0 153837.5 10040.0 153772.5 ;
      RECT  9480.0 155182.5 10040.0 155117.5 ;
      RECT  10107.5 154987.5 10172.5 155182.5 ;
      RECT  10107.5 154147.5 10172.5 153772.5 ;
      RECT  10487.5 154147.5 10552.5 153772.5 ;
      RECT  10657.5 153990.0 10722.5 153805.0 ;
      RECT  10657.5 155150.0 10722.5 154965.0 ;
      RECT  10107.5 154147.5 10172.5 154012.5 ;
      RECT  10297.5 154147.5 10362.5 154012.5 ;
      RECT  10297.5 154147.5 10362.5 154012.5 ;
      RECT  10107.5 154147.5 10172.5 154012.5 ;
      RECT  10297.5 154147.5 10362.5 154012.5 ;
      RECT  10487.5 154147.5 10552.5 154012.5 ;
      RECT  10487.5 154147.5 10552.5 154012.5 ;
      RECT  10297.5 154147.5 10362.5 154012.5 ;
      RECT  10107.5 154987.5 10172.5 154852.5 ;
      RECT  10297.5 154987.5 10362.5 154852.5 ;
      RECT  10297.5 154987.5 10362.5 154852.5 ;
      RECT  10107.5 154987.5 10172.5 154852.5 ;
      RECT  10297.5 154987.5 10362.5 154852.5 ;
      RECT  10487.5 154987.5 10552.5 154852.5 ;
      RECT  10487.5 154987.5 10552.5 154852.5 ;
      RECT  10297.5 154987.5 10362.5 154852.5 ;
      RECT  10657.5 154057.5 10722.5 153922.5 ;
      RECT  10657.5 155032.5 10722.5 154897.5 ;
      RECT  10492.5 154757.5 10357.5 154692.5 ;
      RECT  10235.0 154542.5 10100.0 154477.5 ;
      RECT  10297.5 154147.5 10362.5 154012.5 ;
      RECT  10487.5 154987.5 10552.5 154852.5 ;
      RECT  10587.5 154542.5 10452.5 154477.5 ;
      RECT  10100.0 154542.5 10235.0 154477.5 ;
      RECT  10357.5 154757.5 10492.5 154692.5 ;
      RECT  10452.5 154542.5 10587.5 154477.5 ;
      RECT  10040.0 153837.5 10960.0 153772.5 ;
      RECT  10040.0 155182.5 10960.0 155117.5 ;
      RECT  11387.5 153990.0 11452.5 153805.0 ;
      RECT  11387.5 155150.0 11452.5 154965.0 ;
      RECT  11027.5 155032.5 11092.5 155182.5 ;
      RECT  11027.5 154147.5 11092.5 153772.5 ;
      RECT  11217.5 155032.5 11282.5 154147.5 ;
      RECT  11027.5 154147.5 11092.5 154012.5 ;
      RECT  11217.5 154147.5 11282.5 154012.5 ;
      RECT  11217.5 154147.5 11282.5 154012.5 ;
      RECT  11027.5 154147.5 11092.5 154012.5 ;
      RECT  11027.5 155032.5 11092.5 154897.5 ;
      RECT  11217.5 155032.5 11282.5 154897.5 ;
      RECT  11217.5 155032.5 11282.5 154897.5 ;
      RECT  11027.5 155032.5 11092.5 154897.5 ;
      RECT  11387.5 154057.5 11452.5 153922.5 ;
      RECT  11387.5 155032.5 11452.5 154897.5 ;
      RECT  11085.0 154590.0 11150.0 154455.0 ;
      RECT  11085.0 154590.0 11150.0 154455.0 ;
      RECT  11250.0 154555.0 11315.0 154490.0 ;
      RECT  10960.0 153837.5 11520.0 153772.5 ;
      RECT  10960.0 155182.5 11520.0 155117.5 ;
      RECT  9222.5 154455.0 9287.5 154590.0 ;
      RECT  9362.5 154727.5 9427.5 154862.5 ;
      RECT  10357.5 154692.5 10222.5 154757.5 ;
      RECT  9907.5 156310.0 9972.5 156495.0 ;
      RECT  9907.5 155150.0 9972.5 155335.0 ;
      RECT  9547.5 155267.5 9612.5 155117.5 ;
      RECT  9547.5 156152.5 9612.5 156527.5 ;
      RECT  9737.5 155267.5 9802.5 156152.5 ;
      RECT  9547.5 156152.5 9612.5 156287.5 ;
      RECT  9737.5 156152.5 9802.5 156287.5 ;
      RECT  9737.5 156152.5 9802.5 156287.5 ;
      RECT  9547.5 156152.5 9612.5 156287.5 ;
      RECT  9547.5 155267.5 9612.5 155402.5 ;
      RECT  9737.5 155267.5 9802.5 155402.5 ;
      RECT  9737.5 155267.5 9802.5 155402.5 ;
      RECT  9547.5 155267.5 9612.5 155402.5 ;
      RECT  9907.5 156242.5 9972.5 156377.5 ;
      RECT  9907.5 155267.5 9972.5 155402.5 ;
      RECT  9605.0 155710.0 9670.0 155845.0 ;
      RECT  9605.0 155710.0 9670.0 155845.0 ;
      RECT  9770.0 155745.0 9835.0 155810.0 ;
      RECT  9480.0 156462.5 10040.0 156527.5 ;
      RECT  9480.0 155117.5 10040.0 155182.5 ;
      RECT  10107.5 155312.5 10172.5 155117.5 ;
      RECT  10107.5 156152.5 10172.5 156527.5 ;
      RECT  10487.5 156152.5 10552.5 156527.5 ;
      RECT  10657.5 156310.0 10722.5 156495.0 ;
      RECT  10657.5 155150.0 10722.5 155335.0 ;
      RECT  10107.5 156152.5 10172.5 156287.5 ;
      RECT  10297.5 156152.5 10362.5 156287.5 ;
      RECT  10297.5 156152.5 10362.5 156287.5 ;
      RECT  10107.5 156152.5 10172.5 156287.5 ;
      RECT  10297.5 156152.5 10362.5 156287.5 ;
      RECT  10487.5 156152.5 10552.5 156287.5 ;
      RECT  10487.5 156152.5 10552.5 156287.5 ;
      RECT  10297.5 156152.5 10362.5 156287.5 ;
      RECT  10107.5 155312.5 10172.5 155447.5 ;
      RECT  10297.5 155312.5 10362.5 155447.5 ;
      RECT  10297.5 155312.5 10362.5 155447.5 ;
      RECT  10107.5 155312.5 10172.5 155447.5 ;
      RECT  10297.5 155312.5 10362.5 155447.5 ;
      RECT  10487.5 155312.5 10552.5 155447.5 ;
      RECT  10487.5 155312.5 10552.5 155447.5 ;
      RECT  10297.5 155312.5 10362.5 155447.5 ;
      RECT  10657.5 156242.5 10722.5 156377.5 ;
      RECT  10657.5 155267.5 10722.5 155402.5 ;
      RECT  10492.5 155542.5 10357.5 155607.5 ;
      RECT  10235.0 155757.5 10100.0 155822.5 ;
      RECT  10297.5 156152.5 10362.5 156287.5 ;
      RECT  10487.5 155312.5 10552.5 155447.5 ;
      RECT  10587.5 155757.5 10452.5 155822.5 ;
      RECT  10100.0 155757.5 10235.0 155822.5 ;
      RECT  10357.5 155542.5 10492.5 155607.5 ;
      RECT  10452.5 155757.5 10587.5 155822.5 ;
      RECT  10040.0 156462.5 10960.0 156527.5 ;
      RECT  10040.0 155117.5 10960.0 155182.5 ;
      RECT  11387.5 156310.0 11452.5 156495.0 ;
      RECT  11387.5 155150.0 11452.5 155335.0 ;
      RECT  11027.5 155267.5 11092.5 155117.5 ;
      RECT  11027.5 156152.5 11092.5 156527.5 ;
      RECT  11217.5 155267.5 11282.5 156152.5 ;
      RECT  11027.5 156152.5 11092.5 156287.5 ;
      RECT  11217.5 156152.5 11282.5 156287.5 ;
      RECT  11217.5 156152.5 11282.5 156287.5 ;
      RECT  11027.5 156152.5 11092.5 156287.5 ;
      RECT  11027.5 155267.5 11092.5 155402.5 ;
      RECT  11217.5 155267.5 11282.5 155402.5 ;
      RECT  11217.5 155267.5 11282.5 155402.5 ;
      RECT  11027.5 155267.5 11092.5 155402.5 ;
      RECT  11387.5 156242.5 11452.5 156377.5 ;
      RECT  11387.5 155267.5 11452.5 155402.5 ;
      RECT  11085.0 155710.0 11150.0 155845.0 ;
      RECT  11085.0 155710.0 11150.0 155845.0 ;
      RECT  11250.0 155745.0 11315.0 155810.0 ;
      RECT  10960.0 156462.5 11520.0 156527.5 ;
      RECT  10960.0 155117.5 11520.0 155182.5 ;
      RECT  9222.5 155710.0 9287.5 155845.0 ;
      RECT  9362.5 155437.5 9427.5 155572.5 ;
      RECT  10357.5 155542.5 10222.5 155607.5 ;
      RECT  9907.5 156680.0 9972.5 156495.0 ;
      RECT  9907.5 157840.0 9972.5 157655.0 ;
      RECT  9547.5 157722.5 9612.5 157872.5 ;
      RECT  9547.5 156837.5 9612.5 156462.5 ;
      RECT  9737.5 157722.5 9802.5 156837.5 ;
      RECT  9547.5 156837.5 9612.5 156702.5 ;
      RECT  9737.5 156837.5 9802.5 156702.5 ;
      RECT  9737.5 156837.5 9802.5 156702.5 ;
      RECT  9547.5 156837.5 9612.5 156702.5 ;
      RECT  9547.5 157722.5 9612.5 157587.5 ;
      RECT  9737.5 157722.5 9802.5 157587.5 ;
      RECT  9737.5 157722.5 9802.5 157587.5 ;
      RECT  9547.5 157722.5 9612.5 157587.5 ;
      RECT  9907.5 156747.5 9972.5 156612.5 ;
      RECT  9907.5 157722.5 9972.5 157587.5 ;
      RECT  9605.0 157280.0 9670.0 157145.0 ;
      RECT  9605.0 157280.0 9670.0 157145.0 ;
      RECT  9770.0 157245.0 9835.0 157180.0 ;
      RECT  9480.0 156527.5 10040.0 156462.5 ;
      RECT  9480.0 157872.5 10040.0 157807.5 ;
      RECT  10107.5 157677.5 10172.5 157872.5 ;
      RECT  10107.5 156837.5 10172.5 156462.5 ;
      RECT  10487.5 156837.5 10552.5 156462.5 ;
      RECT  10657.5 156680.0 10722.5 156495.0 ;
      RECT  10657.5 157840.0 10722.5 157655.0 ;
      RECT  10107.5 156837.5 10172.5 156702.5 ;
      RECT  10297.5 156837.5 10362.5 156702.5 ;
      RECT  10297.5 156837.5 10362.5 156702.5 ;
      RECT  10107.5 156837.5 10172.5 156702.5 ;
      RECT  10297.5 156837.5 10362.5 156702.5 ;
      RECT  10487.5 156837.5 10552.5 156702.5 ;
      RECT  10487.5 156837.5 10552.5 156702.5 ;
      RECT  10297.5 156837.5 10362.5 156702.5 ;
      RECT  10107.5 157677.5 10172.5 157542.5 ;
      RECT  10297.5 157677.5 10362.5 157542.5 ;
      RECT  10297.5 157677.5 10362.5 157542.5 ;
      RECT  10107.5 157677.5 10172.5 157542.5 ;
      RECT  10297.5 157677.5 10362.5 157542.5 ;
      RECT  10487.5 157677.5 10552.5 157542.5 ;
      RECT  10487.5 157677.5 10552.5 157542.5 ;
      RECT  10297.5 157677.5 10362.5 157542.5 ;
      RECT  10657.5 156747.5 10722.5 156612.5 ;
      RECT  10657.5 157722.5 10722.5 157587.5 ;
      RECT  10492.5 157447.5 10357.5 157382.5 ;
      RECT  10235.0 157232.5 10100.0 157167.5 ;
      RECT  10297.5 156837.5 10362.5 156702.5 ;
      RECT  10487.5 157677.5 10552.5 157542.5 ;
      RECT  10587.5 157232.5 10452.5 157167.5 ;
      RECT  10100.0 157232.5 10235.0 157167.5 ;
      RECT  10357.5 157447.5 10492.5 157382.5 ;
      RECT  10452.5 157232.5 10587.5 157167.5 ;
      RECT  10040.0 156527.5 10960.0 156462.5 ;
      RECT  10040.0 157872.5 10960.0 157807.5 ;
      RECT  11387.5 156680.0 11452.5 156495.0 ;
      RECT  11387.5 157840.0 11452.5 157655.0 ;
      RECT  11027.5 157722.5 11092.5 157872.5 ;
      RECT  11027.5 156837.5 11092.5 156462.5 ;
      RECT  11217.5 157722.5 11282.5 156837.5 ;
      RECT  11027.5 156837.5 11092.5 156702.5 ;
      RECT  11217.5 156837.5 11282.5 156702.5 ;
      RECT  11217.5 156837.5 11282.5 156702.5 ;
      RECT  11027.5 156837.5 11092.5 156702.5 ;
      RECT  11027.5 157722.5 11092.5 157587.5 ;
      RECT  11217.5 157722.5 11282.5 157587.5 ;
      RECT  11217.5 157722.5 11282.5 157587.5 ;
      RECT  11027.5 157722.5 11092.5 157587.5 ;
      RECT  11387.5 156747.5 11452.5 156612.5 ;
      RECT  11387.5 157722.5 11452.5 157587.5 ;
      RECT  11085.0 157280.0 11150.0 157145.0 ;
      RECT  11085.0 157280.0 11150.0 157145.0 ;
      RECT  11250.0 157245.0 11315.0 157180.0 ;
      RECT  10960.0 156527.5 11520.0 156462.5 ;
      RECT  10960.0 157872.5 11520.0 157807.5 ;
      RECT  9222.5 157145.0 9287.5 157280.0 ;
      RECT  9362.5 157417.5 9427.5 157552.5 ;
      RECT  10357.5 157382.5 10222.5 157447.5 ;
      RECT  9907.5 159000.0 9972.5 159185.0 ;
      RECT  9907.5 157840.0 9972.5 158025.0 ;
      RECT  9547.5 157957.5 9612.5 157807.5 ;
      RECT  9547.5 158842.5 9612.5 159217.5 ;
      RECT  9737.5 157957.5 9802.5 158842.5 ;
      RECT  9547.5 158842.5 9612.5 158977.5 ;
      RECT  9737.5 158842.5 9802.5 158977.5 ;
      RECT  9737.5 158842.5 9802.5 158977.5 ;
      RECT  9547.5 158842.5 9612.5 158977.5 ;
      RECT  9547.5 157957.5 9612.5 158092.5 ;
      RECT  9737.5 157957.5 9802.5 158092.5 ;
      RECT  9737.5 157957.5 9802.5 158092.5 ;
      RECT  9547.5 157957.5 9612.5 158092.5 ;
      RECT  9907.5 158932.5 9972.5 159067.5 ;
      RECT  9907.5 157957.5 9972.5 158092.5 ;
      RECT  9605.0 158400.0 9670.0 158535.0 ;
      RECT  9605.0 158400.0 9670.0 158535.0 ;
      RECT  9770.0 158435.0 9835.0 158500.0 ;
      RECT  9480.0 159152.5 10040.0 159217.5 ;
      RECT  9480.0 157807.5 10040.0 157872.5 ;
      RECT  10107.5 158002.5 10172.5 157807.5 ;
      RECT  10107.5 158842.5 10172.5 159217.5 ;
      RECT  10487.5 158842.5 10552.5 159217.5 ;
      RECT  10657.5 159000.0 10722.5 159185.0 ;
      RECT  10657.5 157840.0 10722.5 158025.0 ;
      RECT  10107.5 158842.5 10172.5 158977.5 ;
      RECT  10297.5 158842.5 10362.5 158977.5 ;
      RECT  10297.5 158842.5 10362.5 158977.5 ;
      RECT  10107.5 158842.5 10172.5 158977.5 ;
      RECT  10297.5 158842.5 10362.5 158977.5 ;
      RECT  10487.5 158842.5 10552.5 158977.5 ;
      RECT  10487.5 158842.5 10552.5 158977.5 ;
      RECT  10297.5 158842.5 10362.5 158977.5 ;
      RECT  10107.5 158002.5 10172.5 158137.5 ;
      RECT  10297.5 158002.5 10362.5 158137.5 ;
      RECT  10297.5 158002.5 10362.5 158137.5 ;
      RECT  10107.5 158002.5 10172.5 158137.5 ;
      RECT  10297.5 158002.5 10362.5 158137.5 ;
      RECT  10487.5 158002.5 10552.5 158137.5 ;
      RECT  10487.5 158002.5 10552.5 158137.5 ;
      RECT  10297.5 158002.5 10362.5 158137.5 ;
      RECT  10657.5 158932.5 10722.5 159067.5 ;
      RECT  10657.5 157957.5 10722.5 158092.5 ;
      RECT  10492.5 158232.5 10357.5 158297.5 ;
      RECT  10235.0 158447.5 10100.0 158512.5 ;
      RECT  10297.5 158842.5 10362.5 158977.5 ;
      RECT  10487.5 158002.5 10552.5 158137.5 ;
      RECT  10587.5 158447.5 10452.5 158512.5 ;
      RECT  10100.0 158447.5 10235.0 158512.5 ;
      RECT  10357.5 158232.5 10492.5 158297.5 ;
      RECT  10452.5 158447.5 10587.5 158512.5 ;
      RECT  10040.0 159152.5 10960.0 159217.5 ;
      RECT  10040.0 157807.5 10960.0 157872.5 ;
      RECT  11387.5 159000.0 11452.5 159185.0 ;
      RECT  11387.5 157840.0 11452.5 158025.0 ;
      RECT  11027.5 157957.5 11092.5 157807.5 ;
      RECT  11027.5 158842.5 11092.5 159217.5 ;
      RECT  11217.5 157957.5 11282.5 158842.5 ;
      RECT  11027.5 158842.5 11092.5 158977.5 ;
      RECT  11217.5 158842.5 11282.5 158977.5 ;
      RECT  11217.5 158842.5 11282.5 158977.5 ;
      RECT  11027.5 158842.5 11092.5 158977.5 ;
      RECT  11027.5 157957.5 11092.5 158092.5 ;
      RECT  11217.5 157957.5 11282.5 158092.5 ;
      RECT  11217.5 157957.5 11282.5 158092.5 ;
      RECT  11027.5 157957.5 11092.5 158092.5 ;
      RECT  11387.5 158932.5 11452.5 159067.5 ;
      RECT  11387.5 157957.5 11452.5 158092.5 ;
      RECT  11085.0 158400.0 11150.0 158535.0 ;
      RECT  11085.0 158400.0 11150.0 158535.0 ;
      RECT  11250.0 158435.0 11315.0 158500.0 ;
      RECT  10960.0 159152.5 11520.0 159217.5 ;
      RECT  10960.0 157807.5 11520.0 157872.5 ;
      RECT  9222.5 158400.0 9287.5 158535.0 ;
      RECT  9362.5 158127.5 9427.5 158262.5 ;
      RECT  10357.5 158232.5 10222.5 158297.5 ;
      RECT  9907.5 159370.0 9972.5 159185.0 ;
      RECT  9907.5 160530.0 9972.5 160345.0 ;
      RECT  9547.5 160412.5 9612.5 160562.5 ;
      RECT  9547.5 159527.5 9612.5 159152.5 ;
      RECT  9737.5 160412.5 9802.5 159527.5 ;
      RECT  9547.5 159527.5 9612.5 159392.5 ;
      RECT  9737.5 159527.5 9802.5 159392.5 ;
      RECT  9737.5 159527.5 9802.5 159392.5 ;
      RECT  9547.5 159527.5 9612.5 159392.5 ;
      RECT  9547.5 160412.5 9612.5 160277.5 ;
      RECT  9737.5 160412.5 9802.5 160277.5 ;
      RECT  9737.5 160412.5 9802.5 160277.5 ;
      RECT  9547.5 160412.5 9612.5 160277.5 ;
      RECT  9907.5 159437.5 9972.5 159302.5 ;
      RECT  9907.5 160412.5 9972.5 160277.5 ;
      RECT  9605.0 159970.0 9670.0 159835.0 ;
      RECT  9605.0 159970.0 9670.0 159835.0 ;
      RECT  9770.0 159935.0 9835.0 159870.0 ;
      RECT  9480.0 159217.5 10040.0 159152.5 ;
      RECT  9480.0 160562.5 10040.0 160497.5 ;
      RECT  10107.5 160367.5 10172.5 160562.5 ;
      RECT  10107.5 159527.5 10172.5 159152.5 ;
      RECT  10487.5 159527.5 10552.5 159152.5 ;
      RECT  10657.5 159370.0 10722.5 159185.0 ;
      RECT  10657.5 160530.0 10722.5 160345.0 ;
      RECT  10107.5 159527.5 10172.5 159392.5 ;
      RECT  10297.5 159527.5 10362.5 159392.5 ;
      RECT  10297.5 159527.5 10362.5 159392.5 ;
      RECT  10107.5 159527.5 10172.5 159392.5 ;
      RECT  10297.5 159527.5 10362.5 159392.5 ;
      RECT  10487.5 159527.5 10552.5 159392.5 ;
      RECT  10487.5 159527.5 10552.5 159392.5 ;
      RECT  10297.5 159527.5 10362.5 159392.5 ;
      RECT  10107.5 160367.5 10172.5 160232.5 ;
      RECT  10297.5 160367.5 10362.5 160232.5 ;
      RECT  10297.5 160367.5 10362.5 160232.5 ;
      RECT  10107.5 160367.5 10172.5 160232.5 ;
      RECT  10297.5 160367.5 10362.5 160232.5 ;
      RECT  10487.5 160367.5 10552.5 160232.5 ;
      RECT  10487.5 160367.5 10552.5 160232.5 ;
      RECT  10297.5 160367.5 10362.5 160232.5 ;
      RECT  10657.5 159437.5 10722.5 159302.5 ;
      RECT  10657.5 160412.5 10722.5 160277.5 ;
      RECT  10492.5 160137.5 10357.5 160072.5 ;
      RECT  10235.0 159922.5 10100.0 159857.5 ;
      RECT  10297.5 159527.5 10362.5 159392.5 ;
      RECT  10487.5 160367.5 10552.5 160232.5 ;
      RECT  10587.5 159922.5 10452.5 159857.5 ;
      RECT  10100.0 159922.5 10235.0 159857.5 ;
      RECT  10357.5 160137.5 10492.5 160072.5 ;
      RECT  10452.5 159922.5 10587.5 159857.5 ;
      RECT  10040.0 159217.5 10960.0 159152.5 ;
      RECT  10040.0 160562.5 10960.0 160497.5 ;
      RECT  11387.5 159370.0 11452.5 159185.0 ;
      RECT  11387.5 160530.0 11452.5 160345.0 ;
      RECT  11027.5 160412.5 11092.5 160562.5 ;
      RECT  11027.5 159527.5 11092.5 159152.5 ;
      RECT  11217.5 160412.5 11282.5 159527.5 ;
      RECT  11027.5 159527.5 11092.5 159392.5 ;
      RECT  11217.5 159527.5 11282.5 159392.5 ;
      RECT  11217.5 159527.5 11282.5 159392.5 ;
      RECT  11027.5 159527.5 11092.5 159392.5 ;
      RECT  11027.5 160412.5 11092.5 160277.5 ;
      RECT  11217.5 160412.5 11282.5 160277.5 ;
      RECT  11217.5 160412.5 11282.5 160277.5 ;
      RECT  11027.5 160412.5 11092.5 160277.5 ;
      RECT  11387.5 159437.5 11452.5 159302.5 ;
      RECT  11387.5 160412.5 11452.5 160277.5 ;
      RECT  11085.0 159970.0 11150.0 159835.0 ;
      RECT  11085.0 159970.0 11150.0 159835.0 ;
      RECT  11250.0 159935.0 11315.0 159870.0 ;
      RECT  10960.0 159217.5 11520.0 159152.5 ;
      RECT  10960.0 160562.5 11520.0 160497.5 ;
      RECT  9222.5 159835.0 9287.5 159970.0 ;
      RECT  9362.5 160107.5 9427.5 160242.5 ;
      RECT  10357.5 160072.5 10222.5 160137.5 ;
      RECT  9907.5 161690.0 9972.5 161875.0 ;
      RECT  9907.5 160530.0 9972.5 160715.0 ;
      RECT  9547.5 160647.5 9612.5 160497.5 ;
      RECT  9547.5 161532.5 9612.5 161907.5 ;
      RECT  9737.5 160647.5 9802.5 161532.5 ;
      RECT  9547.5 161532.5 9612.5 161667.5 ;
      RECT  9737.5 161532.5 9802.5 161667.5 ;
      RECT  9737.5 161532.5 9802.5 161667.5 ;
      RECT  9547.5 161532.5 9612.5 161667.5 ;
      RECT  9547.5 160647.5 9612.5 160782.5 ;
      RECT  9737.5 160647.5 9802.5 160782.5 ;
      RECT  9737.5 160647.5 9802.5 160782.5 ;
      RECT  9547.5 160647.5 9612.5 160782.5 ;
      RECT  9907.5 161622.5 9972.5 161757.5 ;
      RECT  9907.5 160647.5 9972.5 160782.5 ;
      RECT  9605.0 161090.0 9670.0 161225.0 ;
      RECT  9605.0 161090.0 9670.0 161225.0 ;
      RECT  9770.0 161125.0 9835.0 161190.0 ;
      RECT  9480.0 161842.5 10040.0 161907.5 ;
      RECT  9480.0 160497.5 10040.0 160562.5 ;
      RECT  10107.5 160692.5 10172.5 160497.5 ;
      RECT  10107.5 161532.5 10172.5 161907.5 ;
      RECT  10487.5 161532.5 10552.5 161907.5 ;
      RECT  10657.5 161690.0 10722.5 161875.0 ;
      RECT  10657.5 160530.0 10722.5 160715.0 ;
      RECT  10107.5 161532.5 10172.5 161667.5 ;
      RECT  10297.5 161532.5 10362.5 161667.5 ;
      RECT  10297.5 161532.5 10362.5 161667.5 ;
      RECT  10107.5 161532.5 10172.5 161667.5 ;
      RECT  10297.5 161532.5 10362.5 161667.5 ;
      RECT  10487.5 161532.5 10552.5 161667.5 ;
      RECT  10487.5 161532.5 10552.5 161667.5 ;
      RECT  10297.5 161532.5 10362.5 161667.5 ;
      RECT  10107.5 160692.5 10172.5 160827.5 ;
      RECT  10297.5 160692.5 10362.5 160827.5 ;
      RECT  10297.5 160692.5 10362.5 160827.5 ;
      RECT  10107.5 160692.5 10172.5 160827.5 ;
      RECT  10297.5 160692.5 10362.5 160827.5 ;
      RECT  10487.5 160692.5 10552.5 160827.5 ;
      RECT  10487.5 160692.5 10552.5 160827.5 ;
      RECT  10297.5 160692.5 10362.5 160827.5 ;
      RECT  10657.5 161622.5 10722.5 161757.5 ;
      RECT  10657.5 160647.5 10722.5 160782.5 ;
      RECT  10492.5 160922.5 10357.5 160987.5 ;
      RECT  10235.0 161137.5 10100.0 161202.5 ;
      RECT  10297.5 161532.5 10362.5 161667.5 ;
      RECT  10487.5 160692.5 10552.5 160827.5 ;
      RECT  10587.5 161137.5 10452.5 161202.5 ;
      RECT  10100.0 161137.5 10235.0 161202.5 ;
      RECT  10357.5 160922.5 10492.5 160987.5 ;
      RECT  10452.5 161137.5 10587.5 161202.5 ;
      RECT  10040.0 161842.5 10960.0 161907.5 ;
      RECT  10040.0 160497.5 10960.0 160562.5 ;
      RECT  11387.5 161690.0 11452.5 161875.0 ;
      RECT  11387.5 160530.0 11452.5 160715.0 ;
      RECT  11027.5 160647.5 11092.5 160497.5 ;
      RECT  11027.5 161532.5 11092.5 161907.5 ;
      RECT  11217.5 160647.5 11282.5 161532.5 ;
      RECT  11027.5 161532.5 11092.5 161667.5 ;
      RECT  11217.5 161532.5 11282.5 161667.5 ;
      RECT  11217.5 161532.5 11282.5 161667.5 ;
      RECT  11027.5 161532.5 11092.5 161667.5 ;
      RECT  11027.5 160647.5 11092.5 160782.5 ;
      RECT  11217.5 160647.5 11282.5 160782.5 ;
      RECT  11217.5 160647.5 11282.5 160782.5 ;
      RECT  11027.5 160647.5 11092.5 160782.5 ;
      RECT  11387.5 161622.5 11452.5 161757.5 ;
      RECT  11387.5 160647.5 11452.5 160782.5 ;
      RECT  11085.0 161090.0 11150.0 161225.0 ;
      RECT  11085.0 161090.0 11150.0 161225.0 ;
      RECT  11250.0 161125.0 11315.0 161190.0 ;
      RECT  10960.0 161842.5 11520.0 161907.5 ;
      RECT  10960.0 160497.5 11520.0 160562.5 ;
      RECT  9222.5 161090.0 9287.5 161225.0 ;
      RECT  9362.5 160817.5 9427.5 160952.5 ;
      RECT  10357.5 160922.5 10222.5 160987.5 ;
      RECT  9907.5 162060.0 9972.5 161875.0 ;
      RECT  9907.5 163220.0 9972.5 163035.0 ;
      RECT  9547.5 163102.5 9612.5 163252.5 ;
      RECT  9547.5 162217.5 9612.5 161842.5 ;
      RECT  9737.5 163102.5 9802.5 162217.5 ;
      RECT  9547.5 162217.5 9612.5 162082.5 ;
      RECT  9737.5 162217.5 9802.5 162082.5 ;
      RECT  9737.5 162217.5 9802.5 162082.5 ;
      RECT  9547.5 162217.5 9612.5 162082.5 ;
      RECT  9547.5 163102.5 9612.5 162967.5 ;
      RECT  9737.5 163102.5 9802.5 162967.5 ;
      RECT  9737.5 163102.5 9802.5 162967.5 ;
      RECT  9547.5 163102.5 9612.5 162967.5 ;
      RECT  9907.5 162127.5 9972.5 161992.5 ;
      RECT  9907.5 163102.5 9972.5 162967.5 ;
      RECT  9605.0 162660.0 9670.0 162525.0 ;
      RECT  9605.0 162660.0 9670.0 162525.0 ;
      RECT  9770.0 162625.0 9835.0 162560.0 ;
      RECT  9480.0 161907.5 10040.0 161842.5 ;
      RECT  9480.0 163252.5 10040.0 163187.5 ;
      RECT  10107.5 163057.5 10172.5 163252.5 ;
      RECT  10107.5 162217.5 10172.5 161842.5 ;
      RECT  10487.5 162217.5 10552.5 161842.5 ;
      RECT  10657.5 162060.0 10722.5 161875.0 ;
      RECT  10657.5 163220.0 10722.5 163035.0 ;
      RECT  10107.5 162217.5 10172.5 162082.5 ;
      RECT  10297.5 162217.5 10362.5 162082.5 ;
      RECT  10297.5 162217.5 10362.5 162082.5 ;
      RECT  10107.5 162217.5 10172.5 162082.5 ;
      RECT  10297.5 162217.5 10362.5 162082.5 ;
      RECT  10487.5 162217.5 10552.5 162082.5 ;
      RECT  10487.5 162217.5 10552.5 162082.5 ;
      RECT  10297.5 162217.5 10362.5 162082.5 ;
      RECT  10107.5 163057.5 10172.5 162922.5 ;
      RECT  10297.5 163057.5 10362.5 162922.5 ;
      RECT  10297.5 163057.5 10362.5 162922.5 ;
      RECT  10107.5 163057.5 10172.5 162922.5 ;
      RECT  10297.5 163057.5 10362.5 162922.5 ;
      RECT  10487.5 163057.5 10552.5 162922.5 ;
      RECT  10487.5 163057.5 10552.5 162922.5 ;
      RECT  10297.5 163057.5 10362.5 162922.5 ;
      RECT  10657.5 162127.5 10722.5 161992.5 ;
      RECT  10657.5 163102.5 10722.5 162967.5 ;
      RECT  10492.5 162827.5 10357.5 162762.5 ;
      RECT  10235.0 162612.5 10100.0 162547.5 ;
      RECT  10297.5 162217.5 10362.5 162082.5 ;
      RECT  10487.5 163057.5 10552.5 162922.5 ;
      RECT  10587.5 162612.5 10452.5 162547.5 ;
      RECT  10100.0 162612.5 10235.0 162547.5 ;
      RECT  10357.5 162827.5 10492.5 162762.5 ;
      RECT  10452.5 162612.5 10587.5 162547.5 ;
      RECT  10040.0 161907.5 10960.0 161842.5 ;
      RECT  10040.0 163252.5 10960.0 163187.5 ;
      RECT  11387.5 162060.0 11452.5 161875.0 ;
      RECT  11387.5 163220.0 11452.5 163035.0 ;
      RECT  11027.5 163102.5 11092.5 163252.5 ;
      RECT  11027.5 162217.5 11092.5 161842.5 ;
      RECT  11217.5 163102.5 11282.5 162217.5 ;
      RECT  11027.5 162217.5 11092.5 162082.5 ;
      RECT  11217.5 162217.5 11282.5 162082.5 ;
      RECT  11217.5 162217.5 11282.5 162082.5 ;
      RECT  11027.5 162217.5 11092.5 162082.5 ;
      RECT  11027.5 163102.5 11092.5 162967.5 ;
      RECT  11217.5 163102.5 11282.5 162967.5 ;
      RECT  11217.5 163102.5 11282.5 162967.5 ;
      RECT  11027.5 163102.5 11092.5 162967.5 ;
      RECT  11387.5 162127.5 11452.5 161992.5 ;
      RECT  11387.5 163102.5 11452.5 162967.5 ;
      RECT  11085.0 162660.0 11150.0 162525.0 ;
      RECT  11085.0 162660.0 11150.0 162525.0 ;
      RECT  11250.0 162625.0 11315.0 162560.0 ;
      RECT  10960.0 161907.5 11520.0 161842.5 ;
      RECT  10960.0 163252.5 11520.0 163187.5 ;
      RECT  9222.5 162525.0 9287.5 162660.0 ;
      RECT  9362.5 162797.5 9427.5 162932.5 ;
      RECT  10357.5 162762.5 10222.5 162827.5 ;
      RECT  9907.5 164380.0 9972.5 164565.0 ;
      RECT  9907.5 163220.0 9972.5 163405.0 ;
      RECT  9547.5 163337.5 9612.5 163187.5 ;
      RECT  9547.5 164222.5 9612.5 164597.5 ;
      RECT  9737.5 163337.5 9802.5 164222.5 ;
      RECT  9547.5 164222.5 9612.5 164357.5 ;
      RECT  9737.5 164222.5 9802.5 164357.5 ;
      RECT  9737.5 164222.5 9802.5 164357.5 ;
      RECT  9547.5 164222.5 9612.5 164357.5 ;
      RECT  9547.5 163337.5 9612.5 163472.5 ;
      RECT  9737.5 163337.5 9802.5 163472.5 ;
      RECT  9737.5 163337.5 9802.5 163472.5 ;
      RECT  9547.5 163337.5 9612.5 163472.5 ;
      RECT  9907.5 164312.5 9972.5 164447.5 ;
      RECT  9907.5 163337.5 9972.5 163472.5 ;
      RECT  9605.0 163780.0 9670.0 163915.0 ;
      RECT  9605.0 163780.0 9670.0 163915.0 ;
      RECT  9770.0 163815.0 9835.0 163880.0 ;
      RECT  9480.0 164532.5 10040.0 164597.5 ;
      RECT  9480.0 163187.5 10040.0 163252.5 ;
      RECT  10107.5 163382.5 10172.5 163187.5 ;
      RECT  10107.5 164222.5 10172.5 164597.5 ;
      RECT  10487.5 164222.5 10552.5 164597.5 ;
      RECT  10657.5 164380.0 10722.5 164565.0 ;
      RECT  10657.5 163220.0 10722.5 163405.0 ;
      RECT  10107.5 164222.5 10172.5 164357.5 ;
      RECT  10297.5 164222.5 10362.5 164357.5 ;
      RECT  10297.5 164222.5 10362.5 164357.5 ;
      RECT  10107.5 164222.5 10172.5 164357.5 ;
      RECT  10297.5 164222.5 10362.5 164357.5 ;
      RECT  10487.5 164222.5 10552.5 164357.5 ;
      RECT  10487.5 164222.5 10552.5 164357.5 ;
      RECT  10297.5 164222.5 10362.5 164357.5 ;
      RECT  10107.5 163382.5 10172.5 163517.5 ;
      RECT  10297.5 163382.5 10362.5 163517.5 ;
      RECT  10297.5 163382.5 10362.5 163517.5 ;
      RECT  10107.5 163382.5 10172.5 163517.5 ;
      RECT  10297.5 163382.5 10362.5 163517.5 ;
      RECT  10487.5 163382.5 10552.5 163517.5 ;
      RECT  10487.5 163382.5 10552.5 163517.5 ;
      RECT  10297.5 163382.5 10362.5 163517.5 ;
      RECT  10657.5 164312.5 10722.5 164447.5 ;
      RECT  10657.5 163337.5 10722.5 163472.5 ;
      RECT  10492.5 163612.5 10357.5 163677.5 ;
      RECT  10235.0 163827.5 10100.0 163892.5 ;
      RECT  10297.5 164222.5 10362.5 164357.5 ;
      RECT  10487.5 163382.5 10552.5 163517.5 ;
      RECT  10587.5 163827.5 10452.5 163892.5 ;
      RECT  10100.0 163827.5 10235.0 163892.5 ;
      RECT  10357.5 163612.5 10492.5 163677.5 ;
      RECT  10452.5 163827.5 10587.5 163892.5 ;
      RECT  10040.0 164532.5 10960.0 164597.5 ;
      RECT  10040.0 163187.5 10960.0 163252.5 ;
      RECT  11387.5 164380.0 11452.5 164565.0 ;
      RECT  11387.5 163220.0 11452.5 163405.0 ;
      RECT  11027.5 163337.5 11092.5 163187.5 ;
      RECT  11027.5 164222.5 11092.5 164597.5 ;
      RECT  11217.5 163337.5 11282.5 164222.5 ;
      RECT  11027.5 164222.5 11092.5 164357.5 ;
      RECT  11217.5 164222.5 11282.5 164357.5 ;
      RECT  11217.5 164222.5 11282.5 164357.5 ;
      RECT  11027.5 164222.5 11092.5 164357.5 ;
      RECT  11027.5 163337.5 11092.5 163472.5 ;
      RECT  11217.5 163337.5 11282.5 163472.5 ;
      RECT  11217.5 163337.5 11282.5 163472.5 ;
      RECT  11027.5 163337.5 11092.5 163472.5 ;
      RECT  11387.5 164312.5 11452.5 164447.5 ;
      RECT  11387.5 163337.5 11452.5 163472.5 ;
      RECT  11085.0 163780.0 11150.0 163915.0 ;
      RECT  11085.0 163780.0 11150.0 163915.0 ;
      RECT  11250.0 163815.0 11315.0 163880.0 ;
      RECT  10960.0 164532.5 11520.0 164597.5 ;
      RECT  10960.0 163187.5 11520.0 163252.5 ;
      RECT  9222.5 163780.0 9287.5 163915.0 ;
      RECT  9362.5 163507.5 9427.5 163642.5 ;
      RECT  10357.5 163612.5 10222.5 163677.5 ;
      RECT  9907.5 164750.0 9972.5 164565.0 ;
      RECT  9907.5 165910.0 9972.5 165725.0 ;
      RECT  9547.5 165792.5 9612.5 165942.5 ;
      RECT  9547.5 164907.5 9612.5 164532.5 ;
      RECT  9737.5 165792.5 9802.5 164907.5 ;
      RECT  9547.5 164907.5 9612.5 164772.5 ;
      RECT  9737.5 164907.5 9802.5 164772.5 ;
      RECT  9737.5 164907.5 9802.5 164772.5 ;
      RECT  9547.5 164907.5 9612.5 164772.5 ;
      RECT  9547.5 165792.5 9612.5 165657.5 ;
      RECT  9737.5 165792.5 9802.5 165657.5 ;
      RECT  9737.5 165792.5 9802.5 165657.5 ;
      RECT  9547.5 165792.5 9612.5 165657.5 ;
      RECT  9907.5 164817.5 9972.5 164682.5 ;
      RECT  9907.5 165792.5 9972.5 165657.5 ;
      RECT  9605.0 165350.0 9670.0 165215.0 ;
      RECT  9605.0 165350.0 9670.0 165215.0 ;
      RECT  9770.0 165315.0 9835.0 165250.0 ;
      RECT  9480.0 164597.5 10040.0 164532.5 ;
      RECT  9480.0 165942.5 10040.0 165877.5 ;
      RECT  10107.5 165747.5 10172.5 165942.5 ;
      RECT  10107.5 164907.5 10172.5 164532.5 ;
      RECT  10487.5 164907.5 10552.5 164532.5 ;
      RECT  10657.5 164750.0 10722.5 164565.0 ;
      RECT  10657.5 165910.0 10722.5 165725.0 ;
      RECT  10107.5 164907.5 10172.5 164772.5 ;
      RECT  10297.5 164907.5 10362.5 164772.5 ;
      RECT  10297.5 164907.5 10362.5 164772.5 ;
      RECT  10107.5 164907.5 10172.5 164772.5 ;
      RECT  10297.5 164907.5 10362.5 164772.5 ;
      RECT  10487.5 164907.5 10552.5 164772.5 ;
      RECT  10487.5 164907.5 10552.5 164772.5 ;
      RECT  10297.5 164907.5 10362.5 164772.5 ;
      RECT  10107.5 165747.5 10172.5 165612.5 ;
      RECT  10297.5 165747.5 10362.5 165612.5 ;
      RECT  10297.5 165747.5 10362.5 165612.5 ;
      RECT  10107.5 165747.5 10172.5 165612.5 ;
      RECT  10297.5 165747.5 10362.5 165612.5 ;
      RECT  10487.5 165747.5 10552.5 165612.5 ;
      RECT  10487.5 165747.5 10552.5 165612.5 ;
      RECT  10297.5 165747.5 10362.5 165612.5 ;
      RECT  10657.5 164817.5 10722.5 164682.5 ;
      RECT  10657.5 165792.5 10722.5 165657.5 ;
      RECT  10492.5 165517.5 10357.5 165452.5 ;
      RECT  10235.0 165302.5 10100.0 165237.5 ;
      RECT  10297.5 164907.5 10362.5 164772.5 ;
      RECT  10487.5 165747.5 10552.5 165612.5 ;
      RECT  10587.5 165302.5 10452.5 165237.5 ;
      RECT  10100.0 165302.5 10235.0 165237.5 ;
      RECT  10357.5 165517.5 10492.5 165452.5 ;
      RECT  10452.5 165302.5 10587.5 165237.5 ;
      RECT  10040.0 164597.5 10960.0 164532.5 ;
      RECT  10040.0 165942.5 10960.0 165877.5 ;
      RECT  11387.5 164750.0 11452.5 164565.0 ;
      RECT  11387.5 165910.0 11452.5 165725.0 ;
      RECT  11027.5 165792.5 11092.5 165942.5 ;
      RECT  11027.5 164907.5 11092.5 164532.5 ;
      RECT  11217.5 165792.5 11282.5 164907.5 ;
      RECT  11027.5 164907.5 11092.5 164772.5 ;
      RECT  11217.5 164907.5 11282.5 164772.5 ;
      RECT  11217.5 164907.5 11282.5 164772.5 ;
      RECT  11027.5 164907.5 11092.5 164772.5 ;
      RECT  11027.5 165792.5 11092.5 165657.5 ;
      RECT  11217.5 165792.5 11282.5 165657.5 ;
      RECT  11217.5 165792.5 11282.5 165657.5 ;
      RECT  11027.5 165792.5 11092.5 165657.5 ;
      RECT  11387.5 164817.5 11452.5 164682.5 ;
      RECT  11387.5 165792.5 11452.5 165657.5 ;
      RECT  11085.0 165350.0 11150.0 165215.0 ;
      RECT  11085.0 165350.0 11150.0 165215.0 ;
      RECT  11250.0 165315.0 11315.0 165250.0 ;
      RECT  10960.0 164597.5 11520.0 164532.5 ;
      RECT  10960.0 165942.5 11520.0 165877.5 ;
      RECT  9222.5 165215.0 9287.5 165350.0 ;
      RECT  9362.5 165487.5 9427.5 165622.5 ;
      RECT  10357.5 165452.5 10222.5 165517.5 ;
      RECT  9907.5 167070.0 9972.5 167255.0 ;
      RECT  9907.5 165910.0 9972.5 166095.0 ;
      RECT  9547.5 166027.5 9612.5 165877.5 ;
      RECT  9547.5 166912.5 9612.5 167287.5 ;
      RECT  9737.5 166027.5 9802.5 166912.5 ;
      RECT  9547.5 166912.5 9612.5 167047.5 ;
      RECT  9737.5 166912.5 9802.5 167047.5 ;
      RECT  9737.5 166912.5 9802.5 167047.5 ;
      RECT  9547.5 166912.5 9612.5 167047.5 ;
      RECT  9547.5 166027.5 9612.5 166162.5 ;
      RECT  9737.5 166027.5 9802.5 166162.5 ;
      RECT  9737.5 166027.5 9802.5 166162.5 ;
      RECT  9547.5 166027.5 9612.5 166162.5 ;
      RECT  9907.5 167002.5 9972.5 167137.5 ;
      RECT  9907.5 166027.5 9972.5 166162.5 ;
      RECT  9605.0 166470.0 9670.0 166605.0 ;
      RECT  9605.0 166470.0 9670.0 166605.0 ;
      RECT  9770.0 166505.0 9835.0 166570.0 ;
      RECT  9480.0 167222.5 10040.0 167287.5 ;
      RECT  9480.0 165877.5 10040.0 165942.5 ;
      RECT  10107.5 166072.5 10172.5 165877.5 ;
      RECT  10107.5 166912.5 10172.5 167287.5 ;
      RECT  10487.5 166912.5 10552.5 167287.5 ;
      RECT  10657.5 167070.0 10722.5 167255.0 ;
      RECT  10657.5 165910.0 10722.5 166095.0 ;
      RECT  10107.5 166912.5 10172.5 167047.5 ;
      RECT  10297.5 166912.5 10362.5 167047.5 ;
      RECT  10297.5 166912.5 10362.5 167047.5 ;
      RECT  10107.5 166912.5 10172.5 167047.5 ;
      RECT  10297.5 166912.5 10362.5 167047.5 ;
      RECT  10487.5 166912.5 10552.5 167047.5 ;
      RECT  10487.5 166912.5 10552.5 167047.5 ;
      RECT  10297.5 166912.5 10362.5 167047.5 ;
      RECT  10107.5 166072.5 10172.5 166207.5 ;
      RECT  10297.5 166072.5 10362.5 166207.5 ;
      RECT  10297.5 166072.5 10362.5 166207.5 ;
      RECT  10107.5 166072.5 10172.5 166207.5 ;
      RECT  10297.5 166072.5 10362.5 166207.5 ;
      RECT  10487.5 166072.5 10552.5 166207.5 ;
      RECT  10487.5 166072.5 10552.5 166207.5 ;
      RECT  10297.5 166072.5 10362.5 166207.5 ;
      RECT  10657.5 167002.5 10722.5 167137.5 ;
      RECT  10657.5 166027.5 10722.5 166162.5 ;
      RECT  10492.5 166302.5 10357.5 166367.5 ;
      RECT  10235.0 166517.5 10100.0 166582.5 ;
      RECT  10297.5 166912.5 10362.5 167047.5 ;
      RECT  10487.5 166072.5 10552.5 166207.5 ;
      RECT  10587.5 166517.5 10452.5 166582.5 ;
      RECT  10100.0 166517.5 10235.0 166582.5 ;
      RECT  10357.5 166302.5 10492.5 166367.5 ;
      RECT  10452.5 166517.5 10587.5 166582.5 ;
      RECT  10040.0 167222.5 10960.0 167287.5 ;
      RECT  10040.0 165877.5 10960.0 165942.5 ;
      RECT  11387.5 167070.0 11452.5 167255.0 ;
      RECT  11387.5 165910.0 11452.5 166095.0 ;
      RECT  11027.5 166027.5 11092.5 165877.5 ;
      RECT  11027.5 166912.5 11092.5 167287.5 ;
      RECT  11217.5 166027.5 11282.5 166912.5 ;
      RECT  11027.5 166912.5 11092.5 167047.5 ;
      RECT  11217.5 166912.5 11282.5 167047.5 ;
      RECT  11217.5 166912.5 11282.5 167047.5 ;
      RECT  11027.5 166912.5 11092.5 167047.5 ;
      RECT  11027.5 166027.5 11092.5 166162.5 ;
      RECT  11217.5 166027.5 11282.5 166162.5 ;
      RECT  11217.5 166027.5 11282.5 166162.5 ;
      RECT  11027.5 166027.5 11092.5 166162.5 ;
      RECT  11387.5 167002.5 11452.5 167137.5 ;
      RECT  11387.5 166027.5 11452.5 166162.5 ;
      RECT  11085.0 166470.0 11150.0 166605.0 ;
      RECT  11085.0 166470.0 11150.0 166605.0 ;
      RECT  11250.0 166505.0 11315.0 166570.0 ;
      RECT  10960.0 167222.5 11520.0 167287.5 ;
      RECT  10960.0 165877.5 11520.0 165942.5 ;
      RECT  9222.5 166470.0 9287.5 166605.0 ;
      RECT  9362.5 166197.5 9427.5 166332.5 ;
      RECT  10357.5 166302.5 10222.5 166367.5 ;
      RECT  9907.5 167440.0 9972.5 167255.0 ;
      RECT  9907.5 168600.0 9972.5 168415.0 ;
      RECT  9547.5 168482.5 9612.5 168632.5 ;
      RECT  9547.5 167597.5 9612.5 167222.5 ;
      RECT  9737.5 168482.5 9802.5 167597.5 ;
      RECT  9547.5 167597.5 9612.5 167462.5 ;
      RECT  9737.5 167597.5 9802.5 167462.5 ;
      RECT  9737.5 167597.5 9802.5 167462.5 ;
      RECT  9547.5 167597.5 9612.5 167462.5 ;
      RECT  9547.5 168482.5 9612.5 168347.5 ;
      RECT  9737.5 168482.5 9802.5 168347.5 ;
      RECT  9737.5 168482.5 9802.5 168347.5 ;
      RECT  9547.5 168482.5 9612.5 168347.5 ;
      RECT  9907.5 167507.5 9972.5 167372.5 ;
      RECT  9907.5 168482.5 9972.5 168347.5 ;
      RECT  9605.0 168040.0 9670.0 167905.0 ;
      RECT  9605.0 168040.0 9670.0 167905.0 ;
      RECT  9770.0 168005.0 9835.0 167940.0 ;
      RECT  9480.0 167287.5 10040.0 167222.5 ;
      RECT  9480.0 168632.5 10040.0 168567.5 ;
      RECT  10107.5 168437.5 10172.5 168632.5 ;
      RECT  10107.5 167597.5 10172.5 167222.5 ;
      RECT  10487.5 167597.5 10552.5 167222.5 ;
      RECT  10657.5 167440.0 10722.5 167255.0 ;
      RECT  10657.5 168600.0 10722.5 168415.0 ;
      RECT  10107.5 167597.5 10172.5 167462.5 ;
      RECT  10297.5 167597.5 10362.5 167462.5 ;
      RECT  10297.5 167597.5 10362.5 167462.5 ;
      RECT  10107.5 167597.5 10172.5 167462.5 ;
      RECT  10297.5 167597.5 10362.5 167462.5 ;
      RECT  10487.5 167597.5 10552.5 167462.5 ;
      RECT  10487.5 167597.5 10552.5 167462.5 ;
      RECT  10297.5 167597.5 10362.5 167462.5 ;
      RECT  10107.5 168437.5 10172.5 168302.5 ;
      RECT  10297.5 168437.5 10362.5 168302.5 ;
      RECT  10297.5 168437.5 10362.5 168302.5 ;
      RECT  10107.5 168437.5 10172.5 168302.5 ;
      RECT  10297.5 168437.5 10362.5 168302.5 ;
      RECT  10487.5 168437.5 10552.5 168302.5 ;
      RECT  10487.5 168437.5 10552.5 168302.5 ;
      RECT  10297.5 168437.5 10362.5 168302.5 ;
      RECT  10657.5 167507.5 10722.5 167372.5 ;
      RECT  10657.5 168482.5 10722.5 168347.5 ;
      RECT  10492.5 168207.5 10357.5 168142.5 ;
      RECT  10235.0 167992.5 10100.0 167927.5 ;
      RECT  10297.5 167597.5 10362.5 167462.5 ;
      RECT  10487.5 168437.5 10552.5 168302.5 ;
      RECT  10587.5 167992.5 10452.5 167927.5 ;
      RECT  10100.0 167992.5 10235.0 167927.5 ;
      RECT  10357.5 168207.5 10492.5 168142.5 ;
      RECT  10452.5 167992.5 10587.5 167927.5 ;
      RECT  10040.0 167287.5 10960.0 167222.5 ;
      RECT  10040.0 168632.5 10960.0 168567.5 ;
      RECT  11387.5 167440.0 11452.5 167255.0 ;
      RECT  11387.5 168600.0 11452.5 168415.0 ;
      RECT  11027.5 168482.5 11092.5 168632.5 ;
      RECT  11027.5 167597.5 11092.5 167222.5 ;
      RECT  11217.5 168482.5 11282.5 167597.5 ;
      RECT  11027.5 167597.5 11092.5 167462.5 ;
      RECT  11217.5 167597.5 11282.5 167462.5 ;
      RECT  11217.5 167597.5 11282.5 167462.5 ;
      RECT  11027.5 167597.5 11092.5 167462.5 ;
      RECT  11027.5 168482.5 11092.5 168347.5 ;
      RECT  11217.5 168482.5 11282.5 168347.5 ;
      RECT  11217.5 168482.5 11282.5 168347.5 ;
      RECT  11027.5 168482.5 11092.5 168347.5 ;
      RECT  11387.5 167507.5 11452.5 167372.5 ;
      RECT  11387.5 168482.5 11452.5 168347.5 ;
      RECT  11085.0 168040.0 11150.0 167905.0 ;
      RECT  11085.0 168040.0 11150.0 167905.0 ;
      RECT  11250.0 168005.0 11315.0 167940.0 ;
      RECT  10960.0 167287.5 11520.0 167222.5 ;
      RECT  10960.0 168632.5 11520.0 168567.5 ;
      RECT  9222.5 167905.0 9287.5 168040.0 ;
      RECT  9362.5 168177.5 9427.5 168312.5 ;
      RECT  10357.5 168142.5 10222.5 168207.5 ;
      RECT  9907.5 169760.0 9972.5 169945.0 ;
      RECT  9907.5 168600.0 9972.5 168785.0 ;
      RECT  9547.5 168717.5 9612.5 168567.5 ;
      RECT  9547.5 169602.5 9612.5 169977.5 ;
      RECT  9737.5 168717.5 9802.5 169602.5 ;
      RECT  9547.5 169602.5 9612.5 169737.5 ;
      RECT  9737.5 169602.5 9802.5 169737.5 ;
      RECT  9737.5 169602.5 9802.5 169737.5 ;
      RECT  9547.5 169602.5 9612.5 169737.5 ;
      RECT  9547.5 168717.5 9612.5 168852.5 ;
      RECT  9737.5 168717.5 9802.5 168852.5 ;
      RECT  9737.5 168717.5 9802.5 168852.5 ;
      RECT  9547.5 168717.5 9612.5 168852.5 ;
      RECT  9907.5 169692.5 9972.5 169827.5 ;
      RECT  9907.5 168717.5 9972.5 168852.5 ;
      RECT  9605.0 169160.0 9670.0 169295.0 ;
      RECT  9605.0 169160.0 9670.0 169295.0 ;
      RECT  9770.0 169195.0 9835.0 169260.0 ;
      RECT  9480.0 169912.5 10040.0 169977.5 ;
      RECT  9480.0 168567.5 10040.0 168632.5 ;
      RECT  10107.5 168762.5 10172.5 168567.5 ;
      RECT  10107.5 169602.5 10172.5 169977.5 ;
      RECT  10487.5 169602.5 10552.5 169977.5 ;
      RECT  10657.5 169760.0 10722.5 169945.0 ;
      RECT  10657.5 168600.0 10722.5 168785.0 ;
      RECT  10107.5 169602.5 10172.5 169737.5 ;
      RECT  10297.5 169602.5 10362.5 169737.5 ;
      RECT  10297.5 169602.5 10362.5 169737.5 ;
      RECT  10107.5 169602.5 10172.5 169737.5 ;
      RECT  10297.5 169602.5 10362.5 169737.5 ;
      RECT  10487.5 169602.5 10552.5 169737.5 ;
      RECT  10487.5 169602.5 10552.5 169737.5 ;
      RECT  10297.5 169602.5 10362.5 169737.5 ;
      RECT  10107.5 168762.5 10172.5 168897.5 ;
      RECT  10297.5 168762.5 10362.5 168897.5 ;
      RECT  10297.5 168762.5 10362.5 168897.5 ;
      RECT  10107.5 168762.5 10172.5 168897.5 ;
      RECT  10297.5 168762.5 10362.5 168897.5 ;
      RECT  10487.5 168762.5 10552.5 168897.5 ;
      RECT  10487.5 168762.5 10552.5 168897.5 ;
      RECT  10297.5 168762.5 10362.5 168897.5 ;
      RECT  10657.5 169692.5 10722.5 169827.5 ;
      RECT  10657.5 168717.5 10722.5 168852.5 ;
      RECT  10492.5 168992.5 10357.5 169057.5 ;
      RECT  10235.0 169207.5 10100.0 169272.5 ;
      RECT  10297.5 169602.5 10362.5 169737.5 ;
      RECT  10487.5 168762.5 10552.5 168897.5 ;
      RECT  10587.5 169207.5 10452.5 169272.5 ;
      RECT  10100.0 169207.5 10235.0 169272.5 ;
      RECT  10357.5 168992.5 10492.5 169057.5 ;
      RECT  10452.5 169207.5 10587.5 169272.5 ;
      RECT  10040.0 169912.5 10960.0 169977.5 ;
      RECT  10040.0 168567.5 10960.0 168632.5 ;
      RECT  11387.5 169760.0 11452.5 169945.0 ;
      RECT  11387.5 168600.0 11452.5 168785.0 ;
      RECT  11027.5 168717.5 11092.5 168567.5 ;
      RECT  11027.5 169602.5 11092.5 169977.5 ;
      RECT  11217.5 168717.5 11282.5 169602.5 ;
      RECT  11027.5 169602.5 11092.5 169737.5 ;
      RECT  11217.5 169602.5 11282.5 169737.5 ;
      RECT  11217.5 169602.5 11282.5 169737.5 ;
      RECT  11027.5 169602.5 11092.5 169737.5 ;
      RECT  11027.5 168717.5 11092.5 168852.5 ;
      RECT  11217.5 168717.5 11282.5 168852.5 ;
      RECT  11217.5 168717.5 11282.5 168852.5 ;
      RECT  11027.5 168717.5 11092.5 168852.5 ;
      RECT  11387.5 169692.5 11452.5 169827.5 ;
      RECT  11387.5 168717.5 11452.5 168852.5 ;
      RECT  11085.0 169160.0 11150.0 169295.0 ;
      RECT  11085.0 169160.0 11150.0 169295.0 ;
      RECT  11250.0 169195.0 11315.0 169260.0 ;
      RECT  10960.0 169912.5 11520.0 169977.5 ;
      RECT  10960.0 168567.5 11520.0 168632.5 ;
      RECT  9222.5 169160.0 9287.5 169295.0 ;
      RECT  9362.5 168887.5 9427.5 169022.5 ;
      RECT  10357.5 168992.5 10222.5 169057.5 ;
      RECT  9907.5 170130.0 9972.5 169945.0 ;
      RECT  9907.5 171290.0 9972.5 171105.0 ;
      RECT  9547.5 171172.5 9612.5 171322.5 ;
      RECT  9547.5 170287.5 9612.5 169912.5 ;
      RECT  9737.5 171172.5 9802.5 170287.5 ;
      RECT  9547.5 170287.5 9612.5 170152.5 ;
      RECT  9737.5 170287.5 9802.5 170152.5 ;
      RECT  9737.5 170287.5 9802.5 170152.5 ;
      RECT  9547.5 170287.5 9612.5 170152.5 ;
      RECT  9547.5 171172.5 9612.5 171037.5 ;
      RECT  9737.5 171172.5 9802.5 171037.5 ;
      RECT  9737.5 171172.5 9802.5 171037.5 ;
      RECT  9547.5 171172.5 9612.5 171037.5 ;
      RECT  9907.5 170197.5 9972.5 170062.5 ;
      RECT  9907.5 171172.5 9972.5 171037.5 ;
      RECT  9605.0 170730.0 9670.0 170595.0 ;
      RECT  9605.0 170730.0 9670.0 170595.0 ;
      RECT  9770.0 170695.0 9835.0 170630.0 ;
      RECT  9480.0 169977.5 10040.0 169912.5 ;
      RECT  9480.0 171322.5 10040.0 171257.5 ;
      RECT  10107.5 171127.5 10172.5 171322.5 ;
      RECT  10107.5 170287.5 10172.5 169912.5 ;
      RECT  10487.5 170287.5 10552.5 169912.5 ;
      RECT  10657.5 170130.0 10722.5 169945.0 ;
      RECT  10657.5 171290.0 10722.5 171105.0 ;
      RECT  10107.5 170287.5 10172.5 170152.5 ;
      RECT  10297.5 170287.5 10362.5 170152.5 ;
      RECT  10297.5 170287.5 10362.5 170152.5 ;
      RECT  10107.5 170287.5 10172.5 170152.5 ;
      RECT  10297.5 170287.5 10362.5 170152.5 ;
      RECT  10487.5 170287.5 10552.5 170152.5 ;
      RECT  10487.5 170287.5 10552.5 170152.5 ;
      RECT  10297.5 170287.5 10362.5 170152.5 ;
      RECT  10107.5 171127.5 10172.5 170992.5 ;
      RECT  10297.5 171127.5 10362.5 170992.5 ;
      RECT  10297.5 171127.5 10362.5 170992.5 ;
      RECT  10107.5 171127.5 10172.5 170992.5 ;
      RECT  10297.5 171127.5 10362.5 170992.5 ;
      RECT  10487.5 171127.5 10552.5 170992.5 ;
      RECT  10487.5 171127.5 10552.5 170992.5 ;
      RECT  10297.5 171127.5 10362.5 170992.5 ;
      RECT  10657.5 170197.5 10722.5 170062.5 ;
      RECT  10657.5 171172.5 10722.5 171037.5 ;
      RECT  10492.5 170897.5 10357.5 170832.5 ;
      RECT  10235.0 170682.5 10100.0 170617.5 ;
      RECT  10297.5 170287.5 10362.5 170152.5 ;
      RECT  10487.5 171127.5 10552.5 170992.5 ;
      RECT  10587.5 170682.5 10452.5 170617.5 ;
      RECT  10100.0 170682.5 10235.0 170617.5 ;
      RECT  10357.5 170897.5 10492.5 170832.5 ;
      RECT  10452.5 170682.5 10587.5 170617.5 ;
      RECT  10040.0 169977.5 10960.0 169912.5 ;
      RECT  10040.0 171322.5 10960.0 171257.5 ;
      RECT  11387.5 170130.0 11452.5 169945.0 ;
      RECT  11387.5 171290.0 11452.5 171105.0 ;
      RECT  11027.5 171172.5 11092.5 171322.5 ;
      RECT  11027.5 170287.5 11092.5 169912.5 ;
      RECT  11217.5 171172.5 11282.5 170287.5 ;
      RECT  11027.5 170287.5 11092.5 170152.5 ;
      RECT  11217.5 170287.5 11282.5 170152.5 ;
      RECT  11217.5 170287.5 11282.5 170152.5 ;
      RECT  11027.5 170287.5 11092.5 170152.5 ;
      RECT  11027.5 171172.5 11092.5 171037.5 ;
      RECT  11217.5 171172.5 11282.5 171037.5 ;
      RECT  11217.5 171172.5 11282.5 171037.5 ;
      RECT  11027.5 171172.5 11092.5 171037.5 ;
      RECT  11387.5 170197.5 11452.5 170062.5 ;
      RECT  11387.5 171172.5 11452.5 171037.5 ;
      RECT  11085.0 170730.0 11150.0 170595.0 ;
      RECT  11085.0 170730.0 11150.0 170595.0 ;
      RECT  11250.0 170695.0 11315.0 170630.0 ;
      RECT  10960.0 169977.5 11520.0 169912.5 ;
      RECT  10960.0 171322.5 11520.0 171257.5 ;
      RECT  9222.5 170595.0 9287.5 170730.0 ;
      RECT  9362.5 170867.5 9427.5 171002.5 ;
      RECT  10357.5 170832.5 10222.5 170897.5 ;
      RECT  9907.5 172450.0 9972.5 172635.0 ;
      RECT  9907.5 171290.0 9972.5 171475.0 ;
      RECT  9547.5 171407.5 9612.5 171257.5 ;
      RECT  9547.5 172292.5 9612.5 172667.5 ;
      RECT  9737.5 171407.5 9802.5 172292.5 ;
      RECT  9547.5 172292.5 9612.5 172427.5 ;
      RECT  9737.5 172292.5 9802.5 172427.5 ;
      RECT  9737.5 172292.5 9802.5 172427.5 ;
      RECT  9547.5 172292.5 9612.5 172427.5 ;
      RECT  9547.5 171407.5 9612.5 171542.5 ;
      RECT  9737.5 171407.5 9802.5 171542.5 ;
      RECT  9737.5 171407.5 9802.5 171542.5 ;
      RECT  9547.5 171407.5 9612.5 171542.5 ;
      RECT  9907.5 172382.5 9972.5 172517.5 ;
      RECT  9907.5 171407.5 9972.5 171542.5 ;
      RECT  9605.0 171850.0 9670.0 171985.0 ;
      RECT  9605.0 171850.0 9670.0 171985.0 ;
      RECT  9770.0 171885.0 9835.0 171950.0 ;
      RECT  9480.0 172602.5 10040.0 172667.5 ;
      RECT  9480.0 171257.5 10040.0 171322.5 ;
      RECT  10107.5 171452.5 10172.5 171257.5 ;
      RECT  10107.5 172292.5 10172.5 172667.5 ;
      RECT  10487.5 172292.5 10552.5 172667.5 ;
      RECT  10657.5 172450.0 10722.5 172635.0 ;
      RECT  10657.5 171290.0 10722.5 171475.0 ;
      RECT  10107.5 172292.5 10172.5 172427.5 ;
      RECT  10297.5 172292.5 10362.5 172427.5 ;
      RECT  10297.5 172292.5 10362.5 172427.5 ;
      RECT  10107.5 172292.5 10172.5 172427.5 ;
      RECT  10297.5 172292.5 10362.5 172427.5 ;
      RECT  10487.5 172292.5 10552.5 172427.5 ;
      RECT  10487.5 172292.5 10552.5 172427.5 ;
      RECT  10297.5 172292.5 10362.5 172427.5 ;
      RECT  10107.5 171452.5 10172.5 171587.5 ;
      RECT  10297.5 171452.5 10362.5 171587.5 ;
      RECT  10297.5 171452.5 10362.5 171587.5 ;
      RECT  10107.5 171452.5 10172.5 171587.5 ;
      RECT  10297.5 171452.5 10362.5 171587.5 ;
      RECT  10487.5 171452.5 10552.5 171587.5 ;
      RECT  10487.5 171452.5 10552.5 171587.5 ;
      RECT  10297.5 171452.5 10362.5 171587.5 ;
      RECT  10657.5 172382.5 10722.5 172517.5 ;
      RECT  10657.5 171407.5 10722.5 171542.5 ;
      RECT  10492.5 171682.5 10357.5 171747.5 ;
      RECT  10235.0 171897.5 10100.0 171962.5 ;
      RECT  10297.5 172292.5 10362.5 172427.5 ;
      RECT  10487.5 171452.5 10552.5 171587.5 ;
      RECT  10587.5 171897.5 10452.5 171962.5 ;
      RECT  10100.0 171897.5 10235.0 171962.5 ;
      RECT  10357.5 171682.5 10492.5 171747.5 ;
      RECT  10452.5 171897.5 10587.5 171962.5 ;
      RECT  10040.0 172602.5 10960.0 172667.5 ;
      RECT  10040.0 171257.5 10960.0 171322.5 ;
      RECT  11387.5 172450.0 11452.5 172635.0 ;
      RECT  11387.5 171290.0 11452.5 171475.0 ;
      RECT  11027.5 171407.5 11092.5 171257.5 ;
      RECT  11027.5 172292.5 11092.5 172667.5 ;
      RECT  11217.5 171407.5 11282.5 172292.5 ;
      RECT  11027.5 172292.5 11092.5 172427.5 ;
      RECT  11217.5 172292.5 11282.5 172427.5 ;
      RECT  11217.5 172292.5 11282.5 172427.5 ;
      RECT  11027.5 172292.5 11092.5 172427.5 ;
      RECT  11027.5 171407.5 11092.5 171542.5 ;
      RECT  11217.5 171407.5 11282.5 171542.5 ;
      RECT  11217.5 171407.5 11282.5 171542.5 ;
      RECT  11027.5 171407.5 11092.5 171542.5 ;
      RECT  11387.5 172382.5 11452.5 172517.5 ;
      RECT  11387.5 171407.5 11452.5 171542.5 ;
      RECT  11085.0 171850.0 11150.0 171985.0 ;
      RECT  11085.0 171850.0 11150.0 171985.0 ;
      RECT  11250.0 171885.0 11315.0 171950.0 ;
      RECT  10960.0 172602.5 11520.0 172667.5 ;
      RECT  10960.0 171257.5 11520.0 171322.5 ;
      RECT  9222.5 171850.0 9287.5 171985.0 ;
      RECT  9362.5 171577.5 9427.5 171712.5 ;
      RECT  10357.5 171682.5 10222.5 171747.5 ;
      RECT  9907.5 172820.0 9972.5 172635.0 ;
      RECT  9907.5 173980.0 9972.5 173795.0 ;
      RECT  9547.5 173862.5 9612.5 174012.5 ;
      RECT  9547.5 172977.5 9612.5 172602.5 ;
      RECT  9737.5 173862.5 9802.5 172977.5 ;
      RECT  9547.5 172977.5 9612.5 172842.5 ;
      RECT  9737.5 172977.5 9802.5 172842.5 ;
      RECT  9737.5 172977.5 9802.5 172842.5 ;
      RECT  9547.5 172977.5 9612.5 172842.5 ;
      RECT  9547.5 173862.5 9612.5 173727.5 ;
      RECT  9737.5 173862.5 9802.5 173727.5 ;
      RECT  9737.5 173862.5 9802.5 173727.5 ;
      RECT  9547.5 173862.5 9612.5 173727.5 ;
      RECT  9907.5 172887.5 9972.5 172752.5 ;
      RECT  9907.5 173862.5 9972.5 173727.5 ;
      RECT  9605.0 173420.0 9670.0 173285.0 ;
      RECT  9605.0 173420.0 9670.0 173285.0 ;
      RECT  9770.0 173385.0 9835.0 173320.0 ;
      RECT  9480.0 172667.5 10040.0 172602.5 ;
      RECT  9480.0 174012.5 10040.0 173947.5 ;
      RECT  10107.5 173817.5 10172.5 174012.5 ;
      RECT  10107.5 172977.5 10172.5 172602.5 ;
      RECT  10487.5 172977.5 10552.5 172602.5 ;
      RECT  10657.5 172820.0 10722.5 172635.0 ;
      RECT  10657.5 173980.0 10722.5 173795.0 ;
      RECT  10107.5 172977.5 10172.5 172842.5 ;
      RECT  10297.5 172977.5 10362.5 172842.5 ;
      RECT  10297.5 172977.5 10362.5 172842.5 ;
      RECT  10107.5 172977.5 10172.5 172842.5 ;
      RECT  10297.5 172977.5 10362.5 172842.5 ;
      RECT  10487.5 172977.5 10552.5 172842.5 ;
      RECT  10487.5 172977.5 10552.5 172842.5 ;
      RECT  10297.5 172977.5 10362.5 172842.5 ;
      RECT  10107.5 173817.5 10172.5 173682.5 ;
      RECT  10297.5 173817.5 10362.5 173682.5 ;
      RECT  10297.5 173817.5 10362.5 173682.5 ;
      RECT  10107.5 173817.5 10172.5 173682.5 ;
      RECT  10297.5 173817.5 10362.5 173682.5 ;
      RECT  10487.5 173817.5 10552.5 173682.5 ;
      RECT  10487.5 173817.5 10552.5 173682.5 ;
      RECT  10297.5 173817.5 10362.5 173682.5 ;
      RECT  10657.5 172887.5 10722.5 172752.5 ;
      RECT  10657.5 173862.5 10722.5 173727.5 ;
      RECT  10492.5 173587.5 10357.5 173522.5 ;
      RECT  10235.0 173372.5 10100.0 173307.5 ;
      RECT  10297.5 172977.5 10362.5 172842.5 ;
      RECT  10487.5 173817.5 10552.5 173682.5 ;
      RECT  10587.5 173372.5 10452.5 173307.5 ;
      RECT  10100.0 173372.5 10235.0 173307.5 ;
      RECT  10357.5 173587.5 10492.5 173522.5 ;
      RECT  10452.5 173372.5 10587.5 173307.5 ;
      RECT  10040.0 172667.5 10960.0 172602.5 ;
      RECT  10040.0 174012.5 10960.0 173947.5 ;
      RECT  11387.5 172820.0 11452.5 172635.0 ;
      RECT  11387.5 173980.0 11452.5 173795.0 ;
      RECT  11027.5 173862.5 11092.5 174012.5 ;
      RECT  11027.5 172977.5 11092.5 172602.5 ;
      RECT  11217.5 173862.5 11282.5 172977.5 ;
      RECT  11027.5 172977.5 11092.5 172842.5 ;
      RECT  11217.5 172977.5 11282.5 172842.5 ;
      RECT  11217.5 172977.5 11282.5 172842.5 ;
      RECT  11027.5 172977.5 11092.5 172842.5 ;
      RECT  11027.5 173862.5 11092.5 173727.5 ;
      RECT  11217.5 173862.5 11282.5 173727.5 ;
      RECT  11217.5 173862.5 11282.5 173727.5 ;
      RECT  11027.5 173862.5 11092.5 173727.5 ;
      RECT  11387.5 172887.5 11452.5 172752.5 ;
      RECT  11387.5 173862.5 11452.5 173727.5 ;
      RECT  11085.0 173420.0 11150.0 173285.0 ;
      RECT  11085.0 173420.0 11150.0 173285.0 ;
      RECT  11250.0 173385.0 11315.0 173320.0 ;
      RECT  10960.0 172667.5 11520.0 172602.5 ;
      RECT  10960.0 174012.5 11520.0 173947.5 ;
      RECT  9222.5 173285.0 9287.5 173420.0 ;
      RECT  9362.5 173557.5 9427.5 173692.5 ;
      RECT  10357.5 173522.5 10222.5 173587.5 ;
      RECT  9907.5 175140.0 9972.5 175325.0 ;
      RECT  9907.5 173980.0 9972.5 174165.0 ;
      RECT  9547.5 174097.5 9612.5 173947.5 ;
      RECT  9547.5 174982.5 9612.5 175357.5 ;
      RECT  9737.5 174097.5 9802.5 174982.5 ;
      RECT  9547.5 174982.5 9612.5 175117.5 ;
      RECT  9737.5 174982.5 9802.5 175117.5 ;
      RECT  9737.5 174982.5 9802.5 175117.5 ;
      RECT  9547.5 174982.5 9612.5 175117.5 ;
      RECT  9547.5 174097.5 9612.5 174232.5 ;
      RECT  9737.5 174097.5 9802.5 174232.5 ;
      RECT  9737.5 174097.5 9802.5 174232.5 ;
      RECT  9547.5 174097.5 9612.5 174232.5 ;
      RECT  9907.5 175072.5 9972.5 175207.5 ;
      RECT  9907.5 174097.5 9972.5 174232.5 ;
      RECT  9605.0 174540.0 9670.0 174675.0 ;
      RECT  9605.0 174540.0 9670.0 174675.0 ;
      RECT  9770.0 174575.0 9835.0 174640.0 ;
      RECT  9480.0 175292.5 10040.0 175357.5 ;
      RECT  9480.0 173947.5 10040.0 174012.5 ;
      RECT  10107.5 174142.5 10172.5 173947.5 ;
      RECT  10107.5 174982.5 10172.5 175357.5 ;
      RECT  10487.5 174982.5 10552.5 175357.5 ;
      RECT  10657.5 175140.0 10722.5 175325.0 ;
      RECT  10657.5 173980.0 10722.5 174165.0 ;
      RECT  10107.5 174982.5 10172.5 175117.5 ;
      RECT  10297.5 174982.5 10362.5 175117.5 ;
      RECT  10297.5 174982.5 10362.5 175117.5 ;
      RECT  10107.5 174982.5 10172.5 175117.5 ;
      RECT  10297.5 174982.5 10362.5 175117.5 ;
      RECT  10487.5 174982.5 10552.5 175117.5 ;
      RECT  10487.5 174982.5 10552.5 175117.5 ;
      RECT  10297.5 174982.5 10362.5 175117.5 ;
      RECT  10107.5 174142.5 10172.5 174277.5 ;
      RECT  10297.5 174142.5 10362.5 174277.5 ;
      RECT  10297.5 174142.5 10362.5 174277.5 ;
      RECT  10107.5 174142.5 10172.5 174277.5 ;
      RECT  10297.5 174142.5 10362.5 174277.5 ;
      RECT  10487.5 174142.5 10552.5 174277.5 ;
      RECT  10487.5 174142.5 10552.5 174277.5 ;
      RECT  10297.5 174142.5 10362.5 174277.5 ;
      RECT  10657.5 175072.5 10722.5 175207.5 ;
      RECT  10657.5 174097.5 10722.5 174232.5 ;
      RECT  10492.5 174372.5 10357.5 174437.5 ;
      RECT  10235.0 174587.5 10100.0 174652.5 ;
      RECT  10297.5 174982.5 10362.5 175117.5 ;
      RECT  10487.5 174142.5 10552.5 174277.5 ;
      RECT  10587.5 174587.5 10452.5 174652.5 ;
      RECT  10100.0 174587.5 10235.0 174652.5 ;
      RECT  10357.5 174372.5 10492.5 174437.5 ;
      RECT  10452.5 174587.5 10587.5 174652.5 ;
      RECT  10040.0 175292.5 10960.0 175357.5 ;
      RECT  10040.0 173947.5 10960.0 174012.5 ;
      RECT  11387.5 175140.0 11452.5 175325.0 ;
      RECT  11387.5 173980.0 11452.5 174165.0 ;
      RECT  11027.5 174097.5 11092.5 173947.5 ;
      RECT  11027.5 174982.5 11092.5 175357.5 ;
      RECT  11217.5 174097.5 11282.5 174982.5 ;
      RECT  11027.5 174982.5 11092.5 175117.5 ;
      RECT  11217.5 174982.5 11282.5 175117.5 ;
      RECT  11217.5 174982.5 11282.5 175117.5 ;
      RECT  11027.5 174982.5 11092.5 175117.5 ;
      RECT  11027.5 174097.5 11092.5 174232.5 ;
      RECT  11217.5 174097.5 11282.5 174232.5 ;
      RECT  11217.5 174097.5 11282.5 174232.5 ;
      RECT  11027.5 174097.5 11092.5 174232.5 ;
      RECT  11387.5 175072.5 11452.5 175207.5 ;
      RECT  11387.5 174097.5 11452.5 174232.5 ;
      RECT  11085.0 174540.0 11150.0 174675.0 ;
      RECT  11085.0 174540.0 11150.0 174675.0 ;
      RECT  11250.0 174575.0 11315.0 174640.0 ;
      RECT  10960.0 175292.5 11520.0 175357.5 ;
      RECT  10960.0 173947.5 11520.0 174012.5 ;
      RECT  9222.5 174540.0 9287.5 174675.0 ;
      RECT  9362.5 174267.5 9427.5 174402.5 ;
      RECT  10357.5 174372.5 10222.5 174437.5 ;
      RECT  9907.5 175510.0 9972.5 175325.0 ;
      RECT  9907.5 176670.0 9972.5 176485.0 ;
      RECT  9547.5 176552.5 9612.5 176702.5 ;
      RECT  9547.5 175667.5 9612.5 175292.5 ;
      RECT  9737.5 176552.5 9802.5 175667.5 ;
      RECT  9547.5 175667.5 9612.5 175532.5 ;
      RECT  9737.5 175667.5 9802.5 175532.5 ;
      RECT  9737.5 175667.5 9802.5 175532.5 ;
      RECT  9547.5 175667.5 9612.5 175532.5 ;
      RECT  9547.5 176552.5 9612.5 176417.5 ;
      RECT  9737.5 176552.5 9802.5 176417.5 ;
      RECT  9737.5 176552.5 9802.5 176417.5 ;
      RECT  9547.5 176552.5 9612.5 176417.5 ;
      RECT  9907.5 175577.5 9972.5 175442.5 ;
      RECT  9907.5 176552.5 9972.5 176417.5 ;
      RECT  9605.0 176110.0 9670.0 175975.0 ;
      RECT  9605.0 176110.0 9670.0 175975.0 ;
      RECT  9770.0 176075.0 9835.0 176010.0 ;
      RECT  9480.0 175357.5 10040.0 175292.5 ;
      RECT  9480.0 176702.5 10040.0 176637.5 ;
      RECT  10107.5 176507.5 10172.5 176702.5 ;
      RECT  10107.5 175667.5 10172.5 175292.5 ;
      RECT  10487.5 175667.5 10552.5 175292.5 ;
      RECT  10657.5 175510.0 10722.5 175325.0 ;
      RECT  10657.5 176670.0 10722.5 176485.0 ;
      RECT  10107.5 175667.5 10172.5 175532.5 ;
      RECT  10297.5 175667.5 10362.5 175532.5 ;
      RECT  10297.5 175667.5 10362.5 175532.5 ;
      RECT  10107.5 175667.5 10172.5 175532.5 ;
      RECT  10297.5 175667.5 10362.5 175532.5 ;
      RECT  10487.5 175667.5 10552.5 175532.5 ;
      RECT  10487.5 175667.5 10552.5 175532.5 ;
      RECT  10297.5 175667.5 10362.5 175532.5 ;
      RECT  10107.5 176507.5 10172.5 176372.5 ;
      RECT  10297.5 176507.5 10362.5 176372.5 ;
      RECT  10297.5 176507.5 10362.5 176372.5 ;
      RECT  10107.5 176507.5 10172.5 176372.5 ;
      RECT  10297.5 176507.5 10362.5 176372.5 ;
      RECT  10487.5 176507.5 10552.5 176372.5 ;
      RECT  10487.5 176507.5 10552.5 176372.5 ;
      RECT  10297.5 176507.5 10362.5 176372.5 ;
      RECT  10657.5 175577.5 10722.5 175442.5 ;
      RECT  10657.5 176552.5 10722.5 176417.5 ;
      RECT  10492.5 176277.5 10357.5 176212.5 ;
      RECT  10235.0 176062.5 10100.0 175997.5 ;
      RECT  10297.5 175667.5 10362.5 175532.5 ;
      RECT  10487.5 176507.5 10552.5 176372.5 ;
      RECT  10587.5 176062.5 10452.5 175997.5 ;
      RECT  10100.0 176062.5 10235.0 175997.5 ;
      RECT  10357.5 176277.5 10492.5 176212.5 ;
      RECT  10452.5 176062.5 10587.5 175997.5 ;
      RECT  10040.0 175357.5 10960.0 175292.5 ;
      RECT  10040.0 176702.5 10960.0 176637.5 ;
      RECT  11387.5 175510.0 11452.5 175325.0 ;
      RECT  11387.5 176670.0 11452.5 176485.0 ;
      RECT  11027.5 176552.5 11092.5 176702.5 ;
      RECT  11027.5 175667.5 11092.5 175292.5 ;
      RECT  11217.5 176552.5 11282.5 175667.5 ;
      RECT  11027.5 175667.5 11092.5 175532.5 ;
      RECT  11217.5 175667.5 11282.5 175532.5 ;
      RECT  11217.5 175667.5 11282.5 175532.5 ;
      RECT  11027.5 175667.5 11092.5 175532.5 ;
      RECT  11027.5 176552.5 11092.5 176417.5 ;
      RECT  11217.5 176552.5 11282.5 176417.5 ;
      RECT  11217.5 176552.5 11282.5 176417.5 ;
      RECT  11027.5 176552.5 11092.5 176417.5 ;
      RECT  11387.5 175577.5 11452.5 175442.5 ;
      RECT  11387.5 176552.5 11452.5 176417.5 ;
      RECT  11085.0 176110.0 11150.0 175975.0 ;
      RECT  11085.0 176110.0 11150.0 175975.0 ;
      RECT  11250.0 176075.0 11315.0 176010.0 ;
      RECT  10960.0 175357.5 11520.0 175292.5 ;
      RECT  10960.0 176702.5 11520.0 176637.5 ;
      RECT  9222.5 175975.0 9287.5 176110.0 ;
      RECT  9362.5 176247.5 9427.5 176382.5 ;
      RECT  10357.5 176212.5 10222.5 176277.5 ;
      RECT  9907.5 177830.0 9972.5 178015.0 ;
      RECT  9907.5 176670.0 9972.5 176855.0 ;
      RECT  9547.5 176787.5 9612.5 176637.5 ;
      RECT  9547.5 177672.5 9612.5 178047.5 ;
      RECT  9737.5 176787.5 9802.5 177672.5 ;
      RECT  9547.5 177672.5 9612.5 177807.5 ;
      RECT  9737.5 177672.5 9802.5 177807.5 ;
      RECT  9737.5 177672.5 9802.5 177807.5 ;
      RECT  9547.5 177672.5 9612.5 177807.5 ;
      RECT  9547.5 176787.5 9612.5 176922.5 ;
      RECT  9737.5 176787.5 9802.5 176922.5 ;
      RECT  9737.5 176787.5 9802.5 176922.5 ;
      RECT  9547.5 176787.5 9612.5 176922.5 ;
      RECT  9907.5 177762.5 9972.5 177897.5 ;
      RECT  9907.5 176787.5 9972.5 176922.5 ;
      RECT  9605.0 177230.0 9670.0 177365.0 ;
      RECT  9605.0 177230.0 9670.0 177365.0 ;
      RECT  9770.0 177265.0 9835.0 177330.0 ;
      RECT  9480.0 177982.5 10040.0 178047.5 ;
      RECT  9480.0 176637.5 10040.0 176702.5 ;
      RECT  10107.5 176832.5 10172.5 176637.5 ;
      RECT  10107.5 177672.5 10172.5 178047.5 ;
      RECT  10487.5 177672.5 10552.5 178047.5 ;
      RECT  10657.5 177830.0 10722.5 178015.0 ;
      RECT  10657.5 176670.0 10722.5 176855.0 ;
      RECT  10107.5 177672.5 10172.5 177807.5 ;
      RECT  10297.5 177672.5 10362.5 177807.5 ;
      RECT  10297.5 177672.5 10362.5 177807.5 ;
      RECT  10107.5 177672.5 10172.5 177807.5 ;
      RECT  10297.5 177672.5 10362.5 177807.5 ;
      RECT  10487.5 177672.5 10552.5 177807.5 ;
      RECT  10487.5 177672.5 10552.5 177807.5 ;
      RECT  10297.5 177672.5 10362.5 177807.5 ;
      RECT  10107.5 176832.5 10172.5 176967.5 ;
      RECT  10297.5 176832.5 10362.5 176967.5 ;
      RECT  10297.5 176832.5 10362.5 176967.5 ;
      RECT  10107.5 176832.5 10172.5 176967.5 ;
      RECT  10297.5 176832.5 10362.5 176967.5 ;
      RECT  10487.5 176832.5 10552.5 176967.5 ;
      RECT  10487.5 176832.5 10552.5 176967.5 ;
      RECT  10297.5 176832.5 10362.5 176967.5 ;
      RECT  10657.5 177762.5 10722.5 177897.5 ;
      RECT  10657.5 176787.5 10722.5 176922.5 ;
      RECT  10492.5 177062.5 10357.5 177127.5 ;
      RECT  10235.0 177277.5 10100.0 177342.5 ;
      RECT  10297.5 177672.5 10362.5 177807.5 ;
      RECT  10487.5 176832.5 10552.5 176967.5 ;
      RECT  10587.5 177277.5 10452.5 177342.5 ;
      RECT  10100.0 177277.5 10235.0 177342.5 ;
      RECT  10357.5 177062.5 10492.5 177127.5 ;
      RECT  10452.5 177277.5 10587.5 177342.5 ;
      RECT  10040.0 177982.5 10960.0 178047.5 ;
      RECT  10040.0 176637.5 10960.0 176702.5 ;
      RECT  11387.5 177830.0 11452.5 178015.0 ;
      RECT  11387.5 176670.0 11452.5 176855.0 ;
      RECT  11027.5 176787.5 11092.5 176637.5 ;
      RECT  11027.5 177672.5 11092.5 178047.5 ;
      RECT  11217.5 176787.5 11282.5 177672.5 ;
      RECT  11027.5 177672.5 11092.5 177807.5 ;
      RECT  11217.5 177672.5 11282.5 177807.5 ;
      RECT  11217.5 177672.5 11282.5 177807.5 ;
      RECT  11027.5 177672.5 11092.5 177807.5 ;
      RECT  11027.5 176787.5 11092.5 176922.5 ;
      RECT  11217.5 176787.5 11282.5 176922.5 ;
      RECT  11217.5 176787.5 11282.5 176922.5 ;
      RECT  11027.5 176787.5 11092.5 176922.5 ;
      RECT  11387.5 177762.5 11452.5 177897.5 ;
      RECT  11387.5 176787.5 11452.5 176922.5 ;
      RECT  11085.0 177230.0 11150.0 177365.0 ;
      RECT  11085.0 177230.0 11150.0 177365.0 ;
      RECT  11250.0 177265.0 11315.0 177330.0 ;
      RECT  10960.0 177982.5 11520.0 178047.5 ;
      RECT  10960.0 176637.5 11520.0 176702.5 ;
      RECT  9222.5 177230.0 9287.5 177365.0 ;
      RECT  9362.5 176957.5 9427.5 177092.5 ;
      RECT  10357.5 177062.5 10222.5 177127.5 ;
      RECT  9907.5 178200.0 9972.5 178015.0 ;
      RECT  9907.5 179360.0 9972.5 179175.0 ;
      RECT  9547.5 179242.5 9612.5 179392.5 ;
      RECT  9547.5 178357.5 9612.5 177982.5 ;
      RECT  9737.5 179242.5 9802.5 178357.5 ;
      RECT  9547.5 178357.5 9612.5 178222.5 ;
      RECT  9737.5 178357.5 9802.5 178222.5 ;
      RECT  9737.5 178357.5 9802.5 178222.5 ;
      RECT  9547.5 178357.5 9612.5 178222.5 ;
      RECT  9547.5 179242.5 9612.5 179107.5 ;
      RECT  9737.5 179242.5 9802.5 179107.5 ;
      RECT  9737.5 179242.5 9802.5 179107.5 ;
      RECT  9547.5 179242.5 9612.5 179107.5 ;
      RECT  9907.5 178267.5 9972.5 178132.5 ;
      RECT  9907.5 179242.5 9972.5 179107.5 ;
      RECT  9605.0 178800.0 9670.0 178665.0 ;
      RECT  9605.0 178800.0 9670.0 178665.0 ;
      RECT  9770.0 178765.0 9835.0 178700.0 ;
      RECT  9480.0 178047.5 10040.0 177982.5 ;
      RECT  9480.0 179392.5 10040.0 179327.5 ;
      RECT  10107.5 179197.5 10172.5 179392.5 ;
      RECT  10107.5 178357.5 10172.5 177982.5 ;
      RECT  10487.5 178357.5 10552.5 177982.5 ;
      RECT  10657.5 178200.0 10722.5 178015.0 ;
      RECT  10657.5 179360.0 10722.5 179175.0 ;
      RECT  10107.5 178357.5 10172.5 178222.5 ;
      RECT  10297.5 178357.5 10362.5 178222.5 ;
      RECT  10297.5 178357.5 10362.5 178222.5 ;
      RECT  10107.5 178357.5 10172.5 178222.5 ;
      RECT  10297.5 178357.5 10362.5 178222.5 ;
      RECT  10487.5 178357.5 10552.5 178222.5 ;
      RECT  10487.5 178357.5 10552.5 178222.5 ;
      RECT  10297.5 178357.5 10362.5 178222.5 ;
      RECT  10107.5 179197.5 10172.5 179062.5 ;
      RECT  10297.5 179197.5 10362.5 179062.5 ;
      RECT  10297.5 179197.5 10362.5 179062.5 ;
      RECT  10107.5 179197.5 10172.5 179062.5 ;
      RECT  10297.5 179197.5 10362.5 179062.5 ;
      RECT  10487.5 179197.5 10552.5 179062.5 ;
      RECT  10487.5 179197.5 10552.5 179062.5 ;
      RECT  10297.5 179197.5 10362.5 179062.5 ;
      RECT  10657.5 178267.5 10722.5 178132.5 ;
      RECT  10657.5 179242.5 10722.5 179107.5 ;
      RECT  10492.5 178967.5 10357.5 178902.5 ;
      RECT  10235.0 178752.5 10100.0 178687.5 ;
      RECT  10297.5 178357.5 10362.5 178222.5 ;
      RECT  10487.5 179197.5 10552.5 179062.5 ;
      RECT  10587.5 178752.5 10452.5 178687.5 ;
      RECT  10100.0 178752.5 10235.0 178687.5 ;
      RECT  10357.5 178967.5 10492.5 178902.5 ;
      RECT  10452.5 178752.5 10587.5 178687.5 ;
      RECT  10040.0 178047.5 10960.0 177982.5 ;
      RECT  10040.0 179392.5 10960.0 179327.5 ;
      RECT  11387.5 178200.0 11452.5 178015.0 ;
      RECT  11387.5 179360.0 11452.5 179175.0 ;
      RECT  11027.5 179242.5 11092.5 179392.5 ;
      RECT  11027.5 178357.5 11092.5 177982.5 ;
      RECT  11217.5 179242.5 11282.5 178357.5 ;
      RECT  11027.5 178357.5 11092.5 178222.5 ;
      RECT  11217.5 178357.5 11282.5 178222.5 ;
      RECT  11217.5 178357.5 11282.5 178222.5 ;
      RECT  11027.5 178357.5 11092.5 178222.5 ;
      RECT  11027.5 179242.5 11092.5 179107.5 ;
      RECT  11217.5 179242.5 11282.5 179107.5 ;
      RECT  11217.5 179242.5 11282.5 179107.5 ;
      RECT  11027.5 179242.5 11092.5 179107.5 ;
      RECT  11387.5 178267.5 11452.5 178132.5 ;
      RECT  11387.5 179242.5 11452.5 179107.5 ;
      RECT  11085.0 178800.0 11150.0 178665.0 ;
      RECT  11085.0 178800.0 11150.0 178665.0 ;
      RECT  11250.0 178765.0 11315.0 178700.0 ;
      RECT  10960.0 178047.5 11520.0 177982.5 ;
      RECT  10960.0 179392.5 11520.0 179327.5 ;
      RECT  9222.5 178665.0 9287.5 178800.0 ;
      RECT  9362.5 178937.5 9427.5 179072.5 ;
      RECT  10357.5 178902.5 10222.5 178967.5 ;
      RECT  9907.5 180520.0 9972.5 180705.0 ;
      RECT  9907.5 179360.0 9972.5 179545.0 ;
      RECT  9547.5 179477.5 9612.5 179327.5 ;
      RECT  9547.5 180362.5 9612.5 180737.5 ;
      RECT  9737.5 179477.5 9802.5 180362.5 ;
      RECT  9547.5 180362.5 9612.5 180497.5 ;
      RECT  9737.5 180362.5 9802.5 180497.5 ;
      RECT  9737.5 180362.5 9802.5 180497.5 ;
      RECT  9547.5 180362.5 9612.5 180497.5 ;
      RECT  9547.5 179477.5 9612.5 179612.5 ;
      RECT  9737.5 179477.5 9802.5 179612.5 ;
      RECT  9737.5 179477.5 9802.5 179612.5 ;
      RECT  9547.5 179477.5 9612.5 179612.5 ;
      RECT  9907.5 180452.5 9972.5 180587.5 ;
      RECT  9907.5 179477.5 9972.5 179612.5 ;
      RECT  9605.0 179920.0 9670.0 180055.0 ;
      RECT  9605.0 179920.0 9670.0 180055.0 ;
      RECT  9770.0 179955.0 9835.0 180020.0 ;
      RECT  9480.0 180672.5 10040.0 180737.5 ;
      RECT  9480.0 179327.5 10040.0 179392.5 ;
      RECT  10107.5 179522.5 10172.5 179327.5 ;
      RECT  10107.5 180362.5 10172.5 180737.5 ;
      RECT  10487.5 180362.5 10552.5 180737.5 ;
      RECT  10657.5 180520.0 10722.5 180705.0 ;
      RECT  10657.5 179360.0 10722.5 179545.0 ;
      RECT  10107.5 180362.5 10172.5 180497.5 ;
      RECT  10297.5 180362.5 10362.5 180497.5 ;
      RECT  10297.5 180362.5 10362.5 180497.5 ;
      RECT  10107.5 180362.5 10172.5 180497.5 ;
      RECT  10297.5 180362.5 10362.5 180497.5 ;
      RECT  10487.5 180362.5 10552.5 180497.5 ;
      RECT  10487.5 180362.5 10552.5 180497.5 ;
      RECT  10297.5 180362.5 10362.5 180497.5 ;
      RECT  10107.5 179522.5 10172.5 179657.5 ;
      RECT  10297.5 179522.5 10362.5 179657.5 ;
      RECT  10297.5 179522.5 10362.5 179657.5 ;
      RECT  10107.5 179522.5 10172.5 179657.5 ;
      RECT  10297.5 179522.5 10362.5 179657.5 ;
      RECT  10487.5 179522.5 10552.5 179657.5 ;
      RECT  10487.5 179522.5 10552.5 179657.5 ;
      RECT  10297.5 179522.5 10362.5 179657.5 ;
      RECT  10657.5 180452.5 10722.5 180587.5 ;
      RECT  10657.5 179477.5 10722.5 179612.5 ;
      RECT  10492.5 179752.5 10357.5 179817.5 ;
      RECT  10235.0 179967.5 10100.0 180032.5 ;
      RECT  10297.5 180362.5 10362.5 180497.5 ;
      RECT  10487.5 179522.5 10552.5 179657.5 ;
      RECT  10587.5 179967.5 10452.5 180032.5 ;
      RECT  10100.0 179967.5 10235.0 180032.5 ;
      RECT  10357.5 179752.5 10492.5 179817.5 ;
      RECT  10452.5 179967.5 10587.5 180032.5 ;
      RECT  10040.0 180672.5 10960.0 180737.5 ;
      RECT  10040.0 179327.5 10960.0 179392.5 ;
      RECT  11387.5 180520.0 11452.5 180705.0 ;
      RECT  11387.5 179360.0 11452.5 179545.0 ;
      RECT  11027.5 179477.5 11092.5 179327.5 ;
      RECT  11027.5 180362.5 11092.5 180737.5 ;
      RECT  11217.5 179477.5 11282.5 180362.5 ;
      RECT  11027.5 180362.5 11092.5 180497.5 ;
      RECT  11217.5 180362.5 11282.5 180497.5 ;
      RECT  11217.5 180362.5 11282.5 180497.5 ;
      RECT  11027.5 180362.5 11092.5 180497.5 ;
      RECT  11027.5 179477.5 11092.5 179612.5 ;
      RECT  11217.5 179477.5 11282.5 179612.5 ;
      RECT  11217.5 179477.5 11282.5 179612.5 ;
      RECT  11027.5 179477.5 11092.5 179612.5 ;
      RECT  11387.5 180452.5 11452.5 180587.5 ;
      RECT  11387.5 179477.5 11452.5 179612.5 ;
      RECT  11085.0 179920.0 11150.0 180055.0 ;
      RECT  11085.0 179920.0 11150.0 180055.0 ;
      RECT  11250.0 179955.0 11315.0 180020.0 ;
      RECT  10960.0 180672.5 11520.0 180737.5 ;
      RECT  10960.0 179327.5 11520.0 179392.5 ;
      RECT  9222.5 179920.0 9287.5 180055.0 ;
      RECT  9362.5 179647.5 9427.5 179782.5 ;
      RECT  10357.5 179752.5 10222.5 179817.5 ;
      RECT  9907.5 180890.0 9972.5 180705.0 ;
      RECT  9907.5 182050.0 9972.5 181865.0 ;
      RECT  9547.5 181932.5 9612.5 182082.5 ;
      RECT  9547.5 181047.5 9612.5 180672.5 ;
      RECT  9737.5 181932.5 9802.5 181047.5 ;
      RECT  9547.5 181047.5 9612.5 180912.5 ;
      RECT  9737.5 181047.5 9802.5 180912.5 ;
      RECT  9737.5 181047.5 9802.5 180912.5 ;
      RECT  9547.5 181047.5 9612.5 180912.5 ;
      RECT  9547.5 181932.5 9612.5 181797.5 ;
      RECT  9737.5 181932.5 9802.5 181797.5 ;
      RECT  9737.5 181932.5 9802.5 181797.5 ;
      RECT  9547.5 181932.5 9612.5 181797.5 ;
      RECT  9907.5 180957.5 9972.5 180822.5 ;
      RECT  9907.5 181932.5 9972.5 181797.5 ;
      RECT  9605.0 181490.0 9670.0 181355.0 ;
      RECT  9605.0 181490.0 9670.0 181355.0 ;
      RECT  9770.0 181455.0 9835.0 181390.0 ;
      RECT  9480.0 180737.5 10040.0 180672.5 ;
      RECT  9480.0 182082.5 10040.0 182017.5 ;
      RECT  10107.5 181887.5 10172.5 182082.5 ;
      RECT  10107.5 181047.5 10172.5 180672.5 ;
      RECT  10487.5 181047.5 10552.5 180672.5 ;
      RECT  10657.5 180890.0 10722.5 180705.0 ;
      RECT  10657.5 182050.0 10722.5 181865.0 ;
      RECT  10107.5 181047.5 10172.5 180912.5 ;
      RECT  10297.5 181047.5 10362.5 180912.5 ;
      RECT  10297.5 181047.5 10362.5 180912.5 ;
      RECT  10107.5 181047.5 10172.5 180912.5 ;
      RECT  10297.5 181047.5 10362.5 180912.5 ;
      RECT  10487.5 181047.5 10552.5 180912.5 ;
      RECT  10487.5 181047.5 10552.5 180912.5 ;
      RECT  10297.5 181047.5 10362.5 180912.5 ;
      RECT  10107.5 181887.5 10172.5 181752.5 ;
      RECT  10297.5 181887.5 10362.5 181752.5 ;
      RECT  10297.5 181887.5 10362.5 181752.5 ;
      RECT  10107.5 181887.5 10172.5 181752.5 ;
      RECT  10297.5 181887.5 10362.5 181752.5 ;
      RECT  10487.5 181887.5 10552.5 181752.5 ;
      RECT  10487.5 181887.5 10552.5 181752.5 ;
      RECT  10297.5 181887.5 10362.5 181752.5 ;
      RECT  10657.5 180957.5 10722.5 180822.5 ;
      RECT  10657.5 181932.5 10722.5 181797.5 ;
      RECT  10492.5 181657.5 10357.5 181592.5 ;
      RECT  10235.0 181442.5 10100.0 181377.5 ;
      RECT  10297.5 181047.5 10362.5 180912.5 ;
      RECT  10487.5 181887.5 10552.5 181752.5 ;
      RECT  10587.5 181442.5 10452.5 181377.5 ;
      RECT  10100.0 181442.5 10235.0 181377.5 ;
      RECT  10357.5 181657.5 10492.5 181592.5 ;
      RECT  10452.5 181442.5 10587.5 181377.5 ;
      RECT  10040.0 180737.5 10960.0 180672.5 ;
      RECT  10040.0 182082.5 10960.0 182017.5 ;
      RECT  11387.5 180890.0 11452.5 180705.0 ;
      RECT  11387.5 182050.0 11452.5 181865.0 ;
      RECT  11027.5 181932.5 11092.5 182082.5 ;
      RECT  11027.5 181047.5 11092.5 180672.5 ;
      RECT  11217.5 181932.5 11282.5 181047.5 ;
      RECT  11027.5 181047.5 11092.5 180912.5 ;
      RECT  11217.5 181047.5 11282.5 180912.5 ;
      RECT  11217.5 181047.5 11282.5 180912.5 ;
      RECT  11027.5 181047.5 11092.5 180912.5 ;
      RECT  11027.5 181932.5 11092.5 181797.5 ;
      RECT  11217.5 181932.5 11282.5 181797.5 ;
      RECT  11217.5 181932.5 11282.5 181797.5 ;
      RECT  11027.5 181932.5 11092.5 181797.5 ;
      RECT  11387.5 180957.5 11452.5 180822.5 ;
      RECT  11387.5 181932.5 11452.5 181797.5 ;
      RECT  11085.0 181490.0 11150.0 181355.0 ;
      RECT  11085.0 181490.0 11150.0 181355.0 ;
      RECT  11250.0 181455.0 11315.0 181390.0 ;
      RECT  10960.0 180737.5 11520.0 180672.5 ;
      RECT  10960.0 182082.5 11520.0 182017.5 ;
      RECT  9222.5 181355.0 9287.5 181490.0 ;
      RECT  9362.5 181627.5 9427.5 181762.5 ;
      RECT  10357.5 181592.5 10222.5 181657.5 ;
      RECT  9907.5 183210.0 9972.5 183395.0 ;
      RECT  9907.5 182050.0 9972.5 182235.0 ;
      RECT  9547.5 182167.5 9612.5 182017.5 ;
      RECT  9547.5 183052.5 9612.5 183427.5 ;
      RECT  9737.5 182167.5 9802.5 183052.5 ;
      RECT  9547.5 183052.5 9612.5 183187.5 ;
      RECT  9737.5 183052.5 9802.5 183187.5 ;
      RECT  9737.5 183052.5 9802.5 183187.5 ;
      RECT  9547.5 183052.5 9612.5 183187.5 ;
      RECT  9547.5 182167.5 9612.5 182302.5 ;
      RECT  9737.5 182167.5 9802.5 182302.5 ;
      RECT  9737.5 182167.5 9802.5 182302.5 ;
      RECT  9547.5 182167.5 9612.5 182302.5 ;
      RECT  9907.5 183142.5 9972.5 183277.5 ;
      RECT  9907.5 182167.5 9972.5 182302.5 ;
      RECT  9605.0 182610.0 9670.0 182745.0 ;
      RECT  9605.0 182610.0 9670.0 182745.0 ;
      RECT  9770.0 182645.0 9835.0 182710.0 ;
      RECT  9480.0 183362.5 10040.0 183427.5 ;
      RECT  9480.0 182017.5 10040.0 182082.5 ;
      RECT  10107.5 182212.5 10172.5 182017.5 ;
      RECT  10107.5 183052.5 10172.5 183427.5 ;
      RECT  10487.5 183052.5 10552.5 183427.5 ;
      RECT  10657.5 183210.0 10722.5 183395.0 ;
      RECT  10657.5 182050.0 10722.5 182235.0 ;
      RECT  10107.5 183052.5 10172.5 183187.5 ;
      RECT  10297.5 183052.5 10362.5 183187.5 ;
      RECT  10297.5 183052.5 10362.5 183187.5 ;
      RECT  10107.5 183052.5 10172.5 183187.5 ;
      RECT  10297.5 183052.5 10362.5 183187.5 ;
      RECT  10487.5 183052.5 10552.5 183187.5 ;
      RECT  10487.5 183052.5 10552.5 183187.5 ;
      RECT  10297.5 183052.5 10362.5 183187.5 ;
      RECT  10107.5 182212.5 10172.5 182347.5 ;
      RECT  10297.5 182212.5 10362.5 182347.5 ;
      RECT  10297.5 182212.5 10362.5 182347.5 ;
      RECT  10107.5 182212.5 10172.5 182347.5 ;
      RECT  10297.5 182212.5 10362.5 182347.5 ;
      RECT  10487.5 182212.5 10552.5 182347.5 ;
      RECT  10487.5 182212.5 10552.5 182347.5 ;
      RECT  10297.5 182212.5 10362.5 182347.5 ;
      RECT  10657.5 183142.5 10722.5 183277.5 ;
      RECT  10657.5 182167.5 10722.5 182302.5 ;
      RECT  10492.5 182442.5 10357.5 182507.5 ;
      RECT  10235.0 182657.5 10100.0 182722.5 ;
      RECT  10297.5 183052.5 10362.5 183187.5 ;
      RECT  10487.5 182212.5 10552.5 182347.5 ;
      RECT  10587.5 182657.5 10452.5 182722.5 ;
      RECT  10100.0 182657.5 10235.0 182722.5 ;
      RECT  10357.5 182442.5 10492.5 182507.5 ;
      RECT  10452.5 182657.5 10587.5 182722.5 ;
      RECT  10040.0 183362.5 10960.0 183427.5 ;
      RECT  10040.0 182017.5 10960.0 182082.5 ;
      RECT  11387.5 183210.0 11452.5 183395.0 ;
      RECT  11387.5 182050.0 11452.5 182235.0 ;
      RECT  11027.5 182167.5 11092.5 182017.5 ;
      RECT  11027.5 183052.5 11092.5 183427.5 ;
      RECT  11217.5 182167.5 11282.5 183052.5 ;
      RECT  11027.5 183052.5 11092.5 183187.5 ;
      RECT  11217.5 183052.5 11282.5 183187.5 ;
      RECT  11217.5 183052.5 11282.5 183187.5 ;
      RECT  11027.5 183052.5 11092.5 183187.5 ;
      RECT  11027.5 182167.5 11092.5 182302.5 ;
      RECT  11217.5 182167.5 11282.5 182302.5 ;
      RECT  11217.5 182167.5 11282.5 182302.5 ;
      RECT  11027.5 182167.5 11092.5 182302.5 ;
      RECT  11387.5 183142.5 11452.5 183277.5 ;
      RECT  11387.5 182167.5 11452.5 182302.5 ;
      RECT  11085.0 182610.0 11150.0 182745.0 ;
      RECT  11085.0 182610.0 11150.0 182745.0 ;
      RECT  11250.0 182645.0 11315.0 182710.0 ;
      RECT  10960.0 183362.5 11520.0 183427.5 ;
      RECT  10960.0 182017.5 11520.0 182082.5 ;
      RECT  9222.5 182610.0 9287.5 182745.0 ;
      RECT  9362.5 182337.5 9427.5 182472.5 ;
      RECT  10357.5 182442.5 10222.5 182507.5 ;
      RECT  9907.5 183580.0 9972.5 183395.0 ;
      RECT  9907.5 184740.0 9972.5 184555.0 ;
      RECT  9547.5 184622.5 9612.5 184772.5 ;
      RECT  9547.5 183737.5 9612.5 183362.5 ;
      RECT  9737.5 184622.5 9802.5 183737.5 ;
      RECT  9547.5 183737.5 9612.5 183602.5 ;
      RECT  9737.5 183737.5 9802.5 183602.5 ;
      RECT  9737.5 183737.5 9802.5 183602.5 ;
      RECT  9547.5 183737.5 9612.5 183602.5 ;
      RECT  9547.5 184622.5 9612.5 184487.5 ;
      RECT  9737.5 184622.5 9802.5 184487.5 ;
      RECT  9737.5 184622.5 9802.5 184487.5 ;
      RECT  9547.5 184622.5 9612.5 184487.5 ;
      RECT  9907.5 183647.5 9972.5 183512.5 ;
      RECT  9907.5 184622.5 9972.5 184487.5 ;
      RECT  9605.0 184180.0 9670.0 184045.0 ;
      RECT  9605.0 184180.0 9670.0 184045.0 ;
      RECT  9770.0 184145.0 9835.0 184080.0 ;
      RECT  9480.0 183427.5 10040.0 183362.5 ;
      RECT  9480.0 184772.5 10040.0 184707.5 ;
      RECT  10107.5 184577.5 10172.5 184772.5 ;
      RECT  10107.5 183737.5 10172.5 183362.5 ;
      RECT  10487.5 183737.5 10552.5 183362.5 ;
      RECT  10657.5 183580.0 10722.5 183395.0 ;
      RECT  10657.5 184740.0 10722.5 184555.0 ;
      RECT  10107.5 183737.5 10172.5 183602.5 ;
      RECT  10297.5 183737.5 10362.5 183602.5 ;
      RECT  10297.5 183737.5 10362.5 183602.5 ;
      RECT  10107.5 183737.5 10172.5 183602.5 ;
      RECT  10297.5 183737.5 10362.5 183602.5 ;
      RECT  10487.5 183737.5 10552.5 183602.5 ;
      RECT  10487.5 183737.5 10552.5 183602.5 ;
      RECT  10297.5 183737.5 10362.5 183602.5 ;
      RECT  10107.5 184577.5 10172.5 184442.5 ;
      RECT  10297.5 184577.5 10362.5 184442.5 ;
      RECT  10297.5 184577.5 10362.5 184442.5 ;
      RECT  10107.5 184577.5 10172.5 184442.5 ;
      RECT  10297.5 184577.5 10362.5 184442.5 ;
      RECT  10487.5 184577.5 10552.5 184442.5 ;
      RECT  10487.5 184577.5 10552.5 184442.5 ;
      RECT  10297.5 184577.5 10362.5 184442.5 ;
      RECT  10657.5 183647.5 10722.5 183512.5 ;
      RECT  10657.5 184622.5 10722.5 184487.5 ;
      RECT  10492.5 184347.5 10357.5 184282.5 ;
      RECT  10235.0 184132.5 10100.0 184067.5 ;
      RECT  10297.5 183737.5 10362.5 183602.5 ;
      RECT  10487.5 184577.5 10552.5 184442.5 ;
      RECT  10587.5 184132.5 10452.5 184067.5 ;
      RECT  10100.0 184132.5 10235.0 184067.5 ;
      RECT  10357.5 184347.5 10492.5 184282.5 ;
      RECT  10452.5 184132.5 10587.5 184067.5 ;
      RECT  10040.0 183427.5 10960.0 183362.5 ;
      RECT  10040.0 184772.5 10960.0 184707.5 ;
      RECT  11387.5 183580.0 11452.5 183395.0 ;
      RECT  11387.5 184740.0 11452.5 184555.0 ;
      RECT  11027.5 184622.5 11092.5 184772.5 ;
      RECT  11027.5 183737.5 11092.5 183362.5 ;
      RECT  11217.5 184622.5 11282.5 183737.5 ;
      RECT  11027.5 183737.5 11092.5 183602.5 ;
      RECT  11217.5 183737.5 11282.5 183602.5 ;
      RECT  11217.5 183737.5 11282.5 183602.5 ;
      RECT  11027.5 183737.5 11092.5 183602.5 ;
      RECT  11027.5 184622.5 11092.5 184487.5 ;
      RECT  11217.5 184622.5 11282.5 184487.5 ;
      RECT  11217.5 184622.5 11282.5 184487.5 ;
      RECT  11027.5 184622.5 11092.5 184487.5 ;
      RECT  11387.5 183647.5 11452.5 183512.5 ;
      RECT  11387.5 184622.5 11452.5 184487.5 ;
      RECT  11085.0 184180.0 11150.0 184045.0 ;
      RECT  11085.0 184180.0 11150.0 184045.0 ;
      RECT  11250.0 184145.0 11315.0 184080.0 ;
      RECT  10960.0 183427.5 11520.0 183362.5 ;
      RECT  10960.0 184772.5 11520.0 184707.5 ;
      RECT  9222.5 184045.0 9287.5 184180.0 ;
      RECT  9362.5 184317.5 9427.5 184452.5 ;
      RECT  10357.5 184282.5 10222.5 184347.5 ;
      RECT  9907.5 185900.0 9972.5 186085.0 ;
      RECT  9907.5 184740.0 9972.5 184925.0 ;
      RECT  9547.5 184857.5 9612.5 184707.5 ;
      RECT  9547.5 185742.5 9612.5 186117.5 ;
      RECT  9737.5 184857.5 9802.5 185742.5 ;
      RECT  9547.5 185742.5 9612.5 185877.5 ;
      RECT  9737.5 185742.5 9802.5 185877.5 ;
      RECT  9737.5 185742.5 9802.5 185877.5 ;
      RECT  9547.5 185742.5 9612.5 185877.5 ;
      RECT  9547.5 184857.5 9612.5 184992.5 ;
      RECT  9737.5 184857.5 9802.5 184992.5 ;
      RECT  9737.5 184857.5 9802.5 184992.5 ;
      RECT  9547.5 184857.5 9612.5 184992.5 ;
      RECT  9907.5 185832.5 9972.5 185967.5 ;
      RECT  9907.5 184857.5 9972.5 184992.5 ;
      RECT  9605.0 185300.0 9670.0 185435.0 ;
      RECT  9605.0 185300.0 9670.0 185435.0 ;
      RECT  9770.0 185335.0 9835.0 185400.0 ;
      RECT  9480.0 186052.5 10040.0 186117.5 ;
      RECT  9480.0 184707.5 10040.0 184772.5 ;
      RECT  10107.5 184902.5 10172.5 184707.5 ;
      RECT  10107.5 185742.5 10172.5 186117.5 ;
      RECT  10487.5 185742.5 10552.5 186117.5 ;
      RECT  10657.5 185900.0 10722.5 186085.0 ;
      RECT  10657.5 184740.0 10722.5 184925.0 ;
      RECT  10107.5 185742.5 10172.5 185877.5 ;
      RECT  10297.5 185742.5 10362.5 185877.5 ;
      RECT  10297.5 185742.5 10362.5 185877.5 ;
      RECT  10107.5 185742.5 10172.5 185877.5 ;
      RECT  10297.5 185742.5 10362.5 185877.5 ;
      RECT  10487.5 185742.5 10552.5 185877.5 ;
      RECT  10487.5 185742.5 10552.5 185877.5 ;
      RECT  10297.5 185742.5 10362.5 185877.5 ;
      RECT  10107.5 184902.5 10172.5 185037.5 ;
      RECT  10297.5 184902.5 10362.5 185037.5 ;
      RECT  10297.5 184902.5 10362.5 185037.5 ;
      RECT  10107.5 184902.5 10172.5 185037.5 ;
      RECT  10297.5 184902.5 10362.5 185037.5 ;
      RECT  10487.5 184902.5 10552.5 185037.5 ;
      RECT  10487.5 184902.5 10552.5 185037.5 ;
      RECT  10297.5 184902.5 10362.5 185037.5 ;
      RECT  10657.5 185832.5 10722.5 185967.5 ;
      RECT  10657.5 184857.5 10722.5 184992.5 ;
      RECT  10492.5 185132.5 10357.5 185197.5 ;
      RECT  10235.0 185347.5 10100.0 185412.5 ;
      RECT  10297.5 185742.5 10362.5 185877.5 ;
      RECT  10487.5 184902.5 10552.5 185037.5 ;
      RECT  10587.5 185347.5 10452.5 185412.5 ;
      RECT  10100.0 185347.5 10235.0 185412.5 ;
      RECT  10357.5 185132.5 10492.5 185197.5 ;
      RECT  10452.5 185347.5 10587.5 185412.5 ;
      RECT  10040.0 186052.5 10960.0 186117.5 ;
      RECT  10040.0 184707.5 10960.0 184772.5 ;
      RECT  11387.5 185900.0 11452.5 186085.0 ;
      RECT  11387.5 184740.0 11452.5 184925.0 ;
      RECT  11027.5 184857.5 11092.5 184707.5 ;
      RECT  11027.5 185742.5 11092.5 186117.5 ;
      RECT  11217.5 184857.5 11282.5 185742.5 ;
      RECT  11027.5 185742.5 11092.5 185877.5 ;
      RECT  11217.5 185742.5 11282.5 185877.5 ;
      RECT  11217.5 185742.5 11282.5 185877.5 ;
      RECT  11027.5 185742.5 11092.5 185877.5 ;
      RECT  11027.5 184857.5 11092.5 184992.5 ;
      RECT  11217.5 184857.5 11282.5 184992.5 ;
      RECT  11217.5 184857.5 11282.5 184992.5 ;
      RECT  11027.5 184857.5 11092.5 184992.5 ;
      RECT  11387.5 185832.5 11452.5 185967.5 ;
      RECT  11387.5 184857.5 11452.5 184992.5 ;
      RECT  11085.0 185300.0 11150.0 185435.0 ;
      RECT  11085.0 185300.0 11150.0 185435.0 ;
      RECT  11250.0 185335.0 11315.0 185400.0 ;
      RECT  10960.0 186052.5 11520.0 186117.5 ;
      RECT  10960.0 184707.5 11520.0 184772.5 ;
      RECT  9222.5 185300.0 9287.5 185435.0 ;
      RECT  9362.5 185027.5 9427.5 185162.5 ;
      RECT  10357.5 185132.5 10222.5 185197.5 ;
      RECT  9907.5 186270.0 9972.5 186085.0 ;
      RECT  9907.5 187430.0 9972.5 187245.0 ;
      RECT  9547.5 187312.5 9612.5 187462.5 ;
      RECT  9547.5 186427.5 9612.5 186052.5 ;
      RECT  9737.5 187312.5 9802.5 186427.5 ;
      RECT  9547.5 186427.5 9612.5 186292.5 ;
      RECT  9737.5 186427.5 9802.5 186292.5 ;
      RECT  9737.5 186427.5 9802.5 186292.5 ;
      RECT  9547.5 186427.5 9612.5 186292.5 ;
      RECT  9547.5 187312.5 9612.5 187177.5 ;
      RECT  9737.5 187312.5 9802.5 187177.5 ;
      RECT  9737.5 187312.5 9802.5 187177.5 ;
      RECT  9547.5 187312.5 9612.5 187177.5 ;
      RECT  9907.5 186337.5 9972.5 186202.5 ;
      RECT  9907.5 187312.5 9972.5 187177.5 ;
      RECT  9605.0 186870.0 9670.0 186735.0 ;
      RECT  9605.0 186870.0 9670.0 186735.0 ;
      RECT  9770.0 186835.0 9835.0 186770.0 ;
      RECT  9480.0 186117.5 10040.0 186052.5 ;
      RECT  9480.0 187462.5 10040.0 187397.5 ;
      RECT  10107.5 187267.5 10172.5 187462.5 ;
      RECT  10107.5 186427.5 10172.5 186052.5 ;
      RECT  10487.5 186427.5 10552.5 186052.5 ;
      RECT  10657.5 186270.0 10722.5 186085.0 ;
      RECT  10657.5 187430.0 10722.5 187245.0 ;
      RECT  10107.5 186427.5 10172.5 186292.5 ;
      RECT  10297.5 186427.5 10362.5 186292.5 ;
      RECT  10297.5 186427.5 10362.5 186292.5 ;
      RECT  10107.5 186427.5 10172.5 186292.5 ;
      RECT  10297.5 186427.5 10362.5 186292.5 ;
      RECT  10487.5 186427.5 10552.5 186292.5 ;
      RECT  10487.5 186427.5 10552.5 186292.5 ;
      RECT  10297.5 186427.5 10362.5 186292.5 ;
      RECT  10107.5 187267.5 10172.5 187132.5 ;
      RECT  10297.5 187267.5 10362.5 187132.5 ;
      RECT  10297.5 187267.5 10362.5 187132.5 ;
      RECT  10107.5 187267.5 10172.5 187132.5 ;
      RECT  10297.5 187267.5 10362.5 187132.5 ;
      RECT  10487.5 187267.5 10552.5 187132.5 ;
      RECT  10487.5 187267.5 10552.5 187132.5 ;
      RECT  10297.5 187267.5 10362.5 187132.5 ;
      RECT  10657.5 186337.5 10722.5 186202.5 ;
      RECT  10657.5 187312.5 10722.5 187177.5 ;
      RECT  10492.5 187037.5 10357.5 186972.5 ;
      RECT  10235.0 186822.5 10100.0 186757.5 ;
      RECT  10297.5 186427.5 10362.5 186292.5 ;
      RECT  10487.5 187267.5 10552.5 187132.5 ;
      RECT  10587.5 186822.5 10452.5 186757.5 ;
      RECT  10100.0 186822.5 10235.0 186757.5 ;
      RECT  10357.5 187037.5 10492.5 186972.5 ;
      RECT  10452.5 186822.5 10587.5 186757.5 ;
      RECT  10040.0 186117.5 10960.0 186052.5 ;
      RECT  10040.0 187462.5 10960.0 187397.5 ;
      RECT  11387.5 186270.0 11452.5 186085.0 ;
      RECT  11387.5 187430.0 11452.5 187245.0 ;
      RECT  11027.5 187312.5 11092.5 187462.5 ;
      RECT  11027.5 186427.5 11092.5 186052.5 ;
      RECT  11217.5 187312.5 11282.5 186427.5 ;
      RECT  11027.5 186427.5 11092.5 186292.5 ;
      RECT  11217.5 186427.5 11282.5 186292.5 ;
      RECT  11217.5 186427.5 11282.5 186292.5 ;
      RECT  11027.5 186427.5 11092.5 186292.5 ;
      RECT  11027.5 187312.5 11092.5 187177.5 ;
      RECT  11217.5 187312.5 11282.5 187177.5 ;
      RECT  11217.5 187312.5 11282.5 187177.5 ;
      RECT  11027.5 187312.5 11092.5 187177.5 ;
      RECT  11387.5 186337.5 11452.5 186202.5 ;
      RECT  11387.5 187312.5 11452.5 187177.5 ;
      RECT  11085.0 186870.0 11150.0 186735.0 ;
      RECT  11085.0 186870.0 11150.0 186735.0 ;
      RECT  11250.0 186835.0 11315.0 186770.0 ;
      RECT  10960.0 186117.5 11520.0 186052.5 ;
      RECT  10960.0 187462.5 11520.0 187397.5 ;
      RECT  9222.5 186735.0 9287.5 186870.0 ;
      RECT  9362.5 187007.5 9427.5 187142.5 ;
      RECT  10357.5 186972.5 10222.5 187037.5 ;
      RECT  9907.5 188590.0 9972.5 188775.0 ;
      RECT  9907.5 187430.0 9972.5 187615.0 ;
      RECT  9547.5 187547.5 9612.5 187397.5 ;
      RECT  9547.5 188432.5 9612.5 188807.5 ;
      RECT  9737.5 187547.5 9802.5 188432.5 ;
      RECT  9547.5 188432.5 9612.5 188567.5 ;
      RECT  9737.5 188432.5 9802.5 188567.5 ;
      RECT  9737.5 188432.5 9802.5 188567.5 ;
      RECT  9547.5 188432.5 9612.5 188567.5 ;
      RECT  9547.5 187547.5 9612.5 187682.5 ;
      RECT  9737.5 187547.5 9802.5 187682.5 ;
      RECT  9737.5 187547.5 9802.5 187682.5 ;
      RECT  9547.5 187547.5 9612.5 187682.5 ;
      RECT  9907.5 188522.5 9972.5 188657.5 ;
      RECT  9907.5 187547.5 9972.5 187682.5 ;
      RECT  9605.0 187990.0 9670.0 188125.0 ;
      RECT  9605.0 187990.0 9670.0 188125.0 ;
      RECT  9770.0 188025.0 9835.0 188090.0 ;
      RECT  9480.0 188742.5 10040.0 188807.5 ;
      RECT  9480.0 187397.5 10040.0 187462.5 ;
      RECT  10107.5 187592.5 10172.5 187397.5 ;
      RECT  10107.5 188432.5 10172.5 188807.5 ;
      RECT  10487.5 188432.5 10552.5 188807.5 ;
      RECT  10657.5 188590.0 10722.5 188775.0 ;
      RECT  10657.5 187430.0 10722.5 187615.0 ;
      RECT  10107.5 188432.5 10172.5 188567.5 ;
      RECT  10297.5 188432.5 10362.5 188567.5 ;
      RECT  10297.5 188432.5 10362.5 188567.5 ;
      RECT  10107.5 188432.5 10172.5 188567.5 ;
      RECT  10297.5 188432.5 10362.5 188567.5 ;
      RECT  10487.5 188432.5 10552.5 188567.5 ;
      RECT  10487.5 188432.5 10552.5 188567.5 ;
      RECT  10297.5 188432.5 10362.5 188567.5 ;
      RECT  10107.5 187592.5 10172.5 187727.5 ;
      RECT  10297.5 187592.5 10362.5 187727.5 ;
      RECT  10297.5 187592.5 10362.5 187727.5 ;
      RECT  10107.5 187592.5 10172.5 187727.5 ;
      RECT  10297.5 187592.5 10362.5 187727.5 ;
      RECT  10487.5 187592.5 10552.5 187727.5 ;
      RECT  10487.5 187592.5 10552.5 187727.5 ;
      RECT  10297.5 187592.5 10362.5 187727.5 ;
      RECT  10657.5 188522.5 10722.5 188657.5 ;
      RECT  10657.5 187547.5 10722.5 187682.5 ;
      RECT  10492.5 187822.5 10357.5 187887.5 ;
      RECT  10235.0 188037.5 10100.0 188102.5 ;
      RECT  10297.5 188432.5 10362.5 188567.5 ;
      RECT  10487.5 187592.5 10552.5 187727.5 ;
      RECT  10587.5 188037.5 10452.5 188102.5 ;
      RECT  10100.0 188037.5 10235.0 188102.5 ;
      RECT  10357.5 187822.5 10492.5 187887.5 ;
      RECT  10452.5 188037.5 10587.5 188102.5 ;
      RECT  10040.0 188742.5 10960.0 188807.5 ;
      RECT  10040.0 187397.5 10960.0 187462.5 ;
      RECT  11387.5 188590.0 11452.5 188775.0 ;
      RECT  11387.5 187430.0 11452.5 187615.0 ;
      RECT  11027.5 187547.5 11092.5 187397.5 ;
      RECT  11027.5 188432.5 11092.5 188807.5 ;
      RECT  11217.5 187547.5 11282.5 188432.5 ;
      RECT  11027.5 188432.5 11092.5 188567.5 ;
      RECT  11217.5 188432.5 11282.5 188567.5 ;
      RECT  11217.5 188432.5 11282.5 188567.5 ;
      RECT  11027.5 188432.5 11092.5 188567.5 ;
      RECT  11027.5 187547.5 11092.5 187682.5 ;
      RECT  11217.5 187547.5 11282.5 187682.5 ;
      RECT  11217.5 187547.5 11282.5 187682.5 ;
      RECT  11027.5 187547.5 11092.5 187682.5 ;
      RECT  11387.5 188522.5 11452.5 188657.5 ;
      RECT  11387.5 187547.5 11452.5 187682.5 ;
      RECT  11085.0 187990.0 11150.0 188125.0 ;
      RECT  11085.0 187990.0 11150.0 188125.0 ;
      RECT  11250.0 188025.0 11315.0 188090.0 ;
      RECT  10960.0 188742.5 11520.0 188807.5 ;
      RECT  10960.0 187397.5 11520.0 187462.5 ;
      RECT  9222.5 187990.0 9287.5 188125.0 ;
      RECT  9362.5 187717.5 9427.5 187852.5 ;
      RECT  10357.5 187822.5 10222.5 187887.5 ;
      RECT  9907.5 188960.0 9972.5 188775.0 ;
      RECT  9907.5 190120.0 9972.5 189935.0 ;
      RECT  9547.5 190002.5 9612.5 190152.5 ;
      RECT  9547.5 189117.5 9612.5 188742.5 ;
      RECT  9737.5 190002.5 9802.5 189117.5 ;
      RECT  9547.5 189117.5 9612.5 188982.5 ;
      RECT  9737.5 189117.5 9802.5 188982.5 ;
      RECT  9737.5 189117.5 9802.5 188982.5 ;
      RECT  9547.5 189117.5 9612.5 188982.5 ;
      RECT  9547.5 190002.5 9612.5 189867.5 ;
      RECT  9737.5 190002.5 9802.5 189867.5 ;
      RECT  9737.5 190002.5 9802.5 189867.5 ;
      RECT  9547.5 190002.5 9612.5 189867.5 ;
      RECT  9907.5 189027.5 9972.5 188892.5 ;
      RECT  9907.5 190002.5 9972.5 189867.5 ;
      RECT  9605.0 189560.0 9670.0 189425.0 ;
      RECT  9605.0 189560.0 9670.0 189425.0 ;
      RECT  9770.0 189525.0 9835.0 189460.0 ;
      RECT  9480.0 188807.5 10040.0 188742.5 ;
      RECT  9480.0 190152.5 10040.0 190087.5 ;
      RECT  10107.5 189957.5 10172.5 190152.5 ;
      RECT  10107.5 189117.5 10172.5 188742.5 ;
      RECT  10487.5 189117.5 10552.5 188742.5 ;
      RECT  10657.5 188960.0 10722.5 188775.0 ;
      RECT  10657.5 190120.0 10722.5 189935.0 ;
      RECT  10107.5 189117.5 10172.5 188982.5 ;
      RECT  10297.5 189117.5 10362.5 188982.5 ;
      RECT  10297.5 189117.5 10362.5 188982.5 ;
      RECT  10107.5 189117.5 10172.5 188982.5 ;
      RECT  10297.5 189117.5 10362.5 188982.5 ;
      RECT  10487.5 189117.5 10552.5 188982.5 ;
      RECT  10487.5 189117.5 10552.5 188982.5 ;
      RECT  10297.5 189117.5 10362.5 188982.5 ;
      RECT  10107.5 189957.5 10172.5 189822.5 ;
      RECT  10297.5 189957.5 10362.5 189822.5 ;
      RECT  10297.5 189957.5 10362.5 189822.5 ;
      RECT  10107.5 189957.5 10172.5 189822.5 ;
      RECT  10297.5 189957.5 10362.5 189822.5 ;
      RECT  10487.5 189957.5 10552.5 189822.5 ;
      RECT  10487.5 189957.5 10552.5 189822.5 ;
      RECT  10297.5 189957.5 10362.5 189822.5 ;
      RECT  10657.5 189027.5 10722.5 188892.5 ;
      RECT  10657.5 190002.5 10722.5 189867.5 ;
      RECT  10492.5 189727.5 10357.5 189662.5 ;
      RECT  10235.0 189512.5 10100.0 189447.5 ;
      RECT  10297.5 189117.5 10362.5 188982.5 ;
      RECT  10487.5 189957.5 10552.5 189822.5 ;
      RECT  10587.5 189512.5 10452.5 189447.5 ;
      RECT  10100.0 189512.5 10235.0 189447.5 ;
      RECT  10357.5 189727.5 10492.5 189662.5 ;
      RECT  10452.5 189512.5 10587.5 189447.5 ;
      RECT  10040.0 188807.5 10960.0 188742.5 ;
      RECT  10040.0 190152.5 10960.0 190087.5 ;
      RECT  11387.5 188960.0 11452.5 188775.0 ;
      RECT  11387.5 190120.0 11452.5 189935.0 ;
      RECT  11027.5 190002.5 11092.5 190152.5 ;
      RECT  11027.5 189117.5 11092.5 188742.5 ;
      RECT  11217.5 190002.5 11282.5 189117.5 ;
      RECT  11027.5 189117.5 11092.5 188982.5 ;
      RECT  11217.5 189117.5 11282.5 188982.5 ;
      RECT  11217.5 189117.5 11282.5 188982.5 ;
      RECT  11027.5 189117.5 11092.5 188982.5 ;
      RECT  11027.5 190002.5 11092.5 189867.5 ;
      RECT  11217.5 190002.5 11282.5 189867.5 ;
      RECT  11217.5 190002.5 11282.5 189867.5 ;
      RECT  11027.5 190002.5 11092.5 189867.5 ;
      RECT  11387.5 189027.5 11452.5 188892.5 ;
      RECT  11387.5 190002.5 11452.5 189867.5 ;
      RECT  11085.0 189560.0 11150.0 189425.0 ;
      RECT  11085.0 189560.0 11150.0 189425.0 ;
      RECT  11250.0 189525.0 11315.0 189460.0 ;
      RECT  10960.0 188807.5 11520.0 188742.5 ;
      RECT  10960.0 190152.5 11520.0 190087.5 ;
      RECT  9222.5 189425.0 9287.5 189560.0 ;
      RECT  9362.5 189697.5 9427.5 189832.5 ;
      RECT  10357.5 189662.5 10222.5 189727.5 ;
      RECT  9907.5 191280.0 9972.5 191465.0 ;
      RECT  9907.5 190120.0 9972.5 190305.0 ;
      RECT  9547.5 190237.5 9612.5 190087.5 ;
      RECT  9547.5 191122.5 9612.5 191497.5 ;
      RECT  9737.5 190237.5 9802.5 191122.5 ;
      RECT  9547.5 191122.5 9612.5 191257.5 ;
      RECT  9737.5 191122.5 9802.5 191257.5 ;
      RECT  9737.5 191122.5 9802.5 191257.5 ;
      RECT  9547.5 191122.5 9612.5 191257.5 ;
      RECT  9547.5 190237.5 9612.5 190372.5 ;
      RECT  9737.5 190237.5 9802.5 190372.5 ;
      RECT  9737.5 190237.5 9802.5 190372.5 ;
      RECT  9547.5 190237.5 9612.5 190372.5 ;
      RECT  9907.5 191212.5 9972.5 191347.5 ;
      RECT  9907.5 190237.5 9972.5 190372.5 ;
      RECT  9605.0 190680.0 9670.0 190815.0 ;
      RECT  9605.0 190680.0 9670.0 190815.0 ;
      RECT  9770.0 190715.0 9835.0 190780.0 ;
      RECT  9480.0 191432.5 10040.0 191497.5 ;
      RECT  9480.0 190087.5 10040.0 190152.5 ;
      RECT  10107.5 190282.5 10172.5 190087.5 ;
      RECT  10107.5 191122.5 10172.5 191497.5 ;
      RECT  10487.5 191122.5 10552.5 191497.5 ;
      RECT  10657.5 191280.0 10722.5 191465.0 ;
      RECT  10657.5 190120.0 10722.5 190305.0 ;
      RECT  10107.5 191122.5 10172.5 191257.5 ;
      RECT  10297.5 191122.5 10362.5 191257.5 ;
      RECT  10297.5 191122.5 10362.5 191257.5 ;
      RECT  10107.5 191122.5 10172.5 191257.5 ;
      RECT  10297.5 191122.5 10362.5 191257.5 ;
      RECT  10487.5 191122.5 10552.5 191257.5 ;
      RECT  10487.5 191122.5 10552.5 191257.5 ;
      RECT  10297.5 191122.5 10362.5 191257.5 ;
      RECT  10107.5 190282.5 10172.5 190417.5 ;
      RECT  10297.5 190282.5 10362.5 190417.5 ;
      RECT  10297.5 190282.5 10362.5 190417.5 ;
      RECT  10107.5 190282.5 10172.5 190417.5 ;
      RECT  10297.5 190282.5 10362.5 190417.5 ;
      RECT  10487.5 190282.5 10552.5 190417.5 ;
      RECT  10487.5 190282.5 10552.5 190417.5 ;
      RECT  10297.5 190282.5 10362.5 190417.5 ;
      RECT  10657.5 191212.5 10722.5 191347.5 ;
      RECT  10657.5 190237.5 10722.5 190372.5 ;
      RECT  10492.5 190512.5 10357.5 190577.5 ;
      RECT  10235.0 190727.5 10100.0 190792.5 ;
      RECT  10297.5 191122.5 10362.5 191257.5 ;
      RECT  10487.5 190282.5 10552.5 190417.5 ;
      RECT  10587.5 190727.5 10452.5 190792.5 ;
      RECT  10100.0 190727.5 10235.0 190792.5 ;
      RECT  10357.5 190512.5 10492.5 190577.5 ;
      RECT  10452.5 190727.5 10587.5 190792.5 ;
      RECT  10040.0 191432.5 10960.0 191497.5 ;
      RECT  10040.0 190087.5 10960.0 190152.5 ;
      RECT  11387.5 191280.0 11452.5 191465.0 ;
      RECT  11387.5 190120.0 11452.5 190305.0 ;
      RECT  11027.5 190237.5 11092.5 190087.5 ;
      RECT  11027.5 191122.5 11092.5 191497.5 ;
      RECT  11217.5 190237.5 11282.5 191122.5 ;
      RECT  11027.5 191122.5 11092.5 191257.5 ;
      RECT  11217.5 191122.5 11282.5 191257.5 ;
      RECT  11217.5 191122.5 11282.5 191257.5 ;
      RECT  11027.5 191122.5 11092.5 191257.5 ;
      RECT  11027.5 190237.5 11092.5 190372.5 ;
      RECT  11217.5 190237.5 11282.5 190372.5 ;
      RECT  11217.5 190237.5 11282.5 190372.5 ;
      RECT  11027.5 190237.5 11092.5 190372.5 ;
      RECT  11387.5 191212.5 11452.5 191347.5 ;
      RECT  11387.5 190237.5 11452.5 190372.5 ;
      RECT  11085.0 190680.0 11150.0 190815.0 ;
      RECT  11085.0 190680.0 11150.0 190815.0 ;
      RECT  11250.0 190715.0 11315.0 190780.0 ;
      RECT  10960.0 191432.5 11520.0 191497.5 ;
      RECT  10960.0 190087.5 11520.0 190152.5 ;
      RECT  9222.5 190680.0 9287.5 190815.0 ;
      RECT  9362.5 190407.5 9427.5 190542.5 ;
      RECT  10357.5 190512.5 10222.5 190577.5 ;
      RECT  9907.5 191650.0 9972.5 191465.0 ;
      RECT  9907.5 192810.0 9972.5 192625.0 ;
      RECT  9547.5 192692.5 9612.5 192842.5 ;
      RECT  9547.5 191807.5 9612.5 191432.5 ;
      RECT  9737.5 192692.5 9802.5 191807.5 ;
      RECT  9547.5 191807.5 9612.5 191672.5 ;
      RECT  9737.5 191807.5 9802.5 191672.5 ;
      RECT  9737.5 191807.5 9802.5 191672.5 ;
      RECT  9547.5 191807.5 9612.5 191672.5 ;
      RECT  9547.5 192692.5 9612.5 192557.5 ;
      RECT  9737.5 192692.5 9802.5 192557.5 ;
      RECT  9737.5 192692.5 9802.5 192557.5 ;
      RECT  9547.5 192692.5 9612.5 192557.5 ;
      RECT  9907.5 191717.5 9972.5 191582.5 ;
      RECT  9907.5 192692.5 9972.5 192557.5 ;
      RECT  9605.0 192250.0 9670.0 192115.0 ;
      RECT  9605.0 192250.0 9670.0 192115.0 ;
      RECT  9770.0 192215.0 9835.0 192150.0 ;
      RECT  9480.0 191497.5 10040.0 191432.5 ;
      RECT  9480.0 192842.5 10040.0 192777.5 ;
      RECT  10107.5 192647.5 10172.5 192842.5 ;
      RECT  10107.5 191807.5 10172.5 191432.5 ;
      RECT  10487.5 191807.5 10552.5 191432.5 ;
      RECT  10657.5 191650.0 10722.5 191465.0 ;
      RECT  10657.5 192810.0 10722.5 192625.0 ;
      RECT  10107.5 191807.5 10172.5 191672.5 ;
      RECT  10297.5 191807.5 10362.5 191672.5 ;
      RECT  10297.5 191807.5 10362.5 191672.5 ;
      RECT  10107.5 191807.5 10172.5 191672.5 ;
      RECT  10297.5 191807.5 10362.5 191672.5 ;
      RECT  10487.5 191807.5 10552.5 191672.5 ;
      RECT  10487.5 191807.5 10552.5 191672.5 ;
      RECT  10297.5 191807.5 10362.5 191672.5 ;
      RECT  10107.5 192647.5 10172.5 192512.5 ;
      RECT  10297.5 192647.5 10362.5 192512.5 ;
      RECT  10297.5 192647.5 10362.5 192512.5 ;
      RECT  10107.5 192647.5 10172.5 192512.5 ;
      RECT  10297.5 192647.5 10362.5 192512.5 ;
      RECT  10487.5 192647.5 10552.5 192512.5 ;
      RECT  10487.5 192647.5 10552.5 192512.5 ;
      RECT  10297.5 192647.5 10362.5 192512.5 ;
      RECT  10657.5 191717.5 10722.5 191582.5 ;
      RECT  10657.5 192692.5 10722.5 192557.5 ;
      RECT  10492.5 192417.5 10357.5 192352.5 ;
      RECT  10235.0 192202.5 10100.0 192137.5 ;
      RECT  10297.5 191807.5 10362.5 191672.5 ;
      RECT  10487.5 192647.5 10552.5 192512.5 ;
      RECT  10587.5 192202.5 10452.5 192137.5 ;
      RECT  10100.0 192202.5 10235.0 192137.5 ;
      RECT  10357.5 192417.5 10492.5 192352.5 ;
      RECT  10452.5 192202.5 10587.5 192137.5 ;
      RECT  10040.0 191497.5 10960.0 191432.5 ;
      RECT  10040.0 192842.5 10960.0 192777.5 ;
      RECT  11387.5 191650.0 11452.5 191465.0 ;
      RECT  11387.5 192810.0 11452.5 192625.0 ;
      RECT  11027.5 192692.5 11092.5 192842.5 ;
      RECT  11027.5 191807.5 11092.5 191432.5 ;
      RECT  11217.5 192692.5 11282.5 191807.5 ;
      RECT  11027.5 191807.5 11092.5 191672.5 ;
      RECT  11217.5 191807.5 11282.5 191672.5 ;
      RECT  11217.5 191807.5 11282.5 191672.5 ;
      RECT  11027.5 191807.5 11092.5 191672.5 ;
      RECT  11027.5 192692.5 11092.5 192557.5 ;
      RECT  11217.5 192692.5 11282.5 192557.5 ;
      RECT  11217.5 192692.5 11282.5 192557.5 ;
      RECT  11027.5 192692.5 11092.5 192557.5 ;
      RECT  11387.5 191717.5 11452.5 191582.5 ;
      RECT  11387.5 192692.5 11452.5 192557.5 ;
      RECT  11085.0 192250.0 11150.0 192115.0 ;
      RECT  11085.0 192250.0 11150.0 192115.0 ;
      RECT  11250.0 192215.0 11315.0 192150.0 ;
      RECT  10960.0 191497.5 11520.0 191432.5 ;
      RECT  10960.0 192842.5 11520.0 192777.5 ;
      RECT  9222.5 192115.0 9287.5 192250.0 ;
      RECT  9362.5 192387.5 9427.5 192522.5 ;
      RECT  10357.5 192352.5 10222.5 192417.5 ;
      RECT  9907.5 193970.0 9972.5 194155.0 ;
      RECT  9907.5 192810.0 9972.5 192995.0 ;
      RECT  9547.5 192927.5 9612.5 192777.5 ;
      RECT  9547.5 193812.5 9612.5 194187.5 ;
      RECT  9737.5 192927.5 9802.5 193812.5 ;
      RECT  9547.5 193812.5 9612.5 193947.5 ;
      RECT  9737.5 193812.5 9802.5 193947.5 ;
      RECT  9737.5 193812.5 9802.5 193947.5 ;
      RECT  9547.5 193812.5 9612.5 193947.5 ;
      RECT  9547.5 192927.5 9612.5 193062.5 ;
      RECT  9737.5 192927.5 9802.5 193062.5 ;
      RECT  9737.5 192927.5 9802.5 193062.5 ;
      RECT  9547.5 192927.5 9612.5 193062.5 ;
      RECT  9907.5 193902.5 9972.5 194037.5 ;
      RECT  9907.5 192927.5 9972.5 193062.5 ;
      RECT  9605.0 193370.0 9670.0 193505.0 ;
      RECT  9605.0 193370.0 9670.0 193505.0 ;
      RECT  9770.0 193405.0 9835.0 193470.0 ;
      RECT  9480.0 194122.5 10040.0 194187.5 ;
      RECT  9480.0 192777.5 10040.0 192842.5 ;
      RECT  10107.5 192972.5 10172.5 192777.5 ;
      RECT  10107.5 193812.5 10172.5 194187.5 ;
      RECT  10487.5 193812.5 10552.5 194187.5 ;
      RECT  10657.5 193970.0 10722.5 194155.0 ;
      RECT  10657.5 192810.0 10722.5 192995.0 ;
      RECT  10107.5 193812.5 10172.5 193947.5 ;
      RECT  10297.5 193812.5 10362.5 193947.5 ;
      RECT  10297.5 193812.5 10362.5 193947.5 ;
      RECT  10107.5 193812.5 10172.5 193947.5 ;
      RECT  10297.5 193812.5 10362.5 193947.5 ;
      RECT  10487.5 193812.5 10552.5 193947.5 ;
      RECT  10487.5 193812.5 10552.5 193947.5 ;
      RECT  10297.5 193812.5 10362.5 193947.5 ;
      RECT  10107.5 192972.5 10172.5 193107.5 ;
      RECT  10297.5 192972.5 10362.5 193107.5 ;
      RECT  10297.5 192972.5 10362.5 193107.5 ;
      RECT  10107.5 192972.5 10172.5 193107.5 ;
      RECT  10297.5 192972.5 10362.5 193107.5 ;
      RECT  10487.5 192972.5 10552.5 193107.5 ;
      RECT  10487.5 192972.5 10552.5 193107.5 ;
      RECT  10297.5 192972.5 10362.5 193107.5 ;
      RECT  10657.5 193902.5 10722.5 194037.5 ;
      RECT  10657.5 192927.5 10722.5 193062.5 ;
      RECT  10492.5 193202.5 10357.5 193267.5 ;
      RECT  10235.0 193417.5 10100.0 193482.5 ;
      RECT  10297.5 193812.5 10362.5 193947.5 ;
      RECT  10487.5 192972.5 10552.5 193107.5 ;
      RECT  10587.5 193417.5 10452.5 193482.5 ;
      RECT  10100.0 193417.5 10235.0 193482.5 ;
      RECT  10357.5 193202.5 10492.5 193267.5 ;
      RECT  10452.5 193417.5 10587.5 193482.5 ;
      RECT  10040.0 194122.5 10960.0 194187.5 ;
      RECT  10040.0 192777.5 10960.0 192842.5 ;
      RECT  11387.5 193970.0 11452.5 194155.0 ;
      RECT  11387.5 192810.0 11452.5 192995.0 ;
      RECT  11027.5 192927.5 11092.5 192777.5 ;
      RECT  11027.5 193812.5 11092.5 194187.5 ;
      RECT  11217.5 192927.5 11282.5 193812.5 ;
      RECT  11027.5 193812.5 11092.5 193947.5 ;
      RECT  11217.5 193812.5 11282.5 193947.5 ;
      RECT  11217.5 193812.5 11282.5 193947.5 ;
      RECT  11027.5 193812.5 11092.5 193947.5 ;
      RECT  11027.5 192927.5 11092.5 193062.5 ;
      RECT  11217.5 192927.5 11282.5 193062.5 ;
      RECT  11217.5 192927.5 11282.5 193062.5 ;
      RECT  11027.5 192927.5 11092.5 193062.5 ;
      RECT  11387.5 193902.5 11452.5 194037.5 ;
      RECT  11387.5 192927.5 11452.5 193062.5 ;
      RECT  11085.0 193370.0 11150.0 193505.0 ;
      RECT  11085.0 193370.0 11150.0 193505.0 ;
      RECT  11250.0 193405.0 11315.0 193470.0 ;
      RECT  10960.0 194122.5 11520.0 194187.5 ;
      RECT  10960.0 192777.5 11520.0 192842.5 ;
      RECT  9222.5 193370.0 9287.5 193505.0 ;
      RECT  9362.5 193097.5 9427.5 193232.5 ;
      RECT  10357.5 193202.5 10222.5 193267.5 ;
      RECT  9907.5 194340.0 9972.5 194155.0 ;
      RECT  9907.5 195500.0 9972.5 195315.0 ;
      RECT  9547.5 195382.5 9612.5 195532.5 ;
      RECT  9547.5 194497.5 9612.5 194122.5 ;
      RECT  9737.5 195382.5 9802.5 194497.5 ;
      RECT  9547.5 194497.5 9612.5 194362.5 ;
      RECT  9737.5 194497.5 9802.5 194362.5 ;
      RECT  9737.5 194497.5 9802.5 194362.5 ;
      RECT  9547.5 194497.5 9612.5 194362.5 ;
      RECT  9547.5 195382.5 9612.5 195247.5 ;
      RECT  9737.5 195382.5 9802.5 195247.5 ;
      RECT  9737.5 195382.5 9802.5 195247.5 ;
      RECT  9547.5 195382.5 9612.5 195247.5 ;
      RECT  9907.5 194407.5 9972.5 194272.5 ;
      RECT  9907.5 195382.5 9972.5 195247.5 ;
      RECT  9605.0 194940.0 9670.0 194805.0 ;
      RECT  9605.0 194940.0 9670.0 194805.0 ;
      RECT  9770.0 194905.0 9835.0 194840.0 ;
      RECT  9480.0 194187.5 10040.0 194122.5 ;
      RECT  9480.0 195532.5 10040.0 195467.5 ;
      RECT  10107.5 195337.5 10172.5 195532.5 ;
      RECT  10107.5 194497.5 10172.5 194122.5 ;
      RECT  10487.5 194497.5 10552.5 194122.5 ;
      RECT  10657.5 194340.0 10722.5 194155.0 ;
      RECT  10657.5 195500.0 10722.5 195315.0 ;
      RECT  10107.5 194497.5 10172.5 194362.5 ;
      RECT  10297.5 194497.5 10362.5 194362.5 ;
      RECT  10297.5 194497.5 10362.5 194362.5 ;
      RECT  10107.5 194497.5 10172.5 194362.5 ;
      RECT  10297.5 194497.5 10362.5 194362.5 ;
      RECT  10487.5 194497.5 10552.5 194362.5 ;
      RECT  10487.5 194497.5 10552.5 194362.5 ;
      RECT  10297.5 194497.5 10362.5 194362.5 ;
      RECT  10107.5 195337.5 10172.5 195202.5 ;
      RECT  10297.5 195337.5 10362.5 195202.5 ;
      RECT  10297.5 195337.5 10362.5 195202.5 ;
      RECT  10107.5 195337.5 10172.5 195202.5 ;
      RECT  10297.5 195337.5 10362.5 195202.5 ;
      RECT  10487.5 195337.5 10552.5 195202.5 ;
      RECT  10487.5 195337.5 10552.5 195202.5 ;
      RECT  10297.5 195337.5 10362.5 195202.5 ;
      RECT  10657.5 194407.5 10722.5 194272.5 ;
      RECT  10657.5 195382.5 10722.5 195247.5 ;
      RECT  10492.5 195107.5 10357.5 195042.5 ;
      RECT  10235.0 194892.5 10100.0 194827.5 ;
      RECT  10297.5 194497.5 10362.5 194362.5 ;
      RECT  10487.5 195337.5 10552.5 195202.5 ;
      RECT  10587.5 194892.5 10452.5 194827.5 ;
      RECT  10100.0 194892.5 10235.0 194827.5 ;
      RECT  10357.5 195107.5 10492.5 195042.5 ;
      RECT  10452.5 194892.5 10587.5 194827.5 ;
      RECT  10040.0 194187.5 10960.0 194122.5 ;
      RECT  10040.0 195532.5 10960.0 195467.5 ;
      RECT  11387.5 194340.0 11452.5 194155.0 ;
      RECT  11387.5 195500.0 11452.5 195315.0 ;
      RECT  11027.5 195382.5 11092.5 195532.5 ;
      RECT  11027.5 194497.5 11092.5 194122.5 ;
      RECT  11217.5 195382.5 11282.5 194497.5 ;
      RECT  11027.5 194497.5 11092.5 194362.5 ;
      RECT  11217.5 194497.5 11282.5 194362.5 ;
      RECT  11217.5 194497.5 11282.5 194362.5 ;
      RECT  11027.5 194497.5 11092.5 194362.5 ;
      RECT  11027.5 195382.5 11092.5 195247.5 ;
      RECT  11217.5 195382.5 11282.5 195247.5 ;
      RECT  11217.5 195382.5 11282.5 195247.5 ;
      RECT  11027.5 195382.5 11092.5 195247.5 ;
      RECT  11387.5 194407.5 11452.5 194272.5 ;
      RECT  11387.5 195382.5 11452.5 195247.5 ;
      RECT  11085.0 194940.0 11150.0 194805.0 ;
      RECT  11085.0 194940.0 11150.0 194805.0 ;
      RECT  11250.0 194905.0 11315.0 194840.0 ;
      RECT  10960.0 194187.5 11520.0 194122.5 ;
      RECT  10960.0 195532.5 11520.0 195467.5 ;
      RECT  9222.5 194805.0 9287.5 194940.0 ;
      RECT  9362.5 195077.5 9427.5 195212.5 ;
      RECT  10357.5 195042.5 10222.5 195107.5 ;
      RECT  9907.5 196660.0 9972.5 196845.0 ;
      RECT  9907.5 195500.0 9972.5 195685.0 ;
      RECT  9547.5 195617.5 9612.5 195467.5 ;
      RECT  9547.5 196502.5 9612.5 196877.5 ;
      RECT  9737.5 195617.5 9802.5 196502.5 ;
      RECT  9547.5 196502.5 9612.5 196637.5 ;
      RECT  9737.5 196502.5 9802.5 196637.5 ;
      RECT  9737.5 196502.5 9802.5 196637.5 ;
      RECT  9547.5 196502.5 9612.5 196637.5 ;
      RECT  9547.5 195617.5 9612.5 195752.5 ;
      RECT  9737.5 195617.5 9802.5 195752.5 ;
      RECT  9737.5 195617.5 9802.5 195752.5 ;
      RECT  9547.5 195617.5 9612.5 195752.5 ;
      RECT  9907.5 196592.5 9972.5 196727.5 ;
      RECT  9907.5 195617.5 9972.5 195752.5 ;
      RECT  9605.0 196060.0 9670.0 196195.0 ;
      RECT  9605.0 196060.0 9670.0 196195.0 ;
      RECT  9770.0 196095.0 9835.0 196160.0 ;
      RECT  9480.0 196812.5 10040.0 196877.5 ;
      RECT  9480.0 195467.5 10040.0 195532.5 ;
      RECT  10107.5 195662.5 10172.5 195467.5 ;
      RECT  10107.5 196502.5 10172.5 196877.5 ;
      RECT  10487.5 196502.5 10552.5 196877.5 ;
      RECT  10657.5 196660.0 10722.5 196845.0 ;
      RECT  10657.5 195500.0 10722.5 195685.0 ;
      RECT  10107.5 196502.5 10172.5 196637.5 ;
      RECT  10297.5 196502.5 10362.5 196637.5 ;
      RECT  10297.5 196502.5 10362.5 196637.5 ;
      RECT  10107.5 196502.5 10172.5 196637.5 ;
      RECT  10297.5 196502.5 10362.5 196637.5 ;
      RECT  10487.5 196502.5 10552.5 196637.5 ;
      RECT  10487.5 196502.5 10552.5 196637.5 ;
      RECT  10297.5 196502.5 10362.5 196637.5 ;
      RECT  10107.5 195662.5 10172.5 195797.5 ;
      RECT  10297.5 195662.5 10362.5 195797.5 ;
      RECT  10297.5 195662.5 10362.5 195797.5 ;
      RECT  10107.5 195662.5 10172.5 195797.5 ;
      RECT  10297.5 195662.5 10362.5 195797.5 ;
      RECT  10487.5 195662.5 10552.5 195797.5 ;
      RECT  10487.5 195662.5 10552.5 195797.5 ;
      RECT  10297.5 195662.5 10362.5 195797.5 ;
      RECT  10657.5 196592.5 10722.5 196727.5 ;
      RECT  10657.5 195617.5 10722.5 195752.5 ;
      RECT  10492.5 195892.5 10357.5 195957.5 ;
      RECT  10235.0 196107.5 10100.0 196172.5 ;
      RECT  10297.5 196502.5 10362.5 196637.5 ;
      RECT  10487.5 195662.5 10552.5 195797.5 ;
      RECT  10587.5 196107.5 10452.5 196172.5 ;
      RECT  10100.0 196107.5 10235.0 196172.5 ;
      RECT  10357.5 195892.5 10492.5 195957.5 ;
      RECT  10452.5 196107.5 10587.5 196172.5 ;
      RECT  10040.0 196812.5 10960.0 196877.5 ;
      RECT  10040.0 195467.5 10960.0 195532.5 ;
      RECT  11387.5 196660.0 11452.5 196845.0 ;
      RECT  11387.5 195500.0 11452.5 195685.0 ;
      RECT  11027.5 195617.5 11092.5 195467.5 ;
      RECT  11027.5 196502.5 11092.5 196877.5 ;
      RECT  11217.5 195617.5 11282.5 196502.5 ;
      RECT  11027.5 196502.5 11092.5 196637.5 ;
      RECT  11217.5 196502.5 11282.5 196637.5 ;
      RECT  11217.5 196502.5 11282.5 196637.5 ;
      RECT  11027.5 196502.5 11092.5 196637.5 ;
      RECT  11027.5 195617.5 11092.5 195752.5 ;
      RECT  11217.5 195617.5 11282.5 195752.5 ;
      RECT  11217.5 195617.5 11282.5 195752.5 ;
      RECT  11027.5 195617.5 11092.5 195752.5 ;
      RECT  11387.5 196592.5 11452.5 196727.5 ;
      RECT  11387.5 195617.5 11452.5 195752.5 ;
      RECT  11085.0 196060.0 11150.0 196195.0 ;
      RECT  11085.0 196060.0 11150.0 196195.0 ;
      RECT  11250.0 196095.0 11315.0 196160.0 ;
      RECT  10960.0 196812.5 11520.0 196877.5 ;
      RECT  10960.0 195467.5 11520.0 195532.5 ;
      RECT  9222.5 196060.0 9287.5 196195.0 ;
      RECT  9362.5 195787.5 9427.5 195922.5 ;
      RECT  10357.5 195892.5 10222.5 195957.5 ;
      RECT  9907.5 197030.0 9972.5 196845.0 ;
      RECT  9907.5 198190.0 9972.5 198005.0 ;
      RECT  9547.5 198072.5 9612.5 198222.5 ;
      RECT  9547.5 197187.5 9612.5 196812.5 ;
      RECT  9737.5 198072.5 9802.5 197187.5 ;
      RECT  9547.5 197187.5 9612.5 197052.5 ;
      RECT  9737.5 197187.5 9802.5 197052.5 ;
      RECT  9737.5 197187.5 9802.5 197052.5 ;
      RECT  9547.5 197187.5 9612.5 197052.5 ;
      RECT  9547.5 198072.5 9612.5 197937.5 ;
      RECT  9737.5 198072.5 9802.5 197937.5 ;
      RECT  9737.5 198072.5 9802.5 197937.5 ;
      RECT  9547.5 198072.5 9612.5 197937.5 ;
      RECT  9907.5 197097.5 9972.5 196962.5 ;
      RECT  9907.5 198072.5 9972.5 197937.5 ;
      RECT  9605.0 197630.0 9670.0 197495.0 ;
      RECT  9605.0 197630.0 9670.0 197495.0 ;
      RECT  9770.0 197595.0 9835.0 197530.0 ;
      RECT  9480.0 196877.5 10040.0 196812.5 ;
      RECT  9480.0 198222.5 10040.0 198157.5 ;
      RECT  10107.5 198027.5 10172.5 198222.5 ;
      RECT  10107.5 197187.5 10172.5 196812.5 ;
      RECT  10487.5 197187.5 10552.5 196812.5 ;
      RECT  10657.5 197030.0 10722.5 196845.0 ;
      RECT  10657.5 198190.0 10722.5 198005.0 ;
      RECT  10107.5 197187.5 10172.5 197052.5 ;
      RECT  10297.5 197187.5 10362.5 197052.5 ;
      RECT  10297.5 197187.5 10362.5 197052.5 ;
      RECT  10107.5 197187.5 10172.5 197052.5 ;
      RECT  10297.5 197187.5 10362.5 197052.5 ;
      RECT  10487.5 197187.5 10552.5 197052.5 ;
      RECT  10487.5 197187.5 10552.5 197052.5 ;
      RECT  10297.5 197187.5 10362.5 197052.5 ;
      RECT  10107.5 198027.5 10172.5 197892.5 ;
      RECT  10297.5 198027.5 10362.5 197892.5 ;
      RECT  10297.5 198027.5 10362.5 197892.5 ;
      RECT  10107.5 198027.5 10172.5 197892.5 ;
      RECT  10297.5 198027.5 10362.5 197892.5 ;
      RECT  10487.5 198027.5 10552.5 197892.5 ;
      RECT  10487.5 198027.5 10552.5 197892.5 ;
      RECT  10297.5 198027.5 10362.5 197892.5 ;
      RECT  10657.5 197097.5 10722.5 196962.5 ;
      RECT  10657.5 198072.5 10722.5 197937.5 ;
      RECT  10492.5 197797.5 10357.5 197732.5 ;
      RECT  10235.0 197582.5 10100.0 197517.5 ;
      RECT  10297.5 197187.5 10362.5 197052.5 ;
      RECT  10487.5 198027.5 10552.5 197892.5 ;
      RECT  10587.5 197582.5 10452.5 197517.5 ;
      RECT  10100.0 197582.5 10235.0 197517.5 ;
      RECT  10357.5 197797.5 10492.5 197732.5 ;
      RECT  10452.5 197582.5 10587.5 197517.5 ;
      RECT  10040.0 196877.5 10960.0 196812.5 ;
      RECT  10040.0 198222.5 10960.0 198157.5 ;
      RECT  11387.5 197030.0 11452.5 196845.0 ;
      RECT  11387.5 198190.0 11452.5 198005.0 ;
      RECT  11027.5 198072.5 11092.5 198222.5 ;
      RECT  11027.5 197187.5 11092.5 196812.5 ;
      RECT  11217.5 198072.5 11282.5 197187.5 ;
      RECT  11027.5 197187.5 11092.5 197052.5 ;
      RECT  11217.5 197187.5 11282.5 197052.5 ;
      RECT  11217.5 197187.5 11282.5 197052.5 ;
      RECT  11027.5 197187.5 11092.5 197052.5 ;
      RECT  11027.5 198072.5 11092.5 197937.5 ;
      RECT  11217.5 198072.5 11282.5 197937.5 ;
      RECT  11217.5 198072.5 11282.5 197937.5 ;
      RECT  11027.5 198072.5 11092.5 197937.5 ;
      RECT  11387.5 197097.5 11452.5 196962.5 ;
      RECT  11387.5 198072.5 11452.5 197937.5 ;
      RECT  11085.0 197630.0 11150.0 197495.0 ;
      RECT  11085.0 197630.0 11150.0 197495.0 ;
      RECT  11250.0 197595.0 11315.0 197530.0 ;
      RECT  10960.0 196877.5 11520.0 196812.5 ;
      RECT  10960.0 198222.5 11520.0 198157.5 ;
      RECT  9222.5 197495.0 9287.5 197630.0 ;
      RECT  9362.5 197767.5 9427.5 197902.5 ;
      RECT  10357.5 197732.5 10222.5 197797.5 ;
      RECT  9907.5 199350.0 9972.5 199535.0 ;
      RECT  9907.5 198190.0 9972.5 198375.0 ;
      RECT  9547.5 198307.5 9612.5 198157.5 ;
      RECT  9547.5 199192.5 9612.5 199567.5 ;
      RECT  9737.5 198307.5 9802.5 199192.5 ;
      RECT  9547.5 199192.5 9612.5 199327.5 ;
      RECT  9737.5 199192.5 9802.5 199327.5 ;
      RECT  9737.5 199192.5 9802.5 199327.5 ;
      RECT  9547.5 199192.5 9612.5 199327.5 ;
      RECT  9547.5 198307.5 9612.5 198442.5 ;
      RECT  9737.5 198307.5 9802.5 198442.5 ;
      RECT  9737.5 198307.5 9802.5 198442.5 ;
      RECT  9547.5 198307.5 9612.5 198442.5 ;
      RECT  9907.5 199282.5 9972.5 199417.5 ;
      RECT  9907.5 198307.5 9972.5 198442.5 ;
      RECT  9605.0 198750.0 9670.0 198885.0 ;
      RECT  9605.0 198750.0 9670.0 198885.0 ;
      RECT  9770.0 198785.0 9835.0 198850.0 ;
      RECT  9480.0 199502.5 10040.0 199567.5 ;
      RECT  9480.0 198157.5 10040.0 198222.5 ;
      RECT  10107.5 198352.5 10172.5 198157.5 ;
      RECT  10107.5 199192.5 10172.5 199567.5 ;
      RECT  10487.5 199192.5 10552.5 199567.5 ;
      RECT  10657.5 199350.0 10722.5 199535.0 ;
      RECT  10657.5 198190.0 10722.5 198375.0 ;
      RECT  10107.5 199192.5 10172.5 199327.5 ;
      RECT  10297.5 199192.5 10362.5 199327.5 ;
      RECT  10297.5 199192.5 10362.5 199327.5 ;
      RECT  10107.5 199192.5 10172.5 199327.5 ;
      RECT  10297.5 199192.5 10362.5 199327.5 ;
      RECT  10487.5 199192.5 10552.5 199327.5 ;
      RECT  10487.5 199192.5 10552.5 199327.5 ;
      RECT  10297.5 199192.5 10362.5 199327.5 ;
      RECT  10107.5 198352.5 10172.5 198487.5 ;
      RECT  10297.5 198352.5 10362.5 198487.5 ;
      RECT  10297.5 198352.5 10362.5 198487.5 ;
      RECT  10107.5 198352.5 10172.5 198487.5 ;
      RECT  10297.5 198352.5 10362.5 198487.5 ;
      RECT  10487.5 198352.5 10552.5 198487.5 ;
      RECT  10487.5 198352.5 10552.5 198487.5 ;
      RECT  10297.5 198352.5 10362.5 198487.5 ;
      RECT  10657.5 199282.5 10722.5 199417.5 ;
      RECT  10657.5 198307.5 10722.5 198442.5 ;
      RECT  10492.5 198582.5 10357.5 198647.5 ;
      RECT  10235.0 198797.5 10100.0 198862.5 ;
      RECT  10297.5 199192.5 10362.5 199327.5 ;
      RECT  10487.5 198352.5 10552.5 198487.5 ;
      RECT  10587.5 198797.5 10452.5 198862.5 ;
      RECT  10100.0 198797.5 10235.0 198862.5 ;
      RECT  10357.5 198582.5 10492.5 198647.5 ;
      RECT  10452.5 198797.5 10587.5 198862.5 ;
      RECT  10040.0 199502.5 10960.0 199567.5 ;
      RECT  10040.0 198157.5 10960.0 198222.5 ;
      RECT  11387.5 199350.0 11452.5 199535.0 ;
      RECT  11387.5 198190.0 11452.5 198375.0 ;
      RECT  11027.5 198307.5 11092.5 198157.5 ;
      RECT  11027.5 199192.5 11092.5 199567.5 ;
      RECT  11217.5 198307.5 11282.5 199192.5 ;
      RECT  11027.5 199192.5 11092.5 199327.5 ;
      RECT  11217.5 199192.5 11282.5 199327.5 ;
      RECT  11217.5 199192.5 11282.5 199327.5 ;
      RECT  11027.5 199192.5 11092.5 199327.5 ;
      RECT  11027.5 198307.5 11092.5 198442.5 ;
      RECT  11217.5 198307.5 11282.5 198442.5 ;
      RECT  11217.5 198307.5 11282.5 198442.5 ;
      RECT  11027.5 198307.5 11092.5 198442.5 ;
      RECT  11387.5 199282.5 11452.5 199417.5 ;
      RECT  11387.5 198307.5 11452.5 198442.5 ;
      RECT  11085.0 198750.0 11150.0 198885.0 ;
      RECT  11085.0 198750.0 11150.0 198885.0 ;
      RECT  11250.0 198785.0 11315.0 198850.0 ;
      RECT  10960.0 199502.5 11520.0 199567.5 ;
      RECT  10960.0 198157.5 11520.0 198222.5 ;
      RECT  9222.5 198750.0 9287.5 198885.0 ;
      RECT  9362.5 198477.5 9427.5 198612.5 ;
      RECT  10357.5 198582.5 10222.5 198647.5 ;
      RECT  9907.5 199720.0 9972.5 199535.0 ;
      RECT  9907.5 200880.0 9972.5 200695.0 ;
      RECT  9547.5 200762.5 9612.5 200912.5 ;
      RECT  9547.5 199877.5 9612.5 199502.5 ;
      RECT  9737.5 200762.5 9802.5 199877.5 ;
      RECT  9547.5 199877.5 9612.5 199742.5 ;
      RECT  9737.5 199877.5 9802.5 199742.5 ;
      RECT  9737.5 199877.5 9802.5 199742.5 ;
      RECT  9547.5 199877.5 9612.5 199742.5 ;
      RECT  9547.5 200762.5 9612.5 200627.5 ;
      RECT  9737.5 200762.5 9802.5 200627.5 ;
      RECT  9737.5 200762.5 9802.5 200627.5 ;
      RECT  9547.5 200762.5 9612.5 200627.5 ;
      RECT  9907.5 199787.5 9972.5 199652.5 ;
      RECT  9907.5 200762.5 9972.5 200627.5 ;
      RECT  9605.0 200320.0 9670.0 200185.0 ;
      RECT  9605.0 200320.0 9670.0 200185.0 ;
      RECT  9770.0 200285.0 9835.0 200220.0 ;
      RECT  9480.0 199567.5 10040.0 199502.5 ;
      RECT  9480.0 200912.5 10040.0 200847.5 ;
      RECT  10107.5 200717.5 10172.5 200912.5 ;
      RECT  10107.5 199877.5 10172.5 199502.5 ;
      RECT  10487.5 199877.5 10552.5 199502.5 ;
      RECT  10657.5 199720.0 10722.5 199535.0 ;
      RECT  10657.5 200880.0 10722.5 200695.0 ;
      RECT  10107.5 199877.5 10172.5 199742.5 ;
      RECT  10297.5 199877.5 10362.5 199742.5 ;
      RECT  10297.5 199877.5 10362.5 199742.5 ;
      RECT  10107.5 199877.5 10172.5 199742.5 ;
      RECT  10297.5 199877.5 10362.5 199742.5 ;
      RECT  10487.5 199877.5 10552.5 199742.5 ;
      RECT  10487.5 199877.5 10552.5 199742.5 ;
      RECT  10297.5 199877.5 10362.5 199742.5 ;
      RECT  10107.5 200717.5 10172.5 200582.5 ;
      RECT  10297.5 200717.5 10362.5 200582.5 ;
      RECT  10297.5 200717.5 10362.5 200582.5 ;
      RECT  10107.5 200717.5 10172.5 200582.5 ;
      RECT  10297.5 200717.5 10362.5 200582.5 ;
      RECT  10487.5 200717.5 10552.5 200582.5 ;
      RECT  10487.5 200717.5 10552.5 200582.5 ;
      RECT  10297.5 200717.5 10362.5 200582.5 ;
      RECT  10657.5 199787.5 10722.5 199652.5 ;
      RECT  10657.5 200762.5 10722.5 200627.5 ;
      RECT  10492.5 200487.5 10357.5 200422.5 ;
      RECT  10235.0 200272.5 10100.0 200207.5 ;
      RECT  10297.5 199877.5 10362.5 199742.5 ;
      RECT  10487.5 200717.5 10552.5 200582.5 ;
      RECT  10587.5 200272.5 10452.5 200207.5 ;
      RECT  10100.0 200272.5 10235.0 200207.5 ;
      RECT  10357.5 200487.5 10492.5 200422.5 ;
      RECT  10452.5 200272.5 10587.5 200207.5 ;
      RECT  10040.0 199567.5 10960.0 199502.5 ;
      RECT  10040.0 200912.5 10960.0 200847.5 ;
      RECT  11387.5 199720.0 11452.5 199535.0 ;
      RECT  11387.5 200880.0 11452.5 200695.0 ;
      RECT  11027.5 200762.5 11092.5 200912.5 ;
      RECT  11027.5 199877.5 11092.5 199502.5 ;
      RECT  11217.5 200762.5 11282.5 199877.5 ;
      RECT  11027.5 199877.5 11092.5 199742.5 ;
      RECT  11217.5 199877.5 11282.5 199742.5 ;
      RECT  11217.5 199877.5 11282.5 199742.5 ;
      RECT  11027.5 199877.5 11092.5 199742.5 ;
      RECT  11027.5 200762.5 11092.5 200627.5 ;
      RECT  11217.5 200762.5 11282.5 200627.5 ;
      RECT  11217.5 200762.5 11282.5 200627.5 ;
      RECT  11027.5 200762.5 11092.5 200627.5 ;
      RECT  11387.5 199787.5 11452.5 199652.5 ;
      RECT  11387.5 200762.5 11452.5 200627.5 ;
      RECT  11085.0 200320.0 11150.0 200185.0 ;
      RECT  11085.0 200320.0 11150.0 200185.0 ;
      RECT  11250.0 200285.0 11315.0 200220.0 ;
      RECT  10960.0 199567.5 11520.0 199502.5 ;
      RECT  10960.0 200912.5 11520.0 200847.5 ;
      RECT  9222.5 200185.0 9287.5 200320.0 ;
      RECT  9362.5 200457.5 9427.5 200592.5 ;
      RECT  10357.5 200422.5 10222.5 200487.5 ;
      RECT  9907.5 202040.0 9972.5 202225.0 ;
      RECT  9907.5 200880.0 9972.5 201065.0 ;
      RECT  9547.5 200997.5 9612.5 200847.5 ;
      RECT  9547.5 201882.5 9612.5 202257.5 ;
      RECT  9737.5 200997.5 9802.5 201882.5 ;
      RECT  9547.5 201882.5 9612.5 202017.5 ;
      RECT  9737.5 201882.5 9802.5 202017.5 ;
      RECT  9737.5 201882.5 9802.5 202017.5 ;
      RECT  9547.5 201882.5 9612.5 202017.5 ;
      RECT  9547.5 200997.5 9612.5 201132.5 ;
      RECT  9737.5 200997.5 9802.5 201132.5 ;
      RECT  9737.5 200997.5 9802.5 201132.5 ;
      RECT  9547.5 200997.5 9612.5 201132.5 ;
      RECT  9907.5 201972.5 9972.5 202107.5 ;
      RECT  9907.5 200997.5 9972.5 201132.5 ;
      RECT  9605.0 201440.0 9670.0 201575.0 ;
      RECT  9605.0 201440.0 9670.0 201575.0 ;
      RECT  9770.0 201475.0 9835.0 201540.0 ;
      RECT  9480.0 202192.5 10040.0 202257.5 ;
      RECT  9480.0 200847.5 10040.0 200912.5 ;
      RECT  10107.5 201042.5 10172.5 200847.5 ;
      RECT  10107.5 201882.5 10172.5 202257.5 ;
      RECT  10487.5 201882.5 10552.5 202257.5 ;
      RECT  10657.5 202040.0 10722.5 202225.0 ;
      RECT  10657.5 200880.0 10722.5 201065.0 ;
      RECT  10107.5 201882.5 10172.5 202017.5 ;
      RECT  10297.5 201882.5 10362.5 202017.5 ;
      RECT  10297.5 201882.5 10362.5 202017.5 ;
      RECT  10107.5 201882.5 10172.5 202017.5 ;
      RECT  10297.5 201882.5 10362.5 202017.5 ;
      RECT  10487.5 201882.5 10552.5 202017.5 ;
      RECT  10487.5 201882.5 10552.5 202017.5 ;
      RECT  10297.5 201882.5 10362.5 202017.5 ;
      RECT  10107.5 201042.5 10172.5 201177.5 ;
      RECT  10297.5 201042.5 10362.5 201177.5 ;
      RECT  10297.5 201042.5 10362.5 201177.5 ;
      RECT  10107.5 201042.5 10172.5 201177.5 ;
      RECT  10297.5 201042.5 10362.5 201177.5 ;
      RECT  10487.5 201042.5 10552.5 201177.5 ;
      RECT  10487.5 201042.5 10552.5 201177.5 ;
      RECT  10297.5 201042.5 10362.5 201177.5 ;
      RECT  10657.5 201972.5 10722.5 202107.5 ;
      RECT  10657.5 200997.5 10722.5 201132.5 ;
      RECT  10492.5 201272.5 10357.5 201337.5 ;
      RECT  10235.0 201487.5 10100.0 201552.5 ;
      RECT  10297.5 201882.5 10362.5 202017.5 ;
      RECT  10487.5 201042.5 10552.5 201177.5 ;
      RECT  10587.5 201487.5 10452.5 201552.5 ;
      RECT  10100.0 201487.5 10235.0 201552.5 ;
      RECT  10357.5 201272.5 10492.5 201337.5 ;
      RECT  10452.5 201487.5 10587.5 201552.5 ;
      RECT  10040.0 202192.5 10960.0 202257.5 ;
      RECT  10040.0 200847.5 10960.0 200912.5 ;
      RECT  11387.5 202040.0 11452.5 202225.0 ;
      RECT  11387.5 200880.0 11452.5 201065.0 ;
      RECT  11027.5 200997.5 11092.5 200847.5 ;
      RECT  11027.5 201882.5 11092.5 202257.5 ;
      RECT  11217.5 200997.5 11282.5 201882.5 ;
      RECT  11027.5 201882.5 11092.5 202017.5 ;
      RECT  11217.5 201882.5 11282.5 202017.5 ;
      RECT  11217.5 201882.5 11282.5 202017.5 ;
      RECT  11027.5 201882.5 11092.5 202017.5 ;
      RECT  11027.5 200997.5 11092.5 201132.5 ;
      RECT  11217.5 200997.5 11282.5 201132.5 ;
      RECT  11217.5 200997.5 11282.5 201132.5 ;
      RECT  11027.5 200997.5 11092.5 201132.5 ;
      RECT  11387.5 201972.5 11452.5 202107.5 ;
      RECT  11387.5 200997.5 11452.5 201132.5 ;
      RECT  11085.0 201440.0 11150.0 201575.0 ;
      RECT  11085.0 201440.0 11150.0 201575.0 ;
      RECT  11250.0 201475.0 11315.0 201540.0 ;
      RECT  10960.0 202192.5 11520.0 202257.5 ;
      RECT  10960.0 200847.5 11520.0 200912.5 ;
      RECT  9222.5 201440.0 9287.5 201575.0 ;
      RECT  9362.5 201167.5 9427.5 201302.5 ;
      RECT  10357.5 201272.5 10222.5 201337.5 ;
      RECT  9907.5 202410.0 9972.5 202225.0 ;
      RECT  9907.5 203570.0 9972.5 203385.0 ;
      RECT  9547.5 203452.5 9612.5 203602.5 ;
      RECT  9547.5 202567.5 9612.5 202192.5 ;
      RECT  9737.5 203452.5 9802.5 202567.5 ;
      RECT  9547.5 202567.5 9612.5 202432.5 ;
      RECT  9737.5 202567.5 9802.5 202432.5 ;
      RECT  9737.5 202567.5 9802.5 202432.5 ;
      RECT  9547.5 202567.5 9612.5 202432.5 ;
      RECT  9547.5 203452.5 9612.5 203317.5 ;
      RECT  9737.5 203452.5 9802.5 203317.5 ;
      RECT  9737.5 203452.5 9802.5 203317.5 ;
      RECT  9547.5 203452.5 9612.5 203317.5 ;
      RECT  9907.5 202477.5 9972.5 202342.5 ;
      RECT  9907.5 203452.5 9972.5 203317.5 ;
      RECT  9605.0 203010.0 9670.0 202875.0 ;
      RECT  9605.0 203010.0 9670.0 202875.0 ;
      RECT  9770.0 202975.0 9835.0 202910.0 ;
      RECT  9480.0 202257.5 10040.0 202192.5 ;
      RECT  9480.0 203602.5 10040.0 203537.5 ;
      RECT  10107.5 203407.5 10172.5 203602.5 ;
      RECT  10107.5 202567.5 10172.5 202192.5 ;
      RECT  10487.5 202567.5 10552.5 202192.5 ;
      RECT  10657.5 202410.0 10722.5 202225.0 ;
      RECT  10657.5 203570.0 10722.5 203385.0 ;
      RECT  10107.5 202567.5 10172.5 202432.5 ;
      RECT  10297.5 202567.5 10362.5 202432.5 ;
      RECT  10297.5 202567.5 10362.5 202432.5 ;
      RECT  10107.5 202567.5 10172.5 202432.5 ;
      RECT  10297.5 202567.5 10362.5 202432.5 ;
      RECT  10487.5 202567.5 10552.5 202432.5 ;
      RECT  10487.5 202567.5 10552.5 202432.5 ;
      RECT  10297.5 202567.5 10362.5 202432.5 ;
      RECT  10107.5 203407.5 10172.5 203272.5 ;
      RECT  10297.5 203407.5 10362.5 203272.5 ;
      RECT  10297.5 203407.5 10362.5 203272.5 ;
      RECT  10107.5 203407.5 10172.5 203272.5 ;
      RECT  10297.5 203407.5 10362.5 203272.5 ;
      RECT  10487.5 203407.5 10552.5 203272.5 ;
      RECT  10487.5 203407.5 10552.5 203272.5 ;
      RECT  10297.5 203407.5 10362.5 203272.5 ;
      RECT  10657.5 202477.5 10722.5 202342.5 ;
      RECT  10657.5 203452.5 10722.5 203317.5 ;
      RECT  10492.5 203177.5 10357.5 203112.5 ;
      RECT  10235.0 202962.5 10100.0 202897.5 ;
      RECT  10297.5 202567.5 10362.5 202432.5 ;
      RECT  10487.5 203407.5 10552.5 203272.5 ;
      RECT  10587.5 202962.5 10452.5 202897.5 ;
      RECT  10100.0 202962.5 10235.0 202897.5 ;
      RECT  10357.5 203177.5 10492.5 203112.5 ;
      RECT  10452.5 202962.5 10587.5 202897.5 ;
      RECT  10040.0 202257.5 10960.0 202192.5 ;
      RECT  10040.0 203602.5 10960.0 203537.5 ;
      RECT  11387.5 202410.0 11452.5 202225.0 ;
      RECT  11387.5 203570.0 11452.5 203385.0 ;
      RECT  11027.5 203452.5 11092.5 203602.5 ;
      RECT  11027.5 202567.5 11092.5 202192.5 ;
      RECT  11217.5 203452.5 11282.5 202567.5 ;
      RECT  11027.5 202567.5 11092.5 202432.5 ;
      RECT  11217.5 202567.5 11282.5 202432.5 ;
      RECT  11217.5 202567.5 11282.5 202432.5 ;
      RECT  11027.5 202567.5 11092.5 202432.5 ;
      RECT  11027.5 203452.5 11092.5 203317.5 ;
      RECT  11217.5 203452.5 11282.5 203317.5 ;
      RECT  11217.5 203452.5 11282.5 203317.5 ;
      RECT  11027.5 203452.5 11092.5 203317.5 ;
      RECT  11387.5 202477.5 11452.5 202342.5 ;
      RECT  11387.5 203452.5 11452.5 203317.5 ;
      RECT  11085.0 203010.0 11150.0 202875.0 ;
      RECT  11085.0 203010.0 11150.0 202875.0 ;
      RECT  11250.0 202975.0 11315.0 202910.0 ;
      RECT  10960.0 202257.5 11520.0 202192.5 ;
      RECT  10960.0 203602.5 11520.0 203537.5 ;
      RECT  9222.5 202875.0 9287.5 203010.0 ;
      RECT  9362.5 203147.5 9427.5 203282.5 ;
      RECT  10357.5 203112.5 10222.5 203177.5 ;
      RECT  9907.5 204730.0 9972.5 204915.0 ;
      RECT  9907.5 203570.0 9972.5 203755.0 ;
      RECT  9547.5 203687.5 9612.5 203537.5 ;
      RECT  9547.5 204572.5 9612.5 204947.5 ;
      RECT  9737.5 203687.5 9802.5 204572.5 ;
      RECT  9547.5 204572.5 9612.5 204707.5 ;
      RECT  9737.5 204572.5 9802.5 204707.5 ;
      RECT  9737.5 204572.5 9802.5 204707.5 ;
      RECT  9547.5 204572.5 9612.5 204707.5 ;
      RECT  9547.5 203687.5 9612.5 203822.5 ;
      RECT  9737.5 203687.5 9802.5 203822.5 ;
      RECT  9737.5 203687.5 9802.5 203822.5 ;
      RECT  9547.5 203687.5 9612.5 203822.5 ;
      RECT  9907.5 204662.5 9972.5 204797.5 ;
      RECT  9907.5 203687.5 9972.5 203822.5 ;
      RECT  9605.0 204130.0 9670.0 204265.0 ;
      RECT  9605.0 204130.0 9670.0 204265.0 ;
      RECT  9770.0 204165.0 9835.0 204230.0 ;
      RECT  9480.0 204882.5 10040.0 204947.5 ;
      RECT  9480.0 203537.5 10040.0 203602.5 ;
      RECT  10107.5 203732.5 10172.5 203537.5 ;
      RECT  10107.5 204572.5 10172.5 204947.5 ;
      RECT  10487.5 204572.5 10552.5 204947.5 ;
      RECT  10657.5 204730.0 10722.5 204915.0 ;
      RECT  10657.5 203570.0 10722.5 203755.0 ;
      RECT  10107.5 204572.5 10172.5 204707.5 ;
      RECT  10297.5 204572.5 10362.5 204707.5 ;
      RECT  10297.5 204572.5 10362.5 204707.5 ;
      RECT  10107.5 204572.5 10172.5 204707.5 ;
      RECT  10297.5 204572.5 10362.5 204707.5 ;
      RECT  10487.5 204572.5 10552.5 204707.5 ;
      RECT  10487.5 204572.5 10552.5 204707.5 ;
      RECT  10297.5 204572.5 10362.5 204707.5 ;
      RECT  10107.5 203732.5 10172.5 203867.5 ;
      RECT  10297.5 203732.5 10362.5 203867.5 ;
      RECT  10297.5 203732.5 10362.5 203867.5 ;
      RECT  10107.5 203732.5 10172.5 203867.5 ;
      RECT  10297.5 203732.5 10362.5 203867.5 ;
      RECT  10487.5 203732.5 10552.5 203867.5 ;
      RECT  10487.5 203732.5 10552.5 203867.5 ;
      RECT  10297.5 203732.5 10362.5 203867.5 ;
      RECT  10657.5 204662.5 10722.5 204797.5 ;
      RECT  10657.5 203687.5 10722.5 203822.5 ;
      RECT  10492.5 203962.5 10357.5 204027.5 ;
      RECT  10235.0 204177.5 10100.0 204242.5 ;
      RECT  10297.5 204572.5 10362.5 204707.5 ;
      RECT  10487.5 203732.5 10552.5 203867.5 ;
      RECT  10587.5 204177.5 10452.5 204242.5 ;
      RECT  10100.0 204177.5 10235.0 204242.5 ;
      RECT  10357.5 203962.5 10492.5 204027.5 ;
      RECT  10452.5 204177.5 10587.5 204242.5 ;
      RECT  10040.0 204882.5 10960.0 204947.5 ;
      RECT  10040.0 203537.5 10960.0 203602.5 ;
      RECT  11387.5 204730.0 11452.5 204915.0 ;
      RECT  11387.5 203570.0 11452.5 203755.0 ;
      RECT  11027.5 203687.5 11092.5 203537.5 ;
      RECT  11027.5 204572.5 11092.5 204947.5 ;
      RECT  11217.5 203687.5 11282.5 204572.5 ;
      RECT  11027.5 204572.5 11092.5 204707.5 ;
      RECT  11217.5 204572.5 11282.5 204707.5 ;
      RECT  11217.5 204572.5 11282.5 204707.5 ;
      RECT  11027.5 204572.5 11092.5 204707.5 ;
      RECT  11027.5 203687.5 11092.5 203822.5 ;
      RECT  11217.5 203687.5 11282.5 203822.5 ;
      RECT  11217.5 203687.5 11282.5 203822.5 ;
      RECT  11027.5 203687.5 11092.5 203822.5 ;
      RECT  11387.5 204662.5 11452.5 204797.5 ;
      RECT  11387.5 203687.5 11452.5 203822.5 ;
      RECT  11085.0 204130.0 11150.0 204265.0 ;
      RECT  11085.0 204130.0 11150.0 204265.0 ;
      RECT  11250.0 204165.0 11315.0 204230.0 ;
      RECT  10960.0 204882.5 11520.0 204947.5 ;
      RECT  10960.0 203537.5 11520.0 203602.5 ;
      RECT  9222.5 204130.0 9287.5 204265.0 ;
      RECT  9362.5 203857.5 9427.5 203992.5 ;
      RECT  10357.5 203962.5 10222.5 204027.5 ;
      RECT  9907.5 205100.0 9972.5 204915.0 ;
      RECT  9907.5 206260.0 9972.5 206075.0 ;
      RECT  9547.5 206142.5 9612.5 206292.5 ;
      RECT  9547.5 205257.5 9612.5 204882.5 ;
      RECT  9737.5 206142.5 9802.5 205257.5 ;
      RECT  9547.5 205257.5 9612.5 205122.5 ;
      RECT  9737.5 205257.5 9802.5 205122.5 ;
      RECT  9737.5 205257.5 9802.5 205122.5 ;
      RECT  9547.5 205257.5 9612.5 205122.5 ;
      RECT  9547.5 206142.5 9612.5 206007.5 ;
      RECT  9737.5 206142.5 9802.5 206007.5 ;
      RECT  9737.5 206142.5 9802.5 206007.5 ;
      RECT  9547.5 206142.5 9612.5 206007.5 ;
      RECT  9907.5 205167.5 9972.5 205032.5 ;
      RECT  9907.5 206142.5 9972.5 206007.5 ;
      RECT  9605.0 205700.0 9670.0 205565.0 ;
      RECT  9605.0 205700.0 9670.0 205565.0 ;
      RECT  9770.0 205665.0 9835.0 205600.0 ;
      RECT  9480.0 204947.5 10040.0 204882.5 ;
      RECT  9480.0 206292.5 10040.0 206227.5 ;
      RECT  10107.5 206097.5 10172.5 206292.5 ;
      RECT  10107.5 205257.5 10172.5 204882.5 ;
      RECT  10487.5 205257.5 10552.5 204882.5 ;
      RECT  10657.5 205100.0 10722.5 204915.0 ;
      RECT  10657.5 206260.0 10722.5 206075.0 ;
      RECT  10107.5 205257.5 10172.5 205122.5 ;
      RECT  10297.5 205257.5 10362.5 205122.5 ;
      RECT  10297.5 205257.5 10362.5 205122.5 ;
      RECT  10107.5 205257.5 10172.5 205122.5 ;
      RECT  10297.5 205257.5 10362.5 205122.5 ;
      RECT  10487.5 205257.5 10552.5 205122.5 ;
      RECT  10487.5 205257.5 10552.5 205122.5 ;
      RECT  10297.5 205257.5 10362.5 205122.5 ;
      RECT  10107.5 206097.5 10172.5 205962.5 ;
      RECT  10297.5 206097.5 10362.5 205962.5 ;
      RECT  10297.5 206097.5 10362.5 205962.5 ;
      RECT  10107.5 206097.5 10172.5 205962.5 ;
      RECT  10297.5 206097.5 10362.5 205962.5 ;
      RECT  10487.5 206097.5 10552.5 205962.5 ;
      RECT  10487.5 206097.5 10552.5 205962.5 ;
      RECT  10297.5 206097.5 10362.5 205962.5 ;
      RECT  10657.5 205167.5 10722.5 205032.5 ;
      RECT  10657.5 206142.5 10722.5 206007.5 ;
      RECT  10492.5 205867.5 10357.5 205802.5 ;
      RECT  10235.0 205652.5 10100.0 205587.5 ;
      RECT  10297.5 205257.5 10362.5 205122.5 ;
      RECT  10487.5 206097.5 10552.5 205962.5 ;
      RECT  10587.5 205652.5 10452.5 205587.5 ;
      RECT  10100.0 205652.5 10235.0 205587.5 ;
      RECT  10357.5 205867.5 10492.5 205802.5 ;
      RECT  10452.5 205652.5 10587.5 205587.5 ;
      RECT  10040.0 204947.5 10960.0 204882.5 ;
      RECT  10040.0 206292.5 10960.0 206227.5 ;
      RECT  11387.5 205100.0 11452.5 204915.0 ;
      RECT  11387.5 206260.0 11452.5 206075.0 ;
      RECT  11027.5 206142.5 11092.5 206292.5 ;
      RECT  11027.5 205257.5 11092.5 204882.5 ;
      RECT  11217.5 206142.5 11282.5 205257.5 ;
      RECT  11027.5 205257.5 11092.5 205122.5 ;
      RECT  11217.5 205257.5 11282.5 205122.5 ;
      RECT  11217.5 205257.5 11282.5 205122.5 ;
      RECT  11027.5 205257.5 11092.5 205122.5 ;
      RECT  11027.5 206142.5 11092.5 206007.5 ;
      RECT  11217.5 206142.5 11282.5 206007.5 ;
      RECT  11217.5 206142.5 11282.5 206007.5 ;
      RECT  11027.5 206142.5 11092.5 206007.5 ;
      RECT  11387.5 205167.5 11452.5 205032.5 ;
      RECT  11387.5 206142.5 11452.5 206007.5 ;
      RECT  11085.0 205700.0 11150.0 205565.0 ;
      RECT  11085.0 205700.0 11150.0 205565.0 ;
      RECT  11250.0 205665.0 11315.0 205600.0 ;
      RECT  10960.0 204947.5 11520.0 204882.5 ;
      RECT  10960.0 206292.5 11520.0 206227.5 ;
      RECT  9222.5 205565.0 9287.5 205700.0 ;
      RECT  9362.5 205837.5 9427.5 205972.5 ;
      RECT  10357.5 205802.5 10222.5 205867.5 ;
      RECT  9025.0 34422.5 9395.0 34487.5 ;
      RECT  9025.0 36402.5 9395.0 36467.5 ;
      RECT  9025.0 37112.5 9395.0 37177.5 ;
      RECT  9025.0 39092.5 9395.0 39157.5 ;
      RECT  9025.0 39802.5 9395.0 39867.5 ;
      RECT  9025.0 41782.5 9395.0 41847.5 ;
      RECT  9025.0 42492.5 9395.0 42557.5 ;
      RECT  9025.0 44472.5 9395.0 44537.5 ;
      RECT  9025.0 45182.5 9395.0 45247.5 ;
      RECT  9025.0 47162.5 9395.0 47227.5 ;
      RECT  9025.0 47872.5 9395.0 47937.5 ;
      RECT  9025.0 49852.5 9395.0 49917.5 ;
      RECT  9025.0 50562.5 9395.0 50627.5 ;
      RECT  9025.0 52542.5 9395.0 52607.5 ;
      RECT  9025.0 53252.5 9395.0 53317.5 ;
      RECT  9025.0 55232.5 9395.0 55297.5 ;
      RECT  9025.0 55942.5 9395.0 56007.5 ;
      RECT  9025.0 57922.5 9395.0 57987.5 ;
      RECT  9025.0 58632.5 9395.0 58697.5 ;
      RECT  9025.0 60612.5 9395.0 60677.5 ;
      RECT  9025.0 61322.5 9395.0 61387.5 ;
      RECT  9025.0 63302.5 9395.0 63367.5 ;
      RECT  9025.0 64012.5 9395.0 64077.5 ;
      RECT  9025.0 65992.5 9395.0 66057.5 ;
      RECT  9025.0 66702.5 9395.0 66767.5 ;
      RECT  9025.0 68682.5 9395.0 68747.5 ;
      RECT  9025.0 69392.5 9395.0 69457.5 ;
      RECT  9025.0 71372.5 9395.0 71437.5 ;
      RECT  9025.0 72082.5 9395.0 72147.5 ;
      RECT  9025.0 74062.5 9395.0 74127.5 ;
      RECT  9025.0 74772.5 9395.0 74837.5 ;
      RECT  9025.0 76752.5 9395.0 76817.5 ;
      RECT  9025.0 77462.5 9395.0 77527.5 ;
      RECT  9025.0 79442.5 9395.0 79507.5 ;
      RECT  9025.0 80152.5 9395.0 80217.5 ;
      RECT  9025.0 82132.5 9395.0 82197.5 ;
      RECT  9025.0 82842.5 9395.0 82907.5 ;
      RECT  9025.0 84822.5 9395.0 84887.5 ;
      RECT  9025.0 85532.5 9395.0 85597.5 ;
      RECT  9025.0 87512.5 9395.0 87577.5 ;
      RECT  9025.0 88222.5 9395.0 88287.5 ;
      RECT  9025.0 90202.5 9395.0 90267.5 ;
      RECT  9025.0 90912.5 9395.0 90977.5 ;
      RECT  9025.0 92892.5 9395.0 92957.5 ;
      RECT  9025.0 93602.5 9395.0 93667.5 ;
      RECT  9025.0 95582.5 9395.0 95647.5 ;
      RECT  9025.0 96292.5 9395.0 96357.5 ;
      RECT  9025.0 98272.5 9395.0 98337.5 ;
      RECT  9025.0 98982.5 9395.0 99047.5 ;
      RECT  9025.0 100962.5 9395.0 101027.5 ;
      RECT  9025.0 101672.5 9395.0 101737.5 ;
      RECT  9025.0 103652.5 9395.0 103717.5 ;
      RECT  9025.0 104362.5 9395.0 104427.5 ;
      RECT  9025.0 106342.5 9395.0 106407.5 ;
      RECT  9025.0 107052.5 9395.0 107117.5 ;
      RECT  9025.0 109032.5 9395.0 109097.5 ;
      RECT  9025.0 109742.5 9395.0 109807.5 ;
      RECT  9025.0 111722.5 9395.0 111787.5 ;
      RECT  9025.0 112432.5 9395.0 112497.5 ;
      RECT  9025.0 114412.5 9395.0 114477.5 ;
      RECT  9025.0 115122.5 9395.0 115187.5 ;
      RECT  9025.0 117102.5 9395.0 117167.5 ;
      RECT  9025.0 117812.5 9395.0 117877.5 ;
      RECT  9025.0 119792.5 9395.0 119857.5 ;
      RECT  9025.0 120502.5 9395.0 120567.5 ;
      RECT  9025.0 122482.5 9395.0 122547.5 ;
      RECT  9025.0 123192.5 9395.0 123257.5 ;
      RECT  9025.0 125172.5 9395.0 125237.5 ;
      RECT  9025.0 125882.5 9395.0 125947.5 ;
      RECT  9025.0 127862.5 9395.0 127927.5 ;
      RECT  9025.0 128572.5 9395.0 128637.5 ;
      RECT  9025.0 130552.5 9395.0 130617.5 ;
      RECT  9025.0 131262.5 9395.0 131327.5 ;
      RECT  9025.0 133242.5 9395.0 133307.5 ;
      RECT  9025.0 133952.5 9395.0 134017.5 ;
      RECT  9025.0 135932.5 9395.0 135997.5 ;
      RECT  9025.0 136642.5 9395.0 136707.5 ;
      RECT  9025.0 138622.5 9395.0 138687.5 ;
      RECT  9025.0 139332.5 9395.0 139397.5 ;
      RECT  9025.0 141312.5 9395.0 141377.5 ;
      RECT  9025.0 142022.5 9395.0 142087.5 ;
      RECT  9025.0 144002.5 9395.0 144067.5 ;
      RECT  9025.0 144712.5 9395.0 144777.5 ;
      RECT  9025.0 146692.5 9395.0 146757.5 ;
      RECT  9025.0 147402.5 9395.0 147467.5 ;
      RECT  9025.0 149382.5 9395.0 149447.5 ;
      RECT  9025.0 150092.5 9395.0 150157.5 ;
      RECT  9025.0 152072.5 9395.0 152137.5 ;
      RECT  9025.0 152782.5 9395.0 152847.5 ;
      RECT  9025.0 154762.5 9395.0 154827.5 ;
      RECT  9025.0 155472.5 9395.0 155537.5 ;
      RECT  9025.0 157452.5 9395.0 157517.5 ;
      RECT  9025.0 158162.5 9395.0 158227.5 ;
      RECT  9025.0 160142.5 9395.0 160207.5 ;
      RECT  9025.0 160852.5 9395.0 160917.5 ;
      RECT  9025.0 162832.5 9395.0 162897.5 ;
      RECT  9025.0 163542.5 9395.0 163607.5 ;
      RECT  9025.0 165522.5 9395.0 165587.5 ;
      RECT  9025.0 166232.5 9395.0 166297.5 ;
      RECT  9025.0 168212.5 9395.0 168277.5 ;
      RECT  9025.0 168922.5 9395.0 168987.5 ;
      RECT  9025.0 170902.5 9395.0 170967.5 ;
      RECT  9025.0 171612.5 9395.0 171677.5 ;
      RECT  9025.0 173592.5 9395.0 173657.5 ;
      RECT  9025.0 174302.5 9395.0 174367.5 ;
      RECT  9025.0 176282.5 9395.0 176347.5 ;
      RECT  9025.0 176992.5 9395.0 177057.5 ;
      RECT  9025.0 178972.5 9395.0 179037.5 ;
      RECT  9025.0 179682.5 9395.0 179747.5 ;
      RECT  9025.0 181662.5 9395.0 181727.5 ;
      RECT  9025.0 182372.5 9395.0 182437.5 ;
      RECT  9025.0 184352.5 9395.0 184417.5 ;
      RECT  9025.0 185062.5 9395.0 185127.5 ;
      RECT  9025.0 187042.5 9395.0 187107.5 ;
      RECT  9025.0 187752.5 9395.0 187817.5 ;
      RECT  9025.0 189732.5 9395.0 189797.5 ;
      RECT  9025.0 190442.5 9395.0 190507.5 ;
      RECT  9025.0 192422.5 9395.0 192487.5 ;
      RECT  9025.0 193132.5 9395.0 193197.5 ;
      RECT  9025.0 195112.5 9395.0 195177.5 ;
      RECT  9025.0 195822.5 9395.0 195887.5 ;
      RECT  9025.0 197802.5 9395.0 197867.5 ;
      RECT  9025.0 198512.5 9395.0 198577.5 ;
      RECT  9025.0 200492.5 9395.0 200557.5 ;
      RECT  9025.0 201202.5 9395.0 201267.5 ;
      RECT  9025.0 203182.5 9395.0 203247.5 ;
      RECT  9025.0 203892.5 9395.0 203957.5 ;
      RECT  9025.0 205872.5 9395.0 205937.5 ;
      RECT  11250.0 34695.0 11315.0 34760.0 ;
      RECT  11250.0 36130.0 11315.0 36195.0 ;
      RECT  11250.0 37385.0 11315.0 37450.0 ;
      RECT  11250.0 38820.0 11315.0 38885.0 ;
      RECT  11250.0 40075.0 11315.0 40140.0 ;
      RECT  11250.0 41510.0 11315.0 41575.0 ;
      RECT  11250.0 42765.0 11315.0 42830.0 ;
      RECT  11250.0 44200.0 11315.0 44265.0 ;
      RECT  11250.0 45455.0 11315.0 45520.0 ;
      RECT  11250.0 46890.0 11315.0 46955.0 ;
      RECT  11250.0 48145.0 11315.0 48210.0 ;
      RECT  11250.0 49580.0 11315.0 49645.0 ;
      RECT  11250.0 50835.0 11315.0 50900.0 ;
      RECT  11250.0 52270.0 11315.0 52335.0 ;
      RECT  11250.0 53525.0 11315.0 53590.0 ;
      RECT  11250.0 54960.0 11315.0 55025.0 ;
      RECT  11250.0 56215.0 11315.0 56280.0 ;
      RECT  11250.0 57650.0 11315.0 57715.0 ;
      RECT  11250.0 58905.0 11315.0 58970.0 ;
      RECT  11250.0 60340.0 11315.0 60405.0 ;
      RECT  11250.0 61595.0 11315.0 61660.0 ;
      RECT  11250.0 63030.0 11315.0 63095.0 ;
      RECT  11250.0 64285.0 11315.0 64350.0 ;
      RECT  11250.0 65720.0 11315.0 65785.0 ;
      RECT  11250.0 66975.0 11315.0 67040.0 ;
      RECT  11250.0 68410.0 11315.0 68475.0 ;
      RECT  11250.0 69665.0 11315.0 69730.0 ;
      RECT  11250.0 71100.0 11315.0 71165.0 ;
      RECT  11250.0 72355.0 11315.0 72420.0 ;
      RECT  11250.0 73790.0 11315.0 73855.0 ;
      RECT  11250.0 75045.0 11315.0 75110.0 ;
      RECT  11250.0 76480.0 11315.0 76545.0 ;
      RECT  11250.0 77735.0 11315.0 77800.0 ;
      RECT  11250.0 79170.0 11315.0 79235.0 ;
      RECT  11250.0 80425.0 11315.0 80490.0 ;
      RECT  11250.0 81860.0 11315.0 81925.0 ;
      RECT  11250.0 83115.0 11315.0 83180.0 ;
      RECT  11250.0 84550.0 11315.0 84615.0 ;
      RECT  11250.0 85805.0 11315.0 85870.0 ;
      RECT  11250.0 87240.0 11315.0 87305.0 ;
      RECT  11250.0 88495.0 11315.0 88560.0 ;
      RECT  11250.0 89930.0 11315.0 89995.0 ;
      RECT  11250.0 91185.0 11315.0 91250.0 ;
      RECT  11250.0 92620.0 11315.0 92685.0 ;
      RECT  11250.0 93875.0 11315.0 93940.0 ;
      RECT  11250.0 95310.0 11315.0 95375.0 ;
      RECT  11250.0 96565.0 11315.0 96630.0 ;
      RECT  11250.0 98000.0 11315.0 98065.0 ;
      RECT  11250.0 99255.0 11315.0 99320.0 ;
      RECT  11250.0 100690.0 11315.0 100755.0 ;
      RECT  11250.0 101945.0 11315.0 102010.0 ;
      RECT  11250.0 103380.0 11315.0 103445.0 ;
      RECT  11250.0 104635.0 11315.0 104700.0 ;
      RECT  11250.0 106070.0 11315.0 106135.0 ;
      RECT  11250.0 107325.0 11315.0 107390.0 ;
      RECT  11250.0 108760.0 11315.0 108825.0 ;
      RECT  11250.0 110015.0 11315.0 110080.0 ;
      RECT  11250.0 111450.0 11315.0 111515.0 ;
      RECT  11250.0 112705.0 11315.0 112770.0 ;
      RECT  11250.0 114140.0 11315.0 114205.0 ;
      RECT  11250.0 115395.0 11315.0 115460.0 ;
      RECT  11250.0 116830.0 11315.0 116895.0 ;
      RECT  11250.0 118085.0 11315.0 118150.0 ;
      RECT  11250.0 119520.0 11315.0 119585.0 ;
      RECT  11250.0 120775.0 11315.0 120840.0 ;
      RECT  11250.0 122210.0 11315.0 122275.0 ;
      RECT  11250.0 123465.0 11315.0 123530.0 ;
      RECT  11250.0 124900.0 11315.0 124965.0 ;
      RECT  11250.0 126155.0 11315.0 126220.0 ;
      RECT  11250.0 127590.0 11315.0 127655.0 ;
      RECT  11250.0 128845.0 11315.0 128910.0 ;
      RECT  11250.0 130280.0 11315.0 130345.0 ;
      RECT  11250.0 131535.0 11315.0 131600.0 ;
      RECT  11250.0 132970.0 11315.0 133035.0 ;
      RECT  11250.0 134225.0 11315.0 134290.0 ;
      RECT  11250.0 135660.0 11315.0 135725.0 ;
      RECT  11250.0 136915.0 11315.0 136980.0 ;
      RECT  11250.0 138350.0 11315.0 138415.0 ;
      RECT  11250.0 139605.0 11315.0 139670.0 ;
      RECT  11250.0 141040.0 11315.0 141105.0 ;
      RECT  11250.0 142295.0 11315.0 142360.0 ;
      RECT  11250.0 143730.0 11315.0 143795.0 ;
      RECT  11250.0 144985.0 11315.0 145050.0 ;
      RECT  11250.0 146420.0 11315.0 146485.0 ;
      RECT  11250.0 147675.0 11315.0 147740.0 ;
      RECT  11250.0 149110.0 11315.0 149175.0 ;
      RECT  11250.0 150365.0 11315.0 150430.0 ;
      RECT  11250.0 151800.0 11315.0 151865.0 ;
      RECT  11250.0 153055.0 11315.0 153120.0 ;
      RECT  11250.0 154490.0 11315.0 154555.0 ;
      RECT  11250.0 155745.0 11315.0 155810.0 ;
      RECT  11250.0 157180.0 11315.0 157245.0 ;
      RECT  11250.0 158435.0 11315.0 158500.0 ;
      RECT  11250.0 159870.0 11315.0 159935.0 ;
      RECT  11250.0 161125.0 11315.0 161190.0 ;
      RECT  11250.0 162560.0 11315.0 162625.0 ;
      RECT  11250.0 163815.0 11315.0 163880.0 ;
      RECT  11250.0 165250.0 11315.0 165315.0 ;
      RECT  11250.0 166505.0 11315.0 166570.0 ;
      RECT  11250.0 167940.0 11315.0 168005.0 ;
      RECT  11250.0 169195.0 11315.0 169260.0 ;
      RECT  11250.0 170630.0 11315.0 170695.0 ;
      RECT  11250.0 171885.0 11315.0 171950.0 ;
      RECT  11250.0 173320.0 11315.0 173385.0 ;
      RECT  11250.0 174575.0 11315.0 174640.0 ;
      RECT  11250.0 176010.0 11315.0 176075.0 ;
      RECT  11250.0 177265.0 11315.0 177330.0 ;
      RECT  11250.0 178700.0 11315.0 178765.0 ;
      RECT  11250.0 179955.0 11315.0 180020.0 ;
      RECT  11250.0 181390.0 11315.0 181455.0 ;
      RECT  11250.0 182645.0 11315.0 182710.0 ;
      RECT  11250.0 184080.0 11315.0 184145.0 ;
      RECT  11250.0 185335.0 11315.0 185400.0 ;
      RECT  11250.0 186770.0 11315.0 186835.0 ;
      RECT  11250.0 188025.0 11315.0 188090.0 ;
      RECT  11250.0 189460.0 11315.0 189525.0 ;
      RECT  11250.0 190715.0 11315.0 190780.0 ;
      RECT  11250.0 192150.0 11315.0 192215.0 ;
      RECT  11250.0 193405.0 11315.0 193470.0 ;
      RECT  11250.0 194840.0 11315.0 194905.0 ;
      RECT  11250.0 196095.0 11315.0 196160.0 ;
      RECT  11250.0 197530.0 11315.0 197595.0 ;
      RECT  11250.0 198785.0 11315.0 198850.0 ;
      RECT  11250.0 200220.0 11315.0 200285.0 ;
      RECT  11250.0 201475.0 11315.0 201540.0 ;
      RECT  11250.0 202910.0 11315.0 202975.0 ;
      RECT  11250.0 204165.0 11315.0 204230.0 ;
      RECT  11250.0 205600.0 11315.0 205665.0 ;
      RECT  9025.0 35412.5 9480.0 35477.5 ;
      RECT  9025.0 38102.5 9480.0 38167.5 ;
      RECT  9025.0 40792.5 9480.0 40857.5 ;
      RECT  9025.0 43482.5 9480.0 43547.5 ;
      RECT  9025.0 46172.5 9480.0 46237.5 ;
      RECT  9025.0 48862.5 9480.0 48927.5 ;
      RECT  9025.0 51552.5 9480.0 51617.5 ;
      RECT  9025.0 54242.5 9480.0 54307.5 ;
      RECT  9025.0 56932.5 9480.0 56997.5 ;
      RECT  9025.0 59622.5 9480.0 59687.5 ;
      RECT  9025.0 62312.5 9480.0 62377.5 ;
      RECT  9025.0 65002.5 9480.0 65067.5 ;
      RECT  9025.0 67692.5 9480.0 67757.5 ;
      RECT  9025.0 70382.5 9480.0 70447.5 ;
      RECT  9025.0 73072.5 9480.0 73137.5 ;
      RECT  9025.0 75762.5 9480.0 75827.5 ;
      RECT  9025.0 78452.5 9480.0 78517.5 ;
      RECT  9025.0 81142.5 9480.0 81207.5 ;
      RECT  9025.0 83832.5 9480.0 83897.5 ;
      RECT  9025.0 86522.5 9480.0 86587.5 ;
      RECT  9025.0 89212.5 9480.0 89277.5 ;
      RECT  9025.0 91902.5 9480.0 91967.5 ;
      RECT  9025.0 94592.5 9480.0 94657.5 ;
      RECT  9025.0 97282.5 9480.0 97347.5 ;
      RECT  9025.0 99972.5 9480.0 100037.5 ;
      RECT  9025.0 102662.5 9480.0 102727.5 ;
      RECT  9025.0 105352.5 9480.0 105417.5 ;
      RECT  9025.0 108042.5 9480.0 108107.5 ;
      RECT  9025.0 110732.5 9480.0 110797.5 ;
      RECT  9025.0 113422.5 9480.0 113487.5 ;
      RECT  9025.0 116112.5 9480.0 116177.5 ;
      RECT  9025.0 118802.5 9480.0 118867.5 ;
      RECT  9025.0 121492.5 9480.0 121557.5 ;
      RECT  9025.0 124182.5 9480.0 124247.5 ;
      RECT  9025.0 126872.5 9480.0 126937.5 ;
      RECT  9025.0 129562.5 9480.0 129627.5 ;
      RECT  9025.0 132252.5 9480.0 132317.5 ;
      RECT  9025.0 134942.5 9480.0 135007.5 ;
      RECT  9025.0 137632.5 9480.0 137697.5 ;
      RECT  9025.0 140322.5 9480.0 140387.5 ;
      RECT  9025.0 143012.5 9480.0 143077.5 ;
      RECT  9025.0 145702.5 9480.0 145767.5 ;
      RECT  9025.0 148392.5 9480.0 148457.5 ;
      RECT  9025.0 151082.5 9480.0 151147.5 ;
      RECT  9025.0 153772.5 9480.0 153837.5 ;
      RECT  9025.0 156462.5 9480.0 156527.5 ;
      RECT  9025.0 159152.5 9480.0 159217.5 ;
      RECT  9025.0 161842.5 9480.0 161907.5 ;
      RECT  9025.0 164532.5 9480.0 164597.5 ;
      RECT  9025.0 167222.5 9480.0 167287.5 ;
      RECT  9025.0 169912.5 9480.0 169977.5 ;
      RECT  9025.0 172602.5 9480.0 172667.5 ;
      RECT  9025.0 175292.5 9480.0 175357.5 ;
      RECT  9025.0 177982.5 9480.0 178047.5 ;
      RECT  9025.0 180672.5 9480.0 180737.5 ;
      RECT  9025.0 183362.5 9480.0 183427.5 ;
      RECT  9025.0 186052.5 9480.0 186117.5 ;
      RECT  9025.0 188742.5 9480.0 188807.5 ;
      RECT  9025.0 191432.5 9480.0 191497.5 ;
      RECT  9025.0 194122.5 9480.0 194187.5 ;
      RECT  9025.0 196812.5 9480.0 196877.5 ;
      RECT  9025.0 199502.5 9480.0 199567.5 ;
      RECT  9025.0 202192.5 9480.0 202257.5 ;
      RECT  9025.0 204882.5 9480.0 204947.5 ;
      RECT  9025.0 34067.5 9480.0 34132.5 ;
      RECT  9025.0 36757.5 9480.0 36822.5 ;
      RECT  9025.0 39447.5 9480.0 39512.5 ;
      RECT  9025.0 42137.5 9480.0 42202.5 ;
      RECT  9025.0 44827.5 9480.0 44892.5 ;
      RECT  9025.0 47517.5 9480.0 47582.5 ;
      RECT  9025.0 50207.5 9480.0 50272.5 ;
      RECT  9025.0 52897.5 9480.0 52962.5 ;
      RECT  9025.0 55587.5 9480.0 55652.5 ;
      RECT  9025.0 58277.5 9480.0 58342.5 ;
      RECT  9025.0 60967.5 9480.0 61032.5 ;
      RECT  9025.0 63657.5 9480.0 63722.5 ;
      RECT  9025.0 66347.5 9480.0 66412.5 ;
      RECT  9025.0 69037.5 9480.0 69102.5 ;
      RECT  9025.0 71727.5 9480.0 71792.5 ;
      RECT  9025.0 74417.5 9480.0 74482.5 ;
      RECT  9025.0 77107.5 9480.0 77172.5 ;
      RECT  9025.0 79797.5 9480.0 79862.5 ;
      RECT  9025.0 82487.5 9480.0 82552.5 ;
      RECT  9025.0 85177.5 9480.0 85242.5 ;
      RECT  9025.0 87867.5 9480.0 87932.5 ;
      RECT  9025.0 90557.5 9480.0 90622.5 ;
      RECT  9025.0 93247.5 9480.0 93312.5 ;
      RECT  9025.0 95937.5 9480.0 96002.5 ;
      RECT  9025.0 98627.5 9480.0 98692.5 ;
      RECT  9025.0 101317.5 9480.0 101382.5 ;
      RECT  9025.0 104007.5 9480.0 104072.5 ;
      RECT  9025.0 106697.5 9480.0 106762.5 ;
      RECT  9025.0 109387.5 9480.0 109452.5 ;
      RECT  9025.0 112077.5 9480.0 112142.5 ;
      RECT  9025.0 114767.5 9480.0 114832.5 ;
      RECT  9025.0 117457.5 9480.0 117522.5 ;
      RECT  9025.0 120147.5 9480.0 120212.5 ;
      RECT  9025.0 122837.5 9480.0 122902.5 ;
      RECT  9025.0 125527.5 9480.0 125592.5 ;
      RECT  9025.0 128217.5 9480.0 128282.5 ;
      RECT  9025.0 130907.5 9480.0 130972.5 ;
      RECT  9025.0 133597.5 9480.0 133662.5 ;
      RECT  9025.0 136287.5 9480.0 136352.5 ;
      RECT  9025.0 138977.5 9480.0 139042.5 ;
      RECT  9025.0 141667.5 9480.0 141732.5 ;
      RECT  9025.0 144357.5 9480.0 144422.5 ;
      RECT  9025.0 147047.5 9480.0 147112.5 ;
      RECT  9025.0 149737.5 9480.0 149802.5 ;
      RECT  9025.0 152427.5 9480.0 152492.5 ;
      RECT  9025.0 155117.5 9480.0 155182.5 ;
      RECT  9025.0 157807.5 9480.0 157872.5 ;
      RECT  9025.0 160497.5 9480.0 160562.5 ;
      RECT  9025.0 163187.5 9480.0 163252.5 ;
      RECT  9025.0 165877.5 9480.0 165942.5 ;
      RECT  9025.0 168567.5 9480.0 168632.5 ;
      RECT  9025.0 171257.5 9480.0 171322.5 ;
      RECT  9025.0 173947.5 9480.0 174012.5 ;
      RECT  9025.0 176637.5 9480.0 176702.5 ;
      RECT  9025.0 179327.5 9480.0 179392.5 ;
      RECT  9025.0 182017.5 9480.0 182082.5 ;
      RECT  9025.0 184707.5 9480.0 184772.5 ;
      RECT  9025.0 187397.5 9480.0 187462.5 ;
      RECT  9025.0 190087.5 9480.0 190152.5 ;
      RECT  9025.0 192777.5 9480.0 192842.5 ;
      RECT  9025.0 195467.5 9480.0 195532.5 ;
      RECT  9025.0 198157.5 9480.0 198222.5 ;
      RECT  9025.0 200847.5 9480.0 200912.5 ;
      RECT  9025.0 203537.5 9480.0 203602.5 ;
      RECT  9025.0 206227.5 9480.0 206292.5 ;
      RECT  4655.0 12170.0 11095.0 11465.0 ;
      RECT  4655.0 10760.0 11095.0 11465.0 ;
      RECT  4655.0 10760.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 5825.0 ;
      RECT  4860.0 12170.0 4925.0 5825.0 ;
      RECT  7865.0 12170.0 7930.0 5825.0 ;
      RECT  10825.0 12170.0 10890.0 5825.0 ;
      RECT  5875.0 12170.0 5940.0 5825.0 ;
      RECT  8835.0 12170.0 8900.0 5825.0 ;
      RECT  5020.0 12170.0 5085.0 5825.0 ;
      RECT  15102.5 34132.5 15237.5 34067.5 ;
      RECT  15102.5 36822.5 15237.5 36757.5 ;
      RECT  15102.5 39512.5 15237.5 39447.5 ;
      RECT  15102.5 42202.5 15237.5 42137.5 ;
      RECT  15102.5 44892.5 15237.5 44827.5 ;
      RECT  15102.5 47582.5 15237.5 47517.5 ;
      RECT  15102.5 50272.5 15237.5 50207.5 ;
      RECT  15102.5 52962.5 15237.5 52897.5 ;
      RECT  15102.5 55652.5 15237.5 55587.5 ;
      RECT  15102.5 58342.5 15237.5 58277.5 ;
      RECT  15102.5 61032.5 15237.5 60967.5 ;
      RECT  15102.5 63722.5 15237.5 63657.5 ;
      RECT  15102.5 66412.5 15237.5 66347.5 ;
      RECT  15102.5 69102.5 15237.5 69037.5 ;
      RECT  15102.5 71792.5 15237.5 71727.5 ;
      RECT  15102.5 74482.5 15237.5 74417.5 ;
      RECT  15102.5 77172.5 15237.5 77107.5 ;
      RECT  15102.5 79862.5 15237.5 79797.5 ;
      RECT  15102.5 82552.5 15237.5 82487.5 ;
      RECT  15102.5 85242.5 15237.5 85177.5 ;
      RECT  15102.5 87932.5 15237.5 87867.5 ;
      RECT  15102.5 90622.5 15237.5 90557.5 ;
      RECT  15102.5 93312.5 15237.5 93247.5 ;
      RECT  15102.5 96002.5 15237.5 95937.5 ;
      RECT  15102.5 98692.5 15237.5 98627.5 ;
      RECT  15102.5 101382.5 15237.5 101317.5 ;
      RECT  15102.5 104072.5 15237.5 104007.5 ;
      RECT  15102.5 106762.5 15237.5 106697.5 ;
      RECT  15102.5 109452.5 15237.5 109387.5 ;
      RECT  15102.5 112142.5 15237.5 112077.5 ;
      RECT  15102.5 114832.5 15237.5 114767.5 ;
      RECT  15102.5 117522.5 15237.5 117457.5 ;
      RECT  15102.5 120212.5 15237.5 120147.5 ;
      RECT  15102.5 122902.5 15237.5 122837.5 ;
      RECT  15102.5 125592.5 15237.5 125527.5 ;
      RECT  15102.5 128282.5 15237.5 128217.5 ;
      RECT  15102.5 130972.5 15237.5 130907.5 ;
      RECT  15102.5 133662.5 15237.5 133597.5 ;
      RECT  15102.5 136352.5 15237.5 136287.5 ;
      RECT  15102.5 139042.5 15237.5 138977.5 ;
      RECT  15102.5 141732.5 15237.5 141667.5 ;
      RECT  15102.5 144422.5 15237.5 144357.5 ;
      RECT  15102.5 147112.5 15237.5 147047.5 ;
      RECT  15102.5 149802.5 15237.5 149737.5 ;
      RECT  15102.5 152492.5 15237.5 152427.5 ;
      RECT  15102.5 155182.5 15237.5 155117.5 ;
      RECT  15102.5 157872.5 15237.5 157807.5 ;
      RECT  15102.5 160562.5 15237.5 160497.5 ;
      RECT  15102.5 163252.5 15237.5 163187.5 ;
      RECT  15102.5 165942.5 15237.5 165877.5 ;
      RECT  15102.5 168632.5 15237.5 168567.5 ;
      RECT  15102.5 171322.5 15237.5 171257.5 ;
      RECT  15102.5 174012.5 15237.5 173947.5 ;
      RECT  15102.5 176702.5 15237.5 176637.5 ;
      RECT  15102.5 179392.5 15237.5 179327.5 ;
      RECT  15102.5 182082.5 15237.5 182017.5 ;
      RECT  15102.5 184772.5 15237.5 184707.5 ;
      RECT  15102.5 187462.5 15237.5 187397.5 ;
      RECT  15102.5 190152.5 15237.5 190087.5 ;
      RECT  15102.5 192842.5 15237.5 192777.5 ;
      RECT  15102.5 195532.5 15237.5 195467.5 ;
      RECT  15102.5 198222.5 15237.5 198157.5 ;
      RECT  15102.5 200912.5 15237.5 200847.5 ;
      RECT  15102.5 203602.5 15237.5 203537.5 ;
      RECT  15102.5 206292.5 15237.5 206227.5 ;
      RECT  11420.0 12752.5 11285.0 12817.5 ;
      RECT  12745.0 12752.5 12610.0 12817.5 ;
      RECT  11145.0 14097.5 11010.0 14162.5 ;
      RECT  12950.0 14097.5 12815.0 14162.5 ;
      RECT  11420.0 18132.5 11285.0 18197.5 ;
      RECT  13155.0 18132.5 13020.0 18197.5 ;
      RECT  11145.0 19477.5 11010.0 19542.5 ;
      RECT  13360.0 19477.5 13225.0 19542.5 ;
      RECT  12335.0 23512.5 12200.0 23577.5 ;
      RECT  13565.0 23512.5 13430.0 23577.5 ;
      RECT  12060.0 24857.5 11925.0 24922.5 ;
      RECT  13770.0 24857.5 13635.0 24922.5 ;
      RECT  11785.0 26202.5 11650.0 26267.5 ;
      RECT  13975.0 26202.5 13840.0 26267.5 ;
      RECT  12540.0 12547.5 12405.0 12612.5 ;
      RECT  12540.0 15237.5 12405.0 15302.5 ;
      RECT  12540.0 17927.5 12405.0 17992.5 ;
      RECT  12540.0 20617.5 12405.0 20682.5 ;
      RECT  12540.0 23307.5 12405.0 23372.5 ;
      RECT  12540.0 25997.5 12405.0 26062.5 ;
      RECT  12540.0 28687.5 12405.0 28752.5 ;
      RECT  12540.0 31377.5 12405.0 31442.5 ;
      RECT  14180.0 32097.5 14045.0 32162.5 ;
      RECT  14385.0 31957.5 14250.0 32022.5 ;
      RECT  14590.0 31817.5 14455.0 31882.5 ;
      RECT  14795.0 31677.5 14660.0 31742.5 ;
      RECT  14180.0 630.0 14045.0 695.0 ;
      RECT  14385.0 2065.0 14250.0 2130.0 ;
      RECT  14590.0 3320.0 14455.0 3385.0 ;
      RECT  14795.0 4755.0 14660.0 4820.0 ;
      RECT  15102.5 67.5 15237.5 2.5 ;
      RECT  15102.5 2757.5 15237.5 2692.5 ;
      RECT  15102.5 5447.5 15237.5 5382.5 ;
      RECT  11162.5 11785.0 11027.5 11850.0 ;
      RECT  12745.0 11785.0 12610.0 11850.0 ;
      RECT  11162.5 11080.0 11027.5 11145.0 ;
      RECT  12950.0 11080.0 12815.0 11145.0 ;
      RECT  11162.5 10375.0 11027.5 10440.0 ;
      RECT  13155.0 10375.0 13020.0 10440.0 ;
      RECT  11162.5 9670.0 11027.5 9735.0 ;
      RECT  13360.0 9670.0 13225.0 9735.0 ;
      RECT  11162.5 8965.0 11027.5 9030.0 ;
      RECT  13565.0 8965.0 13430.0 9030.0 ;
      RECT  11162.5 8260.0 11027.5 8325.0 ;
      RECT  13770.0 8260.0 13635.0 8325.0 ;
      RECT  11162.5 7555.0 11027.5 7620.0 ;
      RECT  13975.0 7555.0 13840.0 7620.0 ;
      RECT  11230.0 12137.5 11095.0 12202.5 ;
      RECT  15237.5 12137.5 15102.5 12202.5 ;
      RECT  11230.0 11432.5 11095.0 11497.5 ;
      RECT  15237.5 11432.5 15102.5 11497.5 ;
      RECT  11230.0 10727.5 11095.0 10792.5 ;
      RECT  15237.5 10727.5 15102.5 10792.5 ;
      RECT  11230.0 10022.5 11095.0 10087.5 ;
      RECT  15237.5 10022.5 15102.5 10087.5 ;
      RECT  11230.0 9317.5 11095.0 9382.5 ;
      RECT  15237.5 9317.5 15102.5 9382.5 ;
      RECT  11230.0 8612.5 11095.0 8677.5 ;
      RECT  15237.5 8612.5 15102.5 8677.5 ;
      RECT  11230.0 7907.5 11095.0 7972.5 ;
      RECT  15237.5 7907.5 15102.5 7972.5 ;
      RECT  11230.0 7202.5 11095.0 7267.5 ;
      RECT  15237.5 7202.5 15102.5 7267.5 ;
      RECT  11230.0 6497.5 11095.0 6562.5 ;
      RECT  15237.5 6497.5 15102.5 6562.5 ;
      RECT  11230.0 5792.5 11095.0 5857.5 ;
      RECT  15237.5 5792.5 15102.5 5857.5 ;
      RECT  16375.0 15960.0 16240.0 16025.0 ;
      RECT  15965.0 13775.0 15830.0 13840.0 ;
      RECT  16170.0 15322.5 16035.0 15387.5 ;
      RECT  16375.0 207237.5 16240.0 207302.5 ;
      RECT  16580.0 22462.5 16445.0 22527.5 ;
      RECT  16785.0 26487.5 16650.0 26552.5 ;
      RECT  15760.0 12342.5 15625.0 12407.5 ;
      RECT  9322.5 206432.5 9187.5 206497.5 ;
      RECT  15760.0 206432.5 15625.0 206497.5 ;
      RECT  15452.5 15192.5 15317.5 15257.5 ;
      RECT  15452.5 26617.5 15317.5 26682.5 ;
      RECT  15452.5 16120.0 15317.5 16185.0 ;
      RECT  15452.5 23395.0 15317.5 23460.0 ;
      RECT  107630.0 35.0 107980.0 207987.5 ;
      RECT  4175.0 35.0 4525.0 207987.5 ;
      RECT  3455.0 34530.0 3390.0 34595.0 ;
      RECT  3422.5 34530.0 3407.5 34595.0 ;
      RECT  3455.0 34562.5 3390.0 35147.5 ;
      RECT  3455.0 35692.5 3390.0 36087.5 ;
      RECT  3455.0 37012.5 3390.0 37597.5 ;
      RECT  2657.5 37450.0 2280.0 37515.0 ;
      RECT  2657.5 40410.0 2280.0 40475.0 ;
      RECT  2657.5 35460.0 2280.0 35525.0 ;
      RECT  2657.5 38420.0 2280.0 38485.0 ;
      RECT  3440.0 34530.0 3375.0 34595.0 ;
      RECT  3455.0 35660.0 3390.0 35725.0 ;
      RECT  2005.0 46345.0 1940.0 47110.0 ;
      RECT  3455.0 39695.0 3390.0 41125.0 ;
      RECT  2485.0 34445.0 2280.0 34510.0 ;
      RECT  1962.5 41125.0 1897.5 43062.5 ;
      RECT  1747.5 41535.0 1682.5 43320.0 ;
      RECT  3380.0 42560.0 3315.0 43130.0 ;
      RECT  3520.0 42355.0 3455.0 43320.0 ;
      RECT  3660.0 41740.0 3595.0 43510.0 ;
      RECT  3380.0 44070.0 3315.0 44135.0 ;
      RECT  3380.0 43605.0 3315.0 44102.5 ;
      RECT  3407.5 44070.0 3347.5 44135.0 ;
      RECT  3475.0 44235.0 3410.0 44300.0 ;
      RECT  3442.5 44235.0 3407.5 44300.0 ;
      RECT  3475.0 44267.5 3410.0 47807.5 ;
      RECT  690.0 42560.0 625.0 43690.0 ;
      RECT  830.0 41740.0 765.0 43880.0 ;
      RECT  970.0 41945.0 905.0 44070.0 ;
      RECT  690.0 44630.0 625.0 44695.0 ;
      RECT  690.0 44165.0 625.0 44662.5 ;
      RECT  717.5 44630.0 657.5 44695.0 ;
      RECT  750.0 44827.5 685.0 45222.5 ;
      RECT  750.0 45387.5 685.0 45782.5 ;
      RECT  2005.0 46312.5 1940.0 46377.5 ;
      RECT  1972.5 46312.5 1940.0 46377.5 ;
      RECT  2005.0 46220.0 1940.0 46345.0 ;
      RECT  2005.0 45627.5 1940.0 46022.5 ;
      RECT  1962.5 43485.0 1897.5 43855.0 ;
      RECT  2017.5 44560.0 1952.5 45000.0 ;
      RECT  750.0 45947.5 685.0 46185.0 ;
      RECT  2005.0 45225.0 1940.0 45462.5 ;
      RECT  4067.5 34240.0 4002.5 46345.0 ;
      RECT  4067.5 41330.0 4002.5 42935.0 ;
      RECT  2722.5 34240.0 2657.5 46345.0 ;
      RECT  2722.5 42150.0 2657.5 42935.0 ;
      RECT  1377.5 42935.0 1312.5 46345.0 ;
      RECT  1377.5 41330.0 1312.5 42935.0 ;
      RECT  32.5 42935.0 -32.5 46345.0 ;
      RECT  32.5 42150.0 -32.5 42935.0 ;
      RECT  32.5 46312.5 -32.5 46377.5 ;
      RECT  32.5 46140.0 -32.5 46345.0 ;
      RECT  8.881784197e-13 46312.5 -45.0 46377.5 ;
      RECT  165.0 34240.0 870.0 40680.0 ;
      RECT  1575.0 34240.0 870.0 40680.0 ;
      RECT  1575.0 34240.0 2280.0 40680.0 ;
      RECT  165.0 34445.0 2280.0 34510.0 ;
      RECT  165.0 37450.0 2280.0 37515.0 ;
      RECT  165.0 40410.0 2280.0 40475.0 ;
      RECT  165.0 35460.0 2280.0 35525.0 ;
      RECT  165.0 38420.0 2280.0 38485.0 ;
      RECT  165.0 34605.0 2280.0 34670.0 ;
      RECT  2875.0 34857.5 2690.0 34922.5 ;
      RECT  4035.0 34857.5 3850.0 34922.5 ;
      RECT  2832.5 34307.5 2657.5 34752.5 ;
      RECT  3917.5 34497.5 3032.5 34562.5 ;
      RECT  2965.0 34307.5 2800.0 34372.5 ;
      RECT  2965.0 34687.5 2800.0 34752.5 ;
      RECT  3032.5 34307.5 2897.5 34372.5 ;
      RECT  3032.5 34687.5 2897.5 34752.5 ;
      RECT  3032.5 34497.5 2897.5 34562.5 ;
      RECT  3032.5 34497.5 2897.5 34562.5 ;
      RECT  2832.5 34307.5 2767.5 34752.5 ;
      RECT  4015.0 34307.5 3850.0 34372.5 ;
      RECT  4015.0 34687.5 3850.0 34752.5 ;
      RECT  3917.5 34307.5 3782.5 34372.5 ;
      RECT  3917.5 34687.5 3782.5 34752.5 ;
      RECT  3917.5 34497.5 3782.5 34562.5 ;
      RECT  3917.5 34497.5 3782.5 34562.5 ;
      RECT  4047.5 34307.5 3982.5 34752.5 ;
      RECT  2942.5 34857.5 2807.5 34922.5 ;
      RECT  3917.5 34857.5 3782.5 34922.5 ;
      RECT  3475.0 34365.0 3340.0 34430.0 ;
      RECT  3475.0 34365.0 3340.0 34430.0 ;
      RECT  3440.0 34530.0 3375.0 34595.0 ;
      RECT  2722.5 34240.0 2657.5 34990.0 ;
      RECT  4067.5 34240.0 4002.5 34990.0 ;
      RECT  2875.0 35797.5 2690.0 35862.5 ;
      RECT  4035.0 35797.5 3850.0 35862.5 ;
      RECT  2877.5 35057.5 2657.5 35502.5 ;
      RECT  3702.5 35627.5 3207.5 35692.5 ;
      RECT  3010.0 35057.5 2845.0 35122.5 ;
      RECT  3010.0 35437.5 2845.0 35502.5 ;
      RECT  3175.0 35247.5 3010.0 35312.5 ;
      RECT  3175.0 35627.5 3010.0 35692.5 ;
      RECT  3077.5 35057.5 2942.5 35122.5 ;
      RECT  3077.5 35437.5 2942.5 35502.5 ;
      RECT  3077.5 35247.5 2942.5 35312.5 ;
      RECT  3077.5 35627.5 2942.5 35692.5 ;
      RECT  3207.5 35247.5 3142.5 35692.5 ;
      RECT  2877.5 35057.5 2812.5 35502.5 ;
      RECT  4000.0 35057.5 3835.0 35122.5 ;
      RECT  4000.0 35437.5 3835.0 35502.5 ;
      RECT  3835.0 35247.5 3670.0 35312.5 ;
      RECT  3835.0 35627.5 3670.0 35692.5 ;
      RECT  3902.5 35057.5 3767.5 35122.5 ;
      RECT  3902.5 35437.5 3767.5 35502.5 ;
      RECT  3902.5 35247.5 3767.5 35312.5 ;
      RECT  3902.5 35627.5 3767.5 35692.5 ;
      RECT  3702.5 35247.5 3637.5 35692.5 ;
      RECT  4032.5 35057.5 3967.5 35502.5 ;
      RECT  2942.5 35797.5 2807.5 35862.5 ;
      RECT  3917.5 35797.5 3782.5 35862.5 ;
      RECT  3490.0 35115.0 3355.0 35180.0 ;
      RECT  3490.0 35115.0 3355.0 35180.0 ;
      RECT  3455.0 35660.0 3390.0 35725.0 ;
      RECT  2722.5 34990.0 2657.5 35930.0 ;
      RECT  4067.5 34990.0 4002.5 35930.0 ;
      RECT  2875.0 37307.5 2690.0 37372.5 ;
      RECT  4035.0 37307.5 3850.0 37372.5 ;
      RECT  2877.5 35997.5 2657.5 37202.5 ;
      RECT  3702.5 36947.5 3207.5 37012.5 ;
      RECT  3010.0 35997.5 2845.0 36062.5 ;
      RECT  3010.0 36377.5 2845.0 36442.5 ;
      RECT  3010.0 36757.5 2845.0 36822.5 ;
      RECT  3010.0 37137.5 2845.0 37202.5 ;
      RECT  3175.0 36187.5 3010.0 36252.5 ;
      RECT  3175.0 36567.5 3010.0 36632.5 ;
      RECT  3175.0 36947.5 3010.0 37012.5 ;
      RECT  3077.5 35997.5 2942.5 36062.5 ;
      RECT  3077.5 36377.5 2942.5 36442.5 ;
      RECT  3077.5 36757.5 2942.5 36822.5 ;
      RECT  3077.5 37137.5 2942.5 37202.5 ;
      RECT  3077.5 36187.5 2942.5 36252.5 ;
      RECT  3077.5 36567.5 2942.5 36632.5 ;
      RECT  3077.5 36947.5 2942.5 37012.5 ;
      RECT  3207.5 36187.5 3142.5 37012.5 ;
      RECT  2877.5 35997.5 2812.5 37202.5 ;
      RECT  4000.0 35997.5 3835.0 36062.5 ;
      RECT  4000.0 36377.5 3835.0 36442.5 ;
      RECT  4000.0 36757.5 3835.0 36822.5 ;
      RECT  4000.0 37137.5 3835.0 37202.5 ;
      RECT  3835.0 36187.5 3670.0 36252.5 ;
      RECT  3835.0 36567.5 3670.0 36632.5 ;
      RECT  3835.0 36947.5 3670.0 37012.5 ;
      RECT  3902.5 35997.5 3767.5 36062.5 ;
      RECT  3902.5 36377.5 3767.5 36442.5 ;
      RECT  3902.5 36757.5 3767.5 36822.5 ;
      RECT  3902.5 37137.5 3767.5 37202.5 ;
      RECT  3902.5 36187.5 3767.5 36252.5 ;
      RECT  3902.5 36567.5 3767.5 36632.5 ;
      RECT  3902.5 36947.5 3767.5 37012.5 ;
      RECT  3702.5 36187.5 3637.5 37012.5 ;
      RECT  4032.5 35997.5 3967.5 37202.5 ;
      RECT  2942.5 37307.5 2807.5 37372.5 ;
      RECT  3917.5 37307.5 3782.5 37372.5 ;
      RECT  3490.0 36055.0 3355.0 36120.0 ;
      RECT  3490.0 36055.0 3355.0 36120.0 ;
      RECT  3455.0 36980.0 3390.0 37045.0 ;
      RECT  2722.5 35930.0 2657.5 37440.0 ;
      RECT  4067.5 35930.0 4002.5 37440.0 ;
      RECT  2875.0 39957.5 2690.0 40022.5 ;
      RECT  4035.0 39957.5 3850.0 40022.5 ;
      RECT  2877.5 37507.5 2657.5 39852.5 ;
      RECT  3702.5 39597.5 3207.5 39662.5 ;
      RECT  3010.0 37507.5 2845.0 37572.5 ;
      RECT  3010.0 37887.5 2845.0 37952.5 ;
      RECT  3010.0 38267.5 2845.0 38332.5 ;
      RECT  3010.0 38647.5 2845.0 38712.5 ;
      RECT  3010.0 39027.5 2845.0 39092.5 ;
      RECT  3010.0 39407.5 2845.0 39472.5 ;
      RECT  3010.0 39787.5 2845.0 39852.5 ;
      RECT  3175.0 37697.5 3010.0 37762.5 ;
      RECT  3175.0 38077.5 3010.0 38142.5 ;
      RECT  3175.0 38457.5 3010.0 38522.5 ;
      RECT  3175.0 38837.5 3010.0 38902.5 ;
      RECT  3175.0 39217.5 3010.0 39282.5 ;
      RECT  3175.0 39597.5 3010.0 39662.5 ;
      RECT  3077.5 37507.5 2942.5 37572.5 ;
      RECT  3077.5 37887.5 2942.5 37952.5 ;
      RECT  3077.5 38267.5 2942.5 38332.5 ;
      RECT  3077.5 38647.5 2942.5 38712.5 ;
      RECT  3077.5 39027.5 2942.5 39092.5 ;
      RECT  3077.5 39407.5 2942.5 39472.5 ;
      RECT  3077.5 39787.5 2942.5 39852.5 ;
      RECT  3077.5 37697.5 2942.5 37762.5 ;
      RECT  3077.5 38077.5 2942.5 38142.5 ;
      RECT  3077.5 38457.5 2942.5 38522.5 ;
      RECT  3077.5 38837.5 2942.5 38902.5 ;
      RECT  3077.5 39217.5 2942.5 39282.5 ;
      RECT  3077.5 39597.5 2942.5 39662.5 ;
      RECT  3207.5 37697.5 3142.5 39662.5 ;
      RECT  2877.5 37507.5 2812.5 39852.5 ;
      RECT  4000.0 37507.5 3835.0 37572.5 ;
      RECT  4000.0 37887.5 3835.0 37952.5 ;
      RECT  4000.0 38267.5 3835.0 38332.5 ;
      RECT  4000.0 38647.5 3835.0 38712.5 ;
      RECT  4000.0 39027.5 3835.0 39092.5 ;
      RECT  4000.0 39407.5 3835.0 39472.5 ;
      RECT  4000.0 39787.5 3835.0 39852.5 ;
      RECT  3835.0 37697.5 3670.0 37762.5 ;
      RECT  3835.0 38077.5 3670.0 38142.5 ;
      RECT  3835.0 38457.5 3670.0 38522.5 ;
      RECT  3835.0 38837.5 3670.0 38902.5 ;
      RECT  3835.0 39217.5 3670.0 39282.5 ;
      RECT  3835.0 39597.5 3670.0 39662.5 ;
      RECT  3902.5 37507.5 3767.5 37572.5 ;
      RECT  3902.5 37887.5 3767.5 37952.5 ;
      RECT  3902.5 38267.5 3767.5 38332.5 ;
      RECT  3902.5 38647.5 3767.5 38712.5 ;
      RECT  3902.5 39027.5 3767.5 39092.5 ;
      RECT  3902.5 39407.5 3767.5 39472.5 ;
      RECT  3902.5 39787.5 3767.5 39852.5 ;
      RECT  3902.5 37697.5 3767.5 37762.5 ;
      RECT  3902.5 38077.5 3767.5 38142.5 ;
      RECT  3902.5 38457.5 3767.5 38522.5 ;
      RECT  3902.5 38837.5 3767.5 38902.5 ;
      RECT  3902.5 39217.5 3767.5 39282.5 ;
      RECT  3902.5 39597.5 3767.5 39662.5 ;
      RECT  3702.5 37697.5 3637.5 39662.5 ;
      RECT  4032.5 37507.5 3967.5 39852.5 ;
      RECT  2942.5 39957.5 2807.5 40022.5 ;
      RECT  3917.5 39957.5 3782.5 40022.5 ;
      RECT  3490.0 37565.0 3355.0 37630.0 ;
      RECT  3490.0 37565.0 3355.0 37630.0 ;
      RECT  3455.0 39630.0 3390.0 39695.0 ;
      RECT  2722.5 37440.0 2657.5 40090.0 ;
      RECT  4067.5 37440.0 4002.5 40090.0 ;
      RECT  3872.5 43002.5 4067.5 43067.5 ;
      RECT  3032.5 43002.5 2657.5 43067.5 ;
      RECT  3032.5 43382.5 2657.5 43447.5 ;
      RECT  2875.0 43742.5 2690.0 43807.5 ;
      RECT  4035.0 43742.5 3850.0 43807.5 ;
      RECT  3032.5 43002.5 2897.5 43067.5 ;
      RECT  3032.5 43192.5 2897.5 43257.5 ;
      RECT  3032.5 43192.5 2897.5 43257.5 ;
      RECT  3032.5 43002.5 2897.5 43067.5 ;
      RECT  3032.5 43192.5 2897.5 43257.5 ;
      RECT  3032.5 43382.5 2897.5 43447.5 ;
      RECT  3032.5 43382.5 2897.5 43447.5 ;
      RECT  3032.5 43192.5 2897.5 43257.5 ;
      RECT  3032.5 43382.5 2897.5 43447.5 ;
      RECT  3032.5 43572.5 2897.5 43637.5 ;
      RECT  3032.5 43572.5 2897.5 43637.5 ;
      RECT  3032.5 43382.5 2897.5 43447.5 ;
      RECT  3872.5 43002.5 3737.5 43067.5 ;
      RECT  3872.5 43192.5 3737.5 43257.5 ;
      RECT  3872.5 43192.5 3737.5 43257.5 ;
      RECT  3872.5 43002.5 3737.5 43067.5 ;
      RECT  3872.5 43192.5 3737.5 43257.5 ;
      RECT  3872.5 43382.5 3737.5 43447.5 ;
      RECT  3872.5 43382.5 3737.5 43447.5 ;
      RECT  3872.5 43192.5 3737.5 43257.5 ;
      RECT  3872.5 43382.5 3737.5 43447.5 ;
      RECT  3872.5 43572.5 3737.5 43637.5 ;
      RECT  3872.5 43572.5 3737.5 43637.5 ;
      RECT  3872.5 43382.5 3737.5 43447.5 ;
      RECT  2942.5 43742.5 2807.5 43807.5 ;
      RECT  3917.5 43742.5 3782.5 43807.5 ;
      RECT  3660.0 43577.5 3595.0 43442.5 ;
      RECT  3520.0 43387.5 3455.0 43252.5 ;
      RECT  3380.0 43197.5 3315.0 43062.5 ;
      RECT  3032.5 43192.5 2897.5 43257.5 ;
      RECT  3032.5 43572.5 2897.5 43637.5 ;
      RECT  3872.5 43572.5 3737.5 43637.5 ;
      RECT  3415.0 43572.5 3280.0 43637.5 ;
      RECT  3380.0 43062.5 3315.0 43197.5 ;
      RECT  3520.0 43252.5 3455.0 43387.5 ;
      RECT  3660.0 43442.5 3595.0 43577.5 ;
      RECT  3415.0 43572.5 3280.0 43637.5 ;
      RECT  2722.5 42935.0 2657.5 43945.0 ;
      RECT  4067.5 42935.0 4002.5 43945.0 ;
      RECT  2875.0 44372.5 2690.0 44437.5 ;
      RECT  4035.0 44372.5 3850.0 44437.5 ;
      RECT  3917.5 44012.5 4067.5 44077.5 ;
      RECT  3032.5 44012.5 2657.5 44077.5 ;
      RECT  3917.5 44202.5 3032.5 44267.5 ;
      RECT  3032.5 44012.5 2897.5 44077.5 ;
      RECT  3032.5 44202.5 2897.5 44267.5 ;
      RECT  3032.5 44202.5 2897.5 44267.5 ;
      RECT  3032.5 44012.5 2897.5 44077.5 ;
      RECT  3917.5 44012.5 3782.5 44077.5 ;
      RECT  3917.5 44202.5 3782.5 44267.5 ;
      RECT  3917.5 44202.5 3782.5 44267.5 ;
      RECT  3917.5 44012.5 3782.5 44077.5 ;
      RECT  2942.5 44372.5 2807.5 44437.5 ;
      RECT  3917.5 44372.5 3782.5 44437.5 ;
      RECT  3475.0 44070.0 3340.0 44135.0 ;
      RECT  3475.0 44070.0 3340.0 44135.0 ;
      RECT  3440.0 44235.0 3375.0 44300.0 ;
      RECT  2722.5 43945.0 2657.5 44505.0 ;
      RECT  4067.5 43945.0 4002.5 44505.0 ;
      RECT  1462.5 43002.5 1312.5 43067.5 ;
      RECT  1462.5 43382.5 1312.5 43447.5 ;
      RECT  2280.0 43002.5 2722.5 43067.5 ;
      RECT  2505.0 43552.5 2690.0 43617.5 ;
      RECT  1345.0 43552.5 1530.0 43617.5 ;
      RECT  2280.0 43002.5 2415.0 43067.5 ;
      RECT  2280.0 43192.5 2415.0 43257.5 ;
      RECT  2280.0 43192.5 2415.0 43257.5 ;
      RECT  2280.0 43002.5 2415.0 43067.5 ;
      RECT  2280.0 43192.5 2415.0 43257.5 ;
      RECT  2280.0 43382.5 2415.0 43447.5 ;
      RECT  2280.0 43382.5 2415.0 43447.5 ;
      RECT  2280.0 43192.5 2415.0 43257.5 ;
      RECT  1462.5 43002.5 1597.5 43067.5 ;
      RECT  1462.5 43192.5 1597.5 43257.5 ;
      RECT  1462.5 43192.5 1597.5 43257.5 ;
      RECT  1462.5 43002.5 1597.5 43067.5 ;
      RECT  1462.5 43192.5 1597.5 43257.5 ;
      RECT  1462.5 43382.5 1597.5 43447.5 ;
      RECT  1462.5 43382.5 1597.5 43447.5 ;
      RECT  1462.5 43192.5 1597.5 43257.5 ;
      RECT  2437.5 43552.5 2572.5 43617.5 ;
      RECT  1462.5 43552.5 1597.5 43617.5 ;
      RECT  1682.5 43387.5 1747.5 43252.5 ;
      RECT  1897.5 43130.0 1962.5 42995.0 ;
      RECT  2280.0 43382.5 2415.0 43447.5 ;
      RECT  1497.5 43292.5 1562.5 43157.5 ;
      RECT  1897.5 43552.5 1962.5 43417.5 ;
      RECT  1897.5 42995.0 1962.5 43130.0 ;
      RECT  1682.5 43252.5 1747.5 43387.5 ;
      RECT  1897.5 43417.5 1962.5 43552.5 ;
      RECT  2657.5 42935.0 2722.5 43855.0 ;
      RECT  1312.5 42935.0 1377.5 43855.0 ;
      RECT  1507.5 44147.5 1312.5 44212.5 ;
      RECT  2347.5 44147.5 2722.5 44212.5 ;
      RECT  2347.5 44527.5 2722.5 44592.5 ;
      RECT  2505.0 44697.5 2690.0 44762.5 ;
      RECT  1345.0 44697.5 1530.0 44762.5 ;
      RECT  2347.5 44147.5 2482.5 44212.5 ;
      RECT  2347.5 44337.5 2482.5 44402.5 ;
      RECT  2347.5 44337.5 2482.5 44402.5 ;
      RECT  2347.5 44147.5 2482.5 44212.5 ;
      RECT  2347.5 44337.5 2482.5 44402.5 ;
      RECT  2347.5 44527.5 2482.5 44592.5 ;
      RECT  2347.5 44527.5 2482.5 44592.5 ;
      RECT  2347.5 44337.5 2482.5 44402.5 ;
      RECT  1507.5 44147.5 1642.5 44212.5 ;
      RECT  1507.5 44337.5 1642.5 44402.5 ;
      RECT  1507.5 44337.5 1642.5 44402.5 ;
      RECT  1507.5 44147.5 1642.5 44212.5 ;
      RECT  1507.5 44337.5 1642.5 44402.5 ;
      RECT  1507.5 44527.5 1642.5 44592.5 ;
      RECT  1507.5 44527.5 1642.5 44592.5 ;
      RECT  1507.5 44337.5 1642.5 44402.5 ;
      RECT  2437.5 44697.5 2572.5 44762.5 ;
      RECT  1462.5 44697.5 1597.5 44762.5 ;
      RECT  1737.5 44532.5 1802.5 44397.5 ;
      RECT  1952.5 44275.0 2017.5 44140.0 ;
      RECT  2347.5 44337.5 2482.5 44402.5 ;
      RECT  1507.5 44527.5 1642.5 44592.5 ;
      RECT  1952.5 44627.5 2017.5 44492.5 ;
      RECT  1952.5 44140.0 2017.5 44275.0 ;
      RECT  1737.5 44397.5 1802.5 44532.5 ;
      RECT  1952.5 44492.5 2017.5 44627.5 ;
      RECT  2657.5 44080.0 2722.5 45000.0 ;
      RECT  1312.5 44080.0 1377.5 45000.0 ;
      RECT  2505.0 45357.5 2690.0 45292.5 ;
      RECT  1345.0 45357.5 1530.0 45292.5 ;
      RECT  1462.5 45717.5 1312.5 45652.5 ;
      RECT  2347.5 45717.5 2722.5 45652.5 ;
      RECT  1462.5 45527.5 2347.5 45462.5 ;
      RECT  2347.5 45717.5 2482.5 45652.5 ;
      RECT  2347.5 45527.5 2482.5 45462.5 ;
      RECT  2347.5 45527.5 2482.5 45462.5 ;
      RECT  2347.5 45717.5 2482.5 45652.5 ;
      RECT  1462.5 45717.5 1597.5 45652.5 ;
      RECT  1462.5 45527.5 1597.5 45462.5 ;
      RECT  1462.5 45527.5 1597.5 45462.5 ;
      RECT  1462.5 45717.5 1597.5 45652.5 ;
      RECT  2437.5 45357.5 2572.5 45292.5 ;
      RECT  1462.5 45357.5 1597.5 45292.5 ;
      RECT  1905.0 45660.0 2040.0 45595.0 ;
      RECT  1905.0 45660.0 2040.0 45595.0 ;
      RECT  1940.0 45495.0 2005.0 45430.0 ;
      RECT  2657.5 45785.0 2722.5 45225.0 ;
      RECT  1312.5 45785.0 1377.5 45225.0 ;
      RECT  2505.0 45917.5 2690.0 45852.5 ;
      RECT  1345.0 45917.5 1530.0 45852.5 ;
      RECT  1462.5 46277.5 1312.5 46212.5 ;
      RECT  2347.5 46277.5 2722.5 46212.5 ;
      RECT  1462.5 46087.5 2347.5 46022.5 ;
      RECT  2347.5 46277.5 2482.5 46212.5 ;
      RECT  2347.5 46087.5 2482.5 46022.5 ;
      RECT  2347.5 46087.5 2482.5 46022.5 ;
      RECT  2347.5 46277.5 2482.5 46212.5 ;
      RECT  1462.5 46277.5 1597.5 46212.5 ;
      RECT  1462.5 46087.5 1597.5 46022.5 ;
      RECT  1462.5 46087.5 1597.5 46022.5 ;
      RECT  1462.5 46277.5 1597.5 46212.5 ;
      RECT  2437.5 45917.5 2572.5 45852.5 ;
      RECT  1462.5 45917.5 1597.5 45852.5 ;
      RECT  1905.0 46220.0 2040.0 46155.0 ;
      RECT  1905.0 46220.0 2040.0 46155.0 ;
      RECT  1940.0 46055.0 2005.0 45990.0 ;
      RECT  2657.5 46345.0 2722.5 45785.0 ;
      RECT  1312.5 46345.0 1377.5 45785.0 ;
      RECT  1182.5 43562.5 1377.5 43627.5 ;
      RECT  342.5 43562.5 -32.5 43627.5 ;
      RECT  342.5 43942.5 -32.5 44007.5 ;
      RECT  185.0 44302.5 8.881784197e-13 44367.5 ;
      RECT  1345.0 44302.5 1160.0 44367.5 ;
      RECT  342.5 43562.5 207.5 43627.5 ;
      RECT  342.5 43752.5 207.5 43817.5 ;
      RECT  342.5 43752.5 207.5 43817.5 ;
      RECT  342.5 43562.5 207.5 43627.5 ;
      RECT  342.5 43752.5 207.5 43817.5 ;
      RECT  342.5 43942.5 207.5 44007.5 ;
      RECT  342.5 43942.5 207.5 44007.5 ;
      RECT  342.5 43752.5 207.5 43817.5 ;
      RECT  342.5 43942.5 207.5 44007.5 ;
      RECT  342.5 44132.5 207.5 44197.5 ;
      RECT  342.5 44132.5 207.5 44197.5 ;
      RECT  342.5 43942.5 207.5 44007.5 ;
      RECT  1182.5 43562.5 1047.5 43627.5 ;
      RECT  1182.5 43752.5 1047.5 43817.5 ;
      RECT  1182.5 43752.5 1047.5 43817.5 ;
      RECT  1182.5 43562.5 1047.5 43627.5 ;
      RECT  1182.5 43752.5 1047.5 43817.5 ;
      RECT  1182.5 43942.5 1047.5 44007.5 ;
      RECT  1182.5 43942.5 1047.5 44007.5 ;
      RECT  1182.5 43752.5 1047.5 43817.5 ;
      RECT  1182.5 43942.5 1047.5 44007.5 ;
      RECT  1182.5 44132.5 1047.5 44197.5 ;
      RECT  1182.5 44132.5 1047.5 44197.5 ;
      RECT  1182.5 43942.5 1047.5 44007.5 ;
      RECT  252.5 44302.5 117.5 44367.5 ;
      RECT  1227.5 44302.5 1092.5 44367.5 ;
      RECT  970.0 44137.5 905.0 44002.5 ;
      RECT  830.0 43947.5 765.0 43812.5 ;
      RECT  690.0 43757.5 625.0 43622.5 ;
      RECT  342.5 43752.5 207.5 43817.5 ;
      RECT  342.5 44132.5 207.5 44197.5 ;
      RECT  1182.5 44132.5 1047.5 44197.5 ;
      RECT  725.0 44132.5 590.0 44197.5 ;
      RECT  690.0 43622.5 625.0 43757.5 ;
      RECT  830.0 43812.5 765.0 43947.5 ;
      RECT  970.0 44002.5 905.0 44137.5 ;
      RECT  725.0 44132.5 590.0 44197.5 ;
      RECT  32.5 43495.0 -32.5 44505.0 ;
      RECT  1377.5 43495.0 1312.5 44505.0 ;
      RECT  185.0 44932.5 8.881784197e-13 44997.5 ;
      RECT  1345.0 44932.5 1160.0 44997.5 ;
      RECT  1227.5 44572.5 1377.5 44637.5 ;
      RECT  342.5 44572.5 -32.5 44637.5 ;
      RECT  1227.5 44762.5 342.5 44827.5 ;
      RECT  342.5 44572.5 207.5 44637.5 ;
      RECT  342.5 44762.5 207.5 44827.5 ;
      RECT  342.5 44762.5 207.5 44827.5 ;
      RECT  342.5 44572.5 207.5 44637.5 ;
      RECT  1227.5 44572.5 1092.5 44637.5 ;
      RECT  1227.5 44762.5 1092.5 44827.5 ;
      RECT  1227.5 44762.5 1092.5 44827.5 ;
      RECT  1227.5 44572.5 1092.5 44637.5 ;
      RECT  252.5 44932.5 117.5 44997.5 ;
      RECT  1227.5 44932.5 1092.5 44997.5 ;
      RECT  785.0 44630.0 650.0 44695.0 ;
      RECT  785.0 44630.0 650.0 44695.0 ;
      RECT  750.0 44795.0 685.0 44860.0 ;
      RECT  32.5 44505.0 -32.5 45065.0 ;
      RECT  1377.5 44505.0 1312.5 45065.0 ;
      RECT  185.0 45492.5 8.881784197e-13 45557.5 ;
      RECT  1345.0 45492.5 1160.0 45557.5 ;
      RECT  1227.5 45132.5 1377.5 45197.5 ;
      RECT  342.5 45132.5 -32.5 45197.5 ;
      RECT  1227.5 45322.5 342.5 45387.5 ;
      RECT  342.5 45132.5 207.5 45197.5 ;
      RECT  342.5 45322.5 207.5 45387.5 ;
      RECT  342.5 45322.5 207.5 45387.5 ;
      RECT  342.5 45132.5 207.5 45197.5 ;
      RECT  1227.5 45132.5 1092.5 45197.5 ;
      RECT  1227.5 45322.5 1092.5 45387.5 ;
      RECT  1227.5 45322.5 1092.5 45387.5 ;
      RECT  1227.5 45132.5 1092.5 45197.5 ;
      RECT  252.5 45492.5 117.5 45557.5 ;
      RECT  1227.5 45492.5 1092.5 45557.5 ;
      RECT  785.0 45190.0 650.0 45255.0 ;
      RECT  785.0 45190.0 650.0 45255.0 ;
      RECT  750.0 45355.0 685.0 45420.0 ;
      RECT  32.5 45065.0 -32.5 45625.0 ;
      RECT  1377.5 45065.0 1312.5 45625.0 ;
      RECT  185.0 46052.5 8.881784197e-13 46117.5 ;
      RECT  1345.0 46052.5 1160.0 46117.5 ;
      RECT  1227.5 45692.5 1377.5 45757.5 ;
      RECT  342.5 45692.5 -32.5 45757.5 ;
      RECT  1227.5 45882.5 342.5 45947.5 ;
      RECT  342.5 45692.5 207.5 45757.5 ;
      RECT  342.5 45882.5 207.5 45947.5 ;
      RECT  342.5 45882.5 207.5 45947.5 ;
      RECT  342.5 45692.5 207.5 45757.5 ;
      RECT  1227.5 45692.5 1092.5 45757.5 ;
      RECT  1227.5 45882.5 1092.5 45947.5 ;
      RECT  1227.5 45882.5 1092.5 45947.5 ;
      RECT  1227.5 45692.5 1092.5 45757.5 ;
      RECT  252.5 46052.5 117.5 46117.5 ;
      RECT  1227.5 46052.5 1092.5 46117.5 ;
      RECT  785.0 45750.0 650.0 45815.0 ;
      RECT  785.0 45750.0 650.0 45815.0 ;
      RECT  750.0 45915.0 685.0 45980.0 ;
      RECT  32.5 45625.0 -32.5 46185.0 ;
      RECT  1377.5 45625.0 1312.5 46185.0 ;
      RECT  1377.5 53227.5 1312.5 84245.0 ;
      RECT  1312.5 48917.5 1025.0 48982.5 ;
      RECT  1312.5 51327.5 1025.0 51392.5 ;
      RECT  1312.5 51607.5 1025.0 51672.5 ;
      RECT  1312.5 54017.5 1025.0 54082.5 ;
      RECT  1312.5 54297.5 1025.0 54362.5 ;
      RECT  1312.5 56707.5 1025.0 56772.5 ;
      RECT  1312.5 56987.5 1025.0 57052.5 ;
      RECT  1312.5 59397.5 1025.0 59462.5 ;
      RECT  1312.5 59677.5 1025.0 59742.5 ;
      RECT  1312.5 62087.5 1025.0 62152.5 ;
      RECT  1312.5 62367.5 1025.0 62432.5 ;
      RECT  1312.5 64777.5 1025.0 64842.5 ;
      RECT  1312.5 65057.5 1025.0 65122.5 ;
      RECT  1312.5 67467.5 1025.0 67532.5 ;
      RECT  1312.5 67747.5 1025.0 67812.5 ;
      RECT  1312.5 70157.5 1025.0 70222.5 ;
      RECT  1312.5 70437.5 1025.0 70502.5 ;
      RECT  1312.5 72847.5 1025.0 72912.5 ;
      RECT  1312.5 73127.5 1025.0 73192.5 ;
      RECT  1312.5 75537.5 1025.0 75602.5 ;
      RECT  1312.5 75817.5 1025.0 75882.5 ;
      RECT  1312.5 78227.5 1025.0 78292.5 ;
      RECT  1312.5 78507.5 1025.0 78572.5 ;
      RECT  1312.5 80917.5 1025.0 80982.5 ;
      RECT  1312.5 81197.5 1025.0 81262.5 ;
      RECT  1312.5 83607.5 1025.0 83672.5 ;
      RECT  1377.5 46872.5 935.0 46937.5 ;
      RECT  935.0 46872.5 230.0 46937.5 ;
      RECT  20.0 50122.5 935.0 50187.5 ;
      RECT  20.0 52812.5 935.0 52877.5 ;
      RECT  20.0 55502.5 935.0 55567.5 ;
      RECT  20.0 58192.5 935.0 58257.5 ;
      RECT  20.0 60882.5 935.0 60947.5 ;
      RECT  20.0 63572.5 935.0 63637.5 ;
      RECT  20.0 66262.5 935.0 66327.5 ;
      RECT  20.0 68952.5 935.0 69017.5 ;
      RECT  20.0 71642.5 935.0 71707.5 ;
      RECT  20.0 74332.5 935.0 74397.5 ;
      RECT  20.0 77022.5 935.0 77087.5 ;
      RECT  20.0 79712.5 935.0 79777.5 ;
      RECT  20.0 82402.5 935.0 82467.5 ;
      RECT  20.0 47432.5 935.0 47497.5 ;
      RECT  2005.0 48445.0 1940.0 49145.0 ;
      RECT  2005.0 48637.5 1940.0 48702.5 ;
      RECT  2005.0 48445.0 1940.0 48670.0 ;
      RECT  1972.5 48637.5 1025.0 48702.5 ;
      RECT  2690.0 48507.5 2465.0 48572.5 ;
      RECT  2430.0 47637.5 2365.0 47702.5 ;
      RECT  2005.0 47637.5 1940.0 47702.5 ;
      RECT  2430.0 47670.0 2365.0 48317.5 ;
      RECT  2397.5 47637.5 1972.5 47702.5 ;
      RECT  2005.0 47340.0 1940.0 47670.0 ;
      RECT  1972.5 47637.5 1172.5 47702.5 ;
      RECT  1172.5 47040.0 750.0 47105.0 ;
      RECT  2040.0 47275.0 1905.0 47340.0 ;
      RECT  2005.0 49145.0 1940.0 49350.0 ;
      RECT  2505.0 47037.5 2690.0 46972.5 ;
      RECT  1345.0 47037.5 1530.0 46972.5 ;
      RECT  1462.5 47397.5 1312.5 47332.5 ;
      RECT  2347.5 47397.5 2722.5 47332.5 ;
      RECT  1462.5 47207.5 2347.5 47142.5 ;
      RECT  2347.5 47397.5 2482.5 47332.5 ;
      RECT  2347.5 47207.5 2482.5 47142.5 ;
      RECT  2347.5 47207.5 2482.5 47142.5 ;
      RECT  2347.5 47397.5 2482.5 47332.5 ;
      RECT  1462.5 47397.5 1597.5 47332.5 ;
      RECT  1462.5 47207.5 1597.5 47142.5 ;
      RECT  1462.5 47207.5 1597.5 47142.5 ;
      RECT  1462.5 47397.5 1597.5 47332.5 ;
      RECT  2437.5 47037.5 2572.5 46972.5 ;
      RECT  1462.5 47037.5 1597.5 46972.5 ;
      RECT  1905.0 47340.0 2040.0 47275.0 ;
      RECT  1905.0 47340.0 2040.0 47275.0 ;
      RECT  1940.0 47175.0 2005.0 47110.0 ;
      RECT  2657.5 47465.0 2722.5 46905.0 ;
      RECT  1312.5 47465.0 1377.5 46905.0 ;
      RECT  2330.0 48317.5 2465.0 48382.5 ;
      RECT  2330.0 48507.5 2465.0 48572.5 ;
      RECT  2330.0 48507.5 2465.0 48572.5 ;
      RECT  2330.0 48317.5 2465.0 48382.5 ;
      RECT  1312.5 53162.5 1377.5 53227.5 ;
      RECT  4002.5 53162.5 4067.5 53227.5 ;
      RECT  1312.5 53065.0 1377.5 53195.0 ;
      RECT  1345.0 53162.5 4035.0 53227.5 ;
      RECT  4002.5 53065.0 4067.5 53195.0 ;
      RECT  2875.0 49572.5 2690.0 49637.5 ;
      RECT  4035.0 49572.5 3850.0 49637.5 ;
      RECT  3917.5 49212.5 4067.5 49277.5 ;
      RECT  3032.5 49212.5 2657.5 49277.5 ;
      RECT  3917.5 49402.5 3032.5 49467.5 ;
      RECT  3032.5 49212.5 2897.5 49277.5 ;
      RECT  3032.5 49402.5 2897.5 49467.5 ;
      RECT  3032.5 49402.5 2897.5 49467.5 ;
      RECT  3032.5 49212.5 2897.5 49277.5 ;
      RECT  3917.5 49212.5 3782.5 49277.5 ;
      RECT  3917.5 49402.5 3782.5 49467.5 ;
      RECT  3917.5 49402.5 3782.5 49467.5 ;
      RECT  3917.5 49212.5 3782.5 49277.5 ;
      RECT  2942.5 49572.5 2807.5 49637.5 ;
      RECT  3917.5 49572.5 3782.5 49637.5 ;
      RECT  3475.0 49270.0 3340.0 49335.0 ;
      RECT  3475.0 49270.0 3340.0 49335.0 ;
      RECT  3440.0 49435.0 3375.0 49500.0 ;
      RECT  2722.5 49145.0 2657.5 49705.0 ;
      RECT  4067.5 49145.0 4002.5 49705.0 ;
      RECT  2875.0 50132.5 2690.0 50197.5 ;
      RECT  4035.0 50132.5 3850.0 50197.5 ;
      RECT  3917.5 49772.5 4067.5 49837.5 ;
      RECT  3032.5 49772.5 2657.5 49837.5 ;
      RECT  3917.5 49962.5 3032.5 50027.5 ;
      RECT  3032.5 49772.5 2897.5 49837.5 ;
      RECT  3032.5 49962.5 2897.5 50027.5 ;
      RECT  3032.5 49962.5 2897.5 50027.5 ;
      RECT  3032.5 49772.5 2897.5 49837.5 ;
      RECT  3917.5 49772.5 3782.5 49837.5 ;
      RECT  3917.5 49962.5 3782.5 50027.5 ;
      RECT  3917.5 49962.5 3782.5 50027.5 ;
      RECT  3917.5 49772.5 3782.5 49837.5 ;
      RECT  2942.5 50132.5 2807.5 50197.5 ;
      RECT  3917.5 50132.5 3782.5 50197.5 ;
      RECT  3475.0 49830.0 3340.0 49895.0 ;
      RECT  3475.0 49830.0 3340.0 49895.0 ;
      RECT  3440.0 49995.0 3375.0 50060.0 ;
      RECT  2722.5 49705.0 2657.5 50265.0 ;
      RECT  4067.5 49705.0 4002.5 50265.0 ;
      RECT  3340.0 49830.0 3475.0 49895.0 ;
      RECT  2875.0 50692.5 2690.0 50757.5 ;
      RECT  4035.0 50692.5 3850.0 50757.5 ;
      RECT  3917.5 50332.5 4067.5 50397.5 ;
      RECT  3032.5 50332.5 2657.5 50397.5 ;
      RECT  3917.5 50522.5 3032.5 50587.5 ;
      RECT  3032.5 50332.5 2897.5 50397.5 ;
      RECT  3032.5 50522.5 2897.5 50587.5 ;
      RECT  3032.5 50522.5 2897.5 50587.5 ;
      RECT  3032.5 50332.5 2897.5 50397.5 ;
      RECT  3917.5 50332.5 3782.5 50397.5 ;
      RECT  3917.5 50522.5 3782.5 50587.5 ;
      RECT  3917.5 50522.5 3782.5 50587.5 ;
      RECT  3917.5 50332.5 3782.5 50397.5 ;
      RECT  2942.5 50692.5 2807.5 50757.5 ;
      RECT  3917.5 50692.5 3782.5 50757.5 ;
      RECT  3475.0 50390.0 3340.0 50455.0 ;
      RECT  3475.0 50390.0 3340.0 50455.0 ;
      RECT  3440.0 50555.0 3375.0 50620.0 ;
      RECT  2722.5 50265.0 2657.5 50825.0 ;
      RECT  4067.5 50265.0 4002.5 50825.0 ;
      RECT  3340.0 50390.0 3475.0 50455.0 ;
      RECT  2875.0 51252.5 2690.0 51317.5 ;
      RECT  4035.0 51252.5 3850.0 51317.5 ;
      RECT  3917.5 50892.5 4067.5 50957.5 ;
      RECT  3032.5 50892.5 2657.5 50957.5 ;
      RECT  3917.5 51082.5 3032.5 51147.5 ;
      RECT  3032.5 50892.5 2897.5 50957.5 ;
      RECT  3032.5 51082.5 2897.5 51147.5 ;
      RECT  3032.5 51082.5 2897.5 51147.5 ;
      RECT  3032.5 50892.5 2897.5 50957.5 ;
      RECT  3917.5 50892.5 3782.5 50957.5 ;
      RECT  3917.5 51082.5 3782.5 51147.5 ;
      RECT  3917.5 51082.5 3782.5 51147.5 ;
      RECT  3917.5 50892.5 3782.5 50957.5 ;
      RECT  2942.5 51252.5 2807.5 51317.5 ;
      RECT  3917.5 51252.5 3782.5 51317.5 ;
      RECT  3475.0 50950.0 3340.0 51015.0 ;
      RECT  3475.0 50950.0 3340.0 51015.0 ;
      RECT  3440.0 51115.0 3375.0 51180.0 ;
      RECT  2722.5 50825.0 2657.5 51385.0 ;
      RECT  4067.5 50825.0 4002.5 51385.0 ;
      RECT  3340.0 50950.0 3475.0 51015.0 ;
      RECT  2875.0 51812.5 2690.0 51877.5 ;
      RECT  4035.0 51812.5 3850.0 51877.5 ;
      RECT  3917.5 51452.5 4067.5 51517.5 ;
      RECT  3032.5 51452.5 2657.5 51517.5 ;
      RECT  3917.5 51642.5 3032.5 51707.5 ;
      RECT  3032.5 51452.5 2897.5 51517.5 ;
      RECT  3032.5 51642.5 2897.5 51707.5 ;
      RECT  3032.5 51642.5 2897.5 51707.5 ;
      RECT  3032.5 51452.5 2897.5 51517.5 ;
      RECT  3917.5 51452.5 3782.5 51517.5 ;
      RECT  3917.5 51642.5 3782.5 51707.5 ;
      RECT  3917.5 51642.5 3782.5 51707.5 ;
      RECT  3917.5 51452.5 3782.5 51517.5 ;
      RECT  2942.5 51812.5 2807.5 51877.5 ;
      RECT  3917.5 51812.5 3782.5 51877.5 ;
      RECT  3475.0 51510.0 3340.0 51575.0 ;
      RECT  3475.0 51510.0 3340.0 51575.0 ;
      RECT  3440.0 51675.0 3375.0 51740.0 ;
      RECT  2722.5 51385.0 2657.5 51945.0 ;
      RECT  4067.5 51385.0 4002.5 51945.0 ;
      RECT  3340.0 51510.0 3475.0 51575.0 ;
      RECT  2875.0 52372.5 2690.0 52437.5 ;
      RECT  4035.0 52372.5 3850.0 52437.5 ;
      RECT  3917.5 52012.5 4067.5 52077.5 ;
      RECT  3032.5 52012.5 2657.5 52077.5 ;
      RECT  3917.5 52202.5 3032.5 52267.5 ;
      RECT  3032.5 52012.5 2897.5 52077.5 ;
      RECT  3032.5 52202.5 2897.5 52267.5 ;
      RECT  3032.5 52202.5 2897.5 52267.5 ;
      RECT  3032.5 52012.5 2897.5 52077.5 ;
      RECT  3917.5 52012.5 3782.5 52077.5 ;
      RECT  3917.5 52202.5 3782.5 52267.5 ;
      RECT  3917.5 52202.5 3782.5 52267.5 ;
      RECT  3917.5 52012.5 3782.5 52077.5 ;
      RECT  2942.5 52372.5 2807.5 52437.5 ;
      RECT  3917.5 52372.5 3782.5 52437.5 ;
      RECT  3475.0 52070.0 3340.0 52135.0 ;
      RECT  3475.0 52070.0 3340.0 52135.0 ;
      RECT  3440.0 52235.0 3375.0 52300.0 ;
      RECT  2722.5 51945.0 2657.5 52505.0 ;
      RECT  4067.5 51945.0 4002.5 52505.0 ;
      RECT  3340.0 52070.0 3475.0 52135.0 ;
      RECT  2875.0 52932.5 2690.0 52997.5 ;
      RECT  4035.0 52932.5 3850.0 52997.5 ;
      RECT  3917.5 52572.5 4067.5 52637.5 ;
      RECT  3032.5 52572.5 2657.5 52637.5 ;
      RECT  3917.5 52762.5 3032.5 52827.5 ;
      RECT  3032.5 52572.5 2897.5 52637.5 ;
      RECT  3032.5 52762.5 2897.5 52827.5 ;
      RECT  3032.5 52762.5 2897.5 52827.5 ;
      RECT  3032.5 52572.5 2897.5 52637.5 ;
      RECT  3917.5 52572.5 3782.5 52637.5 ;
      RECT  3917.5 52762.5 3782.5 52827.5 ;
      RECT  3917.5 52762.5 3782.5 52827.5 ;
      RECT  3917.5 52572.5 3782.5 52637.5 ;
      RECT  2942.5 52932.5 2807.5 52997.5 ;
      RECT  3917.5 52932.5 3782.5 52997.5 ;
      RECT  3475.0 52630.0 3340.0 52695.0 ;
      RECT  3475.0 52630.0 3340.0 52695.0 ;
      RECT  3440.0 52795.0 3375.0 52860.0 ;
      RECT  2722.5 52505.0 2657.5 53065.0 ;
      RECT  4067.5 52505.0 4002.5 53065.0 ;
      RECT  3340.0 52630.0 3475.0 52695.0 ;
      RECT  2505.0 52077.5 2690.0 52012.5 ;
      RECT  1345.0 52077.5 1530.0 52012.5 ;
      RECT  1462.5 52437.5 1312.5 52372.5 ;
      RECT  2347.5 52437.5 2722.5 52372.5 ;
      RECT  1462.5 52247.5 2347.5 52182.5 ;
      RECT  2347.5 52437.5 2482.5 52372.5 ;
      RECT  2347.5 52247.5 2482.5 52182.5 ;
      RECT  2347.5 52247.5 2482.5 52182.5 ;
      RECT  2347.5 52437.5 2482.5 52372.5 ;
      RECT  1462.5 52437.5 1597.5 52372.5 ;
      RECT  1462.5 52247.5 1597.5 52182.5 ;
      RECT  1462.5 52247.5 1597.5 52182.5 ;
      RECT  1462.5 52437.5 1597.5 52372.5 ;
      RECT  2437.5 52077.5 2572.5 52012.5 ;
      RECT  1462.5 52077.5 1597.5 52012.5 ;
      RECT  1905.0 52380.0 2040.0 52315.0 ;
      RECT  1905.0 52380.0 2040.0 52315.0 ;
      RECT  1940.0 52215.0 2005.0 52150.0 ;
      RECT  2657.5 52505.0 2722.5 51945.0 ;
      RECT  1312.5 52505.0 1377.5 51945.0 ;
      RECT  1905.0 52315.0 2040.0 52380.0 ;
      RECT  2505.0 51517.5 2690.0 51452.5 ;
      RECT  1345.0 51517.5 1530.0 51452.5 ;
      RECT  1462.5 51877.5 1312.5 51812.5 ;
      RECT  2347.5 51877.5 2722.5 51812.5 ;
      RECT  1462.5 51687.5 2347.5 51622.5 ;
      RECT  2347.5 51877.5 2482.5 51812.5 ;
      RECT  2347.5 51687.5 2482.5 51622.5 ;
      RECT  2347.5 51687.5 2482.5 51622.5 ;
      RECT  2347.5 51877.5 2482.5 51812.5 ;
      RECT  1462.5 51877.5 1597.5 51812.5 ;
      RECT  1462.5 51687.5 1597.5 51622.5 ;
      RECT  1462.5 51687.5 1597.5 51622.5 ;
      RECT  1462.5 51877.5 1597.5 51812.5 ;
      RECT  2437.5 51517.5 2572.5 51452.5 ;
      RECT  1462.5 51517.5 1597.5 51452.5 ;
      RECT  1905.0 51820.0 2040.0 51755.0 ;
      RECT  1905.0 51820.0 2040.0 51755.0 ;
      RECT  1940.0 51655.0 2005.0 51590.0 ;
      RECT  2657.5 51945.0 2722.5 51385.0 ;
      RECT  1312.5 51945.0 1377.5 51385.0 ;
      RECT  1905.0 51755.0 2040.0 51820.0 ;
      RECT  2505.0 50957.5 2690.0 50892.5 ;
      RECT  1345.0 50957.5 1530.0 50892.5 ;
      RECT  1462.5 51317.5 1312.5 51252.5 ;
      RECT  2347.5 51317.5 2722.5 51252.5 ;
      RECT  1462.5 51127.5 2347.5 51062.5 ;
      RECT  2347.5 51317.5 2482.5 51252.5 ;
      RECT  2347.5 51127.5 2482.5 51062.5 ;
      RECT  2347.5 51127.5 2482.5 51062.5 ;
      RECT  2347.5 51317.5 2482.5 51252.5 ;
      RECT  1462.5 51317.5 1597.5 51252.5 ;
      RECT  1462.5 51127.5 1597.5 51062.5 ;
      RECT  1462.5 51127.5 1597.5 51062.5 ;
      RECT  1462.5 51317.5 1597.5 51252.5 ;
      RECT  2437.5 50957.5 2572.5 50892.5 ;
      RECT  1462.5 50957.5 1597.5 50892.5 ;
      RECT  1905.0 51260.0 2040.0 51195.0 ;
      RECT  1905.0 51260.0 2040.0 51195.0 ;
      RECT  1940.0 51095.0 2005.0 51030.0 ;
      RECT  2657.5 51385.0 2722.5 50825.0 ;
      RECT  1312.5 51385.0 1377.5 50825.0 ;
      RECT  1905.0 51195.0 2040.0 51260.0 ;
      RECT  2505.0 50397.5 2690.0 50332.5 ;
      RECT  1345.0 50397.5 1530.0 50332.5 ;
      RECT  1462.5 50757.5 1312.5 50692.5 ;
      RECT  2347.5 50757.5 2722.5 50692.5 ;
      RECT  1462.5 50567.5 2347.5 50502.5 ;
      RECT  2347.5 50757.5 2482.5 50692.5 ;
      RECT  2347.5 50567.5 2482.5 50502.5 ;
      RECT  2347.5 50567.5 2482.5 50502.5 ;
      RECT  2347.5 50757.5 2482.5 50692.5 ;
      RECT  1462.5 50757.5 1597.5 50692.5 ;
      RECT  1462.5 50567.5 1597.5 50502.5 ;
      RECT  1462.5 50567.5 1597.5 50502.5 ;
      RECT  1462.5 50757.5 1597.5 50692.5 ;
      RECT  2437.5 50397.5 2572.5 50332.5 ;
      RECT  1462.5 50397.5 1597.5 50332.5 ;
      RECT  1905.0 50700.0 2040.0 50635.0 ;
      RECT  1905.0 50700.0 2040.0 50635.0 ;
      RECT  1940.0 50535.0 2005.0 50470.0 ;
      RECT  2657.5 50825.0 2722.5 50265.0 ;
      RECT  1312.5 50825.0 1377.5 50265.0 ;
      RECT  1905.0 50635.0 2040.0 50700.0 ;
      RECT  2505.0 49837.5 2690.0 49772.5 ;
      RECT  1345.0 49837.5 1530.0 49772.5 ;
      RECT  1462.5 50197.5 1312.5 50132.5 ;
      RECT  2347.5 50197.5 2722.5 50132.5 ;
      RECT  1462.5 50007.5 2347.5 49942.5 ;
      RECT  2347.5 50197.5 2482.5 50132.5 ;
      RECT  2347.5 50007.5 2482.5 49942.5 ;
      RECT  2347.5 50007.5 2482.5 49942.5 ;
      RECT  2347.5 50197.5 2482.5 50132.5 ;
      RECT  1462.5 50197.5 1597.5 50132.5 ;
      RECT  1462.5 50007.5 1597.5 49942.5 ;
      RECT  1462.5 50007.5 1597.5 49942.5 ;
      RECT  1462.5 50197.5 1597.5 50132.5 ;
      RECT  2437.5 49837.5 2572.5 49772.5 ;
      RECT  1462.5 49837.5 1597.5 49772.5 ;
      RECT  1905.0 50140.0 2040.0 50075.0 ;
      RECT  1905.0 50140.0 2040.0 50075.0 ;
      RECT  1940.0 49975.0 2005.0 49910.0 ;
      RECT  2657.5 50265.0 2722.5 49705.0 ;
      RECT  1312.5 50265.0 1377.5 49705.0 ;
      RECT  1905.0 50075.0 2040.0 50140.0 ;
      RECT  2505.0 49277.5 2690.0 49212.5 ;
      RECT  1345.0 49277.5 1530.0 49212.5 ;
      RECT  1462.5 49637.5 1312.5 49572.5 ;
      RECT  2347.5 49637.5 2722.5 49572.5 ;
      RECT  1462.5 49447.5 2347.5 49382.5 ;
      RECT  2347.5 49637.5 2482.5 49572.5 ;
      RECT  2347.5 49447.5 2482.5 49382.5 ;
      RECT  2347.5 49447.5 2482.5 49382.5 ;
      RECT  2347.5 49637.5 2482.5 49572.5 ;
      RECT  1462.5 49637.5 1597.5 49572.5 ;
      RECT  1462.5 49447.5 1597.5 49382.5 ;
      RECT  1462.5 49447.5 1597.5 49382.5 ;
      RECT  1462.5 49637.5 1597.5 49572.5 ;
      RECT  2437.5 49277.5 2572.5 49212.5 ;
      RECT  1462.5 49277.5 1597.5 49212.5 ;
      RECT  1905.0 49580.0 2040.0 49515.0 ;
      RECT  1905.0 49580.0 2040.0 49515.0 ;
      RECT  1940.0 49415.0 2005.0 49350.0 ;
      RECT  2657.5 49705.0 2722.5 49145.0 ;
      RECT  1312.5 49705.0 1377.5 49145.0 ;
      RECT  1905.0 49515.0 2040.0 49580.0 ;
      RECT  3340.0 49435.0 3475.0 49500.0 ;
      RECT  3340.0 51115.0 3475.0 51180.0 ;
      RECT  3340.0 52795.0 3475.0 52860.0 ;
      RECT  1905.0 51030.0 2040.0 51095.0 ;
      RECT  3340.0 49270.0 3475.0 49335.0 ;
      RECT  1940.0 49145.0 2005.0 49350.0 ;
      RECT  2657.5 49145.0 2722.5 53065.0 ;
      RECT  1312.5 49145.0 1377.5 53065.0 ;
      RECT  4002.5 49145.0 4067.5 53065.0 ;
      RECT  935.0 48810.0 225.0 47465.0 ;
      RECT  935.0 48810.0 230.0 50155.0 ;
      RECT  935.0 51500.0 230.0 50155.0 ;
      RECT  935.0 51500.0 230.0 52845.0 ;
      RECT  935.0 54190.0 230.0 52845.0 ;
      RECT  935.0 54190.0 230.0 55535.0 ;
      RECT  935.0 56880.0 230.0 55535.0 ;
      RECT  935.0 56880.0 230.0 58225.0 ;
      RECT  935.0 59570.0 230.0 58225.0 ;
      RECT  935.0 59570.0 230.0 60915.0 ;
      RECT  935.0 62260.0 230.0 60915.0 ;
      RECT  935.0 62260.0 230.0 63605.0 ;
      RECT  935.0 64950.0 230.0 63605.0 ;
      RECT  935.0 64950.0 230.0 66295.0 ;
      RECT  935.0 67640.0 230.0 66295.0 ;
      RECT  935.0 67640.0 230.0 68985.0 ;
      RECT  935.0 70330.0 230.0 68985.0 ;
      RECT  935.0 70330.0 230.0 71675.0 ;
      RECT  935.0 73020.0 230.0 71675.0 ;
      RECT  935.0 73020.0 230.0 74365.0 ;
      RECT  935.0 75710.0 230.0 74365.0 ;
      RECT  935.0 75710.0 230.0 77055.0 ;
      RECT  935.0 78400.0 230.0 77055.0 ;
      RECT  935.0 78400.0 230.0 79745.0 ;
      RECT  935.0 81090.0 230.0 79745.0 ;
      RECT  935.0 81090.0 230.0 82435.0 ;
      RECT  935.0 83780.0 230.0 82435.0 ;
      RECT  1025.0 48917.5 140.0 48982.5 ;
      RECT  1025.0 51327.5 140.0 51392.5 ;
      RECT  1025.0 51607.5 140.0 51672.5 ;
      RECT  1025.0 54017.5 140.0 54082.5 ;
      RECT  1025.0 54297.5 140.0 54362.5 ;
      RECT  1025.0 56707.5 140.0 56772.5 ;
      RECT  1025.0 56987.5 140.0 57052.5 ;
      RECT  1025.0 59397.5 140.0 59462.5 ;
      RECT  1025.0 59677.5 140.0 59742.5 ;
      RECT  1025.0 62087.5 140.0 62152.5 ;
      RECT  1025.0 62367.5 140.0 62432.5 ;
      RECT  1025.0 64777.5 140.0 64842.5 ;
      RECT  1025.0 65057.5 140.0 65122.5 ;
      RECT  1025.0 67467.5 140.0 67532.5 ;
      RECT  1025.0 67747.5 140.0 67812.5 ;
      RECT  1025.0 70157.5 140.0 70222.5 ;
      RECT  1025.0 70437.5 140.0 70502.5 ;
      RECT  1025.0 72847.5 140.0 72912.5 ;
      RECT  1025.0 73127.5 140.0 73192.5 ;
      RECT  1025.0 75537.5 140.0 75602.5 ;
      RECT  1025.0 75817.5 140.0 75882.5 ;
      RECT  1025.0 78227.5 140.0 78292.5 ;
      RECT  1025.0 78507.5 140.0 78572.5 ;
      RECT  1025.0 80917.5 140.0 80982.5 ;
      RECT  1025.0 81197.5 140.0 81262.5 ;
      RECT  1025.0 83607.5 140.0 83672.5 ;
      RECT  1025.0 50122.5 140.0 50187.5 ;
      RECT  1025.0 52812.5 140.0 52877.5 ;
      RECT  1025.0 55502.5 140.0 55567.5 ;
      RECT  1025.0 58192.5 140.0 58257.5 ;
      RECT  1025.0 60882.5 140.0 60947.5 ;
      RECT  1025.0 63572.5 140.0 63637.5 ;
      RECT  1025.0 66262.5 140.0 66327.5 ;
      RECT  1025.0 68952.5 140.0 69017.5 ;
      RECT  1025.0 71642.5 140.0 71707.5 ;
      RECT  1025.0 74332.5 140.0 74397.5 ;
      RECT  1025.0 77022.5 140.0 77087.5 ;
      RECT  1025.0 79712.5 140.0 79777.5 ;
      RECT  1025.0 82402.5 140.0 82467.5 ;
      RECT  1025.0 48777.5 140.0 48842.5 ;
      RECT  1025.0 51467.5 140.0 51532.5 ;
      RECT  1025.0 54157.5 140.0 54222.5 ;
      RECT  1025.0 56847.5 140.0 56912.5 ;
      RECT  1025.0 59537.5 140.0 59602.5 ;
      RECT  1025.0 62227.5 140.0 62292.5 ;
      RECT  1025.0 64917.5 140.0 64982.5 ;
      RECT  1025.0 67607.5 140.0 67672.5 ;
      RECT  1025.0 70297.5 140.0 70362.5 ;
      RECT  1025.0 72987.5 140.0 73052.5 ;
      RECT  1025.0 75677.5 140.0 75742.5 ;
      RECT  1025.0 78367.5 140.0 78432.5 ;
      RECT  1025.0 81057.5 140.0 81122.5 ;
      RECT  1025.0 83747.5 140.0 83812.5 ;
      RECT  1345.0 48882.5 1280.0 49017.5 ;
      RECT  1345.0 51292.5 1280.0 51427.5 ;
      RECT  1345.0 51572.5 1280.0 51707.5 ;
      RECT  1345.0 53982.5 1280.0 54117.5 ;
      RECT  1345.0 54262.5 1280.0 54397.5 ;
      RECT  1345.0 56672.5 1280.0 56807.5 ;
      RECT  1345.0 56952.5 1280.0 57087.5 ;
      RECT  1345.0 59362.5 1280.0 59497.5 ;
      RECT  1345.0 59642.5 1280.0 59777.5 ;
      RECT  1345.0 62052.5 1280.0 62187.5 ;
      RECT  1345.0 62332.5 1280.0 62467.5 ;
      RECT  1345.0 64742.5 1280.0 64877.5 ;
      RECT  1345.0 65022.5 1280.0 65157.5 ;
      RECT  1345.0 67432.5 1280.0 67567.5 ;
      RECT  1345.0 67712.5 1280.0 67847.5 ;
      RECT  1345.0 70122.5 1280.0 70257.5 ;
      RECT  1345.0 70402.5 1280.0 70537.5 ;
      RECT  1345.0 72812.5 1280.0 72947.5 ;
      RECT  1345.0 73092.5 1280.0 73227.5 ;
      RECT  1345.0 75502.5 1280.0 75637.5 ;
      RECT  1345.0 75782.5 1280.0 75917.5 ;
      RECT  1345.0 78192.5 1280.0 78327.5 ;
      RECT  1345.0 78472.5 1280.0 78607.5 ;
      RECT  1345.0 80882.5 1280.0 81017.5 ;
      RECT  1345.0 81162.5 1280.0 81297.5 ;
      RECT  1345.0 83572.5 1280.0 83707.5 ;
      RECT  1342.5 49145.0 1277.5 49280.0 ;
      RECT  1377.5 46770.0 1312.5 46905.0 ;
      RECT  867.5 46872.5 1002.5 46937.5 ;
      RECT  162.5 46872.5 297.5 46937.5 ;
      RECT  2005.0 48377.5 1940.0 48512.5 ;
      RECT  1105.0 47637.5 1240.0 47702.5 ;
      RECT  1105.0 47040.0 1240.0 47105.0 ;
      RECT  682.5 47040.0 817.5 47105.0 ;
      RECT  3475.0 46345.0 3410.0 49270.0 ;
      RECT  2005.0 46345.0 1940.0 47110.0 ;
      RECT  20.0 46345.0 -45.0 83867.5 ;
      RECT  2722.5 46345.0 2657.5 49145.0 ;
      RECT  1377.5 46345.0 1312.5 46905.0 ;
      RECT  4067.5 46345.0 4002.5 49145.0 ;
      RECT  3455.0 41192.5 3390.0 41057.5 ;
      RECT  3455.0 37112.5 3390.0 36977.5 ;
      RECT  2517.5 34545.0 2452.5 34410.0 ;
      RECT  1962.5 41192.5 1897.5 41057.5 ;
      RECT  1747.5 41602.5 1682.5 41467.5 ;
      RECT  2017.5 44140.0 1952.5 44005.0 ;
      RECT  1802.5 44397.5 1737.5 44262.5 ;
      RECT  3380.0 42627.5 3315.0 42492.5 ;
      RECT  3520.0 42422.5 3455.0 42287.5 ;
      RECT  3660.0 41807.5 3595.0 41672.5 ;
      RECT  690.0 42627.5 625.0 42492.5 ;
      RECT  830.0 41807.5 765.0 41672.5 ;
      RECT  970.0 42012.5 905.0 41877.5 ;
      RECT  1997.5 43822.5 1862.5 43887.5 ;
      RECT  2052.5 44967.5 1917.5 45032.5 ;
      RECT  785.0 46152.5 650.0 46217.5 ;
      RECT  2040.0 45192.5 1905.0 45257.5 ;
      RECT  4067.5 41397.5 4002.5 41262.5 ;
      RECT  2722.5 42217.5 2657.5 42082.5 ;
      RECT  1377.5 41397.5 1312.5 41262.5 ;
      RECT  32.5 42217.5 -32.5 42082.5 ;
      RECT  3475.0 34240.0 3340.0 34430.0 ;
      RECT  2722.5 34240.0 2657.5 34305.0 ;
      RECT  4067.5 34240.0 4002.5 34305.0 ;
      RECT  4417.5 42117.5 4282.5 42182.5 ;
   LAYER  metal2 ;
      RECT  16682.5 45020.0 16752.5 45225.0 ;
      RECT  16477.5 45980.0 16547.5 46185.0 ;
      RECT  16067.5 43650.0 16137.5 43855.0 ;
      RECT  15862.5 44795.0 15932.5 45000.0 ;
      RECT  16272.5 42355.0 16342.5 42560.0 ;
      RECT  15657.5 40920.0 15727.5 41125.0 ;
      RECT  4035.0 42115.0 4350.0 42185.0 ;
      RECT  15242.5 41125.0 15312.5 41330.0 ;
      RECT  15657.5 35.0 15727.5 207987.5 ;
      RECT  15862.5 35.0 15932.5 207987.5 ;
      RECT  16067.5 35.0 16137.5 207987.5 ;
      RECT  16272.5 35.0 16342.5 207987.5 ;
      RECT  16477.5 35.0 16547.5 207987.5 ;
      RECT  16682.5 35.0 16752.5 207987.5 ;
      RECT  12642.5 35.0 12712.5 34100.0 ;
      RECT  12847.5 35.0 12917.5 34100.0 ;
      RECT  13052.5 35.0 13122.5 34100.0 ;
      RECT  13257.5 35.0 13327.5 34100.0 ;
      RECT  13462.5 35.0 13532.5 34100.0 ;
      RECT  13667.5 35.0 13737.5 34100.0 ;
      RECT  13872.5 35.0 13942.5 34100.0 ;
      RECT  14077.5 35.0 14147.5 34100.0 ;
      RECT  14282.5 35.0 14352.5 34100.0 ;
      RECT  14487.5 35.0 14557.5 34100.0 ;
      RECT  14692.5 35.0 14762.5 34100.0 ;
      RECT  17345.0 206415.0 17415.0 206820.0 ;
      RECT  17680.0 206415.0 17750.0 206820.0 ;
      RECT  18050.0 206415.0 18120.0 206820.0 ;
      RECT  18385.0 206415.0 18455.0 206820.0 ;
      RECT  18755.0 206415.0 18825.0 206820.0 ;
      RECT  19090.0 206415.0 19160.0 206820.0 ;
      RECT  19460.0 206415.0 19530.0 206820.0 ;
      RECT  19795.0 206415.0 19865.0 206820.0 ;
      RECT  20165.0 206415.0 20235.0 206820.0 ;
      RECT  20500.0 206415.0 20570.0 206820.0 ;
      RECT  20870.0 206415.0 20940.0 206820.0 ;
      RECT  21205.0 206415.0 21275.0 206820.0 ;
      RECT  21575.0 206415.0 21645.0 206820.0 ;
      RECT  21910.0 206415.0 21980.0 206820.0 ;
      RECT  22280.0 206415.0 22350.0 206820.0 ;
      RECT  22615.0 206415.0 22685.0 206820.0 ;
      RECT  22985.0 206415.0 23055.0 206820.0 ;
      RECT  23320.0 206415.0 23390.0 206820.0 ;
      RECT  23690.0 206415.0 23760.0 206820.0 ;
      RECT  24025.0 206415.0 24095.0 206820.0 ;
      RECT  24395.0 206415.0 24465.0 206820.0 ;
      RECT  24730.0 206415.0 24800.0 206820.0 ;
      RECT  25100.0 206415.0 25170.0 206820.0 ;
      RECT  25435.0 206415.0 25505.0 206820.0 ;
      RECT  25805.0 206415.0 25875.0 206820.0 ;
      RECT  26140.0 206415.0 26210.0 206820.0 ;
      RECT  26510.0 206415.0 26580.0 206820.0 ;
      RECT  26845.0 206415.0 26915.0 206820.0 ;
      RECT  27215.0 206415.0 27285.0 206820.0 ;
      RECT  27550.0 206415.0 27620.0 206820.0 ;
      RECT  27920.0 206415.0 27990.0 206820.0 ;
      RECT  28255.0 206415.0 28325.0 206820.0 ;
      RECT  28625.0 206415.0 28695.0 206820.0 ;
      RECT  28960.0 206415.0 29030.0 206820.0 ;
      RECT  29330.0 206415.0 29400.0 206820.0 ;
      RECT  29665.0 206415.0 29735.0 206820.0 ;
      RECT  30035.0 206415.0 30105.0 206820.0 ;
      RECT  30370.0 206415.0 30440.0 206820.0 ;
      RECT  30740.0 206415.0 30810.0 206820.0 ;
      RECT  31075.0 206415.0 31145.0 206820.0 ;
      RECT  31445.0 206415.0 31515.0 206820.0 ;
      RECT  31780.0 206415.0 31850.0 206820.0 ;
      RECT  32150.0 206415.0 32220.0 206820.0 ;
      RECT  32485.0 206415.0 32555.0 206820.0 ;
      RECT  32855.0 206415.0 32925.0 206820.0 ;
      RECT  33190.0 206415.0 33260.0 206820.0 ;
      RECT  33560.0 206415.0 33630.0 206820.0 ;
      RECT  33895.0 206415.0 33965.0 206820.0 ;
      RECT  34265.0 206415.0 34335.0 206820.0 ;
      RECT  34600.0 206415.0 34670.0 206820.0 ;
      RECT  34970.0 206415.0 35040.0 206820.0 ;
      RECT  35305.0 206415.0 35375.0 206820.0 ;
      RECT  35675.0 206415.0 35745.0 206820.0 ;
      RECT  36010.0 206415.0 36080.0 206820.0 ;
      RECT  36380.0 206415.0 36450.0 206820.0 ;
      RECT  36715.0 206415.0 36785.0 206820.0 ;
      RECT  37085.0 206415.0 37155.0 206820.0 ;
      RECT  37420.0 206415.0 37490.0 206820.0 ;
      RECT  37790.0 206415.0 37860.0 206820.0 ;
      RECT  38125.0 206415.0 38195.0 206820.0 ;
      RECT  38495.0 206415.0 38565.0 206820.0 ;
      RECT  38830.0 206415.0 38900.0 206820.0 ;
      RECT  39200.0 206415.0 39270.0 206820.0 ;
      RECT  39535.0 206415.0 39605.0 206820.0 ;
      RECT  39905.0 206415.0 39975.0 206820.0 ;
      RECT  40240.0 206415.0 40310.0 206820.0 ;
      RECT  40610.0 206415.0 40680.0 206820.0 ;
      RECT  40945.0 206415.0 41015.0 206820.0 ;
      RECT  41315.0 206415.0 41385.0 206820.0 ;
      RECT  41650.0 206415.0 41720.0 206820.0 ;
      RECT  42020.0 206415.0 42090.0 206820.0 ;
      RECT  42355.0 206415.0 42425.0 206820.0 ;
      RECT  42725.0 206415.0 42795.0 206820.0 ;
      RECT  43060.0 206415.0 43130.0 206820.0 ;
      RECT  43430.0 206415.0 43500.0 206820.0 ;
      RECT  43765.0 206415.0 43835.0 206820.0 ;
      RECT  44135.0 206415.0 44205.0 206820.0 ;
      RECT  44470.0 206415.0 44540.0 206820.0 ;
      RECT  44840.0 206415.0 44910.0 206820.0 ;
      RECT  45175.0 206415.0 45245.0 206820.0 ;
      RECT  45545.0 206415.0 45615.0 206820.0 ;
      RECT  45880.0 206415.0 45950.0 206820.0 ;
      RECT  46250.0 206415.0 46320.0 206820.0 ;
      RECT  46585.0 206415.0 46655.0 206820.0 ;
      RECT  46955.0 206415.0 47025.0 206820.0 ;
      RECT  47290.0 206415.0 47360.0 206820.0 ;
      RECT  47660.0 206415.0 47730.0 206820.0 ;
      RECT  47995.0 206415.0 48065.0 206820.0 ;
      RECT  48365.0 206415.0 48435.0 206820.0 ;
      RECT  48700.0 206415.0 48770.0 206820.0 ;
      RECT  49070.0 206415.0 49140.0 206820.0 ;
      RECT  49405.0 206415.0 49475.0 206820.0 ;
      RECT  49775.0 206415.0 49845.0 206820.0 ;
      RECT  50110.0 206415.0 50180.0 206820.0 ;
      RECT  50480.0 206415.0 50550.0 206820.0 ;
      RECT  50815.0 206415.0 50885.0 206820.0 ;
      RECT  51185.0 206415.0 51255.0 206820.0 ;
      RECT  51520.0 206415.0 51590.0 206820.0 ;
      RECT  51890.0 206415.0 51960.0 206820.0 ;
      RECT  52225.0 206415.0 52295.0 206820.0 ;
      RECT  52595.0 206415.0 52665.0 206820.0 ;
      RECT  52930.0 206415.0 53000.0 206820.0 ;
      RECT  53300.0 206415.0 53370.0 206820.0 ;
      RECT  53635.0 206415.0 53705.0 206820.0 ;
      RECT  54005.0 206415.0 54075.0 206820.0 ;
      RECT  54340.0 206415.0 54410.0 206820.0 ;
      RECT  54710.0 206415.0 54780.0 206820.0 ;
      RECT  55045.0 206415.0 55115.0 206820.0 ;
      RECT  55415.0 206415.0 55485.0 206820.0 ;
      RECT  55750.0 206415.0 55820.0 206820.0 ;
      RECT  56120.0 206415.0 56190.0 206820.0 ;
      RECT  56455.0 206415.0 56525.0 206820.0 ;
      RECT  56825.0 206415.0 56895.0 206820.0 ;
      RECT  57160.0 206415.0 57230.0 206820.0 ;
      RECT  57530.0 206415.0 57600.0 206820.0 ;
      RECT  57865.0 206415.0 57935.0 206820.0 ;
      RECT  58235.0 206415.0 58305.0 206820.0 ;
      RECT  58570.0 206415.0 58640.0 206820.0 ;
      RECT  58940.0 206415.0 59010.0 206820.0 ;
      RECT  59275.0 206415.0 59345.0 206820.0 ;
      RECT  59645.0 206415.0 59715.0 206820.0 ;
      RECT  59980.0 206415.0 60050.0 206820.0 ;
      RECT  60350.0 206415.0 60420.0 206820.0 ;
      RECT  60685.0 206415.0 60755.0 206820.0 ;
      RECT  61055.0 206415.0 61125.0 206820.0 ;
      RECT  61390.0 206415.0 61460.0 206820.0 ;
      RECT  61760.0 206415.0 61830.0 206820.0 ;
      RECT  62095.0 206415.0 62165.0 206820.0 ;
      RECT  62465.0 206415.0 62535.0 206820.0 ;
      RECT  62800.0 206415.0 62870.0 206820.0 ;
      RECT  63170.0 206415.0 63240.0 206820.0 ;
      RECT  63505.0 206415.0 63575.0 206820.0 ;
      RECT  63875.0 206415.0 63945.0 206820.0 ;
      RECT  64210.0 206415.0 64280.0 206820.0 ;
      RECT  64580.0 206415.0 64650.0 206820.0 ;
      RECT  64915.0 206415.0 64985.0 206820.0 ;
      RECT  65285.0 206415.0 65355.0 206820.0 ;
      RECT  65620.0 206415.0 65690.0 206820.0 ;
      RECT  65990.0 206415.0 66060.0 206820.0 ;
      RECT  66325.0 206415.0 66395.0 206820.0 ;
      RECT  66695.0 206415.0 66765.0 206820.0 ;
      RECT  67030.0 206415.0 67100.0 206820.0 ;
      RECT  67400.0 206415.0 67470.0 206820.0 ;
      RECT  67735.0 206415.0 67805.0 206820.0 ;
      RECT  68105.0 206415.0 68175.0 206820.0 ;
      RECT  68440.0 206415.0 68510.0 206820.0 ;
      RECT  68810.0 206415.0 68880.0 206820.0 ;
      RECT  69145.0 206415.0 69215.0 206820.0 ;
      RECT  69515.0 206415.0 69585.0 206820.0 ;
      RECT  69850.0 206415.0 69920.0 206820.0 ;
      RECT  70220.0 206415.0 70290.0 206820.0 ;
      RECT  70555.0 206415.0 70625.0 206820.0 ;
      RECT  70925.0 206415.0 70995.0 206820.0 ;
      RECT  71260.0 206415.0 71330.0 206820.0 ;
      RECT  71630.0 206415.0 71700.0 206820.0 ;
      RECT  71965.0 206415.0 72035.0 206820.0 ;
      RECT  72335.0 206415.0 72405.0 206820.0 ;
      RECT  72670.0 206415.0 72740.0 206820.0 ;
      RECT  73040.0 206415.0 73110.0 206820.0 ;
      RECT  73375.0 206415.0 73445.0 206820.0 ;
      RECT  73745.0 206415.0 73815.0 206820.0 ;
      RECT  74080.0 206415.0 74150.0 206820.0 ;
      RECT  74450.0 206415.0 74520.0 206820.0 ;
      RECT  74785.0 206415.0 74855.0 206820.0 ;
      RECT  75155.0 206415.0 75225.0 206820.0 ;
      RECT  75490.0 206415.0 75560.0 206820.0 ;
      RECT  75860.0 206415.0 75930.0 206820.0 ;
      RECT  76195.0 206415.0 76265.0 206820.0 ;
      RECT  76565.0 206415.0 76635.0 206820.0 ;
      RECT  76900.0 206415.0 76970.0 206820.0 ;
      RECT  77270.0 206415.0 77340.0 206820.0 ;
      RECT  77605.0 206415.0 77675.0 206820.0 ;
      RECT  77975.0 206415.0 78045.0 206820.0 ;
      RECT  78310.0 206415.0 78380.0 206820.0 ;
      RECT  78680.0 206415.0 78750.0 206820.0 ;
      RECT  79015.0 206415.0 79085.0 206820.0 ;
      RECT  79385.0 206415.0 79455.0 206820.0 ;
      RECT  79720.0 206415.0 79790.0 206820.0 ;
      RECT  80090.0 206415.0 80160.0 206820.0 ;
      RECT  80425.0 206415.0 80495.0 206820.0 ;
      RECT  80795.0 206415.0 80865.0 206820.0 ;
      RECT  81130.0 206415.0 81200.0 206820.0 ;
      RECT  81500.0 206415.0 81570.0 206820.0 ;
      RECT  81835.0 206415.0 81905.0 206820.0 ;
      RECT  82205.0 206415.0 82275.0 206820.0 ;
      RECT  82540.0 206415.0 82610.0 206820.0 ;
      RECT  82910.0 206415.0 82980.0 206820.0 ;
      RECT  83245.0 206415.0 83315.0 206820.0 ;
      RECT  83615.0 206415.0 83685.0 206820.0 ;
      RECT  83950.0 206415.0 84020.0 206820.0 ;
      RECT  84320.0 206415.0 84390.0 206820.0 ;
      RECT  84655.0 206415.0 84725.0 206820.0 ;
      RECT  85025.0 206415.0 85095.0 206820.0 ;
      RECT  85360.0 206415.0 85430.0 206820.0 ;
      RECT  85730.0 206415.0 85800.0 206820.0 ;
      RECT  86065.0 206415.0 86135.0 206820.0 ;
      RECT  86435.0 206415.0 86505.0 206820.0 ;
      RECT  86770.0 206415.0 86840.0 206820.0 ;
      RECT  87140.0 206415.0 87210.0 206820.0 ;
      RECT  87475.0 206415.0 87545.0 206820.0 ;
      RECT  87845.0 206415.0 87915.0 206820.0 ;
      RECT  88180.0 206415.0 88250.0 206820.0 ;
      RECT  88550.0 206415.0 88620.0 206820.0 ;
      RECT  88885.0 206415.0 88955.0 206820.0 ;
      RECT  89255.0 206415.0 89325.0 206820.0 ;
      RECT  89590.0 206415.0 89660.0 206820.0 ;
      RECT  89960.0 206415.0 90030.0 206820.0 ;
      RECT  90295.0 206415.0 90365.0 206820.0 ;
      RECT  90665.0 206415.0 90735.0 206820.0 ;
      RECT  91000.0 206415.0 91070.0 206820.0 ;
      RECT  91370.0 206415.0 91440.0 206820.0 ;
      RECT  91705.0 206415.0 91775.0 206820.0 ;
      RECT  92075.0 206415.0 92145.0 206820.0 ;
      RECT  92410.0 206415.0 92480.0 206820.0 ;
      RECT  92780.0 206415.0 92850.0 206820.0 ;
      RECT  93115.0 206415.0 93185.0 206820.0 ;
      RECT  93485.0 206415.0 93555.0 206820.0 ;
      RECT  93820.0 206415.0 93890.0 206820.0 ;
      RECT  94190.0 206415.0 94260.0 206820.0 ;
      RECT  94525.0 206415.0 94595.0 206820.0 ;
      RECT  94895.0 206415.0 94965.0 206820.0 ;
      RECT  95230.0 206415.0 95300.0 206820.0 ;
      RECT  95600.0 206415.0 95670.0 206820.0 ;
      RECT  95935.0 206415.0 96005.0 206820.0 ;
      RECT  96305.0 206415.0 96375.0 206820.0 ;
      RECT  96640.0 206415.0 96710.0 206820.0 ;
      RECT  97010.0 206415.0 97080.0 206820.0 ;
      RECT  97345.0 206415.0 97415.0 206820.0 ;
      RECT  97715.0 206415.0 97785.0 206820.0 ;
      RECT  98050.0 206415.0 98120.0 206820.0 ;
      RECT  98420.0 206415.0 98490.0 206820.0 ;
      RECT  98755.0 206415.0 98825.0 206820.0 ;
      RECT  99125.0 206415.0 99195.0 206820.0 ;
      RECT  99460.0 206415.0 99530.0 206820.0 ;
      RECT  99830.0 206415.0 99900.0 206820.0 ;
      RECT  100165.0 206415.0 100235.0 206820.0 ;
      RECT  100535.0 206415.0 100605.0 206820.0 ;
      RECT  100870.0 206415.0 100940.0 206820.0 ;
      RECT  101240.0 206415.0 101310.0 206820.0 ;
      RECT  101575.0 206415.0 101645.0 206820.0 ;
      RECT  101945.0 206415.0 102015.0 206820.0 ;
      RECT  102280.0 206415.0 102350.0 206820.0 ;
      RECT  102650.0 206415.0 102720.0 206820.0 ;
      RECT  102985.0 206415.0 103055.0 206820.0 ;
      RECT  103355.0 206415.0 103425.0 206820.0 ;
      RECT  103690.0 206415.0 103760.0 206820.0 ;
      RECT  104060.0 206415.0 104130.0 206820.0 ;
      RECT  104395.0 206415.0 104465.0 206820.0 ;
      RECT  104765.0 206415.0 104835.0 206820.0 ;
      RECT  105100.0 206415.0 105170.0 206820.0 ;
      RECT  105470.0 206415.0 105540.0 206820.0 ;
      RECT  105805.0 206415.0 105875.0 206820.0 ;
      RECT  106175.0 206415.0 106245.0 206820.0 ;
      RECT  106510.0 206415.0 106580.0 206820.0 ;
      RECT  106880.0 206415.0 106950.0 206820.0 ;
      RECT  107215.0 206415.0 107285.0 206820.0 ;
      RECT  17512.5 12605.0 17582.5 12675.0 ;
      RECT  17337.5 12605.0 17547.5 12675.0 ;
      RECT  17512.5 12640.0 17582.5 12780.0 ;
      RECT  20332.5 12605.0 20402.5 12675.0 ;
      RECT  20157.5 12605.0 20367.5 12675.0 ;
      RECT  20332.5 12640.0 20402.5 12780.0 ;
      RECT  23152.5 12605.0 23222.5 12675.0 ;
      RECT  22977.5 12605.0 23187.5 12675.0 ;
      RECT  23152.5 12640.0 23222.5 12780.0 ;
      RECT  25972.5 12605.0 26042.5 12675.0 ;
      RECT  25797.5 12605.0 26007.5 12675.0 ;
      RECT  25972.5 12640.0 26042.5 12780.0 ;
      RECT  28792.5 12605.0 28862.5 12675.0 ;
      RECT  28617.5 12605.0 28827.5 12675.0 ;
      RECT  28792.5 12640.0 28862.5 12780.0 ;
      RECT  31612.5 12605.0 31682.5 12675.0 ;
      RECT  31437.5 12605.0 31647.5 12675.0 ;
      RECT  31612.5 12640.0 31682.5 12780.0 ;
      RECT  34432.5 12605.0 34502.5 12675.0 ;
      RECT  34257.5 12605.0 34467.5 12675.0 ;
      RECT  34432.5 12640.0 34502.5 12780.0 ;
      RECT  37252.5 12605.0 37322.5 12675.0 ;
      RECT  37077.5 12605.0 37287.5 12675.0 ;
      RECT  37252.5 12640.0 37322.5 12780.0 ;
      RECT  40072.5 12605.0 40142.5 12675.0 ;
      RECT  39897.5 12605.0 40107.5 12675.0 ;
      RECT  40072.5 12640.0 40142.5 12780.0 ;
      RECT  42892.5 12605.0 42962.5 12675.0 ;
      RECT  42717.5 12605.0 42927.5 12675.0 ;
      RECT  42892.5 12640.0 42962.5 12780.0 ;
      RECT  45712.5 12605.0 45782.5 12675.0 ;
      RECT  45537.5 12605.0 45747.5 12675.0 ;
      RECT  45712.5 12640.0 45782.5 12780.0 ;
      RECT  48532.5 12605.0 48602.5 12675.0 ;
      RECT  48357.5 12605.0 48567.5 12675.0 ;
      RECT  48532.5 12640.0 48602.5 12780.0 ;
      RECT  51352.5 12605.0 51422.5 12675.0 ;
      RECT  51177.5 12605.0 51387.5 12675.0 ;
      RECT  51352.5 12640.0 51422.5 12780.0 ;
      RECT  54172.5 12605.0 54242.5 12675.0 ;
      RECT  53997.5 12605.0 54207.5 12675.0 ;
      RECT  54172.5 12640.0 54242.5 12780.0 ;
      RECT  56992.5 12605.0 57062.5 12675.0 ;
      RECT  56817.5 12605.0 57027.5 12675.0 ;
      RECT  56992.5 12640.0 57062.5 12780.0 ;
      RECT  59812.5 12605.0 59882.5 12675.0 ;
      RECT  59637.5 12605.0 59847.5 12675.0 ;
      RECT  59812.5 12640.0 59882.5 12780.0 ;
      RECT  62632.5 12605.0 62702.5 12675.0 ;
      RECT  62457.5 12605.0 62667.5 12675.0 ;
      RECT  62632.5 12640.0 62702.5 12780.0 ;
      RECT  65452.5 12605.0 65522.5 12675.0 ;
      RECT  65277.5 12605.0 65487.5 12675.0 ;
      RECT  65452.5 12640.0 65522.5 12780.0 ;
      RECT  68272.5 12605.0 68342.5 12675.0 ;
      RECT  68097.5 12605.0 68307.5 12675.0 ;
      RECT  68272.5 12640.0 68342.5 12780.0 ;
      RECT  71092.5 12605.0 71162.5 12675.0 ;
      RECT  70917.5 12605.0 71127.5 12675.0 ;
      RECT  71092.5 12640.0 71162.5 12780.0 ;
      RECT  73912.5 12605.0 73982.5 12675.0 ;
      RECT  73737.5 12605.0 73947.5 12675.0 ;
      RECT  73912.5 12640.0 73982.5 12780.0 ;
      RECT  76732.5 12605.0 76802.5 12675.0 ;
      RECT  76557.5 12605.0 76767.5 12675.0 ;
      RECT  76732.5 12640.0 76802.5 12780.0 ;
      RECT  79552.5 12605.0 79622.5 12675.0 ;
      RECT  79377.5 12605.0 79587.5 12675.0 ;
      RECT  79552.5 12640.0 79622.5 12780.0 ;
      RECT  82372.5 12605.0 82442.5 12675.0 ;
      RECT  82197.5 12605.0 82407.5 12675.0 ;
      RECT  82372.5 12640.0 82442.5 12780.0 ;
      RECT  85192.5 12605.0 85262.5 12675.0 ;
      RECT  85017.5 12605.0 85227.5 12675.0 ;
      RECT  85192.5 12640.0 85262.5 12780.0 ;
      RECT  88012.5 12605.0 88082.5 12675.0 ;
      RECT  87837.5 12605.0 88047.5 12675.0 ;
      RECT  88012.5 12640.0 88082.5 12780.0 ;
      RECT  90832.5 12605.0 90902.5 12675.0 ;
      RECT  90657.5 12605.0 90867.5 12675.0 ;
      RECT  90832.5 12640.0 90902.5 12780.0 ;
      RECT  93652.5 12605.0 93722.5 12675.0 ;
      RECT  93477.5 12605.0 93687.5 12675.0 ;
      RECT  93652.5 12640.0 93722.5 12780.0 ;
      RECT  96472.5 12605.0 96542.5 12675.0 ;
      RECT  96297.5 12605.0 96507.5 12675.0 ;
      RECT  96472.5 12640.0 96542.5 12780.0 ;
      RECT  99292.5 12605.0 99362.5 12675.0 ;
      RECT  99117.5 12605.0 99327.5 12675.0 ;
      RECT  99292.5 12640.0 99362.5 12780.0 ;
      RECT  102112.5 12605.0 102182.5 12675.0 ;
      RECT  101937.5 12605.0 102147.5 12675.0 ;
      RECT  102112.5 12640.0 102182.5 12780.0 ;
      RECT  104932.5 12605.0 105002.5 12675.0 ;
      RECT  104757.5 12605.0 104967.5 12675.0 ;
      RECT  104932.5 12640.0 105002.5 12780.0 ;
      RECT  9220.0 206260.0 9290.0 206465.0 ;
      RECT  17195.0 34100.0 17900.0 35445.0 ;
      RECT  17195.0 36790.0 17900.0 35445.0 ;
      RECT  17195.0 36790.0 17900.0 38135.0 ;
      RECT  17195.0 39480.0 17900.0 38135.0 ;
      RECT  17195.0 39480.0 17900.0 40825.0 ;
      RECT  17195.0 42170.0 17900.0 40825.0 ;
      RECT  17195.0 42170.0 17900.0 43515.0 ;
      RECT  17195.0 44860.0 17900.0 43515.0 ;
      RECT  17195.0 44860.0 17900.0 46205.0 ;
      RECT  17195.0 47550.0 17900.0 46205.0 ;
      RECT  17195.0 47550.0 17900.0 48895.0 ;
      RECT  17195.0 50240.0 17900.0 48895.0 ;
      RECT  17195.0 50240.0 17900.0 51585.0 ;
      RECT  17195.0 52930.0 17900.0 51585.0 ;
      RECT  17195.0 52930.0 17900.0 54275.0 ;
      RECT  17195.0 55620.0 17900.0 54275.0 ;
      RECT  17195.0 55620.0 17900.0 56965.0 ;
      RECT  17195.0 58310.0 17900.0 56965.0 ;
      RECT  17195.0 58310.0 17900.0 59655.0 ;
      RECT  17195.0 61000.0 17900.0 59655.0 ;
      RECT  17195.0 61000.0 17900.0 62345.0 ;
      RECT  17195.0 63690.0 17900.0 62345.0 ;
      RECT  17195.0 63690.0 17900.0 65035.0 ;
      RECT  17195.0 66380.0 17900.0 65035.0 ;
      RECT  17195.0 66380.0 17900.0 67725.0 ;
      RECT  17195.0 69070.0 17900.0 67725.0 ;
      RECT  17195.0 69070.0 17900.0 70415.0 ;
      RECT  17195.0 71760.0 17900.0 70415.0 ;
      RECT  17195.0 71760.0 17900.0 73105.0 ;
      RECT  17195.0 74450.0 17900.0 73105.0 ;
      RECT  17195.0 74450.0 17900.0 75795.0 ;
      RECT  17195.0 77140.0 17900.0 75795.0 ;
      RECT  17195.0 77140.0 17900.0 78485.0 ;
      RECT  17195.0 79830.0 17900.0 78485.0 ;
      RECT  17195.0 79830.0 17900.0 81175.0 ;
      RECT  17195.0 82520.0 17900.0 81175.0 ;
      RECT  17195.0 82520.0 17900.0 83865.0 ;
      RECT  17195.0 85210.0 17900.0 83865.0 ;
      RECT  17195.0 85210.0 17900.0 86555.0 ;
      RECT  17195.0 87900.0 17900.0 86555.0 ;
      RECT  17195.0 87900.0 17900.0 89245.0 ;
      RECT  17195.0 90590.0 17900.0 89245.0 ;
      RECT  17195.0 90590.0 17900.0 91935.0 ;
      RECT  17195.0 93280.0 17900.0 91935.0 ;
      RECT  17195.0 93280.0 17900.0 94625.0 ;
      RECT  17195.0 95970.0 17900.0 94625.0 ;
      RECT  17195.0 95970.0 17900.0 97315.0 ;
      RECT  17195.0 98660.0 17900.0 97315.0 ;
      RECT  17195.0 98660.0 17900.0 100005.0 ;
      RECT  17195.0 101350.0 17900.0 100005.0 ;
      RECT  17195.0 101350.0 17900.0 102695.0 ;
      RECT  17195.0 104040.0 17900.0 102695.0 ;
      RECT  17195.0 104040.0 17900.0 105385.0 ;
      RECT  17195.0 106730.0 17900.0 105385.0 ;
      RECT  17195.0 106730.0 17900.0 108075.0 ;
      RECT  17195.0 109420.0 17900.0 108075.0 ;
      RECT  17195.0 109420.0 17900.0 110765.0 ;
      RECT  17195.0 112110.0 17900.0 110765.0 ;
      RECT  17195.0 112110.0 17900.0 113455.0 ;
      RECT  17195.0 114800.0 17900.0 113455.0 ;
      RECT  17195.0 114800.0 17900.0 116145.0 ;
      RECT  17195.0 117490.0 17900.0 116145.0 ;
      RECT  17195.0 117490.0 17900.0 118835.0 ;
      RECT  17195.0 120180.0 17900.0 118835.0 ;
      RECT  17195.0 120180.0 17900.0 121525.0 ;
      RECT  17195.0 122870.0 17900.0 121525.0 ;
      RECT  17195.0 122870.0 17900.0 124215.0 ;
      RECT  17195.0 125560.0 17900.0 124215.0 ;
      RECT  17195.0 125560.0 17900.0 126905.0 ;
      RECT  17195.0 128250.0 17900.0 126905.0 ;
      RECT  17195.0 128250.0 17900.0 129595.0 ;
      RECT  17195.0 130940.0 17900.0 129595.0 ;
      RECT  17195.0 130940.0 17900.0 132285.0 ;
      RECT  17195.0 133630.0 17900.0 132285.0 ;
      RECT  17195.0 133630.0 17900.0 134975.0 ;
      RECT  17195.0 136320.0 17900.0 134975.0 ;
      RECT  17195.0 136320.0 17900.0 137665.0 ;
      RECT  17195.0 139010.0 17900.0 137665.0 ;
      RECT  17195.0 139010.0 17900.0 140355.0 ;
      RECT  17195.0 141700.0 17900.0 140355.0 ;
      RECT  17195.0 141700.0 17900.0 143045.0 ;
      RECT  17195.0 144390.0 17900.0 143045.0 ;
      RECT  17195.0 144390.0 17900.0 145735.0 ;
      RECT  17195.0 147080.0 17900.0 145735.0 ;
      RECT  17195.0 147080.0 17900.0 148425.0 ;
      RECT  17195.0 149770.0 17900.0 148425.0 ;
      RECT  17195.0 149770.0 17900.0 151115.0 ;
      RECT  17195.0 152460.0 17900.0 151115.0 ;
      RECT  17195.0 152460.0 17900.0 153805.0 ;
      RECT  17195.0 155150.0 17900.0 153805.0 ;
      RECT  17195.0 155150.0 17900.0 156495.0 ;
      RECT  17195.0 157840.0 17900.0 156495.0 ;
      RECT  17195.0 157840.0 17900.0 159185.0 ;
      RECT  17195.0 160530.0 17900.0 159185.0 ;
      RECT  17195.0 160530.0 17900.0 161875.0 ;
      RECT  17195.0 163220.0 17900.0 161875.0 ;
      RECT  17195.0 163220.0 17900.0 164565.0 ;
      RECT  17195.0 165910.0 17900.0 164565.0 ;
      RECT  17195.0 165910.0 17900.0 167255.0 ;
      RECT  17195.0 168600.0 17900.0 167255.0 ;
      RECT  17195.0 168600.0 17900.0 169945.0 ;
      RECT  17195.0 171290.0 17900.0 169945.0 ;
      RECT  17195.0 171290.0 17900.0 172635.0 ;
      RECT  17195.0 173980.0 17900.0 172635.0 ;
      RECT  17195.0 173980.0 17900.0 175325.0 ;
      RECT  17195.0 176670.0 17900.0 175325.0 ;
      RECT  17195.0 176670.0 17900.0 178015.0 ;
      RECT  17195.0 179360.0 17900.0 178015.0 ;
      RECT  17195.0 179360.0 17900.0 180705.0 ;
      RECT  17195.0 182050.0 17900.0 180705.0 ;
      RECT  17195.0 182050.0 17900.0 183395.0 ;
      RECT  17195.0 184740.0 17900.0 183395.0 ;
      RECT  17195.0 184740.0 17900.0 186085.0 ;
      RECT  17195.0 187430.0 17900.0 186085.0 ;
      RECT  17195.0 187430.0 17900.0 188775.0 ;
      RECT  17195.0 190120.0 17900.0 188775.0 ;
      RECT  17195.0 190120.0 17900.0 191465.0 ;
      RECT  17195.0 192810.0 17900.0 191465.0 ;
      RECT  17195.0 192810.0 17900.0 194155.0 ;
      RECT  17195.0 195500.0 17900.0 194155.0 ;
      RECT  17195.0 195500.0 17900.0 196845.0 ;
      RECT  17195.0 198190.0 17900.0 196845.0 ;
      RECT  17195.0 198190.0 17900.0 199535.0 ;
      RECT  17195.0 200880.0 17900.0 199535.0 ;
      RECT  17195.0 200880.0 17900.0 202225.0 ;
      RECT  17195.0 203570.0 17900.0 202225.0 ;
      RECT  17195.0 203570.0 17900.0 204915.0 ;
      RECT  17195.0 206260.0 17900.0 204915.0 ;
      RECT  17900.0 34100.0 18605.0 35445.0 ;
      RECT  17900.0 36790.0 18605.0 35445.0 ;
      RECT  17900.0 36790.0 18605.0 38135.0 ;
      RECT  17900.0 39480.0 18605.0 38135.0 ;
      RECT  17900.0 39480.0 18605.0 40825.0 ;
      RECT  17900.0 42170.0 18605.0 40825.0 ;
      RECT  17900.0 42170.0 18605.0 43515.0 ;
      RECT  17900.0 44860.0 18605.0 43515.0 ;
      RECT  17900.0 44860.0 18605.0 46205.0 ;
      RECT  17900.0 47550.0 18605.0 46205.0 ;
      RECT  17900.0 47550.0 18605.0 48895.0 ;
      RECT  17900.0 50240.0 18605.0 48895.0 ;
      RECT  17900.0 50240.0 18605.0 51585.0 ;
      RECT  17900.0 52930.0 18605.0 51585.0 ;
      RECT  17900.0 52930.0 18605.0 54275.0 ;
      RECT  17900.0 55620.0 18605.0 54275.0 ;
      RECT  17900.0 55620.0 18605.0 56965.0 ;
      RECT  17900.0 58310.0 18605.0 56965.0 ;
      RECT  17900.0 58310.0 18605.0 59655.0 ;
      RECT  17900.0 61000.0 18605.0 59655.0 ;
      RECT  17900.0 61000.0 18605.0 62345.0 ;
      RECT  17900.0 63690.0 18605.0 62345.0 ;
      RECT  17900.0 63690.0 18605.0 65035.0 ;
      RECT  17900.0 66380.0 18605.0 65035.0 ;
      RECT  17900.0 66380.0 18605.0 67725.0 ;
      RECT  17900.0 69070.0 18605.0 67725.0 ;
      RECT  17900.0 69070.0 18605.0 70415.0 ;
      RECT  17900.0 71760.0 18605.0 70415.0 ;
      RECT  17900.0 71760.0 18605.0 73105.0 ;
      RECT  17900.0 74450.0 18605.0 73105.0 ;
      RECT  17900.0 74450.0 18605.0 75795.0 ;
      RECT  17900.0 77140.0 18605.0 75795.0 ;
      RECT  17900.0 77140.0 18605.0 78485.0 ;
      RECT  17900.0 79830.0 18605.0 78485.0 ;
      RECT  17900.0 79830.0 18605.0 81175.0 ;
      RECT  17900.0 82520.0 18605.0 81175.0 ;
      RECT  17900.0 82520.0 18605.0 83865.0 ;
      RECT  17900.0 85210.0 18605.0 83865.0 ;
      RECT  17900.0 85210.0 18605.0 86555.0 ;
      RECT  17900.0 87900.0 18605.0 86555.0 ;
      RECT  17900.0 87900.0 18605.0 89245.0 ;
      RECT  17900.0 90590.0 18605.0 89245.0 ;
      RECT  17900.0 90590.0 18605.0 91935.0 ;
      RECT  17900.0 93280.0 18605.0 91935.0 ;
      RECT  17900.0 93280.0 18605.0 94625.0 ;
      RECT  17900.0 95970.0 18605.0 94625.0 ;
      RECT  17900.0 95970.0 18605.0 97315.0 ;
      RECT  17900.0 98660.0 18605.0 97315.0 ;
      RECT  17900.0 98660.0 18605.0 100005.0 ;
      RECT  17900.0 101350.0 18605.0 100005.0 ;
      RECT  17900.0 101350.0 18605.0 102695.0 ;
      RECT  17900.0 104040.0 18605.0 102695.0 ;
      RECT  17900.0 104040.0 18605.0 105385.0 ;
      RECT  17900.0 106730.0 18605.0 105385.0 ;
      RECT  17900.0 106730.0 18605.0 108075.0 ;
      RECT  17900.0 109420.0 18605.0 108075.0 ;
      RECT  17900.0 109420.0 18605.0 110765.0 ;
      RECT  17900.0 112110.0 18605.0 110765.0 ;
      RECT  17900.0 112110.0 18605.0 113455.0 ;
      RECT  17900.0 114800.0 18605.0 113455.0 ;
      RECT  17900.0 114800.0 18605.0 116145.0 ;
      RECT  17900.0 117490.0 18605.0 116145.0 ;
      RECT  17900.0 117490.0 18605.0 118835.0 ;
      RECT  17900.0 120180.0 18605.0 118835.0 ;
      RECT  17900.0 120180.0 18605.0 121525.0 ;
      RECT  17900.0 122870.0 18605.0 121525.0 ;
      RECT  17900.0 122870.0 18605.0 124215.0 ;
      RECT  17900.0 125560.0 18605.0 124215.0 ;
      RECT  17900.0 125560.0 18605.0 126905.0 ;
      RECT  17900.0 128250.0 18605.0 126905.0 ;
      RECT  17900.0 128250.0 18605.0 129595.0 ;
      RECT  17900.0 130940.0 18605.0 129595.0 ;
      RECT  17900.0 130940.0 18605.0 132285.0 ;
      RECT  17900.0 133630.0 18605.0 132285.0 ;
      RECT  17900.0 133630.0 18605.0 134975.0 ;
      RECT  17900.0 136320.0 18605.0 134975.0 ;
      RECT  17900.0 136320.0 18605.0 137665.0 ;
      RECT  17900.0 139010.0 18605.0 137665.0 ;
      RECT  17900.0 139010.0 18605.0 140355.0 ;
      RECT  17900.0 141700.0 18605.0 140355.0 ;
      RECT  17900.0 141700.0 18605.0 143045.0 ;
      RECT  17900.0 144390.0 18605.0 143045.0 ;
      RECT  17900.0 144390.0 18605.0 145735.0 ;
      RECT  17900.0 147080.0 18605.0 145735.0 ;
      RECT  17900.0 147080.0 18605.0 148425.0 ;
      RECT  17900.0 149770.0 18605.0 148425.0 ;
      RECT  17900.0 149770.0 18605.0 151115.0 ;
      RECT  17900.0 152460.0 18605.0 151115.0 ;
      RECT  17900.0 152460.0 18605.0 153805.0 ;
      RECT  17900.0 155150.0 18605.0 153805.0 ;
      RECT  17900.0 155150.0 18605.0 156495.0 ;
      RECT  17900.0 157840.0 18605.0 156495.0 ;
      RECT  17900.0 157840.0 18605.0 159185.0 ;
      RECT  17900.0 160530.0 18605.0 159185.0 ;
      RECT  17900.0 160530.0 18605.0 161875.0 ;
      RECT  17900.0 163220.0 18605.0 161875.0 ;
      RECT  17900.0 163220.0 18605.0 164565.0 ;
      RECT  17900.0 165910.0 18605.0 164565.0 ;
      RECT  17900.0 165910.0 18605.0 167255.0 ;
      RECT  17900.0 168600.0 18605.0 167255.0 ;
      RECT  17900.0 168600.0 18605.0 169945.0 ;
      RECT  17900.0 171290.0 18605.0 169945.0 ;
      RECT  17900.0 171290.0 18605.0 172635.0 ;
      RECT  17900.0 173980.0 18605.0 172635.0 ;
      RECT  17900.0 173980.0 18605.0 175325.0 ;
      RECT  17900.0 176670.0 18605.0 175325.0 ;
      RECT  17900.0 176670.0 18605.0 178015.0 ;
      RECT  17900.0 179360.0 18605.0 178015.0 ;
      RECT  17900.0 179360.0 18605.0 180705.0 ;
      RECT  17900.0 182050.0 18605.0 180705.0 ;
      RECT  17900.0 182050.0 18605.0 183395.0 ;
      RECT  17900.0 184740.0 18605.0 183395.0 ;
      RECT  17900.0 184740.0 18605.0 186085.0 ;
      RECT  17900.0 187430.0 18605.0 186085.0 ;
      RECT  17900.0 187430.0 18605.0 188775.0 ;
      RECT  17900.0 190120.0 18605.0 188775.0 ;
      RECT  17900.0 190120.0 18605.0 191465.0 ;
      RECT  17900.0 192810.0 18605.0 191465.0 ;
      RECT  17900.0 192810.0 18605.0 194155.0 ;
      RECT  17900.0 195500.0 18605.0 194155.0 ;
      RECT  17900.0 195500.0 18605.0 196845.0 ;
      RECT  17900.0 198190.0 18605.0 196845.0 ;
      RECT  17900.0 198190.0 18605.0 199535.0 ;
      RECT  17900.0 200880.0 18605.0 199535.0 ;
      RECT  17900.0 200880.0 18605.0 202225.0 ;
      RECT  17900.0 203570.0 18605.0 202225.0 ;
      RECT  17900.0 203570.0 18605.0 204915.0 ;
      RECT  17900.0 206260.0 18605.0 204915.0 ;
      RECT  18605.0 34100.0 19310.0 35445.0 ;
      RECT  18605.0 36790.0 19310.0 35445.0 ;
      RECT  18605.0 36790.0 19310.0 38135.0 ;
      RECT  18605.0 39480.0 19310.0 38135.0 ;
      RECT  18605.0 39480.0 19310.0 40825.0 ;
      RECT  18605.0 42170.0 19310.0 40825.0 ;
      RECT  18605.0 42170.0 19310.0 43515.0 ;
      RECT  18605.0 44860.0 19310.0 43515.0 ;
      RECT  18605.0 44860.0 19310.0 46205.0 ;
      RECT  18605.0 47550.0 19310.0 46205.0 ;
      RECT  18605.0 47550.0 19310.0 48895.0 ;
      RECT  18605.0 50240.0 19310.0 48895.0 ;
      RECT  18605.0 50240.0 19310.0 51585.0 ;
      RECT  18605.0 52930.0 19310.0 51585.0 ;
      RECT  18605.0 52930.0 19310.0 54275.0 ;
      RECT  18605.0 55620.0 19310.0 54275.0 ;
      RECT  18605.0 55620.0 19310.0 56965.0 ;
      RECT  18605.0 58310.0 19310.0 56965.0 ;
      RECT  18605.0 58310.0 19310.0 59655.0 ;
      RECT  18605.0 61000.0 19310.0 59655.0 ;
      RECT  18605.0 61000.0 19310.0 62345.0 ;
      RECT  18605.0 63690.0 19310.0 62345.0 ;
      RECT  18605.0 63690.0 19310.0 65035.0 ;
      RECT  18605.0 66380.0 19310.0 65035.0 ;
      RECT  18605.0 66380.0 19310.0 67725.0 ;
      RECT  18605.0 69070.0 19310.0 67725.0 ;
      RECT  18605.0 69070.0 19310.0 70415.0 ;
      RECT  18605.0 71760.0 19310.0 70415.0 ;
      RECT  18605.0 71760.0 19310.0 73105.0 ;
      RECT  18605.0 74450.0 19310.0 73105.0 ;
      RECT  18605.0 74450.0 19310.0 75795.0 ;
      RECT  18605.0 77140.0 19310.0 75795.0 ;
      RECT  18605.0 77140.0 19310.0 78485.0 ;
      RECT  18605.0 79830.0 19310.0 78485.0 ;
      RECT  18605.0 79830.0 19310.0 81175.0 ;
      RECT  18605.0 82520.0 19310.0 81175.0 ;
      RECT  18605.0 82520.0 19310.0 83865.0 ;
      RECT  18605.0 85210.0 19310.0 83865.0 ;
      RECT  18605.0 85210.0 19310.0 86555.0 ;
      RECT  18605.0 87900.0 19310.0 86555.0 ;
      RECT  18605.0 87900.0 19310.0 89245.0 ;
      RECT  18605.0 90590.0 19310.0 89245.0 ;
      RECT  18605.0 90590.0 19310.0 91935.0 ;
      RECT  18605.0 93280.0 19310.0 91935.0 ;
      RECT  18605.0 93280.0 19310.0 94625.0 ;
      RECT  18605.0 95970.0 19310.0 94625.0 ;
      RECT  18605.0 95970.0 19310.0 97315.0 ;
      RECT  18605.0 98660.0 19310.0 97315.0 ;
      RECT  18605.0 98660.0 19310.0 100005.0 ;
      RECT  18605.0 101350.0 19310.0 100005.0 ;
      RECT  18605.0 101350.0 19310.0 102695.0 ;
      RECT  18605.0 104040.0 19310.0 102695.0 ;
      RECT  18605.0 104040.0 19310.0 105385.0 ;
      RECT  18605.0 106730.0 19310.0 105385.0 ;
      RECT  18605.0 106730.0 19310.0 108075.0 ;
      RECT  18605.0 109420.0 19310.0 108075.0 ;
      RECT  18605.0 109420.0 19310.0 110765.0 ;
      RECT  18605.0 112110.0 19310.0 110765.0 ;
      RECT  18605.0 112110.0 19310.0 113455.0 ;
      RECT  18605.0 114800.0 19310.0 113455.0 ;
      RECT  18605.0 114800.0 19310.0 116145.0 ;
      RECT  18605.0 117490.0 19310.0 116145.0 ;
      RECT  18605.0 117490.0 19310.0 118835.0 ;
      RECT  18605.0 120180.0 19310.0 118835.0 ;
      RECT  18605.0 120180.0 19310.0 121525.0 ;
      RECT  18605.0 122870.0 19310.0 121525.0 ;
      RECT  18605.0 122870.0 19310.0 124215.0 ;
      RECT  18605.0 125560.0 19310.0 124215.0 ;
      RECT  18605.0 125560.0 19310.0 126905.0 ;
      RECT  18605.0 128250.0 19310.0 126905.0 ;
      RECT  18605.0 128250.0 19310.0 129595.0 ;
      RECT  18605.0 130940.0 19310.0 129595.0 ;
      RECT  18605.0 130940.0 19310.0 132285.0 ;
      RECT  18605.0 133630.0 19310.0 132285.0 ;
      RECT  18605.0 133630.0 19310.0 134975.0 ;
      RECT  18605.0 136320.0 19310.0 134975.0 ;
      RECT  18605.0 136320.0 19310.0 137665.0 ;
      RECT  18605.0 139010.0 19310.0 137665.0 ;
      RECT  18605.0 139010.0 19310.0 140355.0 ;
      RECT  18605.0 141700.0 19310.0 140355.0 ;
      RECT  18605.0 141700.0 19310.0 143045.0 ;
      RECT  18605.0 144390.0 19310.0 143045.0 ;
      RECT  18605.0 144390.0 19310.0 145735.0 ;
      RECT  18605.0 147080.0 19310.0 145735.0 ;
      RECT  18605.0 147080.0 19310.0 148425.0 ;
      RECT  18605.0 149770.0 19310.0 148425.0 ;
      RECT  18605.0 149770.0 19310.0 151115.0 ;
      RECT  18605.0 152460.0 19310.0 151115.0 ;
      RECT  18605.0 152460.0 19310.0 153805.0 ;
      RECT  18605.0 155150.0 19310.0 153805.0 ;
      RECT  18605.0 155150.0 19310.0 156495.0 ;
      RECT  18605.0 157840.0 19310.0 156495.0 ;
      RECT  18605.0 157840.0 19310.0 159185.0 ;
      RECT  18605.0 160530.0 19310.0 159185.0 ;
      RECT  18605.0 160530.0 19310.0 161875.0 ;
      RECT  18605.0 163220.0 19310.0 161875.0 ;
      RECT  18605.0 163220.0 19310.0 164565.0 ;
      RECT  18605.0 165910.0 19310.0 164565.0 ;
      RECT  18605.0 165910.0 19310.0 167255.0 ;
      RECT  18605.0 168600.0 19310.0 167255.0 ;
      RECT  18605.0 168600.0 19310.0 169945.0 ;
      RECT  18605.0 171290.0 19310.0 169945.0 ;
      RECT  18605.0 171290.0 19310.0 172635.0 ;
      RECT  18605.0 173980.0 19310.0 172635.0 ;
      RECT  18605.0 173980.0 19310.0 175325.0 ;
      RECT  18605.0 176670.0 19310.0 175325.0 ;
      RECT  18605.0 176670.0 19310.0 178015.0 ;
      RECT  18605.0 179360.0 19310.0 178015.0 ;
      RECT  18605.0 179360.0 19310.0 180705.0 ;
      RECT  18605.0 182050.0 19310.0 180705.0 ;
      RECT  18605.0 182050.0 19310.0 183395.0 ;
      RECT  18605.0 184740.0 19310.0 183395.0 ;
      RECT  18605.0 184740.0 19310.0 186085.0 ;
      RECT  18605.0 187430.0 19310.0 186085.0 ;
      RECT  18605.0 187430.0 19310.0 188775.0 ;
      RECT  18605.0 190120.0 19310.0 188775.0 ;
      RECT  18605.0 190120.0 19310.0 191465.0 ;
      RECT  18605.0 192810.0 19310.0 191465.0 ;
      RECT  18605.0 192810.0 19310.0 194155.0 ;
      RECT  18605.0 195500.0 19310.0 194155.0 ;
      RECT  18605.0 195500.0 19310.0 196845.0 ;
      RECT  18605.0 198190.0 19310.0 196845.0 ;
      RECT  18605.0 198190.0 19310.0 199535.0 ;
      RECT  18605.0 200880.0 19310.0 199535.0 ;
      RECT  18605.0 200880.0 19310.0 202225.0 ;
      RECT  18605.0 203570.0 19310.0 202225.0 ;
      RECT  18605.0 203570.0 19310.0 204915.0 ;
      RECT  18605.0 206260.0 19310.0 204915.0 ;
      RECT  19310.0 34100.0 20015.0 35445.0 ;
      RECT  19310.0 36790.0 20015.0 35445.0 ;
      RECT  19310.0 36790.0 20015.0 38135.0 ;
      RECT  19310.0 39480.0 20015.0 38135.0 ;
      RECT  19310.0 39480.0 20015.0 40825.0 ;
      RECT  19310.0 42170.0 20015.0 40825.0 ;
      RECT  19310.0 42170.0 20015.0 43515.0 ;
      RECT  19310.0 44860.0 20015.0 43515.0 ;
      RECT  19310.0 44860.0 20015.0 46205.0 ;
      RECT  19310.0 47550.0 20015.0 46205.0 ;
      RECT  19310.0 47550.0 20015.0 48895.0 ;
      RECT  19310.0 50240.0 20015.0 48895.0 ;
      RECT  19310.0 50240.0 20015.0 51585.0 ;
      RECT  19310.0 52930.0 20015.0 51585.0 ;
      RECT  19310.0 52930.0 20015.0 54275.0 ;
      RECT  19310.0 55620.0 20015.0 54275.0 ;
      RECT  19310.0 55620.0 20015.0 56965.0 ;
      RECT  19310.0 58310.0 20015.0 56965.0 ;
      RECT  19310.0 58310.0 20015.0 59655.0 ;
      RECT  19310.0 61000.0 20015.0 59655.0 ;
      RECT  19310.0 61000.0 20015.0 62345.0 ;
      RECT  19310.0 63690.0 20015.0 62345.0 ;
      RECT  19310.0 63690.0 20015.0 65035.0 ;
      RECT  19310.0 66380.0 20015.0 65035.0 ;
      RECT  19310.0 66380.0 20015.0 67725.0 ;
      RECT  19310.0 69070.0 20015.0 67725.0 ;
      RECT  19310.0 69070.0 20015.0 70415.0 ;
      RECT  19310.0 71760.0 20015.0 70415.0 ;
      RECT  19310.0 71760.0 20015.0 73105.0 ;
      RECT  19310.0 74450.0 20015.0 73105.0 ;
      RECT  19310.0 74450.0 20015.0 75795.0 ;
      RECT  19310.0 77140.0 20015.0 75795.0 ;
      RECT  19310.0 77140.0 20015.0 78485.0 ;
      RECT  19310.0 79830.0 20015.0 78485.0 ;
      RECT  19310.0 79830.0 20015.0 81175.0 ;
      RECT  19310.0 82520.0 20015.0 81175.0 ;
      RECT  19310.0 82520.0 20015.0 83865.0 ;
      RECT  19310.0 85210.0 20015.0 83865.0 ;
      RECT  19310.0 85210.0 20015.0 86555.0 ;
      RECT  19310.0 87900.0 20015.0 86555.0 ;
      RECT  19310.0 87900.0 20015.0 89245.0 ;
      RECT  19310.0 90590.0 20015.0 89245.0 ;
      RECT  19310.0 90590.0 20015.0 91935.0 ;
      RECT  19310.0 93280.0 20015.0 91935.0 ;
      RECT  19310.0 93280.0 20015.0 94625.0 ;
      RECT  19310.0 95970.0 20015.0 94625.0 ;
      RECT  19310.0 95970.0 20015.0 97315.0 ;
      RECT  19310.0 98660.0 20015.0 97315.0 ;
      RECT  19310.0 98660.0 20015.0 100005.0 ;
      RECT  19310.0 101350.0 20015.0 100005.0 ;
      RECT  19310.0 101350.0 20015.0 102695.0 ;
      RECT  19310.0 104040.0 20015.0 102695.0 ;
      RECT  19310.0 104040.0 20015.0 105385.0 ;
      RECT  19310.0 106730.0 20015.0 105385.0 ;
      RECT  19310.0 106730.0 20015.0 108075.0 ;
      RECT  19310.0 109420.0 20015.0 108075.0 ;
      RECT  19310.0 109420.0 20015.0 110765.0 ;
      RECT  19310.0 112110.0 20015.0 110765.0 ;
      RECT  19310.0 112110.0 20015.0 113455.0 ;
      RECT  19310.0 114800.0 20015.0 113455.0 ;
      RECT  19310.0 114800.0 20015.0 116145.0 ;
      RECT  19310.0 117490.0 20015.0 116145.0 ;
      RECT  19310.0 117490.0 20015.0 118835.0 ;
      RECT  19310.0 120180.0 20015.0 118835.0 ;
      RECT  19310.0 120180.0 20015.0 121525.0 ;
      RECT  19310.0 122870.0 20015.0 121525.0 ;
      RECT  19310.0 122870.0 20015.0 124215.0 ;
      RECT  19310.0 125560.0 20015.0 124215.0 ;
      RECT  19310.0 125560.0 20015.0 126905.0 ;
      RECT  19310.0 128250.0 20015.0 126905.0 ;
      RECT  19310.0 128250.0 20015.0 129595.0 ;
      RECT  19310.0 130940.0 20015.0 129595.0 ;
      RECT  19310.0 130940.0 20015.0 132285.0 ;
      RECT  19310.0 133630.0 20015.0 132285.0 ;
      RECT  19310.0 133630.0 20015.0 134975.0 ;
      RECT  19310.0 136320.0 20015.0 134975.0 ;
      RECT  19310.0 136320.0 20015.0 137665.0 ;
      RECT  19310.0 139010.0 20015.0 137665.0 ;
      RECT  19310.0 139010.0 20015.0 140355.0 ;
      RECT  19310.0 141700.0 20015.0 140355.0 ;
      RECT  19310.0 141700.0 20015.0 143045.0 ;
      RECT  19310.0 144390.0 20015.0 143045.0 ;
      RECT  19310.0 144390.0 20015.0 145735.0 ;
      RECT  19310.0 147080.0 20015.0 145735.0 ;
      RECT  19310.0 147080.0 20015.0 148425.0 ;
      RECT  19310.0 149770.0 20015.0 148425.0 ;
      RECT  19310.0 149770.0 20015.0 151115.0 ;
      RECT  19310.0 152460.0 20015.0 151115.0 ;
      RECT  19310.0 152460.0 20015.0 153805.0 ;
      RECT  19310.0 155150.0 20015.0 153805.0 ;
      RECT  19310.0 155150.0 20015.0 156495.0 ;
      RECT  19310.0 157840.0 20015.0 156495.0 ;
      RECT  19310.0 157840.0 20015.0 159185.0 ;
      RECT  19310.0 160530.0 20015.0 159185.0 ;
      RECT  19310.0 160530.0 20015.0 161875.0 ;
      RECT  19310.0 163220.0 20015.0 161875.0 ;
      RECT  19310.0 163220.0 20015.0 164565.0 ;
      RECT  19310.0 165910.0 20015.0 164565.0 ;
      RECT  19310.0 165910.0 20015.0 167255.0 ;
      RECT  19310.0 168600.0 20015.0 167255.0 ;
      RECT  19310.0 168600.0 20015.0 169945.0 ;
      RECT  19310.0 171290.0 20015.0 169945.0 ;
      RECT  19310.0 171290.0 20015.0 172635.0 ;
      RECT  19310.0 173980.0 20015.0 172635.0 ;
      RECT  19310.0 173980.0 20015.0 175325.0 ;
      RECT  19310.0 176670.0 20015.0 175325.0 ;
      RECT  19310.0 176670.0 20015.0 178015.0 ;
      RECT  19310.0 179360.0 20015.0 178015.0 ;
      RECT  19310.0 179360.0 20015.0 180705.0 ;
      RECT  19310.0 182050.0 20015.0 180705.0 ;
      RECT  19310.0 182050.0 20015.0 183395.0 ;
      RECT  19310.0 184740.0 20015.0 183395.0 ;
      RECT  19310.0 184740.0 20015.0 186085.0 ;
      RECT  19310.0 187430.0 20015.0 186085.0 ;
      RECT  19310.0 187430.0 20015.0 188775.0 ;
      RECT  19310.0 190120.0 20015.0 188775.0 ;
      RECT  19310.0 190120.0 20015.0 191465.0 ;
      RECT  19310.0 192810.0 20015.0 191465.0 ;
      RECT  19310.0 192810.0 20015.0 194155.0 ;
      RECT  19310.0 195500.0 20015.0 194155.0 ;
      RECT  19310.0 195500.0 20015.0 196845.0 ;
      RECT  19310.0 198190.0 20015.0 196845.0 ;
      RECT  19310.0 198190.0 20015.0 199535.0 ;
      RECT  19310.0 200880.0 20015.0 199535.0 ;
      RECT  19310.0 200880.0 20015.0 202225.0 ;
      RECT  19310.0 203570.0 20015.0 202225.0 ;
      RECT  19310.0 203570.0 20015.0 204915.0 ;
      RECT  19310.0 206260.0 20015.0 204915.0 ;
      RECT  20015.0 34100.0 20720.0 35445.0 ;
      RECT  20015.0 36790.0 20720.0 35445.0 ;
      RECT  20015.0 36790.0 20720.0 38135.0 ;
      RECT  20015.0 39480.0 20720.0 38135.0 ;
      RECT  20015.0 39480.0 20720.0 40825.0 ;
      RECT  20015.0 42170.0 20720.0 40825.0 ;
      RECT  20015.0 42170.0 20720.0 43515.0 ;
      RECT  20015.0 44860.0 20720.0 43515.0 ;
      RECT  20015.0 44860.0 20720.0 46205.0 ;
      RECT  20015.0 47550.0 20720.0 46205.0 ;
      RECT  20015.0 47550.0 20720.0 48895.0 ;
      RECT  20015.0 50240.0 20720.0 48895.0 ;
      RECT  20015.0 50240.0 20720.0 51585.0 ;
      RECT  20015.0 52930.0 20720.0 51585.0 ;
      RECT  20015.0 52930.0 20720.0 54275.0 ;
      RECT  20015.0 55620.0 20720.0 54275.0 ;
      RECT  20015.0 55620.0 20720.0 56965.0 ;
      RECT  20015.0 58310.0 20720.0 56965.0 ;
      RECT  20015.0 58310.0 20720.0 59655.0 ;
      RECT  20015.0 61000.0 20720.0 59655.0 ;
      RECT  20015.0 61000.0 20720.0 62345.0 ;
      RECT  20015.0 63690.0 20720.0 62345.0 ;
      RECT  20015.0 63690.0 20720.0 65035.0 ;
      RECT  20015.0 66380.0 20720.0 65035.0 ;
      RECT  20015.0 66380.0 20720.0 67725.0 ;
      RECT  20015.0 69070.0 20720.0 67725.0 ;
      RECT  20015.0 69070.0 20720.0 70415.0 ;
      RECT  20015.0 71760.0 20720.0 70415.0 ;
      RECT  20015.0 71760.0 20720.0 73105.0 ;
      RECT  20015.0 74450.0 20720.0 73105.0 ;
      RECT  20015.0 74450.0 20720.0 75795.0 ;
      RECT  20015.0 77140.0 20720.0 75795.0 ;
      RECT  20015.0 77140.0 20720.0 78485.0 ;
      RECT  20015.0 79830.0 20720.0 78485.0 ;
      RECT  20015.0 79830.0 20720.0 81175.0 ;
      RECT  20015.0 82520.0 20720.0 81175.0 ;
      RECT  20015.0 82520.0 20720.0 83865.0 ;
      RECT  20015.0 85210.0 20720.0 83865.0 ;
      RECT  20015.0 85210.0 20720.0 86555.0 ;
      RECT  20015.0 87900.0 20720.0 86555.0 ;
      RECT  20015.0 87900.0 20720.0 89245.0 ;
      RECT  20015.0 90590.0 20720.0 89245.0 ;
      RECT  20015.0 90590.0 20720.0 91935.0 ;
      RECT  20015.0 93280.0 20720.0 91935.0 ;
      RECT  20015.0 93280.0 20720.0 94625.0 ;
      RECT  20015.0 95970.0 20720.0 94625.0 ;
      RECT  20015.0 95970.0 20720.0 97315.0 ;
      RECT  20015.0 98660.0 20720.0 97315.0 ;
      RECT  20015.0 98660.0 20720.0 100005.0 ;
      RECT  20015.0 101350.0 20720.0 100005.0 ;
      RECT  20015.0 101350.0 20720.0 102695.0 ;
      RECT  20015.0 104040.0 20720.0 102695.0 ;
      RECT  20015.0 104040.0 20720.0 105385.0 ;
      RECT  20015.0 106730.0 20720.0 105385.0 ;
      RECT  20015.0 106730.0 20720.0 108075.0 ;
      RECT  20015.0 109420.0 20720.0 108075.0 ;
      RECT  20015.0 109420.0 20720.0 110765.0 ;
      RECT  20015.0 112110.0 20720.0 110765.0 ;
      RECT  20015.0 112110.0 20720.0 113455.0 ;
      RECT  20015.0 114800.0 20720.0 113455.0 ;
      RECT  20015.0 114800.0 20720.0 116145.0 ;
      RECT  20015.0 117490.0 20720.0 116145.0 ;
      RECT  20015.0 117490.0 20720.0 118835.0 ;
      RECT  20015.0 120180.0 20720.0 118835.0 ;
      RECT  20015.0 120180.0 20720.0 121525.0 ;
      RECT  20015.0 122870.0 20720.0 121525.0 ;
      RECT  20015.0 122870.0 20720.0 124215.0 ;
      RECT  20015.0 125560.0 20720.0 124215.0 ;
      RECT  20015.0 125560.0 20720.0 126905.0 ;
      RECT  20015.0 128250.0 20720.0 126905.0 ;
      RECT  20015.0 128250.0 20720.0 129595.0 ;
      RECT  20015.0 130940.0 20720.0 129595.0 ;
      RECT  20015.0 130940.0 20720.0 132285.0 ;
      RECT  20015.0 133630.0 20720.0 132285.0 ;
      RECT  20015.0 133630.0 20720.0 134975.0 ;
      RECT  20015.0 136320.0 20720.0 134975.0 ;
      RECT  20015.0 136320.0 20720.0 137665.0 ;
      RECT  20015.0 139010.0 20720.0 137665.0 ;
      RECT  20015.0 139010.0 20720.0 140355.0 ;
      RECT  20015.0 141700.0 20720.0 140355.0 ;
      RECT  20015.0 141700.0 20720.0 143045.0 ;
      RECT  20015.0 144390.0 20720.0 143045.0 ;
      RECT  20015.0 144390.0 20720.0 145735.0 ;
      RECT  20015.0 147080.0 20720.0 145735.0 ;
      RECT  20015.0 147080.0 20720.0 148425.0 ;
      RECT  20015.0 149770.0 20720.0 148425.0 ;
      RECT  20015.0 149770.0 20720.0 151115.0 ;
      RECT  20015.0 152460.0 20720.0 151115.0 ;
      RECT  20015.0 152460.0 20720.0 153805.0 ;
      RECT  20015.0 155150.0 20720.0 153805.0 ;
      RECT  20015.0 155150.0 20720.0 156495.0 ;
      RECT  20015.0 157840.0 20720.0 156495.0 ;
      RECT  20015.0 157840.0 20720.0 159185.0 ;
      RECT  20015.0 160530.0 20720.0 159185.0 ;
      RECT  20015.0 160530.0 20720.0 161875.0 ;
      RECT  20015.0 163220.0 20720.0 161875.0 ;
      RECT  20015.0 163220.0 20720.0 164565.0 ;
      RECT  20015.0 165910.0 20720.0 164565.0 ;
      RECT  20015.0 165910.0 20720.0 167255.0 ;
      RECT  20015.0 168600.0 20720.0 167255.0 ;
      RECT  20015.0 168600.0 20720.0 169945.0 ;
      RECT  20015.0 171290.0 20720.0 169945.0 ;
      RECT  20015.0 171290.0 20720.0 172635.0 ;
      RECT  20015.0 173980.0 20720.0 172635.0 ;
      RECT  20015.0 173980.0 20720.0 175325.0 ;
      RECT  20015.0 176670.0 20720.0 175325.0 ;
      RECT  20015.0 176670.0 20720.0 178015.0 ;
      RECT  20015.0 179360.0 20720.0 178015.0 ;
      RECT  20015.0 179360.0 20720.0 180705.0 ;
      RECT  20015.0 182050.0 20720.0 180705.0 ;
      RECT  20015.0 182050.0 20720.0 183395.0 ;
      RECT  20015.0 184740.0 20720.0 183395.0 ;
      RECT  20015.0 184740.0 20720.0 186085.0 ;
      RECT  20015.0 187430.0 20720.0 186085.0 ;
      RECT  20015.0 187430.0 20720.0 188775.0 ;
      RECT  20015.0 190120.0 20720.0 188775.0 ;
      RECT  20015.0 190120.0 20720.0 191465.0 ;
      RECT  20015.0 192810.0 20720.0 191465.0 ;
      RECT  20015.0 192810.0 20720.0 194155.0 ;
      RECT  20015.0 195500.0 20720.0 194155.0 ;
      RECT  20015.0 195500.0 20720.0 196845.0 ;
      RECT  20015.0 198190.0 20720.0 196845.0 ;
      RECT  20015.0 198190.0 20720.0 199535.0 ;
      RECT  20015.0 200880.0 20720.0 199535.0 ;
      RECT  20015.0 200880.0 20720.0 202225.0 ;
      RECT  20015.0 203570.0 20720.0 202225.0 ;
      RECT  20015.0 203570.0 20720.0 204915.0 ;
      RECT  20015.0 206260.0 20720.0 204915.0 ;
      RECT  20720.0 34100.0 21425.0 35445.0 ;
      RECT  20720.0 36790.0 21425.0 35445.0 ;
      RECT  20720.0 36790.0 21425.0 38135.0 ;
      RECT  20720.0 39480.0 21425.0 38135.0 ;
      RECT  20720.0 39480.0 21425.0 40825.0 ;
      RECT  20720.0 42170.0 21425.0 40825.0 ;
      RECT  20720.0 42170.0 21425.0 43515.0 ;
      RECT  20720.0 44860.0 21425.0 43515.0 ;
      RECT  20720.0 44860.0 21425.0 46205.0 ;
      RECT  20720.0 47550.0 21425.0 46205.0 ;
      RECT  20720.0 47550.0 21425.0 48895.0 ;
      RECT  20720.0 50240.0 21425.0 48895.0 ;
      RECT  20720.0 50240.0 21425.0 51585.0 ;
      RECT  20720.0 52930.0 21425.0 51585.0 ;
      RECT  20720.0 52930.0 21425.0 54275.0 ;
      RECT  20720.0 55620.0 21425.0 54275.0 ;
      RECT  20720.0 55620.0 21425.0 56965.0 ;
      RECT  20720.0 58310.0 21425.0 56965.0 ;
      RECT  20720.0 58310.0 21425.0 59655.0 ;
      RECT  20720.0 61000.0 21425.0 59655.0 ;
      RECT  20720.0 61000.0 21425.0 62345.0 ;
      RECT  20720.0 63690.0 21425.0 62345.0 ;
      RECT  20720.0 63690.0 21425.0 65035.0 ;
      RECT  20720.0 66380.0 21425.0 65035.0 ;
      RECT  20720.0 66380.0 21425.0 67725.0 ;
      RECT  20720.0 69070.0 21425.0 67725.0 ;
      RECT  20720.0 69070.0 21425.0 70415.0 ;
      RECT  20720.0 71760.0 21425.0 70415.0 ;
      RECT  20720.0 71760.0 21425.0 73105.0 ;
      RECT  20720.0 74450.0 21425.0 73105.0 ;
      RECT  20720.0 74450.0 21425.0 75795.0 ;
      RECT  20720.0 77140.0 21425.0 75795.0 ;
      RECT  20720.0 77140.0 21425.0 78485.0 ;
      RECT  20720.0 79830.0 21425.0 78485.0 ;
      RECT  20720.0 79830.0 21425.0 81175.0 ;
      RECT  20720.0 82520.0 21425.0 81175.0 ;
      RECT  20720.0 82520.0 21425.0 83865.0 ;
      RECT  20720.0 85210.0 21425.0 83865.0 ;
      RECT  20720.0 85210.0 21425.0 86555.0 ;
      RECT  20720.0 87900.0 21425.0 86555.0 ;
      RECT  20720.0 87900.0 21425.0 89245.0 ;
      RECT  20720.0 90590.0 21425.0 89245.0 ;
      RECT  20720.0 90590.0 21425.0 91935.0 ;
      RECT  20720.0 93280.0 21425.0 91935.0 ;
      RECT  20720.0 93280.0 21425.0 94625.0 ;
      RECT  20720.0 95970.0 21425.0 94625.0 ;
      RECT  20720.0 95970.0 21425.0 97315.0 ;
      RECT  20720.0 98660.0 21425.0 97315.0 ;
      RECT  20720.0 98660.0 21425.0 100005.0 ;
      RECT  20720.0 101350.0 21425.0 100005.0 ;
      RECT  20720.0 101350.0 21425.0 102695.0 ;
      RECT  20720.0 104040.0 21425.0 102695.0 ;
      RECT  20720.0 104040.0 21425.0 105385.0 ;
      RECT  20720.0 106730.0 21425.0 105385.0 ;
      RECT  20720.0 106730.0 21425.0 108075.0 ;
      RECT  20720.0 109420.0 21425.0 108075.0 ;
      RECT  20720.0 109420.0 21425.0 110765.0 ;
      RECT  20720.0 112110.0 21425.0 110765.0 ;
      RECT  20720.0 112110.0 21425.0 113455.0 ;
      RECT  20720.0 114800.0 21425.0 113455.0 ;
      RECT  20720.0 114800.0 21425.0 116145.0 ;
      RECT  20720.0 117490.0 21425.0 116145.0 ;
      RECT  20720.0 117490.0 21425.0 118835.0 ;
      RECT  20720.0 120180.0 21425.0 118835.0 ;
      RECT  20720.0 120180.0 21425.0 121525.0 ;
      RECT  20720.0 122870.0 21425.0 121525.0 ;
      RECT  20720.0 122870.0 21425.0 124215.0 ;
      RECT  20720.0 125560.0 21425.0 124215.0 ;
      RECT  20720.0 125560.0 21425.0 126905.0 ;
      RECT  20720.0 128250.0 21425.0 126905.0 ;
      RECT  20720.0 128250.0 21425.0 129595.0 ;
      RECT  20720.0 130940.0 21425.0 129595.0 ;
      RECT  20720.0 130940.0 21425.0 132285.0 ;
      RECT  20720.0 133630.0 21425.0 132285.0 ;
      RECT  20720.0 133630.0 21425.0 134975.0 ;
      RECT  20720.0 136320.0 21425.0 134975.0 ;
      RECT  20720.0 136320.0 21425.0 137665.0 ;
      RECT  20720.0 139010.0 21425.0 137665.0 ;
      RECT  20720.0 139010.0 21425.0 140355.0 ;
      RECT  20720.0 141700.0 21425.0 140355.0 ;
      RECT  20720.0 141700.0 21425.0 143045.0 ;
      RECT  20720.0 144390.0 21425.0 143045.0 ;
      RECT  20720.0 144390.0 21425.0 145735.0 ;
      RECT  20720.0 147080.0 21425.0 145735.0 ;
      RECT  20720.0 147080.0 21425.0 148425.0 ;
      RECT  20720.0 149770.0 21425.0 148425.0 ;
      RECT  20720.0 149770.0 21425.0 151115.0 ;
      RECT  20720.0 152460.0 21425.0 151115.0 ;
      RECT  20720.0 152460.0 21425.0 153805.0 ;
      RECT  20720.0 155150.0 21425.0 153805.0 ;
      RECT  20720.0 155150.0 21425.0 156495.0 ;
      RECT  20720.0 157840.0 21425.0 156495.0 ;
      RECT  20720.0 157840.0 21425.0 159185.0 ;
      RECT  20720.0 160530.0 21425.0 159185.0 ;
      RECT  20720.0 160530.0 21425.0 161875.0 ;
      RECT  20720.0 163220.0 21425.0 161875.0 ;
      RECT  20720.0 163220.0 21425.0 164565.0 ;
      RECT  20720.0 165910.0 21425.0 164565.0 ;
      RECT  20720.0 165910.0 21425.0 167255.0 ;
      RECT  20720.0 168600.0 21425.0 167255.0 ;
      RECT  20720.0 168600.0 21425.0 169945.0 ;
      RECT  20720.0 171290.0 21425.0 169945.0 ;
      RECT  20720.0 171290.0 21425.0 172635.0 ;
      RECT  20720.0 173980.0 21425.0 172635.0 ;
      RECT  20720.0 173980.0 21425.0 175325.0 ;
      RECT  20720.0 176670.0 21425.0 175325.0 ;
      RECT  20720.0 176670.0 21425.0 178015.0 ;
      RECT  20720.0 179360.0 21425.0 178015.0 ;
      RECT  20720.0 179360.0 21425.0 180705.0 ;
      RECT  20720.0 182050.0 21425.0 180705.0 ;
      RECT  20720.0 182050.0 21425.0 183395.0 ;
      RECT  20720.0 184740.0 21425.0 183395.0 ;
      RECT  20720.0 184740.0 21425.0 186085.0 ;
      RECT  20720.0 187430.0 21425.0 186085.0 ;
      RECT  20720.0 187430.0 21425.0 188775.0 ;
      RECT  20720.0 190120.0 21425.0 188775.0 ;
      RECT  20720.0 190120.0 21425.0 191465.0 ;
      RECT  20720.0 192810.0 21425.0 191465.0 ;
      RECT  20720.0 192810.0 21425.0 194155.0 ;
      RECT  20720.0 195500.0 21425.0 194155.0 ;
      RECT  20720.0 195500.0 21425.0 196845.0 ;
      RECT  20720.0 198190.0 21425.0 196845.0 ;
      RECT  20720.0 198190.0 21425.0 199535.0 ;
      RECT  20720.0 200880.0 21425.0 199535.0 ;
      RECT  20720.0 200880.0 21425.0 202225.0 ;
      RECT  20720.0 203570.0 21425.0 202225.0 ;
      RECT  20720.0 203570.0 21425.0 204915.0 ;
      RECT  20720.0 206260.0 21425.0 204915.0 ;
      RECT  21425.0 34100.0 22130.0 35445.0 ;
      RECT  21425.0 36790.0 22130.0 35445.0 ;
      RECT  21425.0 36790.0 22130.0 38135.0 ;
      RECT  21425.0 39480.0 22130.0 38135.0 ;
      RECT  21425.0 39480.0 22130.0 40825.0 ;
      RECT  21425.0 42170.0 22130.0 40825.0 ;
      RECT  21425.0 42170.0 22130.0 43515.0 ;
      RECT  21425.0 44860.0 22130.0 43515.0 ;
      RECT  21425.0 44860.0 22130.0 46205.0 ;
      RECT  21425.0 47550.0 22130.0 46205.0 ;
      RECT  21425.0 47550.0 22130.0 48895.0 ;
      RECT  21425.0 50240.0 22130.0 48895.0 ;
      RECT  21425.0 50240.0 22130.0 51585.0 ;
      RECT  21425.0 52930.0 22130.0 51585.0 ;
      RECT  21425.0 52930.0 22130.0 54275.0 ;
      RECT  21425.0 55620.0 22130.0 54275.0 ;
      RECT  21425.0 55620.0 22130.0 56965.0 ;
      RECT  21425.0 58310.0 22130.0 56965.0 ;
      RECT  21425.0 58310.0 22130.0 59655.0 ;
      RECT  21425.0 61000.0 22130.0 59655.0 ;
      RECT  21425.0 61000.0 22130.0 62345.0 ;
      RECT  21425.0 63690.0 22130.0 62345.0 ;
      RECT  21425.0 63690.0 22130.0 65035.0 ;
      RECT  21425.0 66380.0 22130.0 65035.0 ;
      RECT  21425.0 66380.0 22130.0 67725.0 ;
      RECT  21425.0 69070.0 22130.0 67725.0 ;
      RECT  21425.0 69070.0 22130.0 70415.0 ;
      RECT  21425.0 71760.0 22130.0 70415.0 ;
      RECT  21425.0 71760.0 22130.0 73105.0 ;
      RECT  21425.0 74450.0 22130.0 73105.0 ;
      RECT  21425.0 74450.0 22130.0 75795.0 ;
      RECT  21425.0 77140.0 22130.0 75795.0 ;
      RECT  21425.0 77140.0 22130.0 78485.0 ;
      RECT  21425.0 79830.0 22130.0 78485.0 ;
      RECT  21425.0 79830.0 22130.0 81175.0 ;
      RECT  21425.0 82520.0 22130.0 81175.0 ;
      RECT  21425.0 82520.0 22130.0 83865.0 ;
      RECT  21425.0 85210.0 22130.0 83865.0 ;
      RECT  21425.0 85210.0 22130.0 86555.0 ;
      RECT  21425.0 87900.0 22130.0 86555.0 ;
      RECT  21425.0 87900.0 22130.0 89245.0 ;
      RECT  21425.0 90590.0 22130.0 89245.0 ;
      RECT  21425.0 90590.0 22130.0 91935.0 ;
      RECT  21425.0 93280.0 22130.0 91935.0 ;
      RECT  21425.0 93280.0 22130.0 94625.0 ;
      RECT  21425.0 95970.0 22130.0 94625.0 ;
      RECT  21425.0 95970.0 22130.0 97315.0 ;
      RECT  21425.0 98660.0 22130.0 97315.0 ;
      RECT  21425.0 98660.0 22130.0 100005.0 ;
      RECT  21425.0 101350.0 22130.0 100005.0 ;
      RECT  21425.0 101350.0 22130.0 102695.0 ;
      RECT  21425.0 104040.0 22130.0 102695.0 ;
      RECT  21425.0 104040.0 22130.0 105385.0 ;
      RECT  21425.0 106730.0 22130.0 105385.0 ;
      RECT  21425.0 106730.0 22130.0 108075.0 ;
      RECT  21425.0 109420.0 22130.0 108075.0 ;
      RECT  21425.0 109420.0 22130.0 110765.0 ;
      RECT  21425.0 112110.0 22130.0 110765.0 ;
      RECT  21425.0 112110.0 22130.0 113455.0 ;
      RECT  21425.0 114800.0 22130.0 113455.0 ;
      RECT  21425.0 114800.0 22130.0 116145.0 ;
      RECT  21425.0 117490.0 22130.0 116145.0 ;
      RECT  21425.0 117490.0 22130.0 118835.0 ;
      RECT  21425.0 120180.0 22130.0 118835.0 ;
      RECT  21425.0 120180.0 22130.0 121525.0 ;
      RECT  21425.0 122870.0 22130.0 121525.0 ;
      RECT  21425.0 122870.0 22130.0 124215.0 ;
      RECT  21425.0 125560.0 22130.0 124215.0 ;
      RECT  21425.0 125560.0 22130.0 126905.0 ;
      RECT  21425.0 128250.0 22130.0 126905.0 ;
      RECT  21425.0 128250.0 22130.0 129595.0 ;
      RECT  21425.0 130940.0 22130.0 129595.0 ;
      RECT  21425.0 130940.0 22130.0 132285.0 ;
      RECT  21425.0 133630.0 22130.0 132285.0 ;
      RECT  21425.0 133630.0 22130.0 134975.0 ;
      RECT  21425.0 136320.0 22130.0 134975.0 ;
      RECT  21425.0 136320.0 22130.0 137665.0 ;
      RECT  21425.0 139010.0 22130.0 137665.0 ;
      RECT  21425.0 139010.0 22130.0 140355.0 ;
      RECT  21425.0 141700.0 22130.0 140355.0 ;
      RECT  21425.0 141700.0 22130.0 143045.0 ;
      RECT  21425.0 144390.0 22130.0 143045.0 ;
      RECT  21425.0 144390.0 22130.0 145735.0 ;
      RECT  21425.0 147080.0 22130.0 145735.0 ;
      RECT  21425.0 147080.0 22130.0 148425.0 ;
      RECT  21425.0 149770.0 22130.0 148425.0 ;
      RECT  21425.0 149770.0 22130.0 151115.0 ;
      RECT  21425.0 152460.0 22130.0 151115.0 ;
      RECT  21425.0 152460.0 22130.0 153805.0 ;
      RECT  21425.0 155150.0 22130.0 153805.0 ;
      RECT  21425.0 155150.0 22130.0 156495.0 ;
      RECT  21425.0 157840.0 22130.0 156495.0 ;
      RECT  21425.0 157840.0 22130.0 159185.0 ;
      RECT  21425.0 160530.0 22130.0 159185.0 ;
      RECT  21425.0 160530.0 22130.0 161875.0 ;
      RECT  21425.0 163220.0 22130.0 161875.0 ;
      RECT  21425.0 163220.0 22130.0 164565.0 ;
      RECT  21425.0 165910.0 22130.0 164565.0 ;
      RECT  21425.0 165910.0 22130.0 167255.0 ;
      RECT  21425.0 168600.0 22130.0 167255.0 ;
      RECT  21425.0 168600.0 22130.0 169945.0 ;
      RECT  21425.0 171290.0 22130.0 169945.0 ;
      RECT  21425.0 171290.0 22130.0 172635.0 ;
      RECT  21425.0 173980.0 22130.0 172635.0 ;
      RECT  21425.0 173980.0 22130.0 175325.0 ;
      RECT  21425.0 176670.0 22130.0 175325.0 ;
      RECT  21425.0 176670.0 22130.0 178015.0 ;
      RECT  21425.0 179360.0 22130.0 178015.0 ;
      RECT  21425.0 179360.0 22130.0 180705.0 ;
      RECT  21425.0 182050.0 22130.0 180705.0 ;
      RECT  21425.0 182050.0 22130.0 183395.0 ;
      RECT  21425.0 184740.0 22130.0 183395.0 ;
      RECT  21425.0 184740.0 22130.0 186085.0 ;
      RECT  21425.0 187430.0 22130.0 186085.0 ;
      RECT  21425.0 187430.0 22130.0 188775.0 ;
      RECT  21425.0 190120.0 22130.0 188775.0 ;
      RECT  21425.0 190120.0 22130.0 191465.0 ;
      RECT  21425.0 192810.0 22130.0 191465.0 ;
      RECT  21425.0 192810.0 22130.0 194155.0 ;
      RECT  21425.0 195500.0 22130.0 194155.0 ;
      RECT  21425.0 195500.0 22130.0 196845.0 ;
      RECT  21425.0 198190.0 22130.0 196845.0 ;
      RECT  21425.0 198190.0 22130.0 199535.0 ;
      RECT  21425.0 200880.0 22130.0 199535.0 ;
      RECT  21425.0 200880.0 22130.0 202225.0 ;
      RECT  21425.0 203570.0 22130.0 202225.0 ;
      RECT  21425.0 203570.0 22130.0 204915.0 ;
      RECT  21425.0 206260.0 22130.0 204915.0 ;
      RECT  22130.0 34100.0 22835.0 35445.0 ;
      RECT  22130.0 36790.0 22835.0 35445.0 ;
      RECT  22130.0 36790.0 22835.0 38135.0 ;
      RECT  22130.0 39480.0 22835.0 38135.0 ;
      RECT  22130.0 39480.0 22835.0 40825.0 ;
      RECT  22130.0 42170.0 22835.0 40825.0 ;
      RECT  22130.0 42170.0 22835.0 43515.0 ;
      RECT  22130.0 44860.0 22835.0 43515.0 ;
      RECT  22130.0 44860.0 22835.0 46205.0 ;
      RECT  22130.0 47550.0 22835.0 46205.0 ;
      RECT  22130.0 47550.0 22835.0 48895.0 ;
      RECT  22130.0 50240.0 22835.0 48895.0 ;
      RECT  22130.0 50240.0 22835.0 51585.0 ;
      RECT  22130.0 52930.0 22835.0 51585.0 ;
      RECT  22130.0 52930.0 22835.0 54275.0 ;
      RECT  22130.0 55620.0 22835.0 54275.0 ;
      RECT  22130.0 55620.0 22835.0 56965.0 ;
      RECT  22130.0 58310.0 22835.0 56965.0 ;
      RECT  22130.0 58310.0 22835.0 59655.0 ;
      RECT  22130.0 61000.0 22835.0 59655.0 ;
      RECT  22130.0 61000.0 22835.0 62345.0 ;
      RECT  22130.0 63690.0 22835.0 62345.0 ;
      RECT  22130.0 63690.0 22835.0 65035.0 ;
      RECT  22130.0 66380.0 22835.0 65035.0 ;
      RECT  22130.0 66380.0 22835.0 67725.0 ;
      RECT  22130.0 69070.0 22835.0 67725.0 ;
      RECT  22130.0 69070.0 22835.0 70415.0 ;
      RECT  22130.0 71760.0 22835.0 70415.0 ;
      RECT  22130.0 71760.0 22835.0 73105.0 ;
      RECT  22130.0 74450.0 22835.0 73105.0 ;
      RECT  22130.0 74450.0 22835.0 75795.0 ;
      RECT  22130.0 77140.0 22835.0 75795.0 ;
      RECT  22130.0 77140.0 22835.0 78485.0 ;
      RECT  22130.0 79830.0 22835.0 78485.0 ;
      RECT  22130.0 79830.0 22835.0 81175.0 ;
      RECT  22130.0 82520.0 22835.0 81175.0 ;
      RECT  22130.0 82520.0 22835.0 83865.0 ;
      RECT  22130.0 85210.0 22835.0 83865.0 ;
      RECT  22130.0 85210.0 22835.0 86555.0 ;
      RECT  22130.0 87900.0 22835.0 86555.0 ;
      RECT  22130.0 87900.0 22835.0 89245.0 ;
      RECT  22130.0 90590.0 22835.0 89245.0 ;
      RECT  22130.0 90590.0 22835.0 91935.0 ;
      RECT  22130.0 93280.0 22835.0 91935.0 ;
      RECT  22130.0 93280.0 22835.0 94625.0 ;
      RECT  22130.0 95970.0 22835.0 94625.0 ;
      RECT  22130.0 95970.0 22835.0 97315.0 ;
      RECT  22130.0 98660.0 22835.0 97315.0 ;
      RECT  22130.0 98660.0 22835.0 100005.0 ;
      RECT  22130.0 101350.0 22835.0 100005.0 ;
      RECT  22130.0 101350.0 22835.0 102695.0 ;
      RECT  22130.0 104040.0 22835.0 102695.0 ;
      RECT  22130.0 104040.0 22835.0 105385.0 ;
      RECT  22130.0 106730.0 22835.0 105385.0 ;
      RECT  22130.0 106730.0 22835.0 108075.0 ;
      RECT  22130.0 109420.0 22835.0 108075.0 ;
      RECT  22130.0 109420.0 22835.0 110765.0 ;
      RECT  22130.0 112110.0 22835.0 110765.0 ;
      RECT  22130.0 112110.0 22835.0 113455.0 ;
      RECT  22130.0 114800.0 22835.0 113455.0 ;
      RECT  22130.0 114800.0 22835.0 116145.0 ;
      RECT  22130.0 117490.0 22835.0 116145.0 ;
      RECT  22130.0 117490.0 22835.0 118835.0 ;
      RECT  22130.0 120180.0 22835.0 118835.0 ;
      RECT  22130.0 120180.0 22835.0 121525.0 ;
      RECT  22130.0 122870.0 22835.0 121525.0 ;
      RECT  22130.0 122870.0 22835.0 124215.0 ;
      RECT  22130.0 125560.0 22835.0 124215.0 ;
      RECT  22130.0 125560.0 22835.0 126905.0 ;
      RECT  22130.0 128250.0 22835.0 126905.0 ;
      RECT  22130.0 128250.0 22835.0 129595.0 ;
      RECT  22130.0 130940.0 22835.0 129595.0 ;
      RECT  22130.0 130940.0 22835.0 132285.0 ;
      RECT  22130.0 133630.0 22835.0 132285.0 ;
      RECT  22130.0 133630.0 22835.0 134975.0 ;
      RECT  22130.0 136320.0 22835.0 134975.0 ;
      RECT  22130.0 136320.0 22835.0 137665.0 ;
      RECT  22130.0 139010.0 22835.0 137665.0 ;
      RECT  22130.0 139010.0 22835.0 140355.0 ;
      RECT  22130.0 141700.0 22835.0 140355.0 ;
      RECT  22130.0 141700.0 22835.0 143045.0 ;
      RECT  22130.0 144390.0 22835.0 143045.0 ;
      RECT  22130.0 144390.0 22835.0 145735.0 ;
      RECT  22130.0 147080.0 22835.0 145735.0 ;
      RECT  22130.0 147080.0 22835.0 148425.0 ;
      RECT  22130.0 149770.0 22835.0 148425.0 ;
      RECT  22130.0 149770.0 22835.0 151115.0 ;
      RECT  22130.0 152460.0 22835.0 151115.0 ;
      RECT  22130.0 152460.0 22835.0 153805.0 ;
      RECT  22130.0 155150.0 22835.0 153805.0 ;
      RECT  22130.0 155150.0 22835.0 156495.0 ;
      RECT  22130.0 157840.0 22835.0 156495.0 ;
      RECT  22130.0 157840.0 22835.0 159185.0 ;
      RECT  22130.0 160530.0 22835.0 159185.0 ;
      RECT  22130.0 160530.0 22835.0 161875.0 ;
      RECT  22130.0 163220.0 22835.0 161875.0 ;
      RECT  22130.0 163220.0 22835.0 164565.0 ;
      RECT  22130.0 165910.0 22835.0 164565.0 ;
      RECT  22130.0 165910.0 22835.0 167255.0 ;
      RECT  22130.0 168600.0 22835.0 167255.0 ;
      RECT  22130.0 168600.0 22835.0 169945.0 ;
      RECT  22130.0 171290.0 22835.0 169945.0 ;
      RECT  22130.0 171290.0 22835.0 172635.0 ;
      RECT  22130.0 173980.0 22835.0 172635.0 ;
      RECT  22130.0 173980.0 22835.0 175325.0 ;
      RECT  22130.0 176670.0 22835.0 175325.0 ;
      RECT  22130.0 176670.0 22835.0 178015.0 ;
      RECT  22130.0 179360.0 22835.0 178015.0 ;
      RECT  22130.0 179360.0 22835.0 180705.0 ;
      RECT  22130.0 182050.0 22835.0 180705.0 ;
      RECT  22130.0 182050.0 22835.0 183395.0 ;
      RECT  22130.0 184740.0 22835.0 183395.0 ;
      RECT  22130.0 184740.0 22835.0 186085.0 ;
      RECT  22130.0 187430.0 22835.0 186085.0 ;
      RECT  22130.0 187430.0 22835.0 188775.0 ;
      RECT  22130.0 190120.0 22835.0 188775.0 ;
      RECT  22130.0 190120.0 22835.0 191465.0 ;
      RECT  22130.0 192810.0 22835.0 191465.0 ;
      RECT  22130.0 192810.0 22835.0 194155.0 ;
      RECT  22130.0 195500.0 22835.0 194155.0 ;
      RECT  22130.0 195500.0 22835.0 196845.0 ;
      RECT  22130.0 198190.0 22835.0 196845.0 ;
      RECT  22130.0 198190.0 22835.0 199535.0 ;
      RECT  22130.0 200880.0 22835.0 199535.0 ;
      RECT  22130.0 200880.0 22835.0 202225.0 ;
      RECT  22130.0 203570.0 22835.0 202225.0 ;
      RECT  22130.0 203570.0 22835.0 204915.0 ;
      RECT  22130.0 206260.0 22835.0 204915.0 ;
      RECT  22835.0 34100.0 23540.0 35445.0 ;
      RECT  22835.0 36790.0 23540.0 35445.0 ;
      RECT  22835.0 36790.0 23540.0 38135.0 ;
      RECT  22835.0 39480.0 23540.0 38135.0 ;
      RECT  22835.0 39480.0 23540.0 40825.0 ;
      RECT  22835.0 42170.0 23540.0 40825.0 ;
      RECT  22835.0 42170.0 23540.0 43515.0 ;
      RECT  22835.0 44860.0 23540.0 43515.0 ;
      RECT  22835.0 44860.0 23540.0 46205.0 ;
      RECT  22835.0 47550.0 23540.0 46205.0 ;
      RECT  22835.0 47550.0 23540.0 48895.0 ;
      RECT  22835.0 50240.0 23540.0 48895.0 ;
      RECT  22835.0 50240.0 23540.0 51585.0 ;
      RECT  22835.0 52930.0 23540.0 51585.0 ;
      RECT  22835.0 52930.0 23540.0 54275.0 ;
      RECT  22835.0 55620.0 23540.0 54275.0 ;
      RECT  22835.0 55620.0 23540.0 56965.0 ;
      RECT  22835.0 58310.0 23540.0 56965.0 ;
      RECT  22835.0 58310.0 23540.0 59655.0 ;
      RECT  22835.0 61000.0 23540.0 59655.0 ;
      RECT  22835.0 61000.0 23540.0 62345.0 ;
      RECT  22835.0 63690.0 23540.0 62345.0 ;
      RECT  22835.0 63690.0 23540.0 65035.0 ;
      RECT  22835.0 66380.0 23540.0 65035.0 ;
      RECT  22835.0 66380.0 23540.0 67725.0 ;
      RECT  22835.0 69070.0 23540.0 67725.0 ;
      RECT  22835.0 69070.0 23540.0 70415.0 ;
      RECT  22835.0 71760.0 23540.0 70415.0 ;
      RECT  22835.0 71760.0 23540.0 73105.0 ;
      RECT  22835.0 74450.0 23540.0 73105.0 ;
      RECT  22835.0 74450.0 23540.0 75795.0 ;
      RECT  22835.0 77140.0 23540.0 75795.0 ;
      RECT  22835.0 77140.0 23540.0 78485.0 ;
      RECT  22835.0 79830.0 23540.0 78485.0 ;
      RECT  22835.0 79830.0 23540.0 81175.0 ;
      RECT  22835.0 82520.0 23540.0 81175.0 ;
      RECT  22835.0 82520.0 23540.0 83865.0 ;
      RECT  22835.0 85210.0 23540.0 83865.0 ;
      RECT  22835.0 85210.0 23540.0 86555.0 ;
      RECT  22835.0 87900.0 23540.0 86555.0 ;
      RECT  22835.0 87900.0 23540.0 89245.0 ;
      RECT  22835.0 90590.0 23540.0 89245.0 ;
      RECT  22835.0 90590.0 23540.0 91935.0 ;
      RECT  22835.0 93280.0 23540.0 91935.0 ;
      RECT  22835.0 93280.0 23540.0 94625.0 ;
      RECT  22835.0 95970.0 23540.0 94625.0 ;
      RECT  22835.0 95970.0 23540.0 97315.0 ;
      RECT  22835.0 98660.0 23540.0 97315.0 ;
      RECT  22835.0 98660.0 23540.0 100005.0 ;
      RECT  22835.0 101350.0 23540.0 100005.0 ;
      RECT  22835.0 101350.0 23540.0 102695.0 ;
      RECT  22835.0 104040.0 23540.0 102695.0 ;
      RECT  22835.0 104040.0 23540.0 105385.0 ;
      RECT  22835.0 106730.0 23540.0 105385.0 ;
      RECT  22835.0 106730.0 23540.0 108075.0 ;
      RECT  22835.0 109420.0 23540.0 108075.0 ;
      RECT  22835.0 109420.0 23540.0 110765.0 ;
      RECT  22835.0 112110.0 23540.0 110765.0 ;
      RECT  22835.0 112110.0 23540.0 113455.0 ;
      RECT  22835.0 114800.0 23540.0 113455.0 ;
      RECT  22835.0 114800.0 23540.0 116145.0 ;
      RECT  22835.0 117490.0 23540.0 116145.0 ;
      RECT  22835.0 117490.0 23540.0 118835.0 ;
      RECT  22835.0 120180.0 23540.0 118835.0 ;
      RECT  22835.0 120180.0 23540.0 121525.0 ;
      RECT  22835.0 122870.0 23540.0 121525.0 ;
      RECT  22835.0 122870.0 23540.0 124215.0 ;
      RECT  22835.0 125560.0 23540.0 124215.0 ;
      RECT  22835.0 125560.0 23540.0 126905.0 ;
      RECT  22835.0 128250.0 23540.0 126905.0 ;
      RECT  22835.0 128250.0 23540.0 129595.0 ;
      RECT  22835.0 130940.0 23540.0 129595.0 ;
      RECT  22835.0 130940.0 23540.0 132285.0 ;
      RECT  22835.0 133630.0 23540.0 132285.0 ;
      RECT  22835.0 133630.0 23540.0 134975.0 ;
      RECT  22835.0 136320.0 23540.0 134975.0 ;
      RECT  22835.0 136320.0 23540.0 137665.0 ;
      RECT  22835.0 139010.0 23540.0 137665.0 ;
      RECT  22835.0 139010.0 23540.0 140355.0 ;
      RECT  22835.0 141700.0 23540.0 140355.0 ;
      RECT  22835.0 141700.0 23540.0 143045.0 ;
      RECT  22835.0 144390.0 23540.0 143045.0 ;
      RECT  22835.0 144390.0 23540.0 145735.0 ;
      RECT  22835.0 147080.0 23540.0 145735.0 ;
      RECT  22835.0 147080.0 23540.0 148425.0 ;
      RECT  22835.0 149770.0 23540.0 148425.0 ;
      RECT  22835.0 149770.0 23540.0 151115.0 ;
      RECT  22835.0 152460.0 23540.0 151115.0 ;
      RECT  22835.0 152460.0 23540.0 153805.0 ;
      RECT  22835.0 155150.0 23540.0 153805.0 ;
      RECT  22835.0 155150.0 23540.0 156495.0 ;
      RECT  22835.0 157840.0 23540.0 156495.0 ;
      RECT  22835.0 157840.0 23540.0 159185.0 ;
      RECT  22835.0 160530.0 23540.0 159185.0 ;
      RECT  22835.0 160530.0 23540.0 161875.0 ;
      RECT  22835.0 163220.0 23540.0 161875.0 ;
      RECT  22835.0 163220.0 23540.0 164565.0 ;
      RECT  22835.0 165910.0 23540.0 164565.0 ;
      RECT  22835.0 165910.0 23540.0 167255.0 ;
      RECT  22835.0 168600.0 23540.0 167255.0 ;
      RECT  22835.0 168600.0 23540.0 169945.0 ;
      RECT  22835.0 171290.0 23540.0 169945.0 ;
      RECT  22835.0 171290.0 23540.0 172635.0 ;
      RECT  22835.0 173980.0 23540.0 172635.0 ;
      RECT  22835.0 173980.0 23540.0 175325.0 ;
      RECT  22835.0 176670.0 23540.0 175325.0 ;
      RECT  22835.0 176670.0 23540.0 178015.0 ;
      RECT  22835.0 179360.0 23540.0 178015.0 ;
      RECT  22835.0 179360.0 23540.0 180705.0 ;
      RECT  22835.0 182050.0 23540.0 180705.0 ;
      RECT  22835.0 182050.0 23540.0 183395.0 ;
      RECT  22835.0 184740.0 23540.0 183395.0 ;
      RECT  22835.0 184740.0 23540.0 186085.0 ;
      RECT  22835.0 187430.0 23540.0 186085.0 ;
      RECT  22835.0 187430.0 23540.0 188775.0 ;
      RECT  22835.0 190120.0 23540.0 188775.0 ;
      RECT  22835.0 190120.0 23540.0 191465.0 ;
      RECT  22835.0 192810.0 23540.0 191465.0 ;
      RECT  22835.0 192810.0 23540.0 194155.0 ;
      RECT  22835.0 195500.0 23540.0 194155.0 ;
      RECT  22835.0 195500.0 23540.0 196845.0 ;
      RECT  22835.0 198190.0 23540.0 196845.0 ;
      RECT  22835.0 198190.0 23540.0 199535.0 ;
      RECT  22835.0 200880.0 23540.0 199535.0 ;
      RECT  22835.0 200880.0 23540.0 202225.0 ;
      RECT  22835.0 203570.0 23540.0 202225.0 ;
      RECT  22835.0 203570.0 23540.0 204915.0 ;
      RECT  22835.0 206260.0 23540.0 204915.0 ;
      RECT  23540.0 34100.0 24245.0 35445.0 ;
      RECT  23540.0 36790.0 24245.0 35445.0 ;
      RECT  23540.0 36790.0 24245.0 38135.0 ;
      RECT  23540.0 39480.0 24245.0 38135.0 ;
      RECT  23540.0 39480.0 24245.0 40825.0 ;
      RECT  23540.0 42170.0 24245.0 40825.0 ;
      RECT  23540.0 42170.0 24245.0 43515.0 ;
      RECT  23540.0 44860.0 24245.0 43515.0 ;
      RECT  23540.0 44860.0 24245.0 46205.0 ;
      RECT  23540.0 47550.0 24245.0 46205.0 ;
      RECT  23540.0 47550.0 24245.0 48895.0 ;
      RECT  23540.0 50240.0 24245.0 48895.0 ;
      RECT  23540.0 50240.0 24245.0 51585.0 ;
      RECT  23540.0 52930.0 24245.0 51585.0 ;
      RECT  23540.0 52930.0 24245.0 54275.0 ;
      RECT  23540.0 55620.0 24245.0 54275.0 ;
      RECT  23540.0 55620.0 24245.0 56965.0 ;
      RECT  23540.0 58310.0 24245.0 56965.0 ;
      RECT  23540.0 58310.0 24245.0 59655.0 ;
      RECT  23540.0 61000.0 24245.0 59655.0 ;
      RECT  23540.0 61000.0 24245.0 62345.0 ;
      RECT  23540.0 63690.0 24245.0 62345.0 ;
      RECT  23540.0 63690.0 24245.0 65035.0 ;
      RECT  23540.0 66380.0 24245.0 65035.0 ;
      RECT  23540.0 66380.0 24245.0 67725.0 ;
      RECT  23540.0 69070.0 24245.0 67725.0 ;
      RECT  23540.0 69070.0 24245.0 70415.0 ;
      RECT  23540.0 71760.0 24245.0 70415.0 ;
      RECT  23540.0 71760.0 24245.0 73105.0 ;
      RECT  23540.0 74450.0 24245.0 73105.0 ;
      RECT  23540.0 74450.0 24245.0 75795.0 ;
      RECT  23540.0 77140.0 24245.0 75795.0 ;
      RECT  23540.0 77140.0 24245.0 78485.0 ;
      RECT  23540.0 79830.0 24245.0 78485.0 ;
      RECT  23540.0 79830.0 24245.0 81175.0 ;
      RECT  23540.0 82520.0 24245.0 81175.0 ;
      RECT  23540.0 82520.0 24245.0 83865.0 ;
      RECT  23540.0 85210.0 24245.0 83865.0 ;
      RECT  23540.0 85210.0 24245.0 86555.0 ;
      RECT  23540.0 87900.0 24245.0 86555.0 ;
      RECT  23540.0 87900.0 24245.0 89245.0 ;
      RECT  23540.0 90590.0 24245.0 89245.0 ;
      RECT  23540.0 90590.0 24245.0 91935.0 ;
      RECT  23540.0 93280.0 24245.0 91935.0 ;
      RECT  23540.0 93280.0 24245.0 94625.0 ;
      RECT  23540.0 95970.0 24245.0 94625.0 ;
      RECT  23540.0 95970.0 24245.0 97315.0 ;
      RECT  23540.0 98660.0 24245.0 97315.0 ;
      RECT  23540.0 98660.0 24245.0 100005.0 ;
      RECT  23540.0 101350.0 24245.0 100005.0 ;
      RECT  23540.0 101350.0 24245.0 102695.0 ;
      RECT  23540.0 104040.0 24245.0 102695.0 ;
      RECT  23540.0 104040.0 24245.0 105385.0 ;
      RECT  23540.0 106730.0 24245.0 105385.0 ;
      RECT  23540.0 106730.0 24245.0 108075.0 ;
      RECT  23540.0 109420.0 24245.0 108075.0 ;
      RECT  23540.0 109420.0 24245.0 110765.0 ;
      RECT  23540.0 112110.0 24245.0 110765.0 ;
      RECT  23540.0 112110.0 24245.0 113455.0 ;
      RECT  23540.0 114800.0 24245.0 113455.0 ;
      RECT  23540.0 114800.0 24245.0 116145.0 ;
      RECT  23540.0 117490.0 24245.0 116145.0 ;
      RECT  23540.0 117490.0 24245.0 118835.0 ;
      RECT  23540.0 120180.0 24245.0 118835.0 ;
      RECT  23540.0 120180.0 24245.0 121525.0 ;
      RECT  23540.0 122870.0 24245.0 121525.0 ;
      RECT  23540.0 122870.0 24245.0 124215.0 ;
      RECT  23540.0 125560.0 24245.0 124215.0 ;
      RECT  23540.0 125560.0 24245.0 126905.0 ;
      RECT  23540.0 128250.0 24245.0 126905.0 ;
      RECT  23540.0 128250.0 24245.0 129595.0 ;
      RECT  23540.0 130940.0 24245.0 129595.0 ;
      RECT  23540.0 130940.0 24245.0 132285.0 ;
      RECT  23540.0 133630.0 24245.0 132285.0 ;
      RECT  23540.0 133630.0 24245.0 134975.0 ;
      RECT  23540.0 136320.0 24245.0 134975.0 ;
      RECT  23540.0 136320.0 24245.0 137665.0 ;
      RECT  23540.0 139010.0 24245.0 137665.0 ;
      RECT  23540.0 139010.0 24245.0 140355.0 ;
      RECT  23540.0 141700.0 24245.0 140355.0 ;
      RECT  23540.0 141700.0 24245.0 143045.0 ;
      RECT  23540.0 144390.0 24245.0 143045.0 ;
      RECT  23540.0 144390.0 24245.0 145735.0 ;
      RECT  23540.0 147080.0 24245.0 145735.0 ;
      RECT  23540.0 147080.0 24245.0 148425.0 ;
      RECT  23540.0 149770.0 24245.0 148425.0 ;
      RECT  23540.0 149770.0 24245.0 151115.0 ;
      RECT  23540.0 152460.0 24245.0 151115.0 ;
      RECT  23540.0 152460.0 24245.0 153805.0 ;
      RECT  23540.0 155150.0 24245.0 153805.0 ;
      RECT  23540.0 155150.0 24245.0 156495.0 ;
      RECT  23540.0 157840.0 24245.0 156495.0 ;
      RECT  23540.0 157840.0 24245.0 159185.0 ;
      RECT  23540.0 160530.0 24245.0 159185.0 ;
      RECT  23540.0 160530.0 24245.0 161875.0 ;
      RECT  23540.0 163220.0 24245.0 161875.0 ;
      RECT  23540.0 163220.0 24245.0 164565.0 ;
      RECT  23540.0 165910.0 24245.0 164565.0 ;
      RECT  23540.0 165910.0 24245.0 167255.0 ;
      RECT  23540.0 168600.0 24245.0 167255.0 ;
      RECT  23540.0 168600.0 24245.0 169945.0 ;
      RECT  23540.0 171290.0 24245.0 169945.0 ;
      RECT  23540.0 171290.0 24245.0 172635.0 ;
      RECT  23540.0 173980.0 24245.0 172635.0 ;
      RECT  23540.0 173980.0 24245.0 175325.0 ;
      RECT  23540.0 176670.0 24245.0 175325.0 ;
      RECT  23540.0 176670.0 24245.0 178015.0 ;
      RECT  23540.0 179360.0 24245.0 178015.0 ;
      RECT  23540.0 179360.0 24245.0 180705.0 ;
      RECT  23540.0 182050.0 24245.0 180705.0 ;
      RECT  23540.0 182050.0 24245.0 183395.0 ;
      RECT  23540.0 184740.0 24245.0 183395.0 ;
      RECT  23540.0 184740.0 24245.0 186085.0 ;
      RECT  23540.0 187430.0 24245.0 186085.0 ;
      RECT  23540.0 187430.0 24245.0 188775.0 ;
      RECT  23540.0 190120.0 24245.0 188775.0 ;
      RECT  23540.0 190120.0 24245.0 191465.0 ;
      RECT  23540.0 192810.0 24245.0 191465.0 ;
      RECT  23540.0 192810.0 24245.0 194155.0 ;
      RECT  23540.0 195500.0 24245.0 194155.0 ;
      RECT  23540.0 195500.0 24245.0 196845.0 ;
      RECT  23540.0 198190.0 24245.0 196845.0 ;
      RECT  23540.0 198190.0 24245.0 199535.0 ;
      RECT  23540.0 200880.0 24245.0 199535.0 ;
      RECT  23540.0 200880.0 24245.0 202225.0 ;
      RECT  23540.0 203570.0 24245.0 202225.0 ;
      RECT  23540.0 203570.0 24245.0 204915.0 ;
      RECT  23540.0 206260.0 24245.0 204915.0 ;
      RECT  24245.0 34100.0 24950.0 35445.0 ;
      RECT  24245.0 36790.0 24950.0 35445.0 ;
      RECT  24245.0 36790.0 24950.0 38135.0 ;
      RECT  24245.0 39480.0 24950.0 38135.0 ;
      RECT  24245.0 39480.0 24950.0 40825.0 ;
      RECT  24245.0 42170.0 24950.0 40825.0 ;
      RECT  24245.0 42170.0 24950.0 43515.0 ;
      RECT  24245.0 44860.0 24950.0 43515.0 ;
      RECT  24245.0 44860.0 24950.0 46205.0 ;
      RECT  24245.0 47550.0 24950.0 46205.0 ;
      RECT  24245.0 47550.0 24950.0 48895.0 ;
      RECT  24245.0 50240.0 24950.0 48895.0 ;
      RECT  24245.0 50240.0 24950.0 51585.0 ;
      RECT  24245.0 52930.0 24950.0 51585.0 ;
      RECT  24245.0 52930.0 24950.0 54275.0 ;
      RECT  24245.0 55620.0 24950.0 54275.0 ;
      RECT  24245.0 55620.0 24950.0 56965.0 ;
      RECT  24245.0 58310.0 24950.0 56965.0 ;
      RECT  24245.0 58310.0 24950.0 59655.0 ;
      RECT  24245.0 61000.0 24950.0 59655.0 ;
      RECT  24245.0 61000.0 24950.0 62345.0 ;
      RECT  24245.0 63690.0 24950.0 62345.0 ;
      RECT  24245.0 63690.0 24950.0 65035.0 ;
      RECT  24245.0 66380.0 24950.0 65035.0 ;
      RECT  24245.0 66380.0 24950.0 67725.0 ;
      RECT  24245.0 69070.0 24950.0 67725.0 ;
      RECT  24245.0 69070.0 24950.0 70415.0 ;
      RECT  24245.0 71760.0 24950.0 70415.0 ;
      RECT  24245.0 71760.0 24950.0 73105.0 ;
      RECT  24245.0 74450.0 24950.0 73105.0 ;
      RECT  24245.0 74450.0 24950.0 75795.0 ;
      RECT  24245.0 77140.0 24950.0 75795.0 ;
      RECT  24245.0 77140.0 24950.0 78485.0 ;
      RECT  24245.0 79830.0 24950.0 78485.0 ;
      RECT  24245.0 79830.0 24950.0 81175.0 ;
      RECT  24245.0 82520.0 24950.0 81175.0 ;
      RECT  24245.0 82520.0 24950.0 83865.0 ;
      RECT  24245.0 85210.0 24950.0 83865.0 ;
      RECT  24245.0 85210.0 24950.0 86555.0 ;
      RECT  24245.0 87900.0 24950.0 86555.0 ;
      RECT  24245.0 87900.0 24950.0 89245.0 ;
      RECT  24245.0 90590.0 24950.0 89245.0 ;
      RECT  24245.0 90590.0 24950.0 91935.0 ;
      RECT  24245.0 93280.0 24950.0 91935.0 ;
      RECT  24245.0 93280.0 24950.0 94625.0 ;
      RECT  24245.0 95970.0 24950.0 94625.0 ;
      RECT  24245.0 95970.0 24950.0 97315.0 ;
      RECT  24245.0 98660.0 24950.0 97315.0 ;
      RECT  24245.0 98660.0 24950.0 100005.0 ;
      RECT  24245.0 101350.0 24950.0 100005.0 ;
      RECT  24245.0 101350.0 24950.0 102695.0 ;
      RECT  24245.0 104040.0 24950.0 102695.0 ;
      RECT  24245.0 104040.0 24950.0 105385.0 ;
      RECT  24245.0 106730.0 24950.0 105385.0 ;
      RECT  24245.0 106730.0 24950.0 108075.0 ;
      RECT  24245.0 109420.0 24950.0 108075.0 ;
      RECT  24245.0 109420.0 24950.0 110765.0 ;
      RECT  24245.0 112110.0 24950.0 110765.0 ;
      RECT  24245.0 112110.0 24950.0 113455.0 ;
      RECT  24245.0 114800.0 24950.0 113455.0 ;
      RECT  24245.0 114800.0 24950.0 116145.0 ;
      RECT  24245.0 117490.0 24950.0 116145.0 ;
      RECT  24245.0 117490.0 24950.0 118835.0 ;
      RECT  24245.0 120180.0 24950.0 118835.0 ;
      RECT  24245.0 120180.0 24950.0 121525.0 ;
      RECT  24245.0 122870.0 24950.0 121525.0 ;
      RECT  24245.0 122870.0 24950.0 124215.0 ;
      RECT  24245.0 125560.0 24950.0 124215.0 ;
      RECT  24245.0 125560.0 24950.0 126905.0 ;
      RECT  24245.0 128250.0 24950.0 126905.0 ;
      RECT  24245.0 128250.0 24950.0 129595.0 ;
      RECT  24245.0 130940.0 24950.0 129595.0 ;
      RECT  24245.0 130940.0 24950.0 132285.0 ;
      RECT  24245.0 133630.0 24950.0 132285.0 ;
      RECT  24245.0 133630.0 24950.0 134975.0 ;
      RECT  24245.0 136320.0 24950.0 134975.0 ;
      RECT  24245.0 136320.0 24950.0 137665.0 ;
      RECT  24245.0 139010.0 24950.0 137665.0 ;
      RECT  24245.0 139010.0 24950.0 140355.0 ;
      RECT  24245.0 141700.0 24950.0 140355.0 ;
      RECT  24245.0 141700.0 24950.0 143045.0 ;
      RECT  24245.0 144390.0 24950.0 143045.0 ;
      RECT  24245.0 144390.0 24950.0 145735.0 ;
      RECT  24245.0 147080.0 24950.0 145735.0 ;
      RECT  24245.0 147080.0 24950.0 148425.0 ;
      RECT  24245.0 149770.0 24950.0 148425.0 ;
      RECT  24245.0 149770.0 24950.0 151115.0 ;
      RECT  24245.0 152460.0 24950.0 151115.0 ;
      RECT  24245.0 152460.0 24950.0 153805.0 ;
      RECT  24245.0 155150.0 24950.0 153805.0 ;
      RECT  24245.0 155150.0 24950.0 156495.0 ;
      RECT  24245.0 157840.0 24950.0 156495.0 ;
      RECT  24245.0 157840.0 24950.0 159185.0 ;
      RECT  24245.0 160530.0 24950.0 159185.0 ;
      RECT  24245.0 160530.0 24950.0 161875.0 ;
      RECT  24245.0 163220.0 24950.0 161875.0 ;
      RECT  24245.0 163220.0 24950.0 164565.0 ;
      RECT  24245.0 165910.0 24950.0 164565.0 ;
      RECT  24245.0 165910.0 24950.0 167255.0 ;
      RECT  24245.0 168600.0 24950.0 167255.0 ;
      RECT  24245.0 168600.0 24950.0 169945.0 ;
      RECT  24245.0 171290.0 24950.0 169945.0 ;
      RECT  24245.0 171290.0 24950.0 172635.0 ;
      RECT  24245.0 173980.0 24950.0 172635.0 ;
      RECT  24245.0 173980.0 24950.0 175325.0 ;
      RECT  24245.0 176670.0 24950.0 175325.0 ;
      RECT  24245.0 176670.0 24950.0 178015.0 ;
      RECT  24245.0 179360.0 24950.0 178015.0 ;
      RECT  24245.0 179360.0 24950.0 180705.0 ;
      RECT  24245.0 182050.0 24950.0 180705.0 ;
      RECT  24245.0 182050.0 24950.0 183395.0 ;
      RECT  24245.0 184740.0 24950.0 183395.0 ;
      RECT  24245.0 184740.0 24950.0 186085.0 ;
      RECT  24245.0 187430.0 24950.0 186085.0 ;
      RECT  24245.0 187430.0 24950.0 188775.0 ;
      RECT  24245.0 190120.0 24950.0 188775.0 ;
      RECT  24245.0 190120.0 24950.0 191465.0 ;
      RECT  24245.0 192810.0 24950.0 191465.0 ;
      RECT  24245.0 192810.0 24950.0 194155.0 ;
      RECT  24245.0 195500.0 24950.0 194155.0 ;
      RECT  24245.0 195500.0 24950.0 196845.0 ;
      RECT  24245.0 198190.0 24950.0 196845.0 ;
      RECT  24245.0 198190.0 24950.0 199535.0 ;
      RECT  24245.0 200880.0 24950.0 199535.0 ;
      RECT  24245.0 200880.0 24950.0 202225.0 ;
      RECT  24245.0 203570.0 24950.0 202225.0 ;
      RECT  24245.0 203570.0 24950.0 204915.0 ;
      RECT  24245.0 206260.0 24950.0 204915.0 ;
      RECT  24950.0 34100.0 25655.0 35445.0 ;
      RECT  24950.0 36790.0 25655.0 35445.0 ;
      RECT  24950.0 36790.0 25655.0 38135.0 ;
      RECT  24950.0 39480.0 25655.0 38135.0 ;
      RECT  24950.0 39480.0 25655.0 40825.0 ;
      RECT  24950.0 42170.0 25655.0 40825.0 ;
      RECT  24950.0 42170.0 25655.0 43515.0 ;
      RECT  24950.0 44860.0 25655.0 43515.0 ;
      RECT  24950.0 44860.0 25655.0 46205.0 ;
      RECT  24950.0 47550.0 25655.0 46205.0 ;
      RECT  24950.0 47550.0 25655.0 48895.0 ;
      RECT  24950.0 50240.0 25655.0 48895.0 ;
      RECT  24950.0 50240.0 25655.0 51585.0 ;
      RECT  24950.0 52930.0 25655.0 51585.0 ;
      RECT  24950.0 52930.0 25655.0 54275.0 ;
      RECT  24950.0 55620.0 25655.0 54275.0 ;
      RECT  24950.0 55620.0 25655.0 56965.0 ;
      RECT  24950.0 58310.0 25655.0 56965.0 ;
      RECT  24950.0 58310.0 25655.0 59655.0 ;
      RECT  24950.0 61000.0 25655.0 59655.0 ;
      RECT  24950.0 61000.0 25655.0 62345.0 ;
      RECT  24950.0 63690.0 25655.0 62345.0 ;
      RECT  24950.0 63690.0 25655.0 65035.0 ;
      RECT  24950.0 66380.0 25655.0 65035.0 ;
      RECT  24950.0 66380.0 25655.0 67725.0 ;
      RECT  24950.0 69070.0 25655.0 67725.0 ;
      RECT  24950.0 69070.0 25655.0 70415.0 ;
      RECT  24950.0 71760.0 25655.0 70415.0 ;
      RECT  24950.0 71760.0 25655.0 73105.0 ;
      RECT  24950.0 74450.0 25655.0 73105.0 ;
      RECT  24950.0 74450.0 25655.0 75795.0 ;
      RECT  24950.0 77140.0 25655.0 75795.0 ;
      RECT  24950.0 77140.0 25655.0 78485.0 ;
      RECT  24950.0 79830.0 25655.0 78485.0 ;
      RECT  24950.0 79830.0 25655.0 81175.0 ;
      RECT  24950.0 82520.0 25655.0 81175.0 ;
      RECT  24950.0 82520.0 25655.0 83865.0 ;
      RECT  24950.0 85210.0 25655.0 83865.0 ;
      RECT  24950.0 85210.0 25655.0 86555.0 ;
      RECT  24950.0 87900.0 25655.0 86555.0 ;
      RECT  24950.0 87900.0 25655.0 89245.0 ;
      RECT  24950.0 90590.0 25655.0 89245.0 ;
      RECT  24950.0 90590.0 25655.0 91935.0 ;
      RECT  24950.0 93280.0 25655.0 91935.0 ;
      RECT  24950.0 93280.0 25655.0 94625.0 ;
      RECT  24950.0 95970.0 25655.0 94625.0 ;
      RECT  24950.0 95970.0 25655.0 97315.0 ;
      RECT  24950.0 98660.0 25655.0 97315.0 ;
      RECT  24950.0 98660.0 25655.0 100005.0 ;
      RECT  24950.0 101350.0 25655.0 100005.0 ;
      RECT  24950.0 101350.0 25655.0 102695.0 ;
      RECT  24950.0 104040.0 25655.0 102695.0 ;
      RECT  24950.0 104040.0 25655.0 105385.0 ;
      RECT  24950.0 106730.0 25655.0 105385.0 ;
      RECT  24950.0 106730.0 25655.0 108075.0 ;
      RECT  24950.0 109420.0 25655.0 108075.0 ;
      RECT  24950.0 109420.0 25655.0 110765.0 ;
      RECT  24950.0 112110.0 25655.0 110765.0 ;
      RECT  24950.0 112110.0 25655.0 113455.0 ;
      RECT  24950.0 114800.0 25655.0 113455.0 ;
      RECT  24950.0 114800.0 25655.0 116145.0 ;
      RECT  24950.0 117490.0 25655.0 116145.0 ;
      RECT  24950.0 117490.0 25655.0 118835.0 ;
      RECT  24950.0 120180.0 25655.0 118835.0 ;
      RECT  24950.0 120180.0 25655.0 121525.0 ;
      RECT  24950.0 122870.0 25655.0 121525.0 ;
      RECT  24950.0 122870.0 25655.0 124215.0 ;
      RECT  24950.0 125560.0 25655.0 124215.0 ;
      RECT  24950.0 125560.0 25655.0 126905.0 ;
      RECT  24950.0 128250.0 25655.0 126905.0 ;
      RECT  24950.0 128250.0 25655.0 129595.0 ;
      RECT  24950.0 130940.0 25655.0 129595.0 ;
      RECT  24950.0 130940.0 25655.0 132285.0 ;
      RECT  24950.0 133630.0 25655.0 132285.0 ;
      RECT  24950.0 133630.0 25655.0 134975.0 ;
      RECT  24950.0 136320.0 25655.0 134975.0 ;
      RECT  24950.0 136320.0 25655.0 137665.0 ;
      RECT  24950.0 139010.0 25655.0 137665.0 ;
      RECT  24950.0 139010.0 25655.0 140355.0 ;
      RECT  24950.0 141700.0 25655.0 140355.0 ;
      RECT  24950.0 141700.0 25655.0 143045.0 ;
      RECT  24950.0 144390.0 25655.0 143045.0 ;
      RECT  24950.0 144390.0 25655.0 145735.0 ;
      RECT  24950.0 147080.0 25655.0 145735.0 ;
      RECT  24950.0 147080.0 25655.0 148425.0 ;
      RECT  24950.0 149770.0 25655.0 148425.0 ;
      RECT  24950.0 149770.0 25655.0 151115.0 ;
      RECT  24950.0 152460.0 25655.0 151115.0 ;
      RECT  24950.0 152460.0 25655.0 153805.0 ;
      RECT  24950.0 155150.0 25655.0 153805.0 ;
      RECT  24950.0 155150.0 25655.0 156495.0 ;
      RECT  24950.0 157840.0 25655.0 156495.0 ;
      RECT  24950.0 157840.0 25655.0 159185.0 ;
      RECT  24950.0 160530.0 25655.0 159185.0 ;
      RECT  24950.0 160530.0 25655.0 161875.0 ;
      RECT  24950.0 163220.0 25655.0 161875.0 ;
      RECT  24950.0 163220.0 25655.0 164565.0 ;
      RECT  24950.0 165910.0 25655.0 164565.0 ;
      RECT  24950.0 165910.0 25655.0 167255.0 ;
      RECT  24950.0 168600.0 25655.0 167255.0 ;
      RECT  24950.0 168600.0 25655.0 169945.0 ;
      RECT  24950.0 171290.0 25655.0 169945.0 ;
      RECT  24950.0 171290.0 25655.0 172635.0 ;
      RECT  24950.0 173980.0 25655.0 172635.0 ;
      RECT  24950.0 173980.0 25655.0 175325.0 ;
      RECT  24950.0 176670.0 25655.0 175325.0 ;
      RECT  24950.0 176670.0 25655.0 178015.0 ;
      RECT  24950.0 179360.0 25655.0 178015.0 ;
      RECT  24950.0 179360.0 25655.0 180705.0 ;
      RECT  24950.0 182050.0 25655.0 180705.0 ;
      RECT  24950.0 182050.0 25655.0 183395.0 ;
      RECT  24950.0 184740.0 25655.0 183395.0 ;
      RECT  24950.0 184740.0 25655.0 186085.0 ;
      RECT  24950.0 187430.0 25655.0 186085.0 ;
      RECT  24950.0 187430.0 25655.0 188775.0 ;
      RECT  24950.0 190120.0 25655.0 188775.0 ;
      RECT  24950.0 190120.0 25655.0 191465.0 ;
      RECT  24950.0 192810.0 25655.0 191465.0 ;
      RECT  24950.0 192810.0 25655.0 194155.0 ;
      RECT  24950.0 195500.0 25655.0 194155.0 ;
      RECT  24950.0 195500.0 25655.0 196845.0 ;
      RECT  24950.0 198190.0 25655.0 196845.0 ;
      RECT  24950.0 198190.0 25655.0 199535.0 ;
      RECT  24950.0 200880.0 25655.0 199535.0 ;
      RECT  24950.0 200880.0 25655.0 202225.0 ;
      RECT  24950.0 203570.0 25655.0 202225.0 ;
      RECT  24950.0 203570.0 25655.0 204915.0 ;
      RECT  24950.0 206260.0 25655.0 204915.0 ;
      RECT  25655.0 34100.0 26360.0 35445.0 ;
      RECT  25655.0 36790.0 26360.0 35445.0 ;
      RECT  25655.0 36790.0 26360.0 38135.0 ;
      RECT  25655.0 39480.0 26360.0 38135.0 ;
      RECT  25655.0 39480.0 26360.0 40825.0 ;
      RECT  25655.0 42170.0 26360.0 40825.0 ;
      RECT  25655.0 42170.0 26360.0 43515.0 ;
      RECT  25655.0 44860.0 26360.0 43515.0 ;
      RECT  25655.0 44860.0 26360.0 46205.0 ;
      RECT  25655.0 47550.0 26360.0 46205.0 ;
      RECT  25655.0 47550.0 26360.0 48895.0 ;
      RECT  25655.0 50240.0 26360.0 48895.0 ;
      RECT  25655.0 50240.0 26360.0 51585.0 ;
      RECT  25655.0 52930.0 26360.0 51585.0 ;
      RECT  25655.0 52930.0 26360.0 54275.0 ;
      RECT  25655.0 55620.0 26360.0 54275.0 ;
      RECT  25655.0 55620.0 26360.0 56965.0 ;
      RECT  25655.0 58310.0 26360.0 56965.0 ;
      RECT  25655.0 58310.0 26360.0 59655.0 ;
      RECT  25655.0 61000.0 26360.0 59655.0 ;
      RECT  25655.0 61000.0 26360.0 62345.0 ;
      RECT  25655.0 63690.0 26360.0 62345.0 ;
      RECT  25655.0 63690.0 26360.0 65035.0 ;
      RECT  25655.0 66380.0 26360.0 65035.0 ;
      RECT  25655.0 66380.0 26360.0 67725.0 ;
      RECT  25655.0 69070.0 26360.0 67725.0 ;
      RECT  25655.0 69070.0 26360.0 70415.0 ;
      RECT  25655.0 71760.0 26360.0 70415.0 ;
      RECT  25655.0 71760.0 26360.0 73105.0 ;
      RECT  25655.0 74450.0 26360.0 73105.0 ;
      RECT  25655.0 74450.0 26360.0 75795.0 ;
      RECT  25655.0 77140.0 26360.0 75795.0 ;
      RECT  25655.0 77140.0 26360.0 78485.0 ;
      RECT  25655.0 79830.0 26360.0 78485.0 ;
      RECT  25655.0 79830.0 26360.0 81175.0 ;
      RECT  25655.0 82520.0 26360.0 81175.0 ;
      RECT  25655.0 82520.0 26360.0 83865.0 ;
      RECT  25655.0 85210.0 26360.0 83865.0 ;
      RECT  25655.0 85210.0 26360.0 86555.0 ;
      RECT  25655.0 87900.0 26360.0 86555.0 ;
      RECT  25655.0 87900.0 26360.0 89245.0 ;
      RECT  25655.0 90590.0 26360.0 89245.0 ;
      RECT  25655.0 90590.0 26360.0 91935.0 ;
      RECT  25655.0 93280.0 26360.0 91935.0 ;
      RECT  25655.0 93280.0 26360.0 94625.0 ;
      RECT  25655.0 95970.0 26360.0 94625.0 ;
      RECT  25655.0 95970.0 26360.0 97315.0 ;
      RECT  25655.0 98660.0 26360.0 97315.0 ;
      RECT  25655.0 98660.0 26360.0 100005.0 ;
      RECT  25655.0 101350.0 26360.0 100005.0 ;
      RECT  25655.0 101350.0 26360.0 102695.0 ;
      RECT  25655.0 104040.0 26360.0 102695.0 ;
      RECT  25655.0 104040.0 26360.0 105385.0 ;
      RECT  25655.0 106730.0 26360.0 105385.0 ;
      RECT  25655.0 106730.0 26360.0 108075.0 ;
      RECT  25655.0 109420.0 26360.0 108075.0 ;
      RECT  25655.0 109420.0 26360.0 110765.0 ;
      RECT  25655.0 112110.0 26360.0 110765.0 ;
      RECT  25655.0 112110.0 26360.0 113455.0 ;
      RECT  25655.0 114800.0 26360.0 113455.0 ;
      RECT  25655.0 114800.0 26360.0 116145.0 ;
      RECT  25655.0 117490.0 26360.0 116145.0 ;
      RECT  25655.0 117490.0 26360.0 118835.0 ;
      RECT  25655.0 120180.0 26360.0 118835.0 ;
      RECT  25655.0 120180.0 26360.0 121525.0 ;
      RECT  25655.0 122870.0 26360.0 121525.0 ;
      RECT  25655.0 122870.0 26360.0 124215.0 ;
      RECT  25655.0 125560.0 26360.0 124215.0 ;
      RECT  25655.0 125560.0 26360.0 126905.0 ;
      RECT  25655.0 128250.0 26360.0 126905.0 ;
      RECT  25655.0 128250.0 26360.0 129595.0 ;
      RECT  25655.0 130940.0 26360.0 129595.0 ;
      RECT  25655.0 130940.0 26360.0 132285.0 ;
      RECT  25655.0 133630.0 26360.0 132285.0 ;
      RECT  25655.0 133630.0 26360.0 134975.0 ;
      RECT  25655.0 136320.0 26360.0 134975.0 ;
      RECT  25655.0 136320.0 26360.0 137665.0 ;
      RECT  25655.0 139010.0 26360.0 137665.0 ;
      RECT  25655.0 139010.0 26360.0 140355.0 ;
      RECT  25655.0 141700.0 26360.0 140355.0 ;
      RECT  25655.0 141700.0 26360.0 143045.0 ;
      RECT  25655.0 144390.0 26360.0 143045.0 ;
      RECT  25655.0 144390.0 26360.0 145735.0 ;
      RECT  25655.0 147080.0 26360.0 145735.0 ;
      RECT  25655.0 147080.0 26360.0 148425.0 ;
      RECT  25655.0 149770.0 26360.0 148425.0 ;
      RECT  25655.0 149770.0 26360.0 151115.0 ;
      RECT  25655.0 152460.0 26360.0 151115.0 ;
      RECT  25655.0 152460.0 26360.0 153805.0 ;
      RECT  25655.0 155150.0 26360.0 153805.0 ;
      RECT  25655.0 155150.0 26360.0 156495.0 ;
      RECT  25655.0 157840.0 26360.0 156495.0 ;
      RECT  25655.0 157840.0 26360.0 159185.0 ;
      RECT  25655.0 160530.0 26360.0 159185.0 ;
      RECT  25655.0 160530.0 26360.0 161875.0 ;
      RECT  25655.0 163220.0 26360.0 161875.0 ;
      RECT  25655.0 163220.0 26360.0 164565.0 ;
      RECT  25655.0 165910.0 26360.0 164565.0 ;
      RECT  25655.0 165910.0 26360.0 167255.0 ;
      RECT  25655.0 168600.0 26360.0 167255.0 ;
      RECT  25655.0 168600.0 26360.0 169945.0 ;
      RECT  25655.0 171290.0 26360.0 169945.0 ;
      RECT  25655.0 171290.0 26360.0 172635.0 ;
      RECT  25655.0 173980.0 26360.0 172635.0 ;
      RECT  25655.0 173980.0 26360.0 175325.0 ;
      RECT  25655.0 176670.0 26360.0 175325.0 ;
      RECT  25655.0 176670.0 26360.0 178015.0 ;
      RECT  25655.0 179360.0 26360.0 178015.0 ;
      RECT  25655.0 179360.0 26360.0 180705.0 ;
      RECT  25655.0 182050.0 26360.0 180705.0 ;
      RECT  25655.0 182050.0 26360.0 183395.0 ;
      RECT  25655.0 184740.0 26360.0 183395.0 ;
      RECT  25655.0 184740.0 26360.0 186085.0 ;
      RECT  25655.0 187430.0 26360.0 186085.0 ;
      RECT  25655.0 187430.0 26360.0 188775.0 ;
      RECT  25655.0 190120.0 26360.0 188775.0 ;
      RECT  25655.0 190120.0 26360.0 191465.0 ;
      RECT  25655.0 192810.0 26360.0 191465.0 ;
      RECT  25655.0 192810.0 26360.0 194155.0 ;
      RECT  25655.0 195500.0 26360.0 194155.0 ;
      RECT  25655.0 195500.0 26360.0 196845.0 ;
      RECT  25655.0 198190.0 26360.0 196845.0 ;
      RECT  25655.0 198190.0 26360.0 199535.0 ;
      RECT  25655.0 200880.0 26360.0 199535.0 ;
      RECT  25655.0 200880.0 26360.0 202225.0 ;
      RECT  25655.0 203570.0 26360.0 202225.0 ;
      RECT  25655.0 203570.0 26360.0 204915.0 ;
      RECT  25655.0 206260.0 26360.0 204915.0 ;
      RECT  26360.0 34100.0 27065.0 35445.0 ;
      RECT  26360.0 36790.0 27065.0 35445.0 ;
      RECT  26360.0 36790.0 27065.0 38135.0 ;
      RECT  26360.0 39480.0 27065.0 38135.0 ;
      RECT  26360.0 39480.0 27065.0 40825.0 ;
      RECT  26360.0 42170.0 27065.0 40825.0 ;
      RECT  26360.0 42170.0 27065.0 43515.0 ;
      RECT  26360.0 44860.0 27065.0 43515.0 ;
      RECT  26360.0 44860.0 27065.0 46205.0 ;
      RECT  26360.0 47550.0 27065.0 46205.0 ;
      RECT  26360.0 47550.0 27065.0 48895.0 ;
      RECT  26360.0 50240.0 27065.0 48895.0 ;
      RECT  26360.0 50240.0 27065.0 51585.0 ;
      RECT  26360.0 52930.0 27065.0 51585.0 ;
      RECT  26360.0 52930.0 27065.0 54275.0 ;
      RECT  26360.0 55620.0 27065.0 54275.0 ;
      RECT  26360.0 55620.0 27065.0 56965.0 ;
      RECT  26360.0 58310.0 27065.0 56965.0 ;
      RECT  26360.0 58310.0 27065.0 59655.0 ;
      RECT  26360.0 61000.0 27065.0 59655.0 ;
      RECT  26360.0 61000.0 27065.0 62345.0 ;
      RECT  26360.0 63690.0 27065.0 62345.0 ;
      RECT  26360.0 63690.0 27065.0 65035.0 ;
      RECT  26360.0 66380.0 27065.0 65035.0 ;
      RECT  26360.0 66380.0 27065.0 67725.0 ;
      RECT  26360.0 69070.0 27065.0 67725.0 ;
      RECT  26360.0 69070.0 27065.0 70415.0 ;
      RECT  26360.0 71760.0 27065.0 70415.0 ;
      RECT  26360.0 71760.0 27065.0 73105.0 ;
      RECT  26360.0 74450.0 27065.0 73105.0 ;
      RECT  26360.0 74450.0 27065.0 75795.0 ;
      RECT  26360.0 77140.0 27065.0 75795.0 ;
      RECT  26360.0 77140.0 27065.0 78485.0 ;
      RECT  26360.0 79830.0 27065.0 78485.0 ;
      RECT  26360.0 79830.0 27065.0 81175.0 ;
      RECT  26360.0 82520.0 27065.0 81175.0 ;
      RECT  26360.0 82520.0 27065.0 83865.0 ;
      RECT  26360.0 85210.0 27065.0 83865.0 ;
      RECT  26360.0 85210.0 27065.0 86555.0 ;
      RECT  26360.0 87900.0 27065.0 86555.0 ;
      RECT  26360.0 87900.0 27065.0 89245.0 ;
      RECT  26360.0 90590.0 27065.0 89245.0 ;
      RECT  26360.0 90590.0 27065.0 91935.0 ;
      RECT  26360.0 93280.0 27065.0 91935.0 ;
      RECT  26360.0 93280.0 27065.0 94625.0 ;
      RECT  26360.0 95970.0 27065.0 94625.0 ;
      RECT  26360.0 95970.0 27065.0 97315.0 ;
      RECT  26360.0 98660.0 27065.0 97315.0 ;
      RECT  26360.0 98660.0 27065.0 100005.0 ;
      RECT  26360.0 101350.0 27065.0 100005.0 ;
      RECT  26360.0 101350.0 27065.0 102695.0 ;
      RECT  26360.0 104040.0 27065.0 102695.0 ;
      RECT  26360.0 104040.0 27065.0 105385.0 ;
      RECT  26360.0 106730.0 27065.0 105385.0 ;
      RECT  26360.0 106730.0 27065.0 108075.0 ;
      RECT  26360.0 109420.0 27065.0 108075.0 ;
      RECT  26360.0 109420.0 27065.0 110765.0 ;
      RECT  26360.0 112110.0 27065.0 110765.0 ;
      RECT  26360.0 112110.0 27065.0 113455.0 ;
      RECT  26360.0 114800.0 27065.0 113455.0 ;
      RECT  26360.0 114800.0 27065.0 116145.0 ;
      RECT  26360.0 117490.0 27065.0 116145.0 ;
      RECT  26360.0 117490.0 27065.0 118835.0 ;
      RECT  26360.0 120180.0 27065.0 118835.0 ;
      RECT  26360.0 120180.0 27065.0 121525.0 ;
      RECT  26360.0 122870.0 27065.0 121525.0 ;
      RECT  26360.0 122870.0 27065.0 124215.0 ;
      RECT  26360.0 125560.0 27065.0 124215.0 ;
      RECT  26360.0 125560.0 27065.0 126905.0 ;
      RECT  26360.0 128250.0 27065.0 126905.0 ;
      RECT  26360.0 128250.0 27065.0 129595.0 ;
      RECT  26360.0 130940.0 27065.0 129595.0 ;
      RECT  26360.0 130940.0 27065.0 132285.0 ;
      RECT  26360.0 133630.0 27065.0 132285.0 ;
      RECT  26360.0 133630.0 27065.0 134975.0 ;
      RECT  26360.0 136320.0 27065.0 134975.0 ;
      RECT  26360.0 136320.0 27065.0 137665.0 ;
      RECT  26360.0 139010.0 27065.0 137665.0 ;
      RECT  26360.0 139010.0 27065.0 140355.0 ;
      RECT  26360.0 141700.0 27065.0 140355.0 ;
      RECT  26360.0 141700.0 27065.0 143045.0 ;
      RECT  26360.0 144390.0 27065.0 143045.0 ;
      RECT  26360.0 144390.0 27065.0 145735.0 ;
      RECT  26360.0 147080.0 27065.0 145735.0 ;
      RECT  26360.0 147080.0 27065.0 148425.0 ;
      RECT  26360.0 149770.0 27065.0 148425.0 ;
      RECT  26360.0 149770.0 27065.0 151115.0 ;
      RECT  26360.0 152460.0 27065.0 151115.0 ;
      RECT  26360.0 152460.0 27065.0 153805.0 ;
      RECT  26360.0 155150.0 27065.0 153805.0 ;
      RECT  26360.0 155150.0 27065.0 156495.0 ;
      RECT  26360.0 157840.0 27065.0 156495.0 ;
      RECT  26360.0 157840.0 27065.0 159185.0 ;
      RECT  26360.0 160530.0 27065.0 159185.0 ;
      RECT  26360.0 160530.0 27065.0 161875.0 ;
      RECT  26360.0 163220.0 27065.0 161875.0 ;
      RECT  26360.0 163220.0 27065.0 164565.0 ;
      RECT  26360.0 165910.0 27065.0 164565.0 ;
      RECT  26360.0 165910.0 27065.0 167255.0 ;
      RECT  26360.0 168600.0 27065.0 167255.0 ;
      RECT  26360.0 168600.0 27065.0 169945.0 ;
      RECT  26360.0 171290.0 27065.0 169945.0 ;
      RECT  26360.0 171290.0 27065.0 172635.0 ;
      RECT  26360.0 173980.0 27065.0 172635.0 ;
      RECT  26360.0 173980.0 27065.0 175325.0 ;
      RECT  26360.0 176670.0 27065.0 175325.0 ;
      RECT  26360.0 176670.0 27065.0 178015.0 ;
      RECT  26360.0 179360.0 27065.0 178015.0 ;
      RECT  26360.0 179360.0 27065.0 180705.0 ;
      RECT  26360.0 182050.0 27065.0 180705.0 ;
      RECT  26360.0 182050.0 27065.0 183395.0 ;
      RECT  26360.0 184740.0 27065.0 183395.0 ;
      RECT  26360.0 184740.0 27065.0 186085.0 ;
      RECT  26360.0 187430.0 27065.0 186085.0 ;
      RECT  26360.0 187430.0 27065.0 188775.0 ;
      RECT  26360.0 190120.0 27065.0 188775.0 ;
      RECT  26360.0 190120.0 27065.0 191465.0 ;
      RECT  26360.0 192810.0 27065.0 191465.0 ;
      RECT  26360.0 192810.0 27065.0 194155.0 ;
      RECT  26360.0 195500.0 27065.0 194155.0 ;
      RECT  26360.0 195500.0 27065.0 196845.0 ;
      RECT  26360.0 198190.0 27065.0 196845.0 ;
      RECT  26360.0 198190.0 27065.0 199535.0 ;
      RECT  26360.0 200880.0 27065.0 199535.0 ;
      RECT  26360.0 200880.0 27065.0 202225.0 ;
      RECT  26360.0 203570.0 27065.0 202225.0 ;
      RECT  26360.0 203570.0 27065.0 204915.0 ;
      RECT  26360.0 206260.0 27065.0 204915.0 ;
      RECT  27065.0 34100.0 27770.0 35445.0 ;
      RECT  27065.0 36790.0 27770.0 35445.0 ;
      RECT  27065.0 36790.0 27770.0 38135.0 ;
      RECT  27065.0 39480.0 27770.0 38135.0 ;
      RECT  27065.0 39480.0 27770.0 40825.0 ;
      RECT  27065.0 42170.0 27770.0 40825.0 ;
      RECT  27065.0 42170.0 27770.0 43515.0 ;
      RECT  27065.0 44860.0 27770.0 43515.0 ;
      RECT  27065.0 44860.0 27770.0 46205.0 ;
      RECT  27065.0 47550.0 27770.0 46205.0 ;
      RECT  27065.0 47550.0 27770.0 48895.0 ;
      RECT  27065.0 50240.0 27770.0 48895.0 ;
      RECT  27065.0 50240.0 27770.0 51585.0 ;
      RECT  27065.0 52930.0 27770.0 51585.0 ;
      RECT  27065.0 52930.0 27770.0 54275.0 ;
      RECT  27065.0 55620.0 27770.0 54275.0 ;
      RECT  27065.0 55620.0 27770.0 56965.0 ;
      RECT  27065.0 58310.0 27770.0 56965.0 ;
      RECT  27065.0 58310.0 27770.0 59655.0 ;
      RECT  27065.0 61000.0 27770.0 59655.0 ;
      RECT  27065.0 61000.0 27770.0 62345.0 ;
      RECT  27065.0 63690.0 27770.0 62345.0 ;
      RECT  27065.0 63690.0 27770.0 65035.0 ;
      RECT  27065.0 66380.0 27770.0 65035.0 ;
      RECT  27065.0 66380.0 27770.0 67725.0 ;
      RECT  27065.0 69070.0 27770.0 67725.0 ;
      RECT  27065.0 69070.0 27770.0 70415.0 ;
      RECT  27065.0 71760.0 27770.0 70415.0 ;
      RECT  27065.0 71760.0 27770.0 73105.0 ;
      RECT  27065.0 74450.0 27770.0 73105.0 ;
      RECT  27065.0 74450.0 27770.0 75795.0 ;
      RECT  27065.0 77140.0 27770.0 75795.0 ;
      RECT  27065.0 77140.0 27770.0 78485.0 ;
      RECT  27065.0 79830.0 27770.0 78485.0 ;
      RECT  27065.0 79830.0 27770.0 81175.0 ;
      RECT  27065.0 82520.0 27770.0 81175.0 ;
      RECT  27065.0 82520.0 27770.0 83865.0 ;
      RECT  27065.0 85210.0 27770.0 83865.0 ;
      RECT  27065.0 85210.0 27770.0 86555.0 ;
      RECT  27065.0 87900.0 27770.0 86555.0 ;
      RECT  27065.0 87900.0 27770.0 89245.0 ;
      RECT  27065.0 90590.0 27770.0 89245.0 ;
      RECT  27065.0 90590.0 27770.0 91935.0 ;
      RECT  27065.0 93280.0 27770.0 91935.0 ;
      RECT  27065.0 93280.0 27770.0 94625.0 ;
      RECT  27065.0 95970.0 27770.0 94625.0 ;
      RECT  27065.0 95970.0 27770.0 97315.0 ;
      RECT  27065.0 98660.0 27770.0 97315.0 ;
      RECT  27065.0 98660.0 27770.0 100005.0 ;
      RECT  27065.0 101350.0 27770.0 100005.0 ;
      RECT  27065.0 101350.0 27770.0 102695.0 ;
      RECT  27065.0 104040.0 27770.0 102695.0 ;
      RECT  27065.0 104040.0 27770.0 105385.0 ;
      RECT  27065.0 106730.0 27770.0 105385.0 ;
      RECT  27065.0 106730.0 27770.0 108075.0 ;
      RECT  27065.0 109420.0 27770.0 108075.0 ;
      RECT  27065.0 109420.0 27770.0 110765.0 ;
      RECT  27065.0 112110.0 27770.0 110765.0 ;
      RECT  27065.0 112110.0 27770.0 113455.0 ;
      RECT  27065.0 114800.0 27770.0 113455.0 ;
      RECT  27065.0 114800.0 27770.0 116145.0 ;
      RECT  27065.0 117490.0 27770.0 116145.0 ;
      RECT  27065.0 117490.0 27770.0 118835.0 ;
      RECT  27065.0 120180.0 27770.0 118835.0 ;
      RECT  27065.0 120180.0 27770.0 121525.0 ;
      RECT  27065.0 122870.0 27770.0 121525.0 ;
      RECT  27065.0 122870.0 27770.0 124215.0 ;
      RECT  27065.0 125560.0 27770.0 124215.0 ;
      RECT  27065.0 125560.0 27770.0 126905.0 ;
      RECT  27065.0 128250.0 27770.0 126905.0 ;
      RECT  27065.0 128250.0 27770.0 129595.0 ;
      RECT  27065.0 130940.0 27770.0 129595.0 ;
      RECT  27065.0 130940.0 27770.0 132285.0 ;
      RECT  27065.0 133630.0 27770.0 132285.0 ;
      RECT  27065.0 133630.0 27770.0 134975.0 ;
      RECT  27065.0 136320.0 27770.0 134975.0 ;
      RECT  27065.0 136320.0 27770.0 137665.0 ;
      RECT  27065.0 139010.0 27770.0 137665.0 ;
      RECT  27065.0 139010.0 27770.0 140355.0 ;
      RECT  27065.0 141700.0 27770.0 140355.0 ;
      RECT  27065.0 141700.0 27770.0 143045.0 ;
      RECT  27065.0 144390.0 27770.0 143045.0 ;
      RECT  27065.0 144390.0 27770.0 145735.0 ;
      RECT  27065.0 147080.0 27770.0 145735.0 ;
      RECT  27065.0 147080.0 27770.0 148425.0 ;
      RECT  27065.0 149770.0 27770.0 148425.0 ;
      RECT  27065.0 149770.0 27770.0 151115.0 ;
      RECT  27065.0 152460.0 27770.0 151115.0 ;
      RECT  27065.0 152460.0 27770.0 153805.0 ;
      RECT  27065.0 155150.0 27770.0 153805.0 ;
      RECT  27065.0 155150.0 27770.0 156495.0 ;
      RECT  27065.0 157840.0 27770.0 156495.0 ;
      RECT  27065.0 157840.0 27770.0 159185.0 ;
      RECT  27065.0 160530.0 27770.0 159185.0 ;
      RECT  27065.0 160530.0 27770.0 161875.0 ;
      RECT  27065.0 163220.0 27770.0 161875.0 ;
      RECT  27065.0 163220.0 27770.0 164565.0 ;
      RECT  27065.0 165910.0 27770.0 164565.0 ;
      RECT  27065.0 165910.0 27770.0 167255.0 ;
      RECT  27065.0 168600.0 27770.0 167255.0 ;
      RECT  27065.0 168600.0 27770.0 169945.0 ;
      RECT  27065.0 171290.0 27770.0 169945.0 ;
      RECT  27065.0 171290.0 27770.0 172635.0 ;
      RECT  27065.0 173980.0 27770.0 172635.0 ;
      RECT  27065.0 173980.0 27770.0 175325.0 ;
      RECT  27065.0 176670.0 27770.0 175325.0 ;
      RECT  27065.0 176670.0 27770.0 178015.0 ;
      RECT  27065.0 179360.0 27770.0 178015.0 ;
      RECT  27065.0 179360.0 27770.0 180705.0 ;
      RECT  27065.0 182050.0 27770.0 180705.0 ;
      RECT  27065.0 182050.0 27770.0 183395.0 ;
      RECT  27065.0 184740.0 27770.0 183395.0 ;
      RECT  27065.0 184740.0 27770.0 186085.0 ;
      RECT  27065.0 187430.0 27770.0 186085.0 ;
      RECT  27065.0 187430.0 27770.0 188775.0 ;
      RECT  27065.0 190120.0 27770.0 188775.0 ;
      RECT  27065.0 190120.0 27770.0 191465.0 ;
      RECT  27065.0 192810.0 27770.0 191465.0 ;
      RECT  27065.0 192810.0 27770.0 194155.0 ;
      RECT  27065.0 195500.0 27770.0 194155.0 ;
      RECT  27065.0 195500.0 27770.0 196845.0 ;
      RECT  27065.0 198190.0 27770.0 196845.0 ;
      RECT  27065.0 198190.0 27770.0 199535.0 ;
      RECT  27065.0 200880.0 27770.0 199535.0 ;
      RECT  27065.0 200880.0 27770.0 202225.0 ;
      RECT  27065.0 203570.0 27770.0 202225.0 ;
      RECT  27065.0 203570.0 27770.0 204915.0 ;
      RECT  27065.0 206260.0 27770.0 204915.0 ;
      RECT  27770.0 34100.0 28475.0 35445.0 ;
      RECT  27770.0 36790.0 28475.0 35445.0 ;
      RECT  27770.0 36790.0 28475.0 38135.0 ;
      RECT  27770.0 39480.0 28475.0 38135.0 ;
      RECT  27770.0 39480.0 28475.0 40825.0 ;
      RECT  27770.0 42170.0 28475.0 40825.0 ;
      RECT  27770.0 42170.0 28475.0 43515.0 ;
      RECT  27770.0 44860.0 28475.0 43515.0 ;
      RECT  27770.0 44860.0 28475.0 46205.0 ;
      RECT  27770.0 47550.0 28475.0 46205.0 ;
      RECT  27770.0 47550.0 28475.0 48895.0 ;
      RECT  27770.0 50240.0 28475.0 48895.0 ;
      RECT  27770.0 50240.0 28475.0 51585.0 ;
      RECT  27770.0 52930.0 28475.0 51585.0 ;
      RECT  27770.0 52930.0 28475.0 54275.0 ;
      RECT  27770.0 55620.0 28475.0 54275.0 ;
      RECT  27770.0 55620.0 28475.0 56965.0 ;
      RECT  27770.0 58310.0 28475.0 56965.0 ;
      RECT  27770.0 58310.0 28475.0 59655.0 ;
      RECT  27770.0 61000.0 28475.0 59655.0 ;
      RECT  27770.0 61000.0 28475.0 62345.0 ;
      RECT  27770.0 63690.0 28475.0 62345.0 ;
      RECT  27770.0 63690.0 28475.0 65035.0 ;
      RECT  27770.0 66380.0 28475.0 65035.0 ;
      RECT  27770.0 66380.0 28475.0 67725.0 ;
      RECT  27770.0 69070.0 28475.0 67725.0 ;
      RECT  27770.0 69070.0 28475.0 70415.0 ;
      RECT  27770.0 71760.0 28475.0 70415.0 ;
      RECT  27770.0 71760.0 28475.0 73105.0 ;
      RECT  27770.0 74450.0 28475.0 73105.0 ;
      RECT  27770.0 74450.0 28475.0 75795.0 ;
      RECT  27770.0 77140.0 28475.0 75795.0 ;
      RECT  27770.0 77140.0 28475.0 78485.0 ;
      RECT  27770.0 79830.0 28475.0 78485.0 ;
      RECT  27770.0 79830.0 28475.0 81175.0 ;
      RECT  27770.0 82520.0 28475.0 81175.0 ;
      RECT  27770.0 82520.0 28475.0 83865.0 ;
      RECT  27770.0 85210.0 28475.0 83865.0 ;
      RECT  27770.0 85210.0 28475.0 86555.0 ;
      RECT  27770.0 87900.0 28475.0 86555.0 ;
      RECT  27770.0 87900.0 28475.0 89245.0 ;
      RECT  27770.0 90590.0 28475.0 89245.0 ;
      RECT  27770.0 90590.0 28475.0 91935.0 ;
      RECT  27770.0 93280.0 28475.0 91935.0 ;
      RECT  27770.0 93280.0 28475.0 94625.0 ;
      RECT  27770.0 95970.0 28475.0 94625.0 ;
      RECT  27770.0 95970.0 28475.0 97315.0 ;
      RECT  27770.0 98660.0 28475.0 97315.0 ;
      RECT  27770.0 98660.0 28475.0 100005.0 ;
      RECT  27770.0 101350.0 28475.0 100005.0 ;
      RECT  27770.0 101350.0 28475.0 102695.0 ;
      RECT  27770.0 104040.0 28475.0 102695.0 ;
      RECT  27770.0 104040.0 28475.0 105385.0 ;
      RECT  27770.0 106730.0 28475.0 105385.0 ;
      RECT  27770.0 106730.0 28475.0 108075.0 ;
      RECT  27770.0 109420.0 28475.0 108075.0 ;
      RECT  27770.0 109420.0 28475.0 110765.0 ;
      RECT  27770.0 112110.0 28475.0 110765.0 ;
      RECT  27770.0 112110.0 28475.0 113455.0 ;
      RECT  27770.0 114800.0 28475.0 113455.0 ;
      RECT  27770.0 114800.0 28475.0 116145.0 ;
      RECT  27770.0 117490.0 28475.0 116145.0 ;
      RECT  27770.0 117490.0 28475.0 118835.0 ;
      RECT  27770.0 120180.0 28475.0 118835.0 ;
      RECT  27770.0 120180.0 28475.0 121525.0 ;
      RECT  27770.0 122870.0 28475.0 121525.0 ;
      RECT  27770.0 122870.0 28475.0 124215.0 ;
      RECT  27770.0 125560.0 28475.0 124215.0 ;
      RECT  27770.0 125560.0 28475.0 126905.0 ;
      RECT  27770.0 128250.0 28475.0 126905.0 ;
      RECT  27770.0 128250.0 28475.0 129595.0 ;
      RECT  27770.0 130940.0 28475.0 129595.0 ;
      RECT  27770.0 130940.0 28475.0 132285.0 ;
      RECT  27770.0 133630.0 28475.0 132285.0 ;
      RECT  27770.0 133630.0 28475.0 134975.0 ;
      RECT  27770.0 136320.0 28475.0 134975.0 ;
      RECT  27770.0 136320.0 28475.0 137665.0 ;
      RECT  27770.0 139010.0 28475.0 137665.0 ;
      RECT  27770.0 139010.0 28475.0 140355.0 ;
      RECT  27770.0 141700.0 28475.0 140355.0 ;
      RECT  27770.0 141700.0 28475.0 143045.0 ;
      RECT  27770.0 144390.0 28475.0 143045.0 ;
      RECT  27770.0 144390.0 28475.0 145735.0 ;
      RECT  27770.0 147080.0 28475.0 145735.0 ;
      RECT  27770.0 147080.0 28475.0 148425.0 ;
      RECT  27770.0 149770.0 28475.0 148425.0 ;
      RECT  27770.0 149770.0 28475.0 151115.0 ;
      RECT  27770.0 152460.0 28475.0 151115.0 ;
      RECT  27770.0 152460.0 28475.0 153805.0 ;
      RECT  27770.0 155150.0 28475.0 153805.0 ;
      RECT  27770.0 155150.0 28475.0 156495.0 ;
      RECT  27770.0 157840.0 28475.0 156495.0 ;
      RECT  27770.0 157840.0 28475.0 159185.0 ;
      RECT  27770.0 160530.0 28475.0 159185.0 ;
      RECT  27770.0 160530.0 28475.0 161875.0 ;
      RECT  27770.0 163220.0 28475.0 161875.0 ;
      RECT  27770.0 163220.0 28475.0 164565.0 ;
      RECT  27770.0 165910.0 28475.0 164565.0 ;
      RECT  27770.0 165910.0 28475.0 167255.0 ;
      RECT  27770.0 168600.0 28475.0 167255.0 ;
      RECT  27770.0 168600.0 28475.0 169945.0 ;
      RECT  27770.0 171290.0 28475.0 169945.0 ;
      RECT  27770.0 171290.0 28475.0 172635.0 ;
      RECT  27770.0 173980.0 28475.0 172635.0 ;
      RECT  27770.0 173980.0 28475.0 175325.0 ;
      RECT  27770.0 176670.0 28475.0 175325.0 ;
      RECT  27770.0 176670.0 28475.0 178015.0 ;
      RECT  27770.0 179360.0 28475.0 178015.0 ;
      RECT  27770.0 179360.0 28475.0 180705.0 ;
      RECT  27770.0 182050.0 28475.0 180705.0 ;
      RECT  27770.0 182050.0 28475.0 183395.0 ;
      RECT  27770.0 184740.0 28475.0 183395.0 ;
      RECT  27770.0 184740.0 28475.0 186085.0 ;
      RECT  27770.0 187430.0 28475.0 186085.0 ;
      RECT  27770.0 187430.0 28475.0 188775.0 ;
      RECT  27770.0 190120.0 28475.0 188775.0 ;
      RECT  27770.0 190120.0 28475.0 191465.0 ;
      RECT  27770.0 192810.0 28475.0 191465.0 ;
      RECT  27770.0 192810.0 28475.0 194155.0 ;
      RECT  27770.0 195500.0 28475.0 194155.0 ;
      RECT  27770.0 195500.0 28475.0 196845.0 ;
      RECT  27770.0 198190.0 28475.0 196845.0 ;
      RECT  27770.0 198190.0 28475.0 199535.0 ;
      RECT  27770.0 200880.0 28475.0 199535.0 ;
      RECT  27770.0 200880.0 28475.0 202225.0 ;
      RECT  27770.0 203570.0 28475.0 202225.0 ;
      RECT  27770.0 203570.0 28475.0 204915.0 ;
      RECT  27770.0 206260.0 28475.0 204915.0 ;
      RECT  28475.0 34100.0 29180.0 35445.0 ;
      RECT  28475.0 36790.0 29180.0 35445.0 ;
      RECT  28475.0 36790.0 29180.0 38135.0 ;
      RECT  28475.0 39480.0 29180.0 38135.0 ;
      RECT  28475.0 39480.0 29180.0 40825.0 ;
      RECT  28475.0 42170.0 29180.0 40825.0 ;
      RECT  28475.0 42170.0 29180.0 43515.0 ;
      RECT  28475.0 44860.0 29180.0 43515.0 ;
      RECT  28475.0 44860.0 29180.0 46205.0 ;
      RECT  28475.0 47550.0 29180.0 46205.0 ;
      RECT  28475.0 47550.0 29180.0 48895.0 ;
      RECT  28475.0 50240.0 29180.0 48895.0 ;
      RECT  28475.0 50240.0 29180.0 51585.0 ;
      RECT  28475.0 52930.0 29180.0 51585.0 ;
      RECT  28475.0 52930.0 29180.0 54275.0 ;
      RECT  28475.0 55620.0 29180.0 54275.0 ;
      RECT  28475.0 55620.0 29180.0 56965.0 ;
      RECT  28475.0 58310.0 29180.0 56965.0 ;
      RECT  28475.0 58310.0 29180.0 59655.0 ;
      RECT  28475.0 61000.0 29180.0 59655.0 ;
      RECT  28475.0 61000.0 29180.0 62345.0 ;
      RECT  28475.0 63690.0 29180.0 62345.0 ;
      RECT  28475.0 63690.0 29180.0 65035.0 ;
      RECT  28475.0 66380.0 29180.0 65035.0 ;
      RECT  28475.0 66380.0 29180.0 67725.0 ;
      RECT  28475.0 69070.0 29180.0 67725.0 ;
      RECT  28475.0 69070.0 29180.0 70415.0 ;
      RECT  28475.0 71760.0 29180.0 70415.0 ;
      RECT  28475.0 71760.0 29180.0 73105.0 ;
      RECT  28475.0 74450.0 29180.0 73105.0 ;
      RECT  28475.0 74450.0 29180.0 75795.0 ;
      RECT  28475.0 77140.0 29180.0 75795.0 ;
      RECT  28475.0 77140.0 29180.0 78485.0 ;
      RECT  28475.0 79830.0 29180.0 78485.0 ;
      RECT  28475.0 79830.0 29180.0 81175.0 ;
      RECT  28475.0 82520.0 29180.0 81175.0 ;
      RECT  28475.0 82520.0 29180.0 83865.0 ;
      RECT  28475.0 85210.0 29180.0 83865.0 ;
      RECT  28475.0 85210.0 29180.0 86555.0 ;
      RECT  28475.0 87900.0 29180.0 86555.0 ;
      RECT  28475.0 87900.0 29180.0 89245.0 ;
      RECT  28475.0 90590.0 29180.0 89245.0 ;
      RECT  28475.0 90590.0 29180.0 91935.0 ;
      RECT  28475.0 93280.0 29180.0 91935.0 ;
      RECT  28475.0 93280.0 29180.0 94625.0 ;
      RECT  28475.0 95970.0 29180.0 94625.0 ;
      RECT  28475.0 95970.0 29180.0 97315.0 ;
      RECT  28475.0 98660.0 29180.0 97315.0 ;
      RECT  28475.0 98660.0 29180.0 100005.0 ;
      RECT  28475.0 101350.0 29180.0 100005.0 ;
      RECT  28475.0 101350.0 29180.0 102695.0 ;
      RECT  28475.0 104040.0 29180.0 102695.0 ;
      RECT  28475.0 104040.0 29180.0 105385.0 ;
      RECT  28475.0 106730.0 29180.0 105385.0 ;
      RECT  28475.0 106730.0 29180.0 108075.0 ;
      RECT  28475.0 109420.0 29180.0 108075.0 ;
      RECT  28475.0 109420.0 29180.0 110765.0 ;
      RECT  28475.0 112110.0 29180.0 110765.0 ;
      RECT  28475.0 112110.0 29180.0 113455.0 ;
      RECT  28475.0 114800.0 29180.0 113455.0 ;
      RECT  28475.0 114800.0 29180.0 116145.0 ;
      RECT  28475.0 117490.0 29180.0 116145.0 ;
      RECT  28475.0 117490.0 29180.0 118835.0 ;
      RECT  28475.0 120180.0 29180.0 118835.0 ;
      RECT  28475.0 120180.0 29180.0 121525.0 ;
      RECT  28475.0 122870.0 29180.0 121525.0 ;
      RECT  28475.0 122870.0 29180.0 124215.0 ;
      RECT  28475.0 125560.0 29180.0 124215.0 ;
      RECT  28475.0 125560.0 29180.0 126905.0 ;
      RECT  28475.0 128250.0 29180.0 126905.0 ;
      RECT  28475.0 128250.0 29180.0 129595.0 ;
      RECT  28475.0 130940.0 29180.0 129595.0 ;
      RECT  28475.0 130940.0 29180.0 132285.0 ;
      RECT  28475.0 133630.0 29180.0 132285.0 ;
      RECT  28475.0 133630.0 29180.0 134975.0 ;
      RECT  28475.0 136320.0 29180.0 134975.0 ;
      RECT  28475.0 136320.0 29180.0 137665.0 ;
      RECT  28475.0 139010.0 29180.0 137665.0 ;
      RECT  28475.0 139010.0 29180.0 140355.0 ;
      RECT  28475.0 141700.0 29180.0 140355.0 ;
      RECT  28475.0 141700.0 29180.0 143045.0 ;
      RECT  28475.0 144390.0 29180.0 143045.0 ;
      RECT  28475.0 144390.0 29180.0 145735.0 ;
      RECT  28475.0 147080.0 29180.0 145735.0 ;
      RECT  28475.0 147080.0 29180.0 148425.0 ;
      RECT  28475.0 149770.0 29180.0 148425.0 ;
      RECT  28475.0 149770.0 29180.0 151115.0 ;
      RECT  28475.0 152460.0 29180.0 151115.0 ;
      RECT  28475.0 152460.0 29180.0 153805.0 ;
      RECT  28475.0 155150.0 29180.0 153805.0 ;
      RECT  28475.0 155150.0 29180.0 156495.0 ;
      RECT  28475.0 157840.0 29180.0 156495.0 ;
      RECT  28475.0 157840.0 29180.0 159185.0 ;
      RECT  28475.0 160530.0 29180.0 159185.0 ;
      RECT  28475.0 160530.0 29180.0 161875.0 ;
      RECT  28475.0 163220.0 29180.0 161875.0 ;
      RECT  28475.0 163220.0 29180.0 164565.0 ;
      RECT  28475.0 165910.0 29180.0 164565.0 ;
      RECT  28475.0 165910.0 29180.0 167255.0 ;
      RECT  28475.0 168600.0 29180.0 167255.0 ;
      RECT  28475.0 168600.0 29180.0 169945.0 ;
      RECT  28475.0 171290.0 29180.0 169945.0 ;
      RECT  28475.0 171290.0 29180.0 172635.0 ;
      RECT  28475.0 173980.0 29180.0 172635.0 ;
      RECT  28475.0 173980.0 29180.0 175325.0 ;
      RECT  28475.0 176670.0 29180.0 175325.0 ;
      RECT  28475.0 176670.0 29180.0 178015.0 ;
      RECT  28475.0 179360.0 29180.0 178015.0 ;
      RECT  28475.0 179360.0 29180.0 180705.0 ;
      RECT  28475.0 182050.0 29180.0 180705.0 ;
      RECT  28475.0 182050.0 29180.0 183395.0 ;
      RECT  28475.0 184740.0 29180.0 183395.0 ;
      RECT  28475.0 184740.0 29180.0 186085.0 ;
      RECT  28475.0 187430.0 29180.0 186085.0 ;
      RECT  28475.0 187430.0 29180.0 188775.0 ;
      RECT  28475.0 190120.0 29180.0 188775.0 ;
      RECT  28475.0 190120.0 29180.0 191465.0 ;
      RECT  28475.0 192810.0 29180.0 191465.0 ;
      RECT  28475.0 192810.0 29180.0 194155.0 ;
      RECT  28475.0 195500.0 29180.0 194155.0 ;
      RECT  28475.0 195500.0 29180.0 196845.0 ;
      RECT  28475.0 198190.0 29180.0 196845.0 ;
      RECT  28475.0 198190.0 29180.0 199535.0 ;
      RECT  28475.0 200880.0 29180.0 199535.0 ;
      RECT  28475.0 200880.0 29180.0 202225.0 ;
      RECT  28475.0 203570.0 29180.0 202225.0 ;
      RECT  28475.0 203570.0 29180.0 204915.0 ;
      RECT  28475.0 206260.0 29180.0 204915.0 ;
      RECT  29180.0 34100.0 29885.0 35445.0 ;
      RECT  29180.0 36790.0 29885.0 35445.0 ;
      RECT  29180.0 36790.0 29885.0 38135.0 ;
      RECT  29180.0 39480.0 29885.0 38135.0 ;
      RECT  29180.0 39480.0 29885.0 40825.0 ;
      RECT  29180.0 42170.0 29885.0 40825.0 ;
      RECT  29180.0 42170.0 29885.0 43515.0 ;
      RECT  29180.0 44860.0 29885.0 43515.0 ;
      RECT  29180.0 44860.0 29885.0 46205.0 ;
      RECT  29180.0 47550.0 29885.0 46205.0 ;
      RECT  29180.0 47550.0 29885.0 48895.0 ;
      RECT  29180.0 50240.0 29885.0 48895.0 ;
      RECT  29180.0 50240.0 29885.0 51585.0 ;
      RECT  29180.0 52930.0 29885.0 51585.0 ;
      RECT  29180.0 52930.0 29885.0 54275.0 ;
      RECT  29180.0 55620.0 29885.0 54275.0 ;
      RECT  29180.0 55620.0 29885.0 56965.0 ;
      RECT  29180.0 58310.0 29885.0 56965.0 ;
      RECT  29180.0 58310.0 29885.0 59655.0 ;
      RECT  29180.0 61000.0 29885.0 59655.0 ;
      RECT  29180.0 61000.0 29885.0 62345.0 ;
      RECT  29180.0 63690.0 29885.0 62345.0 ;
      RECT  29180.0 63690.0 29885.0 65035.0 ;
      RECT  29180.0 66380.0 29885.0 65035.0 ;
      RECT  29180.0 66380.0 29885.0 67725.0 ;
      RECT  29180.0 69070.0 29885.0 67725.0 ;
      RECT  29180.0 69070.0 29885.0 70415.0 ;
      RECT  29180.0 71760.0 29885.0 70415.0 ;
      RECT  29180.0 71760.0 29885.0 73105.0 ;
      RECT  29180.0 74450.0 29885.0 73105.0 ;
      RECT  29180.0 74450.0 29885.0 75795.0 ;
      RECT  29180.0 77140.0 29885.0 75795.0 ;
      RECT  29180.0 77140.0 29885.0 78485.0 ;
      RECT  29180.0 79830.0 29885.0 78485.0 ;
      RECT  29180.0 79830.0 29885.0 81175.0 ;
      RECT  29180.0 82520.0 29885.0 81175.0 ;
      RECT  29180.0 82520.0 29885.0 83865.0 ;
      RECT  29180.0 85210.0 29885.0 83865.0 ;
      RECT  29180.0 85210.0 29885.0 86555.0 ;
      RECT  29180.0 87900.0 29885.0 86555.0 ;
      RECT  29180.0 87900.0 29885.0 89245.0 ;
      RECT  29180.0 90590.0 29885.0 89245.0 ;
      RECT  29180.0 90590.0 29885.0 91935.0 ;
      RECT  29180.0 93280.0 29885.0 91935.0 ;
      RECT  29180.0 93280.0 29885.0 94625.0 ;
      RECT  29180.0 95970.0 29885.0 94625.0 ;
      RECT  29180.0 95970.0 29885.0 97315.0 ;
      RECT  29180.0 98660.0 29885.0 97315.0 ;
      RECT  29180.0 98660.0 29885.0 100005.0 ;
      RECT  29180.0 101350.0 29885.0 100005.0 ;
      RECT  29180.0 101350.0 29885.0 102695.0 ;
      RECT  29180.0 104040.0 29885.0 102695.0 ;
      RECT  29180.0 104040.0 29885.0 105385.0 ;
      RECT  29180.0 106730.0 29885.0 105385.0 ;
      RECT  29180.0 106730.0 29885.0 108075.0 ;
      RECT  29180.0 109420.0 29885.0 108075.0 ;
      RECT  29180.0 109420.0 29885.0 110765.0 ;
      RECT  29180.0 112110.0 29885.0 110765.0 ;
      RECT  29180.0 112110.0 29885.0 113455.0 ;
      RECT  29180.0 114800.0 29885.0 113455.0 ;
      RECT  29180.0 114800.0 29885.0 116145.0 ;
      RECT  29180.0 117490.0 29885.0 116145.0 ;
      RECT  29180.0 117490.0 29885.0 118835.0 ;
      RECT  29180.0 120180.0 29885.0 118835.0 ;
      RECT  29180.0 120180.0 29885.0 121525.0 ;
      RECT  29180.0 122870.0 29885.0 121525.0 ;
      RECT  29180.0 122870.0 29885.0 124215.0 ;
      RECT  29180.0 125560.0 29885.0 124215.0 ;
      RECT  29180.0 125560.0 29885.0 126905.0 ;
      RECT  29180.0 128250.0 29885.0 126905.0 ;
      RECT  29180.0 128250.0 29885.0 129595.0 ;
      RECT  29180.0 130940.0 29885.0 129595.0 ;
      RECT  29180.0 130940.0 29885.0 132285.0 ;
      RECT  29180.0 133630.0 29885.0 132285.0 ;
      RECT  29180.0 133630.0 29885.0 134975.0 ;
      RECT  29180.0 136320.0 29885.0 134975.0 ;
      RECT  29180.0 136320.0 29885.0 137665.0 ;
      RECT  29180.0 139010.0 29885.0 137665.0 ;
      RECT  29180.0 139010.0 29885.0 140355.0 ;
      RECT  29180.0 141700.0 29885.0 140355.0 ;
      RECT  29180.0 141700.0 29885.0 143045.0 ;
      RECT  29180.0 144390.0 29885.0 143045.0 ;
      RECT  29180.0 144390.0 29885.0 145735.0 ;
      RECT  29180.0 147080.0 29885.0 145735.0 ;
      RECT  29180.0 147080.0 29885.0 148425.0 ;
      RECT  29180.0 149770.0 29885.0 148425.0 ;
      RECT  29180.0 149770.0 29885.0 151115.0 ;
      RECT  29180.0 152460.0 29885.0 151115.0 ;
      RECT  29180.0 152460.0 29885.0 153805.0 ;
      RECT  29180.0 155150.0 29885.0 153805.0 ;
      RECT  29180.0 155150.0 29885.0 156495.0 ;
      RECT  29180.0 157840.0 29885.0 156495.0 ;
      RECT  29180.0 157840.0 29885.0 159185.0 ;
      RECT  29180.0 160530.0 29885.0 159185.0 ;
      RECT  29180.0 160530.0 29885.0 161875.0 ;
      RECT  29180.0 163220.0 29885.0 161875.0 ;
      RECT  29180.0 163220.0 29885.0 164565.0 ;
      RECT  29180.0 165910.0 29885.0 164565.0 ;
      RECT  29180.0 165910.0 29885.0 167255.0 ;
      RECT  29180.0 168600.0 29885.0 167255.0 ;
      RECT  29180.0 168600.0 29885.0 169945.0 ;
      RECT  29180.0 171290.0 29885.0 169945.0 ;
      RECT  29180.0 171290.0 29885.0 172635.0 ;
      RECT  29180.0 173980.0 29885.0 172635.0 ;
      RECT  29180.0 173980.0 29885.0 175325.0 ;
      RECT  29180.0 176670.0 29885.0 175325.0 ;
      RECT  29180.0 176670.0 29885.0 178015.0 ;
      RECT  29180.0 179360.0 29885.0 178015.0 ;
      RECT  29180.0 179360.0 29885.0 180705.0 ;
      RECT  29180.0 182050.0 29885.0 180705.0 ;
      RECT  29180.0 182050.0 29885.0 183395.0 ;
      RECT  29180.0 184740.0 29885.0 183395.0 ;
      RECT  29180.0 184740.0 29885.0 186085.0 ;
      RECT  29180.0 187430.0 29885.0 186085.0 ;
      RECT  29180.0 187430.0 29885.0 188775.0 ;
      RECT  29180.0 190120.0 29885.0 188775.0 ;
      RECT  29180.0 190120.0 29885.0 191465.0 ;
      RECT  29180.0 192810.0 29885.0 191465.0 ;
      RECT  29180.0 192810.0 29885.0 194155.0 ;
      RECT  29180.0 195500.0 29885.0 194155.0 ;
      RECT  29180.0 195500.0 29885.0 196845.0 ;
      RECT  29180.0 198190.0 29885.0 196845.0 ;
      RECT  29180.0 198190.0 29885.0 199535.0 ;
      RECT  29180.0 200880.0 29885.0 199535.0 ;
      RECT  29180.0 200880.0 29885.0 202225.0 ;
      RECT  29180.0 203570.0 29885.0 202225.0 ;
      RECT  29180.0 203570.0 29885.0 204915.0 ;
      RECT  29180.0 206260.0 29885.0 204915.0 ;
      RECT  29885.0 34100.0 30590.0 35445.0 ;
      RECT  29885.0 36790.0 30590.0 35445.0 ;
      RECT  29885.0 36790.0 30590.0 38135.0 ;
      RECT  29885.0 39480.0 30590.0 38135.0 ;
      RECT  29885.0 39480.0 30590.0 40825.0 ;
      RECT  29885.0 42170.0 30590.0 40825.0 ;
      RECT  29885.0 42170.0 30590.0 43515.0 ;
      RECT  29885.0 44860.0 30590.0 43515.0 ;
      RECT  29885.0 44860.0 30590.0 46205.0 ;
      RECT  29885.0 47550.0 30590.0 46205.0 ;
      RECT  29885.0 47550.0 30590.0 48895.0 ;
      RECT  29885.0 50240.0 30590.0 48895.0 ;
      RECT  29885.0 50240.0 30590.0 51585.0 ;
      RECT  29885.0 52930.0 30590.0 51585.0 ;
      RECT  29885.0 52930.0 30590.0 54275.0 ;
      RECT  29885.0 55620.0 30590.0 54275.0 ;
      RECT  29885.0 55620.0 30590.0 56965.0 ;
      RECT  29885.0 58310.0 30590.0 56965.0 ;
      RECT  29885.0 58310.0 30590.0 59655.0 ;
      RECT  29885.0 61000.0 30590.0 59655.0 ;
      RECT  29885.0 61000.0 30590.0 62345.0 ;
      RECT  29885.0 63690.0 30590.0 62345.0 ;
      RECT  29885.0 63690.0 30590.0 65035.0 ;
      RECT  29885.0 66380.0 30590.0 65035.0 ;
      RECT  29885.0 66380.0 30590.0 67725.0 ;
      RECT  29885.0 69070.0 30590.0 67725.0 ;
      RECT  29885.0 69070.0 30590.0 70415.0 ;
      RECT  29885.0 71760.0 30590.0 70415.0 ;
      RECT  29885.0 71760.0 30590.0 73105.0 ;
      RECT  29885.0 74450.0 30590.0 73105.0 ;
      RECT  29885.0 74450.0 30590.0 75795.0 ;
      RECT  29885.0 77140.0 30590.0 75795.0 ;
      RECT  29885.0 77140.0 30590.0 78485.0 ;
      RECT  29885.0 79830.0 30590.0 78485.0 ;
      RECT  29885.0 79830.0 30590.0 81175.0 ;
      RECT  29885.0 82520.0 30590.0 81175.0 ;
      RECT  29885.0 82520.0 30590.0 83865.0 ;
      RECT  29885.0 85210.0 30590.0 83865.0 ;
      RECT  29885.0 85210.0 30590.0 86555.0 ;
      RECT  29885.0 87900.0 30590.0 86555.0 ;
      RECT  29885.0 87900.0 30590.0 89245.0 ;
      RECT  29885.0 90590.0 30590.0 89245.0 ;
      RECT  29885.0 90590.0 30590.0 91935.0 ;
      RECT  29885.0 93280.0 30590.0 91935.0 ;
      RECT  29885.0 93280.0 30590.0 94625.0 ;
      RECT  29885.0 95970.0 30590.0 94625.0 ;
      RECT  29885.0 95970.0 30590.0 97315.0 ;
      RECT  29885.0 98660.0 30590.0 97315.0 ;
      RECT  29885.0 98660.0 30590.0 100005.0 ;
      RECT  29885.0 101350.0 30590.0 100005.0 ;
      RECT  29885.0 101350.0 30590.0 102695.0 ;
      RECT  29885.0 104040.0 30590.0 102695.0 ;
      RECT  29885.0 104040.0 30590.0 105385.0 ;
      RECT  29885.0 106730.0 30590.0 105385.0 ;
      RECT  29885.0 106730.0 30590.0 108075.0 ;
      RECT  29885.0 109420.0 30590.0 108075.0 ;
      RECT  29885.0 109420.0 30590.0 110765.0 ;
      RECT  29885.0 112110.0 30590.0 110765.0 ;
      RECT  29885.0 112110.0 30590.0 113455.0 ;
      RECT  29885.0 114800.0 30590.0 113455.0 ;
      RECT  29885.0 114800.0 30590.0 116145.0 ;
      RECT  29885.0 117490.0 30590.0 116145.0 ;
      RECT  29885.0 117490.0 30590.0 118835.0 ;
      RECT  29885.0 120180.0 30590.0 118835.0 ;
      RECT  29885.0 120180.0 30590.0 121525.0 ;
      RECT  29885.0 122870.0 30590.0 121525.0 ;
      RECT  29885.0 122870.0 30590.0 124215.0 ;
      RECT  29885.0 125560.0 30590.0 124215.0 ;
      RECT  29885.0 125560.0 30590.0 126905.0 ;
      RECT  29885.0 128250.0 30590.0 126905.0 ;
      RECT  29885.0 128250.0 30590.0 129595.0 ;
      RECT  29885.0 130940.0 30590.0 129595.0 ;
      RECT  29885.0 130940.0 30590.0 132285.0 ;
      RECT  29885.0 133630.0 30590.0 132285.0 ;
      RECT  29885.0 133630.0 30590.0 134975.0 ;
      RECT  29885.0 136320.0 30590.0 134975.0 ;
      RECT  29885.0 136320.0 30590.0 137665.0 ;
      RECT  29885.0 139010.0 30590.0 137665.0 ;
      RECT  29885.0 139010.0 30590.0 140355.0 ;
      RECT  29885.0 141700.0 30590.0 140355.0 ;
      RECT  29885.0 141700.0 30590.0 143045.0 ;
      RECT  29885.0 144390.0 30590.0 143045.0 ;
      RECT  29885.0 144390.0 30590.0 145735.0 ;
      RECT  29885.0 147080.0 30590.0 145735.0 ;
      RECT  29885.0 147080.0 30590.0 148425.0 ;
      RECT  29885.0 149770.0 30590.0 148425.0 ;
      RECT  29885.0 149770.0 30590.0 151115.0 ;
      RECT  29885.0 152460.0 30590.0 151115.0 ;
      RECT  29885.0 152460.0 30590.0 153805.0 ;
      RECT  29885.0 155150.0 30590.0 153805.0 ;
      RECT  29885.0 155150.0 30590.0 156495.0 ;
      RECT  29885.0 157840.0 30590.0 156495.0 ;
      RECT  29885.0 157840.0 30590.0 159185.0 ;
      RECT  29885.0 160530.0 30590.0 159185.0 ;
      RECT  29885.0 160530.0 30590.0 161875.0 ;
      RECT  29885.0 163220.0 30590.0 161875.0 ;
      RECT  29885.0 163220.0 30590.0 164565.0 ;
      RECT  29885.0 165910.0 30590.0 164565.0 ;
      RECT  29885.0 165910.0 30590.0 167255.0 ;
      RECT  29885.0 168600.0 30590.0 167255.0 ;
      RECT  29885.0 168600.0 30590.0 169945.0 ;
      RECT  29885.0 171290.0 30590.0 169945.0 ;
      RECT  29885.0 171290.0 30590.0 172635.0 ;
      RECT  29885.0 173980.0 30590.0 172635.0 ;
      RECT  29885.0 173980.0 30590.0 175325.0 ;
      RECT  29885.0 176670.0 30590.0 175325.0 ;
      RECT  29885.0 176670.0 30590.0 178015.0 ;
      RECT  29885.0 179360.0 30590.0 178015.0 ;
      RECT  29885.0 179360.0 30590.0 180705.0 ;
      RECT  29885.0 182050.0 30590.0 180705.0 ;
      RECT  29885.0 182050.0 30590.0 183395.0 ;
      RECT  29885.0 184740.0 30590.0 183395.0 ;
      RECT  29885.0 184740.0 30590.0 186085.0 ;
      RECT  29885.0 187430.0 30590.0 186085.0 ;
      RECT  29885.0 187430.0 30590.0 188775.0 ;
      RECT  29885.0 190120.0 30590.0 188775.0 ;
      RECT  29885.0 190120.0 30590.0 191465.0 ;
      RECT  29885.0 192810.0 30590.0 191465.0 ;
      RECT  29885.0 192810.0 30590.0 194155.0 ;
      RECT  29885.0 195500.0 30590.0 194155.0 ;
      RECT  29885.0 195500.0 30590.0 196845.0 ;
      RECT  29885.0 198190.0 30590.0 196845.0 ;
      RECT  29885.0 198190.0 30590.0 199535.0 ;
      RECT  29885.0 200880.0 30590.0 199535.0 ;
      RECT  29885.0 200880.0 30590.0 202225.0 ;
      RECT  29885.0 203570.0 30590.0 202225.0 ;
      RECT  29885.0 203570.0 30590.0 204915.0 ;
      RECT  29885.0 206260.0 30590.0 204915.0 ;
      RECT  30590.0 34100.0 31295.0 35445.0 ;
      RECT  30590.0 36790.0 31295.0 35445.0 ;
      RECT  30590.0 36790.0 31295.0 38135.0 ;
      RECT  30590.0 39480.0 31295.0 38135.0 ;
      RECT  30590.0 39480.0 31295.0 40825.0 ;
      RECT  30590.0 42170.0 31295.0 40825.0 ;
      RECT  30590.0 42170.0 31295.0 43515.0 ;
      RECT  30590.0 44860.0 31295.0 43515.0 ;
      RECT  30590.0 44860.0 31295.0 46205.0 ;
      RECT  30590.0 47550.0 31295.0 46205.0 ;
      RECT  30590.0 47550.0 31295.0 48895.0 ;
      RECT  30590.0 50240.0 31295.0 48895.0 ;
      RECT  30590.0 50240.0 31295.0 51585.0 ;
      RECT  30590.0 52930.0 31295.0 51585.0 ;
      RECT  30590.0 52930.0 31295.0 54275.0 ;
      RECT  30590.0 55620.0 31295.0 54275.0 ;
      RECT  30590.0 55620.0 31295.0 56965.0 ;
      RECT  30590.0 58310.0 31295.0 56965.0 ;
      RECT  30590.0 58310.0 31295.0 59655.0 ;
      RECT  30590.0 61000.0 31295.0 59655.0 ;
      RECT  30590.0 61000.0 31295.0 62345.0 ;
      RECT  30590.0 63690.0 31295.0 62345.0 ;
      RECT  30590.0 63690.0 31295.0 65035.0 ;
      RECT  30590.0 66380.0 31295.0 65035.0 ;
      RECT  30590.0 66380.0 31295.0 67725.0 ;
      RECT  30590.0 69070.0 31295.0 67725.0 ;
      RECT  30590.0 69070.0 31295.0 70415.0 ;
      RECT  30590.0 71760.0 31295.0 70415.0 ;
      RECT  30590.0 71760.0 31295.0 73105.0 ;
      RECT  30590.0 74450.0 31295.0 73105.0 ;
      RECT  30590.0 74450.0 31295.0 75795.0 ;
      RECT  30590.0 77140.0 31295.0 75795.0 ;
      RECT  30590.0 77140.0 31295.0 78485.0 ;
      RECT  30590.0 79830.0 31295.0 78485.0 ;
      RECT  30590.0 79830.0 31295.0 81175.0 ;
      RECT  30590.0 82520.0 31295.0 81175.0 ;
      RECT  30590.0 82520.0 31295.0 83865.0 ;
      RECT  30590.0 85210.0 31295.0 83865.0 ;
      RECT  30590.0 85210.0 31295.0 86555.0 ;
      RECT  30590.0 87900.0 31295.0 86555.0 ;
      RECT  30590.0 87900.0 31295.0 89245.0 ;
      RECT  30590.0 90590.0 31295.0 89245.0 ;
      RECT  30590.0 90590.0 31295.0 91935.0 ;
      RECT  30590.0 93280.0 31295.0 91935.0 ;
      RECT  30590.0 93280.0 31295.0 94625.0 ;
      RECT  30590.0 95970.0 31295.0 94625.0 ;
      RECT  30590.0 95970.0 31295.0 97315.0 ;
      RECT  30590.0 98660.0 31295.0 97315.0 ;
      RECT  30590.0 98660.0 31295.0 100005.0 ;
      RECT  30590.0 101350.0 31295.0 100005.0 ;
      RECT  30590.0 101350.0 31295.0 102695.0 ;
      RECT  30590.0 104040.0 31295.0 102695.0 ;
      RECT  30590.0 104040.0 31295.0 105385.0 ;
      RECT  30590.0 106730.0 31295.0 105385.0 ;
      RECT  30590.0 106730.0 31295.0 108075.0 ;
      RECT  30590.0 109420.0 31295.0 108075.0 ;
      RECT  30590.0 109420.0 31295.0 110765.0 ;
      RECT  30590.0 112110.0 31295.0 110765.0 ;
      RECT  30590.0 112110.0 31295.0 113455.0 ;
      RECT  30590.0 114800.0 31295.0 113455.0 ;
      RECT  30590.0 114800.0 31295.0 116145.0 ;
      RECT  30590.0 117490.0 31295.0 116145.0 ;
      RECT  30590.0 117490.0 31295.0 118835.0 ;
      RECT  30590.0 120180.0 31295.0 118835.0 ;
      RECT  30590.0 120180.0 31295.0 121525.0 ;
      RECT  30590.0 122870.0 31295.0 121525.0 ;
      RECT  30590.0 122870.0 31295.0 124215.0 ;
      RECT  30590.0 125560.0 31295.0 124215.0 ;
      RECT  30590.0 125560.0 31295.0 126905.0 ;
      RECT  30590.0 128250.0 31295.0 126905.0 ;
      RECT  30590.0 128250.0 31295.0 129595.0 ;
      RECT  30590.0 130940.0 31295.0 129595.0 ;
      RECT  30590.0 130940.0 31295.0 132285.0 ;
      RECT  30590.0 133630.0 31295.0 132285.0 ;
      RECT  30590.0 133630.0 31295.0 134975.0 ;
      RECT  30590.0 136320.0 31295.0 134975.0 ;
      RECT  30590.0 136320.0 31295.0 137665.0 ;
      RECT  30590.0 139010.0 31295.0 137665.0 ;
      RECT  30590.0 139010.0 31295.0 140355.0 ;
      RECT  30590.0 141700.0 31295.0 140355.0 ;
      RECT  30590.0 141700.0 31295.0 143045.0 ;
      RECT  30590.0 144390.0 31295.0 143045.0 ;
      RECT  30590.0 144390.0 31295.0 145735.0 ;
      RECT  30590.0 147080.0 31295.0 145735.0 ;
      RECT  30590.0 147080.0 31295.0 148425.0 ;
      RECT  30590.0 149770.0 31295.0 148425.0 ;
      RECT  30590.0 149770.0 31295.0 151115.0 ;
      RECT  30590.0 152460.0 31295.0 151115.0 ;
      RECT  30590.0 152460.0 31295.0 153805.0 ;
      RECT  30590.0 155150.0 31295.0 153805.0 ;
      RECT  30590.0 155150.0 31295.0 156495.0 ;
      RECT  30590.0 157840.0 31295.0 156495.0 ;
      RECT  30590.0 157840.0 31295.0 159185.0 ;
      RECT  30590.0 160530.0 31295.0 159185.0 ;
      RECT  30590.0 160530.0 31295.0 161875.0 ;
      RECT  30590.0 163220.0 31295.0 161875.0 ;
      RECT  30590.0 163220.0 31295.0 164565.0 ;
      RECT  30590.0 165910.0 31295.0 164565.0 ;
      RECT  30590.0 165910.0 31295.0 167255.0 ;
      RECT  30590.0 168600.0 31295.0 167255.0 ;
      RECT  30590.0 168600.0 31295.0 169945.0 ;
      RECT  30590.0 171290.0 31295.0 169945.0 ;
      RECT  30590.0 171290.0 31295.0 172635.0 ;
      RECT  30590.0 173980.0 31295.0 172635.0 ;
      RECT  30590.0 173980.0 31295.0 175325.0 ;
      RECT  30590.0 176670.0 31295.0 175325.0 ;
      RECT  30590.0 176670.0 31295.0 178015.0 ;
      RECT  30590.0 179360.0 31295.0 178015.0 ;
      RECT  30590.0 179360.0 31295.0 180705.0 ;
      RECT  30590.0 182050.0 31295.0 180705.0 ;
      RECT  30590.0 182050.0 31295.0 183395.0 ;
      RECT  30590.0 184740.0 31295.0 183395.0 ;
      RECT  30590.0 184740.0 31295.0 186085.0 ;
      RECT  30590.0 187430.0 31295.0 186085.0 ;
      RECT  30590.0 187430.0 31295.0 188775.0 ;
      RECT  30590.0 190120.0 31295.0 188775.0 ;
      RECT  30590.0 190120.0 31295.0 191465.0 ;
      RECT  30590.0 192810.0 31295.0 191465.0 ;
      RECT  30590.0 192810.0 31295.0 194155.0 ;
      RECT  30590.0 195500.0 31295.0 194155.0 ;
      RECT  30590.0 195500.0 31295.0 196845.0 ;
      RECT  30590.0 198190.0 31295.0 196845.0 ;
      RECT  30590.0 198190.0 31295.0 199535.0 ;
      RECT  30590.0 200880.0 31295.0 199535.0 ;
      RECT  30590.0 200880.0 31295.0 202225.0 ;
      RECT  30590.0 203570.0 31295.0 202225.0 ;
      RECT  30590.0 203570.0 31295.0 204915.0 ;
      RECT  30590.0 206260.0 31295.0 204915.0 ;
      RECT  31295.0 34100.0 32000.0 35445.0 ;
      RECT  31295.0 36790.0 32000.0 35445.0 ;
      RECT  31295.0 36790.0 32000.0 38135.0 ;
      RECT  31295.0 39480.0 32000.0 38135.0 ;
      RECT  31295.0 39480.0 32000.0 40825.0 ;
      RECT  31295.0 42170.0 32000.0 40825.0 ;
      RECT  31295.0 42170.0 32000.0 43515.0 ;
      RECT  31295.0 44860.0 32000.0 43515.0 ;
      RECT  31295.0 44860.0 32000.0 46205.0 ;
      RECT  31295.0 47550.0 32000.0 46205.0 ;
      RECT  31295.0 47550.0 32000.0 48895.0 ;
      RECT  31295.0 50240.0 32000.0 48895.0 ;
      RECT  31295.0 50240.0 32000.0 51585.0 ;
      RECT  31295.0 52930.0 32000.0 51585.0 ;
      RECT  31295.0 52930.0 32000.0 54275.0 ;
      RECT  31295.0 55620.0 32000.0 54275.0 ;
      RECT  31295.0 55620.0 32000.0 56965.0 ;
      RECT  31295.0 58310.0 32000.0 56965.0 ;
      RECT  31295.0 58310.0 32000.0 59655.0 ;
      RECT  31295.0 61000.0 32000.0 59655.0 ;
      RECT  31295.0 61000.0 32000.0 62345.0 ;
      RECT  31295.0 63690.0 32000.0 62345.0 ;
      RECT  31295.0 63690.0 32000.0 65035.0 ;
      RECT  31295.0 66380.0 32000.0 65035.0 ;
      RECT  31295.0 66380.0 32000.0 67725.0 ;
      RECT  31295.0 69070.0 32000.0 67725.0 ;
      RECT  31295.0 69070.0 32000.0 70415.0 ;
      RECT  31295.0 71760.0 32000.0 70415.0 ;
      RECT  31295.0 71760.0 32000.0 73105.0 ;
      RECT  31295.0 74450.0 32000.0 73105.0 ;
      RECT  31295.0 74450.0 32000.0 75795.0 ;
      RECT  31295.0 77140.0 32000.0 75795.0 ;
      RECT  31295.0 77140.0 32000.0 78485.0 ;
      RECT  31295.0 79830.0 32000.0 78485.0 ;
      RECT  31295.0 79830.0 32000.0 81175.0 ;
      RECT  31295.0 82520.0 32000.0 81175.0 ;
      RECT  31295.0 82520.0 32000.0 83865.0 ;
      RECT  31295.0 85210.0 32000.0 83865.0 ;
      RECT  31295.0 85210.0 32000.0 86555.0 ;
      RECT  31295.0 87900.0 32000.0 86555.0 ;
      RECT  31295.0 87900.0 32000.0 89245.0 ;
      RECT  31295.0 90590.0 32000.0 89245.0 ;
      RECT  31295.0 90590.0 32000.0 91935.0 ;
      RECT  31295.0 93280.0 32000.0 91935.0 ;
      RECT  31295.0 93280.0 32000.0 94625.0 ;
      RECT  31295.0 95970.0 32000.0 94625.0 ;
      RECT  31295.0 95970.0 32000.0 97315.0 ;
      RECT  31295.0 98660.0 32000.0 97315.0 ;
      RECT  31295.0 98660.0 32000.0 100005.0 ;
      RECT  31295.0 101350.0 32000.0 100005.0 ;
      RECT  31295.0 101350.0 32000.0 102695.0 ;
      RECT  31295.0 104040.0 32000.0 102695.0 ;
      RECT  31295.0 104040.0 32000.0 105385.0 ;
      RECT  31295.0 106730.0 32000.0 105385.0 ;
      RECT  31295.0 106730.0 32000.0 108075.0 ;
      RECT  31295.0 109420.0 32000.0 108075.0 ;
      RECT  31295.0 109420.0 32000.0 110765.0 ;
      RECT  31295.0 112110.0 32000.0 110765.0 ;
      RECT  31295.0 112110.0 32000.0 113455.0 ;
      RECT  31295.0 114800.0 32000.0 113455.0 ;
      RECT  31295.0 114800.0 32000.0 116145.0 ;
      RECT  31295.0 117490.0 32000.0 116145.0 ;
      RECT  31295.0 117490.0 32000.0 118835.0 ;
      RECT  31295.0 120180.0 32000.0 118835.0 ;
      RECT  31295.0 120180.0 32000.0 121525.0 ;
      RECT  31295.0 122870.0 32000.0 121525.0 ;
      RECT  31295.0 122870.0 32000.0 124215.0 ;
      RECT  31295.0 125560.0 32000.0 124215.0 ;
      RECT  31295.0 125560.0 32000.0 126905.0 ;
      RECT  31295.0 128250.0 32000.0 126905.0 ;
      RECT  31295.0 128250.0 32000.0 129595.0 ;
      RECT  31295.0 130940.0 32000.0 129595.0 ;
      RECT  31295.0 130940.0 32000.0 132285.0 ;
      RECT  31295.0 133630.0 32000.0 132285.0 ;
      RECT  31295.0 133630.0 32000.0 134975.0 ;
      RECT  31295.0 136320.0 32000.0 134975.0 ;
      RECT  31295.0 136320.0 32000.0 137665.0 ;
      RECT  31295.0 139010.0 32000.0 137665.0 ;
      RECT  31295.0 139010.0 32000.0 140355.0 ;
      RECT  31295.0 141700.0 32000.0 140355.0 ;
      RECT  31295.0 141700.0 32000.0 143045.0 ;
      RECT  31295.0 144390.0 32000.0 143045.0 ;
      RECT  31295.0 144390.0 32000.0 145735.0 ;
      RECT  31295.0 147080.0 32000.0 145735.0 ;
      RECT  31295.0 147080.0 32000.0 148425.0 ;
      RECT  31295.0 149770.0 32000.0 148425.0 ;
      RECT  31295.0 149770.0 32000.0 151115.0 ;
      RECT  31295.0 152460.0 32000.0 151115.0 ;
      RECT  31295.0 152460.0 32000.0 153805.0 ;
      RECT  31295.0 155150.0 32000.0 153805.0 ;
      RECT  31295.0 155150.0 32000.0 156495.0 ;
      RECT  31295.0 157840.0 32000.0 156495.0 ;
      RECT  31295.0 157840.0 32000.0 159185.0 ;
      RECT  31295.0 160530.0 32000.0 159185.0 ;
      RECT  31295.0 160530.0 32000.0 161875.0 ;
      RECT  31295.0 163220.0 32000.0 161875.0 ;
      RECT  31295.0 163220.0 32000.0 164565.0 ;
      RECT  31295.0 165910.0 32000.0 164565.0 ;
      RECT  31295.0 165910.0 32000.0 167255.0 ;
      RECT  31295.0 168600.0 32000.0 167255.0 ;
      RECT  31295.0 168600.0 32000.0 169945.0 ;
      RECT  31295.0 171290.0 32000.0 169945.0 ;
      RECT  31295.0 171290.0 32000.0 172635.0 ;
      RECT  31295.0 173980.0 32000.0 172635.0 ;
      RECT  31295.0 173980.0 32000.0 175325.0 ;
      RECT  31295.0 176670.0 32000.0 175325.0 ;
      RECT  31295.0 176670.0 32000.0 178015.0 ;
      RECT  31295.0 179360.0 32000.0 178015.0 ;
      RECT  31295.0 179360.0 32000.0 180705.0 ;
      RECT  31295.0 182050.0 32000.0 180705.0 ;
      RECT  31295.0 182050.0 32000.0 183395.0 ;
      RECT  31295.0 184740.0 32000.0 183395.0 ;
      RECT  31295.0 184740.0 32000.0 186085.0 ;
      RECT  31295.0 187430.0 32000.0 186085.0 ;
      RECT  31295.0 187430.0 32000.0 188775.0 ;
      RECT  31295.0 190120.0 32000.0 188775.0 ;
      RECT  31295.0 190120.0 32000.0 191465.0 ;
      RECT  31295.0 192810.0 32000.0 191465.0 ;
      RECT  31295.0 192810.0 32000.0 194155.0 ;
      RECT  31295.0 195500.0 32000.0 194155.0 ;
      RECT  31295.0 195500.0 32000.0 196845.0 ;
      RECT  31295.0 198190.0 32000.0 196845.0 ;
      RECT  31295.0 198190.0 32000.0 199535.0 ;
      RECT  31295.0 200880.0 32000.0 199535.0 ;
      RECT  31295.0 200880.0 32000.0 202225.0 ;
      RECT  31295.0 203570.0 32000.0 202225.0 ;
      RECT  31295.0 203570.0 32000.0 204915.0 ;
      RECT  31295.0 206260.0 32000.0 204915.0 ;
      RECT  32000.0 34100.0 32705.0 35445.0 ;
      RECT  32000.0 36790.0 32705.0 35445.0 ;
      RECT  32000.0 36790.0 32705.0 38135.0 ;
      RECT  32000.0 39480.0 32705.0 38135.0 ;
      RECT  32000.0 39480.0 32705.0 40825.0 ;
      RECT  32000.0 42170.0 32705.0 40825.0 ;
      RECT  32000.0 42170.0 32705.0 43515.0 ;
      RECT  32000.0 44860.0 32705.0 43515.0 ;
      RECT  32000.0 44860.0 32705.0 46205.0 ;
      RECT  32000.0 47550.0 32705.0 46205.0 ;
      RECT  32000.0 47550.0 32705.0 48895.0 ;
      RECT  32000.0 50240.0 32705.0 48895.0 ;
      RECT  32000.0 50240.0 32705.0 51585.0 ;
      RECT  32000.0 52930.0 32705.0 51585.0 ;
      RECT  32000.0 52930.0 32705.0 54275.0 ;
      RECT  32000.0 55620.0 32705.0 54275.0 ;
      RECT  32000.0 55620.0 32705.0 56965.0 ;
      RECT  32000.0 58310.0 32705.0 56965.0 ;
      RECT  32000.0 58310.0 32705.0 59655.0 ;
      RECT  32000.0 61000.0 32705.0 59655.0 ;
      RECT  32000.0 61000.0 32705.0 62345.0 ;
      RECT  32000.0 63690.0 32705.0 62345.0 ;
      RECT  32000.0 63690.0 32705.0 65035.0 ;
      RECT  32000.0 66380.0 32705.0 65035.0 ;
      RECT  32000.0 66380.0 32705.0 67725.0 ;
      RECT  32000.0 69070.0 32705.0 67725.0 ;
      RECT  32000.0 69070.0 32705.0 70415.0 ;
      RECT  32000.0 71760.0 32705.0 70415.0 ;
      RECT  32000.0 71760.0 32705.0 73105.0 ;
      RECT  32000.0 74450.0 32705.0 73105.0 ;
      RECT  32000.0 74450.0 32705.0 75795.0 ;
      RECT  32000.0 77140.0 32705.0 75795.0 ;
      RECT  32000.0 77140.0 32705.0 78485.0 ;
      RECT  32000.0 79830.0 32705.0 78485.0 ;
      RECT  32000.0 79830.0 32705.0 81175.0 ;
      RECT  32000.0 82520.0 32705.0 81175.0 ;
      RECT  32000.0 82520.0 32705.0 83865.0 ;
      RECT  32000.0 85210.0 32705.0 83865.0 ;
      RECT  32000.0 85210.0 32705.0 86555.0 ;
      RECT  32000.0 87900.0 32705.0 86555.0 ;
      RECT  32000.0 87900.0 32705.0 89245.0 ;
      RECT  32000.0 90590.0 32705.0 89245.0 ;
      RECT  32000.0 90590.0 32705.0 91935.0 ;
      RECT  32000.0 93280.0 32705.0 91935.0 ;
      RECT  32000.0 93280.0 32705.0 94625.0 ;
      RECT  32000.0 95970.0 32705.0 94625.0 ;
      RECT  32000.0 95970.0 32705.0 97315.0 ;
      RECT  32000.0 98660.0 32705.0 97315.0 ;
      RECT  32000.0 98660.0 32705.0 100005.0 ;
      RECT  32000.0 101350.0 32705.0 100005.0 ;
      RECT  32000.0 101350.0 32705.0 102695.0 ;
      RECT  32000.0 104040.0 32705.0 102695.0 ;
      RECT  32000.0 104040.0 32705.0 105385.0 ;
      RECT  32000.0 106730.0 32705.0 105385.0 ;
      RECT  32000.0 106730.0 32705.0 108075.0 ;
      RECT  32000.0 109420.0 32705.0 108075.0 ;
      RECT  32000.0 109420.0 32705.0 110765.0 ;
      RECT  32000.0 112110.0 32705.0 110765.0 ;
      RECT  32000.0 112110.0 32705.0 113455.0 ;
      RECT  32000.0 114800.0 32705.0 113455.0 ;
      RECT  32000.0 114800.0 32705.0 116145.0 ;
      RECT  32000.0 117490.0 32705.0 116145.0 ;
      RECT  32000.0 117490.0 32705.0 118835.0 ;
      RECT  32000.0 120180.0 32705.0 118835.0 ;
      RECT  32000.0 120180.0 32705.0 121525.0 ;
      RECT  32000.0 122870.0 32705.0 121525.0 ;
      RECT  32000.0 122870.0 32705.0 124215.0 ;
      RECT  32000.0 125560.0 32705.0 124215.0 ;
      RECT  32000.0 125560.0 32705.0 126905.0 ;
      RECT  32000.0 128250.0 32705.0 126905.0 ;
      RECT  32000.0 128250.0 32705.0 129595.0 ;
      RECT  32000.0 130940.0 32705.0 129595.0 ;
      RECT  32000.0 130940.0 32705.0 132285.0 ;
      RECT  32000.0 133630.0 32705.0 132285.0 ;
      RECT  32000.0 133630.0 32705.0 134975.0 ;
      RECT  32000.0 136320.0 32705.0 134975.0 ;
      RECT  32000.0 136320.0 32705.0 137665.0 ;
      RECT  32000.0 139010.0 32705.0 137665.0 ;
      RECT  32000.0 139010.0 32705.0 140355.0 ;
      RECT  32000.0 141700.0 32705.0 140355.0 ;
      RECT  32000.0 141700.0 32705.0 143045.0 ;
      RECT  32000.0 144390.0 32705.0 143045.0 ;
      RECT  32000.0 144390.0 32705.0 145735.0 ;
      RECT  32000.0 147080.0 32705.0 145735.0 ;
      RECT  32000.0 147080.0 32705.0 148425.0 ;
      RECT  32000.0 149770.0 32705.0 148425.0 ;
      RECT  32000.0 149770.0 32705.0 151115.0 ;
      RECT  32000.0 152460.0 32705.0 151115.0 ;
      RECT  32000.0 152460.0 32705.0 153805.0 ;
      RECT  32000.0 155150.0 32705.0 153805.0 ;
      RECT  32000.0 155150.0 32705.0 156495.0 ;
      RECT  32000.0 157840.0 32705.0 156495.0 ;
      RECT  32000.0 157840.0 32705.0 159185.0 ;
      RECT  32000.0 160530.0 32705.0 159185.0 ;
      RECT  32000.0 160530.0 32705.0 161875.0 ;
      RECT  32000.0 163220.0 32705.0 161875.0 ;
      RECT  32000.0 163220.0 32705.0 164565.0 ;
      RECT  32000.0 165910.0 32705.0 164565.0 ;
      RECT  32000.0 165910.0 32705.0 167255.0 ;
      RECT  32000.0 168600.0 32705.0 167255.0 ;
      RECT  32000.0 168600.0 32705.0 169945.0 ;
      RECT  32000.0 171290.0 32705.0 169945.0 ;
      RECT  32000.0 171290.0 32705.0 172635.0 ;
      RECT  32000.0 173980.0 32705.0 172635.0 ;
      RECT  32000.0 173980.0 32705.0 175325.0 ;
      RECT  32000.0 176670.0 32705.0 175325.0 ;
      RECT  32000.0 176670.0 32705.0 178015.0 ;
      RECT  32000.0 179360.0 32705.0 178015.0 ;
      RECT  32000.0 179360.0 32705.0 180705.0 ;
      RECT  32000.0 182050.0 32705.0 180705.0 ;
      RECT  32000.0 182050.0 32705.0 183395.0 ;
      RECT  32000.0 184740.0 32705.0 183395.0 ;
      RECT  32000.0 184740.0 32705.0 186085.0 ;
      RECT  32000.0 187430.0 32705.0 186085.0 ;
      RECT  32000.0 187430.0 32705.0 188775.0 ;
      RECT  32000.0 190120.0 32705.0 188775.0 ;
      RECT  32000.0 190120.0 32705.0 191465.0 ;
      RECT  32000.0 192810.0 32705.0 191465.0 ;
      RECT  32000.0 192810.0 32705.0 194155.0 ;
      RECT  32000.0 195500.0 32705.0 194155.0 ;
      RECT  32000.0 195500.0 32705.0 196845.0 ;
      RECT  32000.0 198190.0 32705.0 196845.0 ;
      RECT  32000.0 198190.0 32705.0 199535.0 ;
      RECT  32000.0 200880.0 32705.0 199535.0 ;
      RECT  32000.0 200880.0 32705.0 202225.0 ;
      RECT  32000.0 203570.0 32705.0 202225.0 ;
      RECT  32000.0 203570.0 32705.0 204915.0 ;
      RECT  32000.0 206260.0 32705.0 204915.0 ;
      RECT  32705.0 34100.0 33410.0 35445.0 ;
      RECT  32705.0 36790.0 33410.0 35445.0 ;
      RECT  32705.0 36790.0 33410.0 38135.0 ;
      RECT  32705.0 39480.0 33410.0 38135.0 ;
      RECT  32705.0 39480.0 33410.0 40825.0 ;
      RECT  32705.0 42170.0 33410.0 40825.0 ;
      RECT  32705.0 42170.0 33410.0 43515.0 ;
      RECT  32705.0 44860.0 33410.0 43515.0 ;
      RECT  32705.0 44860.0 33410.0 46205.0 ;
      RECT  32705.0 47550.0 33410.0 46205.0 ;
      RECT  32705.0 47550.0 33410.0 48895.0 ;
      RECT  32705.0 50240.0 33410.0 48895.0 ;
      RECT  32705.0 50240.0 33410.0 51585.0 ;
      RECT  32705.0 52930.0 33410.0 51585.0 ;
      RECT  32705.0 52930.0 33410.0 54275.0 ;
      RECT  32705.0 55620.0 33410.0 54275.0 ;
      RECT  32705.0 55620.0 33410.0 56965.0 ;
      RECT  32705.0 58310.0 33410.0 56965.0 ;
      RECT  32705.0 58310.0 33410.0 59655.0 ;
      RECT  32705.0 61000.0 33410.0 59655.0 ;
      RECT  32705.0 61000.0 33410.0 62345.0 ;
      RECT  32705.0 63690.0 33410.0 62345.0 ;
      RECT  32705.0 63690.0 33410.0 65035.0 ;
      RECT  32705.0 66380.0 33410.0 65035.0 ;
      RECT  32705.0 66380.0 33410.0 67725.0 ;
      RECT  32705.0 69070.0 33410.0 67725.0 ;
      RECT  32705.0 69070.0 33410.0 70415.0 ;
      RECT  32705.0 71760.0 33410.0 70415.0 ;
      RECT  32705.0 71760.0 33410.0 73105.0 ;
      RECT  32705.0 74450.0 33410.0 73105.0 ;
      RECT  32705.0 74450.0 33410.0 75795.0 ;
      RECT  32705.0 77140.0 33410.0 75795.0 ;
      RECT  32705.0 77140.0 33410.0 78485.0 ;
      RECT  32705.0 79830.0 33410.0 78485.0 ;
      RECT  32705.0 79830.0 33410.0 81175.0 ;
      RECT  32705.0 82520.0 33410.0 81175.0 ;
      RECT  32705.0 82520.0 33410.0 83865.0 ;
      RECT  32705.0 85210.0 33410.0 83865.0 ;
      RECT  32705.0 85210.0 33410.0 86555.0 ;
      RECT  32705.0 87900.0 33410.0 86555.0 ;
      RECT  32705.0 87900.0 33410.0 89245.0 ;
      RECT  32705.0 90590.0 33410.0 89245.0 ;
      RECT  32705.0 90590.0 33410.0 91935.0 ;
      RECT  32705.0 93280.0 33410.0 91935.0 ;
      RECT  32705.0 93280.0 33410.0 94625.0 ;
      RECT  32705.0 95970.0 33410.0 94625.0 ;
      RECT  32705.0 95970.0 33410.0 97315.0 ;
      RECT  32705.0 98660.0 33410.0 97315.0 ;
      RECT  32705.0 98660.0 33410.0 100005.0 ;
      RECT  32705.0 101350.0 33410.0 100005.0 ;
      RECT  32705.0 101350.0 33410.0 102695.0 ;
      RECT  32705.0 104040.0 33410.0 102695.0 ;
      RECT  32705.0 104040.0 33410.0 105385.0 ;
      RECT  32705.0 106730.0 33410.0 105385.0 ;
      RECT  32705.0 106730.0 33410.0 108075.0 ;
      RECT  32705.0 109420.0 33410.0 108075.0 ;
      RECT  32705.0 109420.0 33410.0 110765.0 ;
      RECT  32705.0 112110.0 33410.0 110765.0 ;
      RECT  32705.0 112110.0 33410.0 113455.0 ;
      RECT  32705.0 114800.0 33410.0 113455.0 ;
      RECT  32705.0 114800.0 33410.0 116145.0 ;
      RECT  32705.0 117490.0 33410.0 116145.0 ;
      RECT  32705.0 117490.0 33410.0 118835.0 ;
      RECT  32705.0 120180.0 33410.0 118835.0 ;
      RECT  32705.0 120180.0 33410.0 121525.0 ;
      RECT  32705.0 122870.0 33410.0 121525.0 ;
      RECT  32705.0 122870.0 33410.0 124215.0 ;
      RECT  32705.0 125560.0 33410.0 124215.0 ;
      RECT  32705.0 125560.0 33410.0 126905.0 ;
      RECT  32705.0 128250.0 33410.0 126905.0 ;
      RECT  32705.0 128250.0 33410.0 129595.0 ;
      RECT  32705.0 130940.0 33410.0 129595.0 ;
      RECT  32705.0 130940.0 33410.0 132285.0 ;
      RECT  32705.0 133630.0 33410.0 132285.0 ;
      RECT  32705.0 133630.0 33410.0 134975.0 ;
      RECT  32705.0 136320.0 33410.0 134975.0 ;
      RECT  32705.0 136320.0 33410.0 137665.0 ;
      RECT  32705.0 139010.0 33410.0 137665.0 ;
      RECT  32705.0 139010.0 33410.0 140355.0 ;
      RECT  32705.0 141700.0 33410.0 140355.0 ;
      RECT  32705.0 141700.0 33410.0 143045.0 ;
      RECT  32705.0 144390.0 33410.0 143045.0 ;
      RECT  32705.0 144390.0 33410.0 145735.0 ;
      RECT  32705.0 147080.0 33410.0 145735.0 ;
      RECT  32705.0 147080.0 33410.0 148425.0 ;
      RECT  32705.0 149770.0 33410.0 148425.0 ;
      RECT  32705.0 149770.0 33410.0 151115.0 ;
      RECT  32705.0 152460.0 33410.0 151115.0 ;
      RECT  32705.0 152460.0 33410.0 153805.0 ;
      RECT  32705.0 155150.0 33410.0 153805.0 ;
      RECT  32705.0 155150.0 33410.0 156495.0 ;
      RECT  32705.0 157840.0 33410.0 156495.0 ;
      RECT  32705.0 157840.0 33410.0 159185.0 ;
      RECT  32705.0 160530.0 33410.0 159185.0 ;
      RECT  32705.0 160530.0 33410.0 161875.0 ;
      RECT  32705.0 163220.0 33410.0 161875.0 ;
      RECT  32705.0 163220.0 33410.0 164565.0 ;
      RECT  32705.0 165910.0 33410.0 164565.0 ;
      RECT  32705.0 165910.0 33410.0 167255.0 ;
      RECT  32705.0 168600.0 33410.0 167255.0 ;
      RECT  32705.0 168600.0 33410.0 169945.0 ;
      RECT  32705.0 171290.0 33410.0 169945.0 ;
      RECT  32705.0 171290.0 33410.0 172635.0 ;
      RECT  32705.0 173980.0 33410.0 172635.0 ;
      RECT  32705.0 173980.0 33410.0 175325.0 ;
      RECT  32705.0 176670.0 33410.0 175325.0 ;
      RECT  32705.0 176670.0 33410.0 178015.0 ;
      RECT  32705.0 179360.0 33410.0 178015.0 ;
      RECT  32705.0 179360.0 33410.0 180705.0 ;
      RECT  32705.0 182050.0 33410.0 180705.0 ;
      RECT  32705.0 182050.0 33410.0 183395.0 ;
      RECT  32705.0 184740.0 33410.0 183395.0 ;
      RECT  32705.0 184740.0 33410.0 186085.0 ;
      RECT  32705.0 187430.0 33410.0 186085.0 ;
      RECT  32705.0 187430.0 33410.0 188775.0 ;
      RECT  32705.0 190120.0 33410.0 188775.0 ;
      RECT  32705.0 190120.0 33410.0 191465.0 ;
      RECT  32705.0 192810.0 33410.0 191465.0 ;
      RECT  32705.0 192810.0 33410.0 194155.0 ;
      RECT  32705.0 195500.0 33410.0 194155.0 ;
      RECT  32705.0 195500.0 33410.0 196845.0 ;
      RECT  32705.0 198190.0 33410.0 196845.0 ;
      RECT  32705.0 198190.0 33410.0 199535.0 ;
      RECT  32705.0 200880.0 33410.0 199535.0 ;
      RECT  32705.0 200880.0 33410.0 202225.0 ;
      RECT  32705.0 203570.0 33410.0 202225.0 ;
      RECT  32705.0 203570.0 33410.0 204915.0 ;
      RECT  32705.0 206260.0 33410.0 204915.0 ;
      RECT  33410.0 34100.0 34115.0 35445.0 ;
      RECT  33410.0 36790.0 34115.0 35445.0 ;
      RECT  33410.0 36790.0 34115.0 38135.0 ;
      RECT  33410.0 39480.0 34115.0 38135.0 ;
      RECT  33410.0 39480.0 34115.0 40825.0 ;
      RECT  33410.0 42170.0 34115.0 40825.0 ;
      RECT  33410.0 42170.0 34115.0 43515.0 ;
      RECT  33410.0 44860.0 34115.0 43515.0 ;
      RECT  33410.0 44860.0 34115.0 46205.0 ;
      RECT  33410.0 47550.0 34115.0 46205.0 ;
      RECT  33410.0 47550.0 34115.0 48895.0 ;
      RECT  33410.0 50240.0 34115.0 48895.0 ;
      RECT  33410.0 50240.0 34115.0 51585.0 ;
      RECT  33410.0 52930.0 34115.0 51585.0 ;
      RECT  33410.0 52930.0 34115.0 54275.0 ;
      RECT  33410.0 55620.0 34115.0 54275.0 ;
      RECT  33410.0 55620.0 34115.0 56965.0 ;
      RECT  33410.0 58310.0 34115.0 56965.0 ;
      RECT  33410.0 58310.0 34115.0 59655.0 ;
      RECT  33410.0 61000.0 34115.0 59655.0 ;
      RECT  33410.0 61000.0 34115.0 62345.0 ;
      RECT  33410.0 63690.0 34115.0 62345.0 ;
      RECT  33410.0 63690.0 34115.0 65035.0 ;
      RECT  33410.0 66380.0 34115.0 65035.0 ;
      RECT  33410.0 66380.0 34115.0 67725.0 ;
      RECT  33410.0 69070.0 34115.0 67725.0 ;
      RECT  33410.0 69070.0 34115.0 70415.0 ;
      RECT  33410.0 71760.0 34115.0 70415.0 ;
      RECT  33410.0 71760.0 34115.0 73105.0 ;
      RECT  33410.0 74450.0 34115.0 73105.0 ;
      RECT  33410.0 74450.0 34115.0 75795.0 ;
      RECT  33410.0 77140.0 34115.0 75795.0 ;
      RECT  33410.0 77140.0 34115.0 78485.0 ;
      RECT  33410.0 79830.0 34115.0 78485.0 ;
      RECT  33410.0 79830.0 34115.0 81175.0 ;
      RECT  33410.0 82520.0 34115.0 81175.0 ;
      RECT  33410.0 82520.0 34115.0 83865.0 ;
      RECT  33410.0 85210.0 34115.0 83865.0 ;
      RECT  33410.0 85210.0 34115.0 86555.0 ;
      RECT  33410.0 87900.0 34115.0 86555.0 ;
      RECT  33410.0 87900.0 34115.0 89245.0 ;
      RECT  33410.0 90590.0 34115.0 89245.0 ;
      RECT  33410.0 90590.0 34115.0 91935.0 ;
      RECT  33410.0 93280.0 34115.0 91935.0 ;
      RECT  33410.0 93280.0 34115.0 94625.0 ;
      RECT  33410.0 95970.0 34115.0 94625.0 ;
      RECT  33410.0 95970.0 34115.0 97315.0 ;
      RECT  33410.0 98660.0 34115.0 97315.0 ;
      RECT  33410.0 98660.0 34115.0 100005.0 ;
      RECT  33410.0 101350.0 34115.0 100005.0 ;
      RECT  33410.0 101350.0 34115.0 102695.0 ;
      RECT  33410.0 104040.0 34115.0 102695.0 ;
      RECT  33410.0 104040.0 34115.0 105385.0 ;
      RECT  33410.0 106730.0 34115.0 105385.0 ;
      RECT  33410.0 106730.0 34115.0 108075.0 ;
      RECT  33410.0 109420.0 34115.0 108075.0 ;
      RECT  33410.0 109420.0 34115.0 110765.0 ;
      RECT  33410.0 112110.0 34115.0 110765.0 ;
      RECT  33410.0 112110.0 34115.0 113455.0 ;
      RECT  33410.0 114800.0 34115.0 113455.0 ;
      RECT  33410.0 114800.0 34115.0 116145.0 ;
      RECT  33410.0 117490.0 34115.0 116145.0 ;
      RECT  33410.0 117490.0 34115.0 118835.0 ;
      RECT  33410.0 120180.0 34115.0 118835.0 ;
      RECT  33410.0 120180.0 34115.0 121525.0 ;
      RECT  33410.0 122870.0 34115.0 121525.0 ;
      RECT  33410.0 122870.0 34115.0 124215.0 ;
      RECT  33410.0 125560.0 34115.0 124215.0 ;
      RECT  33410.0 125560.0 34115.0 126905.0 ;
      RECT  33410.0 128250.0 34115.0 126905.0 ;
      RECT  33410.0 128250.0 34115.0 129595.0 ;
      RECT  33410.0 130940.0 34115.0 129595.0 ;
      RECT  33410.0 130940.0 34115.0 132285.0 ;
      RECT  33410.0 133630.0 34115.0 132285.0 ;
      RECT  33410.0 133630.0 34115.0 134975.0 ;
      RECT  33410.0 136320.0 34115.0 134975.0 ;
      RECT  33410.0 136320.0 34115.0 137665.0 ;
      RECT  33410.0 139010.0 34115.0 137665.0 ;
      RECT  33410.0 139010.0 34115.0 140355.0 ;
      RECT  33410.0 141700.0 34115.0 140355.0 ;
      RECT  33410.0 141700.0 34115.0 143045.0 ;
      RECT  33410.0 144390.0 34115.0 143045.0 ;
      RECT  33410.0 144390.0 34115.0 145735.0 ;
      RECT  33410.0 147080.0 34115.0 145735.0 ;
      RECT  33410.0 147080.0 34115.0 148425.0 ;
      RECT  33410.0 149770.0 34115.0 148425.0 ;
      RECT  33410.0 149770.0 34115.0 151115.0 ;
      RECT  33410.0 152460.0 34115.0 151115.0 ;
      RECT  33410.0 152460.0 34115.0 153805.0 ;
      RECT  33410.0 155150.0 34115.0 153805.0 ;
      RECT  33410.0 155150.0 34115.0 156495.0 ;
      RECT  33410.0 157840.0 34115.0 156495.0 ;
      RECT  33410.0 157840.0 34115.0 159185.0 ;
      RECT  33410.0 160530.0 34115.0 159185.0 ;
      RECT  33410.0 160530.0 34115.0 161875.0 ;
      RECT  33410.0 163220.0 34115.0 161875.0 ;
      RECT  33410.0 163220.0 34115.0 164565.0 ;
      RECT  33410.0 165910.0 34115.0 164565.0 ;
      RECT  33410.0 165910.0 34115.0 167255.0 ;
      RECT  33410.0 168600.0 34115.0 167255.0 ;
      RECT  33410.0 168600.0 34115.0 169945.0 ;
      RECT  33410.0 171290.0 34115.0 169945.0 ;
      RECT  33410.0 171290.0 34115.0 172635.0 ;
      RECT  33410.0 173980.0 34115.0 172635.0 ;
      RECT  33410.0 173980.0 34115.0 175325.0 ;
      RECT  33410.0 176670.0 34115.0 175325.0 ;
      RECT  33410.0 176670.0 34115.0 178015.0 ;
      RECT  33410.0 179360.0 34115.0 178015.0 ;
      RECT  33410.0 179360.0 34115.0 180705.0 ;
      RECT  33410.0 182050.0 34115.0 180705.0 ;
      RECT  33410.0 182050.0 34115.0 183395.0 ;
      RECT  33410.0 184740.0 34115.0 183395.0 ;
      RECT  33410.0 184740.0 34115.0 186085.0 ;
      RECT  33410.0 187430.0 34115.0 186085.0 ;
      RECT  33410.0 187430.0 34115.0 188775.0 ;
      RECT  33410.0 190120.0 34115.0 188775.0 ;
      RECT  33410.0 190120.0 34115.0 191465.0 ;
      RECT  33410.0 192810.0 34115.0 191465.0 ;
      RECT  33410.0 192810.0 34115.0 194155.0 ;
      RECT  33410.0 195500.0 34115.0 194155.0 ;
      RECT  33410.0 195500.0 34115.0 196845.0 ;
      RECT  33410.0 198190.0 34115.0 196845.0 ;
      RECT  33410.0 198190.0 34115.0 199535.0 ;
      RECT  33410.0 200880.0 34115.0 199535.0 ;
      RECT  33410.0 200880.0 34115.0 202225.0 ;
      RECT  33410.0 203570.0 34115.0 202225.0 ;
      RECT  33410.0 203570.0 34115.0 204915.0 ;
      RECT  33410.0 206260.0 34115.0 204915.0 ;
      RECT  34115.0 34100.0 34820.0 35445.0 ;
      RECT  34115.0 36790.0 34820.0 35445.0 ;
      RECT  34115.0 36790.0 34820.0 38135.0 ;
      RECT  34115.0 39480.0 34820.0 38135.0 ;
      RECT  34115.0 39480.0 34820.0 40825.0 ;
      RECT  34115.0 42170.0 34820.0 40825.0 ;
      RECT  34115.0 42170.0 34820.0 43515.0 ;
      RECT  34115.0 44860.0 34820.0 43515.0 ;
      RECT  34115.0 44860.0 34820.0 46205.0 ;
      RECT  34115.0 47550.0 34820.0 46205.0 ;
      RECT  34115.0 47550.0 34820.0 48895.0 ;
      RECT  34115.0 50240.0 34820.0 48895.0 ;
      RECT  34115.0 50240.0 34820.0 51585.0 ;
      RECT  34115.0 52930.0 34820.0 51585.0 ;
      RECT  34115.0 52930.0 34820.0 54275.0 ;
      RECT  34115.0 55620.0 34820.0 54275.0 ;
      RECT  34115.0 55620.0 34820.0 56965.0 ;
      RECT  34115.0 58310.0 34820.0 56965.0 ;
      RECT  34115.0 58310.0 34820.0 59655.0 ;
      RECT  34115.0 61000.0 34820.0 59655.0 ;
      RECT  34115.0 61000.0 34820.0 62345.0 ;
      RECT  34115.0 63690.0 34820.0 62345.0 ;
      RECT  34115.0 63690.0 34820.0 65035.0 ;
      RECT  34115.0 66380.0 34820.0 65035.0 ;
      RECT  34115.0 66380.0 34820.0 67725.0 ;
      RECT  34115.0 69070.0 34820.0 67725.0 ;
      RECT  34115.0 69070.0 34820.0 70415.0 ;
      RECT  34115.0 71760.0 34820.0 70415.0 ;
      RECT  34115.0 71760.0 34820.0 73105.0 ;
      RECT  34115.0 74450.0 34820.0 73105.0 ;
      RECT  34115.0 74450.0 34820.0 75795.0 ;
      RECT  34115.0 77140.0 34820.0 75795.0 ;
      RECT  34115.0 77140.0 34820.0 78485.0 ;
      RECT  34115.0 79830.0 34820.0 78485.0 ;
      RECT  34115.0 79830.0 34820.0 81175.0 ;
      RECT  34115.0 82520.0 34820.0 81175.0 ;
      RECT  34115.0 82520.0 34820.0 83865.0 ;
      RECT  34115.0 85210.0 34820.0 83865.0 ;
      RECT  34115.0 85210.0 34820.0 86555.0 ;
      RECT  34115.0 87900.0 34820.0 86555.0 ;
      RECT  34115.0 87900.0 34820.0 89245.0 ;
      RECT  34115.0 90590.0 34820.0 89245.0 ;
      RECT  34115.0 90590.0 34820.0 91935.0 ;
      RECT  34115.0 93280.0 34820.0 91935.0 ;
      RECT  34115.0 93280.0 34820.0 94625.0 ;
      RECT  34115.0 95970.0 34820.0 94625.0 ;
      RECT  34115.0 95970.0 34820.0 97315.0 ;
      RECT  34115.0 98660.0 34820.0 97315.0 ;
      RECT  34115.0 98660.0 34820.0 100005.0 ;
      RECT  34115.0 101350.0 34820.0 100005.0 ;
      RECT  34115.0 101350.0 34820.0 102695.0 ;
      RECT  34115.0 104040.0 34820.0 102695.0 ;
      RECT  34115.0 104040.0 34820.0 105385.0 ;
      RECT  34115.0 106730.0 34820.0 105385.0 ;
      RECT  34115.0 106730.0 34820.0 108075.0 ;
      RECT  34115.0 109420.0 34820.0 108075.0 ;
      RECT  34115.0 109420.0 34820.0 110765.0 ;
      RECT  34115.0 112110.0 34820.0 110765.0 ;
      RECT  34115.0 112110.0 34820.0 113455.0 ;
      RECT  34115.0 114800.0 34820.0 113455.0 ;
      RECT  34115.0 114800.0 34820.0 116145.0 ;
      RECT  34115.0 117490.0 34820.0 116145.0 ;
      RECT  34115.0 117490.0 34820.0 118835.0 ;
      RECT  34115.0 120180.0 34820.0 118835.0 ;
      RECT  34115.0 120180.0 34820.0 121525.0 ;
      RECT  34115.0 122870.0 34820.0 121525.0 ;
      RECT  34115.0 122870.0 34820.0 124215.0 ;
      RECT  34115.0 125560.0 34820.0 124215.0 ;
      RECT  34115.0 125560.0 34820.0 126905.0 ;
      RECT  34115.0 128250.0 34820.0 126905.0 ;
      RECT  34115.0 128250.0 34820.0 129595.0 ;
      RECT  34115.0 130940.0 34820.0 129595.0 ;
      RECT  34115.0 130940.0 34820.0 132285.0 ;
      RECT  34115.0 133630.0 34820.0 132285.0 ;
      RECT  34115.0 133630.0 34820.0 134975.0 ;
      RECT  34115.0 136320.0 34820.0 134975.0 ;
      RECT  34115.0 136320.0 34820.0 137665.0 ;
      RECT  34115.0 139010.0 34820.0 137665.0 ;
      RECT  34115.0 139010.0 34820.0 140355.0 ;
      RECT  34115.0 141700.0 34820.0 140355.0 ;
      RECT  34115.0 141700.0 34820.0 143045.0 ;
      RECT  34115.0 144390.0 34820.0 143045.0 ;
      RECT  34115.0 144390.0 34820.0 145735.0 ;
      RECT  34115.0 147080.0 34820.0 145735.0 ;
      RECT  34115.0 147080.0 34820.0 148425.0 ;
      RECT  34115.0 149770.0 34820.0 148425.0 ;
      RECT  34115.0 149770.0 34820.0 151115.0 ;
      RECT  34115.0 152460.0 34820.0 151115.0 ;
      RECT  34115.0 152460.0 34820.0 153805.0 ;
      RECT  34115.0 155150.0 34820.0 153805.0 ;
      RECT  34115.0 155150.0 34820.0 156495.0 ;
      RECT  34115.0 157840.0 34820.0 156495.0 ;
      RECT  34115.0 157840.0 34820.0 159185.0 ;
      RECT  34115.0 160530.0 34820.0 159185.0 ;
      RECT  34115.0 160530.0 34820.0 161875.0 ;
      RECT  34115.0 163220.0 34820.0 161875.0 ;
      RECT  34115.0 163220.0 34820.0 164565.0 ;
      RECT  34115.0 165910.0 34820.0 164565.0 ;
      RECT  34115.0 165910.0 34820.0 167255.0 ;
      RECT  34115.0 168600.0 34820.0 167255.0 ;
      RECT  34115.0 168600.0 34820.0 169945.0 ;
      RECT  34115.0 171290.0 34820.0 169945.0 ;
      RECT  34115.0 171290.0 34820.0 172635.0 ;
      RECT  34115.0 173980.0 34820.0 172635.0 ;
      RECT  34115.0 173980.0 34820.0 175325.0 ;
      RECT  34115.0 176670.0 34820.0 175325.0 ;
      RECT  34115.0 176670.0 34820.0 178015.0 ;
      RECT  34115.0 179360.0 34820.0 178015.0 ;
      RECT  34115.0 179360.0 34820.0 180705.0 ;
      RECT  34115.0 182050.0 34820.0 180705.0 ;
      RECT  34115.0 182050.0 34820.0 183395.0 ;
      RECT  34115.0 184740.0 34820.0 183395.0 ;
      RECT  34115.0 184740.0 34820.0 186085.0 ;
      RECT  34115.0 187430.0 34820.0 186085.0 ;
      RECT  34115.0 187430.0 34820.0 188775.0 ;
      RECT  34115.0 190120.0 34820.0 188775.0 ;
      RECT  34115.0 190120.0 34820.0 191465.0 ;
      RECT  34115.0 192810.0 34820.0 191465.0 ;
      RECT  34115.0 192810.0 34820.0 194155.0 ;
      RECT  34115.0 195500.0 34820.0 194155.0 ;
      RECT  34115.0 195500.0 34820.0 196845.0 ;
      RECT  34115.0 198190.0 34820.0 196845.0 ;
      RECT  34115.0 198190.0 34820.0 199535.0 ;
      RECT  34115.0 200880.0 34820.0 199535.0 ;
      RECT  34115.0 200880.0 34820.0 202225.0 ;
      RECT  34115.0 203570.0 34820.0 202225.0 ;
      RECT  34115.0 203570.0 34820.0 204915.0 ;
      RECT  34115.0 206260.0 34820.0 204915.0 ;
      RECT  34820.0 34100.0 35525.0 35445.0 ;
      RECT  34820.0 36790.0 35525.0 35445.0 ;
      RECT  34820.0 36790.0 35525.0 38135.0 ;
      RECT  34820.0 39480.0 35525.0 38135.0 ;
      RECT  34820.0 39480.0 35525.0 40825.0 ;
      RECT  34820.0 42170.0 35525.0 40825.0 ;
      RECT  34820.0 42170.0 35525.0 43515.0 ;
      RECT  34820.0 44860.0 35525.0 43515.0 ;
      RECT  34820.0 44860.0 35525.0 46205.0 ;
      RECT  34820.0 47550.0 35525.0 46205.0 ;
      RECT  34820.0 47550.0 35525.0 48895.0 ;
      RECT  34820.0 50240.0 35525.0 48895.0 ;
      RECT  34820.0 50240.0 35525.0 51585.0 ;
      RECT  34820.0 52930.0 35525.0 51585.0 ;
      RECT  34820.0 52930.0 35525.0 54275.0 ;
      RECT  34820.0 55620.0 35525.0 54275.0 ;
      RECT  34820.0 55620.0 35525.0 56965.0 ;
      RECT  34820.0 58310.0 35525.0 56965.0 ;
      RECT  34820.0 58310.0 35525.0 59655.0 ;
      RECT  34820.0 61000.0 35525.0 59655.0 ;
      RECT  34820.0 61000.0 35525.0 62345.0 ;
      RECT  34820.0 63690.0 35525.0 62345.0 ;
      RECT  34820.0 63690.0 35525.0 65035.0 ;
      RECT  34820.0 66380.0 35525.0 65035.0 ;
      RECT  34820.0 66380.0 35525.0 67725.0 ;
      RECT  34820.0 69070.0 35525.0 67725.0 ;
      RECT  34820.0 69070.0 35525.0 70415.0 ;
      RECT  34820.0 71760.0 35525.0 70415.0 ;
      RECT  34820.0 71760.0 35525.0 73105.0 ;
      RECT  34820.0 74450.0 35525.0 73105.0 ;
      RECT  34820.0 74450.0 35525.0 75795.0 ;
      RECT  34820.0 77140.0 35525.0 75795.0 ;
      RECT  34820.0 77140.0 35525.0 78485.0 ;
      RECT  34820.0 79830.0 35525.0 78485.0 ;
      RECT  34820.0 79830.0 35525.0 81175.0 ;
      RECT  34820.0 82520.0 35525.0 81175.0 ;
      RECT  34820.0 82520.0 35525.0 83865.0 ;
      RECT  34820.0 85210.0 35525.0 83865.0 ;
      RECT  34820.0 85210.0 35525.0 86555.0 ;
      RECT  34820.0 87900.0 35525.0 86555.0 ;
      RECT  34820.0 87900.0 35525.0 89245.0 ;
      RECT  34820.0 90590.0 35525.0 89245.0 ;
      RECT  34820.0 90590.0 35525.0 91935.0 ;
      RECT  34820.0 93280.0 35525.0 91935.0 ;
      RECT  34820.0 93280.0 35525.0 94625.0 ;
      RECT  34820.0 95970.0 35525.0 94625.0 ;
      RECT  34820.0 95970.0 35525.0 97315.0 ;
      RECT  34820.0 98660.0 35525.0 97315.0 ;
      RECT  34820.0 98660.0 35525.0 100005.0 ;
      RECT  34820.0 101350.0 35525.0 100005.0 ;
      RECT  34820.0 101350.0 35525.0 102695.0 ;
      RECT  34820.0 104040.0 35525.0 102695.0 ;
      RECT  34820.0 104040.0 35525.0 105385.0 ;
      RECT  34820.0 106730.0 35525.0 105385.0 ;
      RECT  34820.0 106730.0 35525.0 108075.0 ;
      RECT  34820.0 109420.0 35525.0 108075.0 ;
      RECT  34820.0 109420.0 35525.0 110765.0 ;
      RECT  34820.0 112110.0 35525.0 110765.0 ;
      RECT  34820.0 112110.0 35525.0 113455.0 ;
      RECT  34820.0 114800.0 35525.0 113455.0 ;
      RECT  34820.0 114800.0 35525.0 116145.0 ;
      RECT  34820.0 117490.0 35525.0 116145.0 ;
      RECT  34820.0 117490.0 35525.0 118835.0 ;
      RECT  34820.0 120180.0 35525.0 118835.0 ;
      RECT  34820.0 120180.0 35525.0 121525.0 ;
      RECT  34820.0 122870.0 35525.0 121525.0 ;
      RECT  34820.0 122870.0 35525.0 124215.0 ;
      RECT  34820.0 125560.0 35525.0 124215.0 ;
      RECT  34820.0 125560.0 35525.0 126905.0 ;
      RECT  34820.0 128250.0 35525.0 126905.0 ;
      RECT  34820.0 128250.0 35525.0 129595.0 ;
      RECT  34820.0 130940.0 35525.0 129595.0 ;
      RECT  34820.0 130940.0 35525.0 132285.0 ;
      RECT  34820.0 133630.0 35525.0 132285.0 ;
      RECT  34820.0 133630.0 35525.0 134975.0 ;
      RECT  34820.0 136320.0 35525.0 134975.0 ;
      RECT  34820.0 136320.0 35525.0 137665.0 ;
      RECT  34820.0 139010.0 35525.0 137665.0 ;
      RECT  34820.0 139010.0 35525.0 140355.0 ;
      RECT  34820.0 141700.0 35525.0 140355.0 ;
      RECT  34820.0 141700.0 35525.0 143045.0 ;
      RECT  34820.0 144390.0 35525.0 143045.0 ;
      RECT  34820.0 144390.0 35525.0 145735.0 ;
      RECT  34820.0 147080.0 35525.0 145735.0 ;
      RECT  34820.0 147080.0 35525.0 148425.0 ;
      RECT  34820.0 149770.0 35525.0 148425.0 ;
      RECT  34820.0 149770.0 35525.0 151115.0 ;
      RECT  34820.0 152460.0 35525.0 151115.0 ;
      RECT  34820.0 152460.0 35525.0 153805.0 ;
      RECT  34820.0 155150.0 35525.0 153805.0 ;
      RECT  34820.0 155150.0 35525.0 156495.0 ;
      RECT  34820.0 157840.0 35525.0 156495.0 ;
      RECT  34820.0 157840.0 35525.0 159185.0 ;
      RECT  34820.0 160530.0 35525.0 159185.0 ;
      RECT  34820.0 160530.0 35525.0 161875.0 ;
      RECT  34820.0 163220.0 35525.0 161875.0 ;
      RECT  34820.0 163220.0 35525.0 164565.0 ;
      RECT  34820.0 165910.0 35525.0 164565.0 ;
      RECT  34820.0 165910.0 35525.0 167255.0 ;
      RECT  34820.0 168600.0 35525.0 167255.0 ;
      RECT  34820.0 168600.0 35525.0 169945.0 ;
      RECT  34820.0 171290.0 35525.0 169945.0 ;
      RECT  34820.0 171290.0 35525.0 172635.0 ;
      RECT  34820.0 173980.0 35525.0 172635.0 ;
      RECT  34820.0 173980.0 35525.0 175325.0 ;
      RECT  34820.0 176670.0 35525.0 175325.0 ;
      RECT  34820.0 176670.0 35525.0 178015.0 ;
      RECT  34820.0 179360.0 35525.0 178015.0 ;
      RECT  34820.0 179360.0 35525.0 180705.0 ;
      RECT  34820.0 182050.0 35525.0 180705.0 ;
      RECT  34820.0 182050.0 35525.0 183395.0 ;
      RECT  34820.0 184740.0 35525.0 183395.0 ;
      RECT  34820.0 184740.0 35525.0 186085.0 ;
      RECT  34820.0 187430.0 35525.0 186085.0 ;
      RECT  34820.0 187430.0 35525.0 188775.0 ;
      RECT  34820.0 190120.0 35525.0 188775.0 ;
      RECT  34820.0 190120.0 35525.0 191465.0 ;
      RECT  34820.0 192810.0 35525.0 191465.0 ;
      RECT  34820.0 192810.0 35525.0 194155.0 ;
      RECT  34820.0 195500.0 35525.0 194155.0 ;
      RECT  34820.0 195500.0 35525.0 196845.0 ;
      RECT  34820.0 198190.0 35525.0 196845.0 ;
      RECT  34820.0 198190.0 35525.0 199535.0 ;
      RECT  34820.0 200880.0 35525.0 199535.0 ;
      RECT  34820.0 200880.0 35525.0 202225.0 ;
      RECT  34820.0 203570.0 35525.0 202225.0 ;
      RECT  34820.0 203570.0 35525.0 204915.0 ;
      RECT  34820.0 206260.0 35525.0 204915.0 ;
      RECT  35525.0 34100.0 36230.0 35445.0 ;
      RECT  35525.0 36790.0 36230.0 35445.0 ;
      RECT  35525.0 36790.0 36230.0 38135.0 ;
      RECT  35525.0 39480.0 36230.0 38135.0 ;
      RECT  35525.0 39480.0 36230.0 40825.0 ;
      RECT  35525.0 42170.0 36230.0 40825.0 ;
      RECT  35525.0 42170.0 36230.0 43515.0 ;
      RECT  35525.0 44860.0 36230.0 43515.0 ;
      RECT  35525.0 44860.0 36230.0 46205.0 ;
      RECT  35525.0 47550.0 36230.0 46205.0 ;
      RECT  35525.0 47550.0 36230.0 48895.0 ;
      RECT  35525.0 50240.0 36230.0 48895.0 ;
      RECT  35525.0 50240.0 36230.0 51585.0 ;
      RECT  35525.0 52930.0 36230.0 51585.0 ;
      RECT  35525.0 52930.0 36230.0 54275.0 ;
      RECT  35525.0 55620.0 36230.0 54275.0 ;
      RECT  35525.0 55620.0 36230.0 56965.0 ;
      RECT  35525.0 58310.0 36230.0 56965.0 ;
      RECT  35525.0 58310.0 36230.0 59655.0 ;
      RECT  35525.0 61000.0 36230.0 59655.0 ;
      RECT  35525.0 61000.0 36230.0 62345.0 ;
      RECT  35525.0 63690.0 36230.0 62345.0 ;
      RECT  35525.0 63690.0 36230.0 65035.0 ;
      RECT  35525.0 66380.0 36230.0 65035.0 ;
      RECT  35525.0 66380.0 36230.0 67725.0 ;
      RECT  35525.0 69070.0 36230.0 67725.0 ;
      RECT  35525.0 69070.0 36230.0 70415.0 ;
      RECT  35525.0 71760.0 36230.0 70415.0 ;
      RECT  35525.0 71760.0 36230.0 73105.0 ;
      RECT  35525.0 74450.0 36230.0 73105.0 ;
      RECT  35525.0 74450.0 36230.0 75795.0 ;
      RECT  35525.0 77140.0 36230.0 75795.0 ;
      RECT  35525.0 77140.0 36230.0 78485.0 ;
      RECT  35525.0 79830.0 36230.0 78485.0 ;
      RECT  35525.0 79830.0 36230.0 81175.0 ;
      RECT  35525.0 82520.0 36230.0 81175.0 ;
      RECT  35525.0 82520.0 36230.0 83865.0 ;
      RECT  35525.0 85210.0 36230.0 83865.0 ;
      RECT  35525.0 85210.0 36230.0 86555.0 ;
      RECT  35525.0 87900.0 36230.0 86555.0 ;
      RECT  35525.0 87900.0 36230.0 89245.0 ;
      RECT  35525.0 90590.0 36230.0 89245.0 ;
      RECT  35525.0 90590.0 36230.0 91935.0 ;
      RECT  35525.0 93280.0 36230.0 91935.0 ;
      RECT  35525.0 93280.0 36230.0 94625.0 ;
      RECT  35525.0 95970.0 36230.0 94625.0 ;
      RECT  35525.0 95970.0 36230.0 97315.0 ;
      RECT  35525.0 98660.0 36230.0 97315.0 ;
      RECT  35525.0 98660.0 36230.0 100005.0 ;
      RECT  35525.0 101350.0 36230.0 100005.0 ;
      RECT  35525.0 101350.0 36230.0 102695.0 ;
      RECT  35525.0 104040.0 36230.0 102695.0 ;
      RECT  35525.0 104040.0 36230.0 105385.0 ;
      RECT  35525.0 106730.0 36230.0 105385.0 ;
      RECT  35525.0 106730.0 36230.0 108075.0 ;
      RECT  35525.0 109420.0 36230.0 108075.0 ;
      RECT  35525.0 109420.0 36230.0 110765.0 ;
      RECT  35525.0 112110.0 36230.0 110765.0 ;
      RECT  35525.0 112110.0 36230.0 113455.0 ;
      RECT  35525.0 114800.0 36230.0 113455.0 ;
      RECT  35525.0 114800.0 36230.0 116145.0 ;
      RECT  35525.0 117490.0 36230.0 116145.0 ;
      RECT  35525.0 117490.0 36230.0 118835.0 ;
      RECT  35525.0 120180.0 36230.0 118835.0 ;
      RECT  35525.0 120180.0 36230.0 121525.0 ;
      RECT  35525.0 122870.0 36230.0 121525.0 ;
      RECT  35525.0 122870.0 36230.0 124215.0 ;
      RECT  35525.0 125560.0 36230.0 124215.0 ;
      RECT  35525.0 125560.0 36230.0 126905.0 ;
      RECT  35525.0 128250.0 36230.0 126905.0 ;
      RECT  35525.0 128250.0 36230.0 129595.0 ;
      RECT  35525.0 130940.0 36230.0 129595.0 ;
      RECT  35525.0 130940.0 36230.0 132285.0 ;
      RECT  35525.0 133630.0 36230.0 132285.0 ;
      RECT  35525.0 133630.0 36230.0 134975.0 ;
      RECT  35525.0 136320.0 36230.0 134975.0 ;
      RECT  35525.0 136320.0 36230.0 137665.0 ;
      RECT  35525.0 139010.0 36230.0 137665.0 ;
      RECT  35525.0 139010.0 36230.0 140355.0 ;
      RECT  35525.0 141700.0 36230.0 140355.0 ;
      RECT  35525.0 141700.0 36230.0 143045.0 ;
      RECT  35525.0 144390.0 36230.0 143045.0 ;
      RECT  35525.0 144390.0 36230.0 145735.0 ;
      RECT  35525.0 147080.0 36230.0 145735.0 ;
      RECT  35525.0 147080.0 36230.0 148425.0 ;
      RECT  35525.0 149770.0 36230.0 148425.0 ;
      RECT  35525.0 149770.0 36230.0 151115.0 ;
      RECT  35525.0 152460.0 36230.0 151115.0 ;
      RECT  35525.0 152460.0 36230.0 153805.0 ;
      RECT  35525.0 155150.0 36230.0 153805.0 ;
      RECT  35525.0 155150.0 36230.0 156495.0 ;
      RECT  35525.0 157840.0 36230.0 156495.0 ;
      RECT  35525.0 157840.0 36230.0 159185.0 ;
      RECT  35525.0 160530.0 36230.0 159185.0 ;
      RECT  35525.0 160530.0 36230.0 161875.0 ;
      RECT  35525.0 163220.0 36230.0 161875.0 ;
      RECT  35525.0 163220.0 36230.0 164565.0 ;
      RECT  35525.0 165910.0 36230.0 164565.0 ;
      RECT  35525.0 165910.0 36230.0 167255.0 ;
      RECT  35525.0 168600.0 36230.0 167255.0 ;
      RECT  35525.0 168600.0 36230.0 169945.0 ;
      RECT  35525.0 171290.0 36230.0 169945.0 ;
      RECT  35525.0 171290.0 36230.0 172635.0 ;
      RECT  35525.0 173980.0 36230.0 172635.0 ;
      RECT  35525.0 173980.0 36230.0 175325.0 ;
      RECT  35525.0 176670.0 36230.0 175325.0 ;
      RECT  35525.0 176670.0 36230.0 178015.0 ;
      RECT  35525.0 179360.0 36230.0 178015.0 ;
      RECT  35525.0 179360.0 36230.0 180705.0 ;
      RECT  35525.0 182050.0 36230.0 180705.0 ;
      RECT  35525.0 182050.0 36230.0 183395.0 ;
      RECT  35525.0 184740.0 36230.0 183395.0 ;
      RECT  35525.0 184740.0 36230.0 186085.0 ;
      RECT  35525.0 187430.0 36230.0 186085.0 ;
      RECT  35525.0 187430.0 36230.0 188775.0 ;
      RECT  35525.0 190120.0 36230.0 188775.0 ;
      RECT  35525.0 190120.0 36230.0 191465.0 ;
      RECT  35525.0 192810.0 36230.0 191465.0 ;
      RECT  35525.0 192810.0 36230.0 194155.0 ;
      RECT  35525.0 195500.0 36230.0 194155.0 ;
      RECT  35525.0 195500.0 36230.0 196845.0 ;
      RECT  35525.0 198190.0 36230.0 196845.0 ;
      RECT  35525.0 198190.0 36230.0 199535.0 ;
      RECT  35525.0 200880.0 36230.0 199535.0 ;
      RECT  35525.0 200880.0 36230.0 202225.0 ;
      RECT  35525.0 203570.0 36230.0 202225.0 ;
      RECT  35525.0 203570.0 36230.0 204915.0 ;
      RECT  35525.0 206260.0 36230.0 204915.0 ;
      RECT  36230.0 34100.0 36935.0 35445.0 ;
      RECT  36230.0 36790.0 36935.0 35445.0 ;
      RECT  36230.0 36790.0 36935.0 38135.0 ;
      RECT  36230.0 39480.0 36935.0 38135.0 ;
      RECT  36230.0 39480.0 36935.0 40825.0 ;
      RECT  36230.0 42170.0 36935.0 40825.0 ;
      RECT  36230.0 42170.0 36935.0 43515.0 ;
      RECT  36230.0 44860.0 36935.0 43515.0 ;
      RECT  36230.0 44860.0 36935.0 46205.0 ;
      RECT  36230.0 47550.0 36935.0 46205.0 ;
      RECT  36230.0 47550.0 36935.0 48895.0 ;
      RECT  36230.0 50240.0 36935.0 48895.0 ;
      RECT  36230.0 50240.0 36935.0 51585.0 ;
      RECT  36230.0 52930.0 36935.0 51585.0 ;
      RECT  36230.0 52930.0 36935.0 54275.0 ;
      RECT  36230.0 55620.0 36935.0 54275.0 ;
      RECT  36230.0 55620.0 36935.0 56965.0 ;
      RECT  36230.0 58310.0 36935.0 56965.0 ;
      RECT  36230.0 58310.0 36935.0 59655.0 ;
      RECT  36230.0 61000.0 36935.0 59655.0 ;
      RECT  36230.0 61000.0 36935.0 62345.0 ;
      RECT  36230.0 63690.0 36935.0 62345.0 ;
      RECT  36230.0 63690.0 36935.0 65035.0 ;
      RECT  36230.0 66380.0 36935.0 65035.0 ;
      RECT  36230.0 66380.0 36935.0 67725.0 ;
      RECT  36230.0 69070.0 36935.0 67725.0 ;
      RECT  36230.0 69070.0 36935.0 70415.0 ;
      RECT  36230.0 71760.0 36935.0 70415.0 ;
      RECT  36230.0 71760.0 36935.0 73105.0 ;
      RECT  36230.0 74450.0 36935.0 73105.0 ;
      RECT  36230.0 74450.0 36935.0 75795.0 ;
      RECT  36230.0 77140.0 36935.0 75795.0 ;
      RECT  36230.0 77140.0 36935.0 78485.0 ;
      RECT  36230.0 79830.0 36935.0 78485.0 ;
      RECT  36230.0 79830.0 36935.0 81175.0 ;
      RECT  36230.0 82520.0 36935.0 81175.0 ;
      RECT  36230.0 82520.0 36935.0 83865.0 ;
      RECT  36230.0 85210.0 36935.0 83865.0 ;
      RECT  36230.0 85210.0 36935.0 86555.0 ;
      RECT  36230.0 87900.0 36935.0 86555.0 ;
      RECT  36230.0 87900.0 36935.0 89245.0 ;
      RECT  36230.0 90590.0 36935.0 89245.0 ;
      RECT  36230.0 90590.0 36935.0 91935.0 ;
      RECT  36230.0 93280.0 36935.0 91935.0 ;
      RECT  36230.0 93280.0 36935.0 94625.0 ;
      RECT  36230.0 95970.0 36935.0 94625.0 ;
      RECT  36230.0 95970.0 36935.0 97315.0 ;
      RECT  36230.0 98660.0 36935.0 97315.0 ;
      RECT  36230.0 98660.0 36935.0 100005.0 ;
      RECT  36230.0 101350.0 36935.0 100005.0 ;
      RECT  36230.0 101350.0 36935.0 102695.0 ;
      RECT  36230.0 104040.0 36935.0 102695.0 ;
      RECT  36230.0 104040.0 36935.0 105385.0 ;
      RECT  36230.0 106730.0 36935.0 105385.0 ;
      RECT  36230.0 106730.0 36935.0 108075.0 ;
      RECT  36230.0 109420.0 36935.0 108075.0 ;
      RECT  36230.0 109420.0 36935.0 110765.0 ;
      RECT  36230.0 112110.0 36935.0 110765.0 ;
      RECT  36230.0 112110.0 36935.0 113455.0 ;
      RECT  36230.0 114800.0 36935.0 113455.0 ;
      RECT  36230.0 114800.0 36935.0 116145.0 ;
      RECT  36230.0 117490.0 36935.0 116145.0 ;
      RECT  36230.0 117490.0 36935.0 118835.0 ;
      RECT  36230.0 120180.0 36935.0 118835.0 ;
      RECT  36230.0 120180.0 36935.0 121525.0 ;
      RECT  36230.0 122870.0 36935.0 121525.0 ;
      RECT  36230.0 122870.0 36935.0 124215.0 ;
      RECT  36230.0 125560.0 36935.0 124215.0 ;
      RECT  36230.0 125560.0 36935.0 126905.0 ;
      RECT  36230.0 128250.0 36935.0 126905.0 ;
      RECT  36230.0 128250.0 36935.0 129595.0 ;
      RECT  36230.0 130940.0 36935.0 129595.0 ;
      RECT  36230.0 130940.0 36935.0 132285.0 ;
      RECT  36230.0 133630.0 36935.0 132285.0 ;
      RECT  36230.0 133630.0 36935.0 134975.0 ;
      RECT  36230.0 136320.0 36935.0 134975.0 ;
      RECT  36230.0 136320.0 36935.0 137665.0 ;
      RECT  36230.0 139010.0 36935.0 137665.0 ;
      RECT  36230.0 139010.0 36935.0 140355.0 ;
      RECT  36230.0 141700.0 36935.0 140355.0 ;
      RECT  36230.0 141700.0 36935.0 143045.0 ;
      RECT  36230.0 144390.0 36935.0 143045.0 ;
      RECT  36230.0 144390.0 36935.0 145735.0 ;
      RECT  36230.0 147080.0 36935.0 145735.0 ;
      RECT  36230.0 147080.0 36935.0 148425.0 ;
      RECT  36230.0 149770.0 36935.0 148425.0 ;
      RECT  36230.0 149770.0 36935.0 151115.0 ;
      RECT  36230.0 152460.0 36935.0 151115.0 ;
      RECT  36230.0 152460.0 36935.0 153805.0 ;
      RECT  36230.0 155150.0 36935.0 153805.0 ;
      RECT  36230.0 155150.0 36935.0 156495.0 ;
      RECT  36230.0 157840.0 36935.0 156495.0 ;
      RECT  36230.0 157840.0 36935.0 159185.0 ;
      RECT  36230.0 160530.0 36935.0 159185.0 ;
      RECT  36230.0 160530.0 36935.0 161875.0 ;
      RECT  36230.0 163220.0 36935.0 161875.0 ;
      RECT  36230.0 163220.0 36935.0 164565.0 ;
      RECT  36230.0 165910.0 36935.0 164565.0 ;
      RECT  36230.0 165910.0 36935.0 167255.0 ;
      RECT  36230.0 168600.0 36935.0 167255.0 ;
      RECT  36230.0 168600.0 36935.0 169945.0 ;
      RECT  36230.0 171290.0 36935.0 169945.0 ;
      RECT  36230.0 171290.0 36935.0 172635.0 ;
      RECT  36230.0 173980.0 36935.0 172635.0 ;
      RECT  36230.0 173980.0 36935.0 175325.0 ;
      RECT  36230.0 176670.0 36935.0 175325.0 ;
      RECT  36230.0 176670.0 36935.0 178015.0 ;
      RECT  36230.0 179360.0 36935.0 178015.0 ;
      RECT  36230.0 179360.0 36935.0 180705.0 ;
      RECT  36230.0 182050.0 36935.0 180705.0 ;
      RECT  36230.0 182050.0 36935.0 183395.0 ;
      RECT  36230.0 184740.0 36935.0 183395.0 ;
      RECT  36230.0 184740.0 36935.0 186085.0 ;
      RECT  36230.0 187430.0 36935.0 186085.0 ;
      RECT  36230.0 187430.0 36935.0 188775.0 ;
      RECT  36230.0 190120.0 36935.0 188775.0 ;
      RECT  36230.0 190120.0 36935.0 191465.0 ;
      RECT  36230.0 192810.0 36935.0 191465.0 ;
      RECT  36230.0 192810.0 36935.0 194155.0 ;
      RECT  36230.0 195500.0 36935.0 194155.0 ;
      RECT  36230.0 195500.0 36935.0 196845.0 ;
      RECT  36230.0 198190.0 36935.0 196845.0 ;
      RECT  36230.0 198190.0 36935.0 199535.0 ;
      RECT  36230.0 200880.0 36935.0 199535.0 ;
      RECT  36230.0 200880.0 36935.0 202225.0 ;
      RECT  36230.0 203570.0 36935.0 202225.0 ;
      RECT  36230.0 203570.0 36935.0 204915.0 ;
      RECT  36230.0 206260.0 36935.0 204915.0 ;
      RECT  36935.0 34100.0 37640.0 35445.0 ;
      RECT  36935.0 36790.0 37640.0 35445.0 ;
      RECT  36935.0 36790.0 37640.0 38135.0 ;
      RECT  36935.0 39480.0 37640.0 38135.0 ;
      RECT  36935.0 39480.0 37640.0 40825.0 ;
      RECT  36935.0 42170.0 37640.0 40825.0 ;
      RECT  36935.0 42170.0 37640.0 43515.0 ;
      RECT  36935.0 44860.0 37640.0 43515.0 ;
      RECT  36935.0 44860.0 37640.0 46205.0 ;
      RECT  36935.0 47550.0 37640.0 46205.0 ;
      RECT  36935.0 47550.0 37640.0 48895.0 ;
      RECT  36935.0 50240.0 37640.0 48895.0 ;
      RECT  36935.0 50240.0 37640.0 51585.0 ;
      RECT  36935.0 52930.0 37640.0 51585.0 ;
      RECT  36935.0 52930.0 37640.0 54275.0 ;
      RECT  36935.0 55620.0 37640.0 54275.0 ;
      RECT  36935.0 55620.0 37640.0 56965.0 ;
      RECT  36935.0 58310.0 37640.0 56965.0 ;
      RECT  36935.0 58310.0 37640.0 59655.0 ;
      RECT  36935.0 61000.0 37640.0 59655.0 ;
      RECT  36935.0 61000.0 37640.0 62345.0 ;
      RECT  36935.0 63690.0 37640.0 62345.0 ;
      RECT  36935.0 63690.0 37640.0 65035.0 ;
      RECT  36935.0 66380.0 37640.0 65035.0 ;
      RECT  36935.0 66380.0 37640.0 67725.0 ;
      RECT  36935.0 69070.0 37640.0 67725.0 ;
      RECT  36935.0 69070.0 37640.0 70415.0 ;
      RECT  36935.0 71760.0 37640.0 70415.0 ;
      RECT  36935.0 71760.0 37640.0 73105.0 ;
      RECT  36935.0 74450.0 37640.0 73105.0 ;
      RECT  36935.0 74450.0 37640.0 75795.0 ;
      RECT  36935.0 77140.0 37640.0 75795.0 ;
      RECT  36935.0 77140.0 37640.0 78485.0 ;
      RECT  36935.0 79830.0 37640.0 78485.0 ;
      RECT  36935.0 79830.0 37640.0 81175.0 ;
      RECT  36935.0 82520.0 37640.0 81175.0 ;
      RECT  36935.0 82520.0 37640.0 83865.0 ;
      RECT  36935.0 85210.0 37640.0 83865.0 ;
      RECT  36935.0 85210.0 37640.0 86555.0 ;
      RECT  36935.0 87900.0 37640.0 86555.0 ;
      RECT  36935.0 87900.0 37640.0 89245.0 ;
      RECT  36935.0 90590.0 37640.0 89245.0 ;
      RECT  36935.0 90590.0 37640.0 91935.0 ;
      RECT  36935.0 93280.0 37640.0 91935.0 ;
      RECT  36935.0 93280.0 37640.0 94625.0 ;
      RECT  36935.0 95970.0 37640.0 94625.0 ;
      RECT  36935.0 95970.0 37640.0 97315.0 ;
      RECT  36935.0 98660.0 37640.0 97315.0 ;
      RECT  36935.0 98660.0 37640.0 100005.0 ;
      RECT  36935.0 101350.0 37640.0 100005.0 ;
      RECT  36935.0 101350.0 37640.0 102695.0 ;
      RECT  36935.0 104040.0 37640.0 102695.0 ;
      RECT  36935.0 104040.0 37640.0 105385.0 ;
      RECT  36935.0 106730.0 37640.0 105385.0 ;
      RECT  36935.0 106730.0 37640.0 108075.0 ;
      RECT  36935.0 109420.0 37640.0 108075.0 ;
      RECT  36935.0 109420.0 37640.0 110765.0 ;
      RECT  36935.0 112110.0 37640.0 110765.0 ;
      RECT  36935.0 112110.0 37640.0 113455.0 ;
      RECT  36935.0 114800.0 37640.0 113455.0 ;
      RECT  36935.0 114800.0 37640.0 116145.0 ;
      RECT  36935.0 117490.0 37640.0 116145.0 ;
      RECT  36935.0 117490.0 37640.0 118835.0 ;
      RECT  36935.0 120180.0 37640.0 118835.0 ;
      RECT  36935.0 120180.0 37640.0 121525.0 ;
      RECT  36935.0 122870.0 37640.0 121525.0 ;
      RECT  36935.0 122870.0 37640.0 124215.0 ;
      RECT  36935.0 125560.0 37640.0 124215.0 ;
      RECT  36935.0 125560.0 37640.0 126905.0 ;
      RECT  36935.0 128250.0 37640.0 126905.0 ;
      RECT  36935.0 128250.0 37640.0 129595.0 ;
      RECT  36935.0 130940.0 37640.0 129595.0 ;
      RECT  36935.0 130940.0 37640.0 132285.0 ;
      RECT  36935.0 133630.0 37640.0 132285.0 ;
      RECT  36935.0 133630.0 37640.0 134975.0 ;
      RECT  36935.0 136320.0 37640.0 134975.0 ;
      RECT  36935.0 136320.0 37640.0 137665.0 ;
      RECT  36935.0 139010.0 37640.0 137665.0 ;
      RECT  36935.0 139010.0 37640.0 140355.0 ;
      RECT  36935.0 141700.0 37640.0 140355.0 ;
      RECT  36935.0 141700.0 37640.0 143045.0 ;
      RECT  36935.0 144390.0 37640.0 143045.0 ;
      RECT  36935.0 144390.0 37640.0 145735.0 ;
      RECT  36935.0 147080.0 37640.0 145735.0 ;
      RECT  36935.0 147080.0 37640.0 148425.0 ;
      RECT  36935.0 149770.0 37640.0 148425.0 ;
      RECT  36935.0 149770.0 37640.0 151115.0 ;
      RECT  36935.0 152460.0 37640.0 151115.0 ;
      RECT  36935.0 152460.0 37640.0 153805.0 ;
      RECT  36935.0 155150.0 37640.0 153805.0 ;
      RECT  36935.0 155150.0 37640.0 156495.0 ;
      RECT  36935.0 157840.0 37640.0 156495.0 ;
      RECT  36935.0 157840.0 37640.0 159185.0 ;
      RECT  36935.0 160530.0 37640.0 159185.0 ;
      RECT  36935.0 160530.0 37640.0 161875.0 ;
      RECT  36935.0 163220.0 37640.0 161875.0 ;
      RECT  36935.0 163220.0 37640.0 164565.0 ;
      RECT  36935.0 165910.0 37640.0 164565.0 ;
      RECT  36935.0 165910.0 37640.0 167255.0 ;
      RECT  36935.0 168600.0 37640.0 167255.0 ;
      RECT  36935.0 168600.0 37640.0 169945.0 ;
      RECT  36935.0 171290.0 37640.0 169945.0 ;
      RECT  36935.0 171290.0 37640.0 172635.0 ;
      RECT  36935.0 173980.0 37640.0 172635.0 ;
      RECT  36935.0 173980.0 37640.0 175325.0 ;
      RECT  36935.0 176670.0 37640.0 175325.0 ;
      RECT  36935.0 176670.0 37640.0 178015.0 ;
      RECT  36935.0 179360.0 37640.0 178015.0 ;
      RECT  36935.0 179360.0 37640.0 180705.0 ;
      RECT  36935.0 182050.0 37640.0 180705.0 ;
      RECT  36935.0 182050.0 37640.0 183395.0 ;
      RECT  36935.0 184740.0 37640.0 183395.0 ;
      RECT  36935.0 184740.0 37640.0 186085.0 ;
      RECT  36935.0 187430.0 37640.0 186085.0 ;
      RECT  36935.0 187430.0 37640.0 188775.0 ;
      RECT  36935.0 190120.0 37640.0 188775.0 ;
      RECT  36935.0 190120.0 37640.0 191465.0 ;
      RECT  36935.0 192810.0 37640.0 191465.0 ;
      RECT  36935.0 192810.0 37640.0 194155.0 ;
      RECT  36935.0 195500.0 37640.0 194155.0 ;
      RECT  36935.0 195500.0 37640.0 196845.0 ;
      RECT  36935.0 198190.0 37640.0 196845.0 ;
      RECT  36935.0 198190.0 37640.0 199535.0 ;
      RECT  36935.0 200880.0 37640.0 199535.0 ;
      RECT  36935.0 200880.0 37640.0 202225.0 ;
      RECT  36935.0 203570.0 37640.0 202225.0 ;
      RECT  36935.0 203570.0 37640.0 204915.0 ;
      RECT  36935.0 206260.0 37640.0 204915.0 ;
      RECT  37640.0 34100.0 38345.0 35445.0 ;
      RECT  37640.0 36790.0 38345.0 35445.0 ;
      RECT  37640.0 36790.0 38345.0 38135.0 ;
      RECT  37640.0 39480.0 38345.0 38135.0 ;
      RECT  37640.0 39480.0 38345.0 40825.0 ;
      RECT  37640.0 42170.0 38345.0 40825.0 ;
      RECT  37640.0 42170.0 38345.0 43515.0 ;
      RECT  37640.0 44860.0 38345.0 43515.0 ;
      RECT  37640.0 44860.0 38345.0 46205.0 ;
      RECT  37640.0 47550.0 38345.0 46205.0 ;
      RECT  37640.0 47550.0 38345.0 48895.0 ;
      RECT  37640.0 50240.0 38345.0 48895.0 ;
      RECT  37640.0 50240.0 38345.0 51585.0 ;
      RECT  37640.0 52930.0 38345.0 51585.0 ;
      RECT  37640.0 52930.0 38345.0 54275.0 ;
      RECT  37640.0 55620.0 38345.0 54275.0 ;
      RECT  37640.0 55620.0 38345.0 56965.0 ;
      RECT  37640.0 58310.0 38345.0 56965.0 ;
      RECT  37640.0 58310.0 38345.0 59655.0 ;
      RECT  37640.0 61000.0 38345.0 59655.0 ;
      RECT  37640.0 61000.0 38345.0 62345.0 ;
      RECT  37640.0 63690.0 38345.0 62345.0 ;
      RECT  37640.0 63690.0 38345.0 65035.0 ;
      RECT  37640.0 66380.0 38345.0 65035.0 ;
      RECT  37640.0 66380.0 38345.0 67725.0 ;
      RECT  37640.0 69070.0 38345.0 67725.0 ;
      RECT  37640.0 69070.0 38345.0 70415.0 ;
      RECT  37640.0 71760.0 38345.0 70415.0 ;
      RECT  37640.0 71760.0 38345.0 73105.0 ;
      RECT  37640.0 74450.0 38345.0 73105.0 ;
      RECT  37640.0 74450.0 38345.0 75795.0 ;
      RECT  37640.0 77140.0 38345.0 75795.0 ;
      RECT  37640.0 77140.0 38345.0 78485.0 ;
      RECT  37640.0 79830.0 38345.0 78485.0 ;
      RECT  37640.0 79830.0 38345.0 81175.0 ;
      RECT  37640.0 82520.0 38345.0 81175.0 ;
      RECT  37640.0 82520.0 38345.0 83865.0 ;
      RECT  37640.0 85210.0 38345.0 83865.0 ;
      RECT  37640.0 85210.0 38345.0 86555.0 ;
      RECT  37640.0 87900.0 38345.0 86555.0 ;
      RECT  37640.0 87900.0 38345.0 89245.0 ;
      RECT  37640.0 90590.0 38345.0 89245.0 ;
      RECT  37640.0 90590.0 38345.0 91935.0 ;
      RECT  37640.0 93280.0 38345.0 91935.0 ;
      RECT  37640.0 93280.0 38345.0 94625.0 ;
      RECT  37640.0 95970.0 38345.0 94625.0 ;
      RECT  37640.0 95970.0 38345.0 97315.0 ;
      RECT  37640.0 98660.0 38345.0 97315.0 ;
      RECT  37640.0 98660.0 38345.0 100005.0 ;
      RECT  37640.0 101350.0 38345.0 100005.0 ;
      RECT  37640.0 101350.0 38345.0 102695.0 ;
      RECT  37640.0 104040.0 38345.0 102695.0 ;
      RECT  37640.0 104040.0 38345.0 105385.0 ;
      RECT  37640.0 106730.0 38345.0 105385.0 ;
      RECT  37640.0 106730.0 38345.0 108075.0 ;
      RECT  37640.0 109420.0 38345.0 108075.0 ;
      RECT  37640.0 109420.0 38345.0 110765.0 ;
      RECT  37640.0 112110.0 38345.0 110765.0 ;
      RECT  37640.0 112110.0 38345.0 113455.0 ;
      RECT  37640.0 114800.0 38345.0 113455.0 ;
      RECT  37640.0 114800.0 38345.0 116145.0 ;
      RECT  37640.0 117490.0 38345.0 116145.0 ;
      RECT  37640.0 117490.0 38345.0 118835.0 ;
      RECT  37640.0 120180.0 38345.0 118835.0 ;
      RECT  37640.0 120180.0 38345.0 121525.0 ;
      RECT  37640.0 122870.0 38345.0 121525.0 ;
      RECT  37640.0 122870.0 38345.0 124215.0 ;
      RECT  37640.0 125560.0 38345.0 124215.0 ;
      RECT  37640.0 125560.0 38345.0 126905.0 ;
      RECT  37640.0 128250.0 38345.0 126905.0 ;
      RECT  37640.0 128250.0 38345.0 129595.0 ;
      RECT  37640.0 130940.0 38345.0 129595.0 ;
      RECT  37640.0 130940.0 38345.0 132285.0 ;
      RECT  37640.0 133630.0 38345.0 132285.0 ;
      RECT  37640.0 133630.0 38345.0 134975.0 ;
      RECT  37640.0 136320.0 38345.0 134975.0 ;
      RECT  37640.0 136320.0 38345.0 137665.0 ;
      RECT  37640.0 139010.0 38345.0 137665.0 ;
      RECT  37640.0 139010.0 38345.0 140355.0 ;
      RECT  37640.0 141700.0 38345.0 140355.0 ;
      RECT  37640.0 141700.0 38345.0 143045.0 ;
      RECT  37640.0 144390.0 38345.0 143045.0 ;
      RECT  37640.0 144390.0 38345.0 145735.0 ;
      RECT  37640.0 147080.0 38345.0 145735.0 ;
      RECT  37640.0 147080.0 38345.0 148425.0 ;
      RECT  37640.0 149770.0 38345.0 148425.0 ;
      RECT  37640.0 149770.0 38345.0 151115.0 ;
      RECT  37640.0 152460.0 38345.0 151115.0 ;
      RECT  37640.0 152460.0 38345.0 153805.0 ;
      RECT  37640.0 155150.0 38345.0 153805.0 ;
      RECT  37640.0 155150.0 38345.0 156495.0 ;
      RECT  37640.0 157840.0 38345.0 156495.0 ;
      RECT  37640.0 157840.0 38345.0 159185.0 ;
      RECT  37640.0 160530.0 38345.0 159185.0 ;
      RECT  37640.0 160530.0 38345.0 161875.0 ;
      RECT  37640.0 163220.0 38345.0 161875.0 ;
      RECT  37640.0 163220.0 38345.0 164565.0 ;
      RECT  37640.0 165910.0 38345.0 164565.0 ;
      RECT  37640.0 165910.0 38345.0 167255.0 ;
      RECT  37640.0 168600.0 38345.0 167255.0 ;
      RECT  37640.0 168600.0 38345.0 169945.0 ;
      RECT  37640.0 171290.0 38345.0 169945.0 ;
      RECT  37640.0 171290.0 38345.0 172635.0 ;
      RECT  37640.0 173980.0 38345.0 172635.0 ;
      RECT  37640.0 173980.0 38345.0 175325.0 ;
      RECT  37640.0 176670.0 38345.0 175325.0 ;
      RECT  37640.0 176670.0 38345.0 178015.0 ;
      RECT  37640.0 179360.0 38345.0 178015.0 ;
      RECT  37640.0 179360.0 38345.0 180705.0 ;
      RECT  37640.0 182050.0 38345.0 180705.0 ;
      RECT  37640.0 182050.0 38345.0 183395.0 ;
      RECT  37640.0 184740.0 38345.0 183395.0 ;
      RECT  37640.0 184740.0 38345.0 186085.0 ;
      RECT  37640.0 187430.0 38345.0 186085.0 ;
      RECT  37640.0 187430.0 38345.0 188775.0 ;
      RECT  37640.0 190120.0 38345.0 188775.0 ;
      RECT  37640.0 190120.0 38345.0 191465.0 ;
      RECT  37640.0 192810.0 38345.0 191465.0 ;
      RECT  37640.0 192810.0 38345.0 194155.0 ;
      RECT  37640.0 195500.0 38345.0 194155.0 ;
      RECT  37640.0 195500.0 38345.0 196845.0 ;
      RECT  37640.0 198190.0 38345.0 196845.0 ;
      RECT  37640.0 198190.0 38345.0 199535.0 ;
      RECT  37640.0 200880.0 38345.0 199535.0 ;
      RECT  37640.0 200880.0 38345.0 202225.0 ;
      RECT  37640.0 203570.0 38345.0 202225.0 ;
      RECT  37640.0 203570.0 38345.0 204915.0 ;
      RECT  37640.0 206260.0 38345.0 204915.0 ;
      RECT  38345.0 34100.0 39050.0 35445.0 ;
      RECT  38345.0 36790.0 39050.0 35445.0 ;
      RECT  38345.0 36790.0 39050.0 38135.0 ;
      RECT  38345.0 39480.0 39050.0 38135.0 ;
      RECT  38345.0 39480.0 39050.0 40825.0 ;
      RECT  38345.0 42170.0 39050.0 40825.0 ;
      RECT  38345.0 42170.0 39050.0 43515.0 ;
      RECT  38345.0 44860.0 39050.0 43515.0 ;
      RECT  38345.0 44860.0 39050.0 46205.0 ;
      RECT  38345.0 47550.0 39050.0 46205.0 ;
      RECT  38345.0 47550.0 39050.0 48895.0 ;
      RECT  38345.0 50240.0 39050.0 48895.0 ;
      RECT  38345.0 50240.0 39050.0 51585.0 ;
      RECT  38345.0 52930.0 39050.0 51585.0 ;
      RECT  38345.0 52930.0 39050.0 54275.0 ;
      RECT  38345.0 55620.0 39050.0 54275.0 ;
      RECT  38345.0 55620.0 39050.0 56965.0 ;
      RECT  38345.0 58310.0 39050.0 56965.0 ;
      RECT  38345.0 58310.0 39050.0 59655.0 ;
      RECT  38345.0 61000.0 39050.0 59655.0 ;
      RECT  38345.0 61000.0 39050.0 62345.0 ;
      RECT  38345.0 63690.0 39050.0 62345.0 ;
      RECT  38345.0 63690.0 39050.0 65035.0 ;
      RECT  38345.0 66380.0 39050.0 65035.0 ;
      RECT  38345.0 66380.0 39050.0 67725.0 ;
      RECT  38345.0 69070.0 39050.0 67725.0 ;
      RECT  38345.0 69070.0 39050.0 70415.0 ;
      RECT  38345.0 71760.0 39050.0 70415.0 ;
      RECT  38345.0 71760.0 39050.0 73105.0 ;
      RECT  38345.0 74450.0 39050.0 73105.0 ;
      RECT  38345.0 74450.0 39050.0 75795.0 ;
      RECT  38345.0 77140.0 39050.0 75795.0 ;
      RECT  38345.0 77140.0 39050.0 78485.0 ;
      RECT  38345.0 79830.0 39050.0 78485.0 ;
      RECT  38345.0 79830.0 39050.0 81175.0 ;
      RECT  38345.0 82520.0 39050.0 81175.0 ;
      RECT  38345.0 82520.0 39050.0 83865.0 ;
      RECT  38345.0 85210.0 39050.0 83865.0 ;
      RECT  38345.0 85210.0 39050.0 86555.0 ;
      RECT  38345.0 87900.0 39050.0 86555.0 ;
      RECT  38345.0 87900.0 39050.0 89245.0 ;
      RECT  38345.0 90590.0 39050.0 89245.0 ;
      RECT  38345.0 90590.0 39050.0 91935.0 ;
      RECT  38345.0 93280.0 39050.0 91935.0 ;
      RECT  38345.0 93280.0 39050.0 94625.0 ;
      RECT  38345.0 95970.0 39050.0 94625.0 ;
      RECT  38345.0 95970.0 39050.0 97315.0 ;
      RECT  38345.0 98660.0 39050.0 97315.0 ;
      RECT  38345.0 98660.0 39050.0 100005.0 ;
      RECT  38345.0 101350.0 39050.0 100005.0 ;
      RECT  38345.0 101350.0 39050.0 102695.0 ;
      RECT  38345.0 104040.0 39050.0 102695.0 ;
      RECT  38345.0 104040.0 39050.0 105385.0 ;
      RECT  38345.0 106730.0 39050.0 105385.0 ;
      RECT  38345.0 106730.0 39050.0 108075.0 ;
      RECT  38345.0 109420.0 39050.0 108075.0 ;
      RECT  38345.0 109420.0 39050.0 110765.0 ;
      RECT  38345.0 112110.0 39050.0 110765.0 ;
      RECT  38345.0 112110.0 39050.0 113455.0 ;
      RECT  38345.0 114800.0 39050.0 113455.0 ;
      RECT  38345.0 114800.0 39050.0 116145.0 ;
      RECT  38345.0 117490.0 39050.0 116145.0 ;
      RECT  38345.0 117490.0 39050.0 118835.0 ;
      RECT  38345.0 120180.0 39050.0 118835.0 ;
      RECT  38345.0 120180.0 39050.0 121525.0 ;
      RECT  38345.0 122870.0 39050.0 121525.0 ;
      RECT  38345.0 122870.0 39050.0 124215.0 ;
      RECT  38345.0 125560.0 39050.0 124215.0 ;
      RECT  38345.0 125560.0 39050.0 126905.0 ;
      RECT  38345.0 128250.0 39050.0 126905.0 ;
      RECT  38345.0 128250.0 39050.0 129595.0 ;
      RECT  38345.0 130940.0 39050.0 129595.0 ;
      RECT  38345.0 130940.0 39050.0 132285.0 ;
      RECT  38345.0 133630.0 39050.0 132285.0 ;
      RECT  38345.0 133630.0 39050.0 134975.0 ;
      RECT  38345.0 136320.0 39050.0 134975.0 ;
      RECT  38345.0 136320.0 39050.0 137665.0 ;
      RECT  38345.0 139010.0 39050.0 137665.0 ;
      RECT  38345.0 139010.0 39050.0 140355.0 ;
      RECT  38345.0 141700.0 39050.0 140355.0 ;
      RECT  38345.0 141700.0 39050.0 143045.0 ;
      RECT  38345.0 144390.0 39050.0 143045.0 ;
      RECT  38345.0 144390.0 39050.0 145735.0 ;
      RECT  38345.0 147080.0 39050.0 145735.0 ;
      RECT  38345.0 147080.0 39050.0 148425.0 ;
      RECT  38345.0 149770.0 39050.0 148425.0 ;
      RECT  38345.0 149770.0 39050.0 151115.0 ;
      RECT  38345.0 152460.0 39050.0 151115.0 ;
      RECT  38345.0 152460.0 39050.0 153805.0 ;
      RECT  38345.0 155150.0 39050.0 153805.0 ;
      RECT  38345.0 155150.0 39050.0 156495.0 ;
      RECT  38345.0 157840.0 39050.0 156495.0 ;
      RECT  38345.0 157840.0 39050.0 159185.0 ;
      RECT  38345.0 160530.0 39050.0 159185.0 ;
      RECT  38345.0 160530.0 39050.0 161875.0 ;
      RECT  38345.0 163220.0 39050.0 161875.0 ;
      RECT  38345.0 163220.0 39050.0 164565.0 ;
      RECT  38345.0 165910.0 39050.0 164565.0 ;
      RECT  38345.0 165910.0 39050.0 167255.0 ;
      RECT  38345.0 168600.0 39050.0 167255.0 ;
      RECT  38345.0 168600.0 39050.0 169945.0 ;
      RECT  38345.0 171290.0 39050.0 169945.0 ;
      RECT  38345.0 171290.0 39050.0 172635.0 ;
      RECT  38345.0 173980.0 39050.0 172635.0 ;
      RECT  38345.0 173980.0 39050.0 175325.0 ;
      RECT  38345.0 176670.0 39050.0 175325.0 ;
      RECT  38345.0 176670.0 39050.0 178015.0 ;
      RECT  38345.0 179360.0 39050.0 178015.0 ;
      RECT  38345.0 179360.0 39050.0 180705.0 ;
      RECT  38345.0 182050.0 39050.0 180705.0 ;
      RECT  38345.0 182050.0 39050.0 183395.0 ;
      RECT  38345.0 184740.0 39050.0 183395.0 ;
      RECT  38345.0 184740.0 39050.0 186085.0 ;
      RECT  38345.0 187430.0 39050.0 186085.0 ;
      RECT  38345.0 187430.0 39050.0 188775.0 ;
      RECT  38345.0 190120.0 39050.0 188775.0 ;
      RECT  38345.0 190120.0 39050.0 191465.0 ;
      RECT  38345.0 192810.0 39050.0 191465.0 ;
      RECT  38345.0 192810.0 39050.0 194155.0 ;
      RECT  38345.0 195500.0 39050.0 194155.0 ;
      RECT  38345.0 195500.0 39050.0 196845.0 ;
      RECT  38345.0 198190.0 39050.0 196845.0 ;
      RECT  38345.0 198190.0 39050.0 199535.0 ;
      RECT  38345.0 200880.0 39050.0 199535.0 ;
      RECT  38345.0 200880.0 39050.0 202225.0 ;
      RECT  38345.0 203570.0 39050.0 202225.0 ;
      RECT  38345.0 203570.0 39050.0 204915.0 ;
      RECT  38345.0 206260.0 39050.0 204915.0 ;
      RECT  39050.0 34100.0 39755.0 35445.0 ;
      RECT  39050.0 36790.0 39755.0 35445.0 ;
      RECT  39050.0 36790.0 39755.0 38135.0 ;
      RECT  39050.0 39480.0 39755.0 38135.0 ;
      RECT  39050.0 39480.0 39755.0 40825.0 ;
      RECT  39050.0 42170.0 39755.0 40825.0 ;
      RECT  39050.0 42170.0 39755.0 43515.0 ;
      RECT  39050.0 44860.0 39755.0 43515.0 ;
      RECT  39050.0 44860.0 39755.0 46205.0 ;
      RECT  39050.0 47550.0 39755.0 46205.0 ;
      RECT  39050.0 47550.0 39755.0 48895.0 ;
      RECT  39050.0 50240.0 39755.0 48895.0 ;
      RECT  39050.0 50240.0 39755.0 51585.0 ;
      RECT  39050.0 52930.0 39755.0 51585.0 ;
      RECT  39050.0 52930.0 39755.0 54275.0 ;
      RECT  39050.0 55620.0 39755.0 54275.0 ;
      RECT  39050.0 55620.0 39755.0 56965.0 ;
      RECT  39050.0 58310.0 39755.0 56965.0 ;
      RECT  39050.0 58310.0 39755.0 59655.0 ;
      RECT  39050.0 61000.0 39755.0 59655.0 ;
      RECT  39050.0 61000.0 39755.0 62345.0 ;
      RECT  39050.0 63690.0 39755.0 62345.0 ;
      RECT  39050.0 63690.0 39755.0 65035.0 ;
      RECT  39050.0 66380.0 39755.0 65035.0 ;
      RECT  39050.0 66380.0 39755.0 67725.0 ;
      RECT  39050.0 69070.0 39755.0 67725.0 ;
      RECT  39050.0 69070.0 39755.0 70415.0 ;
      RECT  39050.0 71760.0 39755.0 70415.0 ;
      RECT  39050.0 71760.0 39755.0 73105.0 ;
      RECT  39050.0 74450.0 39755.0 73105.0 ;
      RECT  39050.0 74450.0 39755.0 75795.0 ;
      RECT  39050.0 77140.0 39755.0 75795.0 ;
      RECT  39050.0 77140.0 39755.0 78485.0 ;
      RECT  39050.0 79830.0 39755.0 78485.0 ;
      RECT  39050.0 79830.0 39755.0 81175.0 ;
      RECT  39050.0 82520.0 39755.0 81175.0 ;
      RECT  39050.0 82520.0 39755.0 83865.0 ;
      RECT  39050.0 85210.0 39755.0 83865.0 ;
      RECT  39050.0 85210.0 39755.0 86555.0 ;
      RECT  39050.0 87900.0 39755.0 86555.0 ;
      RECT  39050.0 87900.0 39755.0 89245.0 ;
      RECT  39050.0 90590.0 39755.0 89245.0 ;
      RECT  39050.0 90590.0 39755.0 91935.0 ;
      RECT  39050.0 93280.0 39755.0 91935.0 ;
      RECT  39050.0 93280.0 39755.0 94625.0 ;
      RECT  39050.0 95970.0 39755.0 94625.0 ;
      RECT  39050.0 95970.0 39755.0 97315.0 ;
      RECT  39050.0 98660.0 39755.0 97315.0 ;
      RECT  39050.0 98660.0 39755.0 100005.0 ;
      RECT  39050.0 101350.0 39755.0 100005.0 ;
      RECT  39050.0 101350.0 39755.0 102695.0 ;
      RECT  39050.0 104040.0 39755.0 102695.0 ;
      RECT  39050.0 104040.0 39755.0 105385.0 ;
      RECT  39050.0 106730.0 39755.0 105385.0 ;
      RECT  39050.0 106730.0 39755.0 108075.0 ;
      RECT  39050.0 109420.0 39755.0 108075.0 ;
      RECT  39050.0 109420.0 39755.0 110765.0 ;
      RECT  39050.0 112110.0 39755.0 110765.0 ;
      RECT  39050.0 112110.0 39755.0 113455.0 ;
      RECT  39050.0 114800.0 39755.0 113455.0 ;
      RECT  39050.0 114800.0 39755.0 116145.0 ;
      RECT  39050.0 117490.0 39755.0 116145.0 ;
      RECT  39050.0 117490.0 39755.0 118835.0 ;
      RECT  39050.0 120180.0 39755.0 118835.0 ;
      RECT  39050.0 120180.0 39755.0 121525.0 ;
      RECT  39050.0 122870.0 39755.0 121525.0 ;
      RECT  39050.0 122870.0 39755.0 124215.0 ;
      RECT  39050.0 125560.0 39755.0 124215.0 ;
      RECT  39050.0 125560.0 39755.0 126905.0 ;
      RECT  39050.0 128250.0 39755.0 126905.0 ;
      RECT  39050.0 128250.0 39755.0 129595.0 ;
      RECT  39050.0 130940.0 39755.0 129595.0 ;
      RECT  39050.0 130940.0 39755.0 132285.0 ;
      RECT  39050.0 133630.0 39755.0 132285.0 ;
      RECT  39050.0 133630.0 39755.0 134975.0 ;
      RECT  39050.0 136320.0 39755.0 134975.0 ;
      RECT  39050.0 136320.0 39755.0 137665.0 ;
      RECT  39050.0 139010.0 39755.0 137665.0 ;
      RECT  39050.0 139010.0 39755.0 140355.0 ;
      RECT  39050.0 141700.0 39755.0 140355.0 ;
      RECT  39050.0 141700.0 39755.0 143045.0 ;
      RECT  39050.0 144390.0 39755.0 143045.0 ;
      RECT  39050.0 144390.0 39755.0 145735.0 ;
      RECT  39050.0 147080.0 39755.0 145735.0 ;
      RECT  39050.0 147080.0 39755.0 148425.0 ;
      RECT  39050.0 149770.0 39755.0 148425.0 ;
      RECT  39050.0 149770.0 39755.0 151115.0 ;
      RECT  39050.0 152460.0 39755.0 151115.0 ;
      RECT  39050.0 152460.0 39755.0 153805.0 ;
      RECT  39050.0 155150.0 39755.0 153805.0 ;
      RECT  39050.0 155150.0 39755.0 156495.0 ;
      RECT  39050.0 157840.0 39755.0 156495.0 ;
      RECT  39050.0 157840.0 39755.0 159185.0 ;
      RECT  39050.0 160530.0 39755.0 159185.0 ;
      RECT  39050.0 160530.0 39755.0 161875.0 ;
      RECT  39050.0 163220.0 39755.0 161875.0 ;
      RECT  39050.0 163220.0 39755.0 164565.0 ;
      RECT  39050.0 165910.0 39755.0 164565.0 ;
      RECT  39050.0 165910.0 39755.0 167255.0 ;
      RECT  39050.0 168600.0 39755.0 167255.0 ;
      RECT  39050.0 168600.0 39755.0 169945.0 ;
      RECT  39050.0 171290.0 39755.0 169945.0 ;
      RECT  39050.0 171290.0 39755.0 172635.0 ;
      RECT  39050.0 173980.0 39755.0 172635.0 ;
      RECT  39050.0 173980.0 39755.0 175325.0 ;
      RECT  39050.0 176670.0 39755.0 175325.0 ;
      RECT  39050.0 176670.0 39755.0 178015.0 ;
      RECT  39050.0 179360.0 39755.0 178015.0 ;
      RECT  39050.0 179360.0 39755.0 180705.0 ;
      RECT  39050.0 182050.0 39755.0 180705.0 ;
      RECT  39050.0 182050.0 39755.0 183395.0 ;
      RECT  39050.0 184740.0 39755.0 183395.0 ;
      RECT  39050.0 184740.0 39755.0 186085.0 ;
      RECT  39050.0 187430.0 39755.0 186085.0 ;
      RECT  39050.0 187430.0 39755.0 188775.0 ;
      RECT  39050.0 190120.0 39755.0 188775.0 ;
      RECT  39050.0 190120.0 39755.0 191465.0 ;
      RECT  39050.0 192810.0 39755.0 191465.0 ;
      RECT  39050.0 192810.0 39755.0 194155.0 ;
      RECT  39050.0 195500.0 39755.0 194155.0 ;
      RECT  39050.0 195500.0 39755.0 196845.0 ;
      RECT  39050.0 198190.0 39755.0 196845.0 ;
      RECT  39050.0 198190.0 39755.0 199535.0 ;
      RECT  39050.0 200880.0 39755.0 199535.0 ;
      RECT  39050.0 200880.0 39755.0 202225.0 ;
      RECT  39050.0 203570.0 39755.0 202225.0 ;
      RECT  39050.0 203570.0 39755.0 204915.0 ;
      RECT  39050.0 206260.0 39755.0 204915.0 ;
      RECT  39755.0 34100.0 40460.0 35445.0 ;
      RECT  39755.0 36790.0 40460.0 35445.0 ;
      RECT  39755.0 36790.0 40460.0 38135.0 ;
      RECT  39755.0 39480.0 40460.0 38135.0 ;
      RECT  39755.0 39480.0 40460.0 40825.0 ;
      RECT  39755.0 42170.0 40460.0 40825.0 ;
      RECT  39755.0 42170.0 40460.0 43515.0 ;
      RECT  39755.0 44860.0 40460.0 43515.0 ;
      RECT  39755.0 44860.0 40460.0 46205.0 ;
      RECT  39755.0 47550.0 40460.0 46205.0 ;
      RECT  39755.0 47550.0 40460.0 48895.0 ;
      RECT  39755.0 50240.0 40460.0 48895.0 ;
      RECT  39755.0 50240.0 40460.0 51585.0 ;
      RECT  39755.0 52930.0 40460.0 51585.0 ;
      RECT  39755.0 52930.0 40460.0 54275.0 ;
      RECT  39755.0 55620.0 40460.0 54275.0 ;
      RECT  39755.0 55620.0 40460.0 56965.0 ;
      RECT  39755.0 58310.0 40460.0 56965.0 ;
      RECT  39755.0 58310.0 40460.0 59655.0 ;
      RECT  39755.0 61000.0 40460.0 59655.0 ;
      RECT  39755.0 61000.0 40460.0 62345.0 ;
      RECT  39755.0 63690.0 40460.0 62345.0 ;
      RECT  39755.0 63690.0 40460.0 65035.0 ;
      RECT  39755.0 66380.0 40460.0 65035.0 ;
      RECT  39755.0 66380.0 40460.0 67725.0 ;
      RECT  39755.0 69070.0 40460.0 67725.0 ;
      RECT  39755.0 69070.0 40460.0 70415.0 ;
      RECT  39755.0 71760.0 40460.0 70415.0 ;
      RECT  39755.0 71760.0 40460.0 73105.0 ;
      RECT  39755.0 74450.0 40460.0 73105.0 ;
      RECT  39755.0 74450.0 40460.0 75795.0 ;
      RECT  39755.0 77140.0 40460.0 75795.0 ;
      RECT  39755.0 77140.0 40460.0 78485.0 ;
      RECT  39755.0 79830.0 40460.0 78485.0 ;
      RECT  39755.0 79830.0 40460.0 81175.0 ;
      RECT  39755.0 82520.0 40460.0 81175.0 ;
      RECT  39755.0 82520.0 40460.0 83865.0 ;
      RECT  39755.0 85210.0 40460.0 83865.0 ;
      RECT  39755.0 85210.0 40460.0 86555.0 ;
      RECT  39755.0 87900.0 40460.0 86555.0 ;
      RECT  39755.0 87900.0 40460.0 89245.0 ;
      RECT  39755.0 90590.0 40460.0 89245.0 ;
      RECT  39755.0 90590.0 40460.0 91935.0 ;
      RECT  39755.0 93280.0 40460.0 91935.0 ;
      RECT  39755.0 93280.0 40460.0 94625.0 ;
      RECT  39755.0 95970.0 40460.0 94625.0 ;
      RECT  39755.0 95970.0 40460.0 97315.0 ;
      RECT  39755.0 98660.0 40460.0 97315.0 ;
      RECT  39755.0 98660.0 40460.0 100005.0 ;
      RECT  39755.0 101350.0 40460.0 100005.0 ;
      RECT  39755.0 101350.0 40460.0 102695.0 ;
      RECT  39755.0 104040.0 40460.0 102695.0 ;
      RECT  39755.0 104040.0 40460.0 105385.0 ;
      RECT  39755.0 106730.0 40460.0 105385.0 ;
      RECT  39755.0 106730.0 40460.0 108075.0 ;
      RECT  39755.0 109420.0 40460.0 108075.0 ;
      RECT  39755.0 109420.0 40460.0 110765.0 ;
      RECT  39755.0 112110.0 40460.0 110765.0 ;
      RECT  39755.0 112110.0 40460.0 113455.0 ;
      RECT  39755.0 114800.0 40460.0 113455.0 ;
      RECT  39755.0 114800.0 40460.0 116145.0 ;
      RECT  39755.0 117490.0 40460.0 116145.0 ;
      RECT  39755.0 117490.0 40460.0 118835.0 ;
      RECT  39755.0 120180.0 40460.0 118835.0 ;
      RECT  39755.0 120180.0 40460.0 121525.0 ;
      RECT  39755.0 122870.0 40460.0 121525.0 ;
      RECT  39755.0 122870.0 40460.0 124215.0 ;
      RECT  39755.0 125560.0 40460.0 124215.0 ;
      RECT  39755.0 125560.0 40460.0 126905.0 ;
      RECT  39755.0 128250.0 40460.0 126905.0 ;
      RECT  39755.0 128250.0 40460.0 129595.0 ;
      RECT  39755.0 130940.0 40460.0 129595.0 ;
      RECT  39755.0 130940.0 40460.0 132285.0 ;
      RECT  39755.0 133630.0 40460.0 132285.0 ;
      RECT  39755.0 133630.0 40460.0 134975.0 ;
      RECT  39755.0 136320.0 40460.0 134975.0 ;
      RECT  39755.0 136320.0 40460.0 137665.0 ;
      RECT  39755.0 139010.0 40460.0 137665.0 ;
      RECT  39755.0 139010.0 40460.0 140355.0 ;
      RECT  39755.0 141700.0 40460.0 140355.0 ;
      RECT  39755.0 141700.0 40460.0 143045.0 ;
      RECT  39755.0 144390.0 40460.0 143045.0 ;
      RECT  39755.0 144390.0 40460.0 145735.0 ;
      RECT  39755.0 147080.0 40460.0 145735.0 ;
      RECT  39755.0 147080.0 40460.0 148425.0 ;
      RECT  39755.0 149770.0 40460.0 148425.0 ;
      RECT  39755.0 149770.0 40460.0 151115.0 ;
      RECT  39755.0 152460.0 40460.0 151115.0 ;
      RECT  39755.0 152460.0 40460.0 153805.0 ;
      RECT  39755.0 155150.0 40460.0 153805.0 ;
      RECT  39755.0 155150.0 40460.0 156495.0 ;
      RECT  39755.0 157840.0 40460.0 156495.0 ;
      RECT  39755.0 157840.0 40460.0 159185.0 ;
      RECT  39755.0 160530.0 40460.0 159185.0 ;
      RECT  39755.0 160530.0 40460.0 161875.0 ;
      RECT  39755.0 163220.0 40460.0 161875.0 ;
      RECT  39755.0 163220.0 40460.0 164565.0 ;
      RECT  39755.0 165910.0 40460.0 164565.0 ;
      RECT  39755.0 165910.0 40460.0 167255.0 ;
      RECT  39755.0 168600.0 40460.0 167255.0 ;
      RECT  39755.0 168600.0 40460.0 169945.0 ;
      RECT  39755.0 171290.0 40460.0 169945.0 ;
      RECT  39755.0 171290.0 40460.0 172635.0 ;
      RECT  39755.0 173980.0 40460.0 172635.0 ;
      RECT  39755.0 173980.0 40460.0 175325.0 ;
      RECT  39755.0 176670.0 40460.0 175325.0 ;
      RECT  39755.0 176670.0 40460.0 178015.0 ;
      RECT  39755.0 179360.0 40460.0 178015.0 ;
      RECT  39755.0 179360.0 40460.0 180705.0 ;
      RECT  39755.0 182050.0 40460.0 180705.0 ;
      RECT  39755.0 182050.0 40460.0 183395.0 ;
      RECT  39755.0 184740.0 40460.0 183395.0 ;
      RECT  39755.0 184740.0 40460.0 186085.0 ;
      RECT  39755.0 187430.0 40460.0 186085.0 ;
      RECT  39755.0 187430.0 40460.0 188775.0 ;
      RECT  39755.0 190120.0 40460.0 188775.0 ;
      RECT  39755.0 190120.0 40460.0 191465.0 ;
      RECT  39755.0 192810.0 40460.0 191465.0 ;
      RECT  39755.0 192810.0 40460.0 194155.0 ;
      RECT  39755.0 195500.0 40460.0 194155.0 ;
      RECT  39755.0 195500.0 40460.0 196845.0 ;
      RECT  39755.0 198190.0 40460.0 196845.0 ;
      RECT  39755.0 198190.0 40460.0 199535.0 ;
      RECT  39755.0 200880.0 40460.0 199535.0 ;
      RECT  39755.0 200880.0 40460.0 202225.0 ;
      RECT  39755.0 203570.0 40460.0 202225.0 ;
      RECT  39755.0 203570.0 40460.0 204915.0 ;
      RECT  39755.0 206260.0 40460.0 204915.0 ;
      RECT  40460.0 34100.0 41165.0 35445.0 ;
      RECT  40460.0 36790.0 41165.0 35445.0 ;
      RECT  40460.0 36790.0 41165.0 38135.0 ;
      RECT  40460.0 39480.0 41165.0 38135.0 ;
      RECT  40460.0 39480.0 41165.0 40825.0 ;
      RECT  40460.0 42170.0 41165.0 40825.0 ;
      RECT  40460.0 42170.0 41165.0 43515.0 ;
      RECT  40460.0 44860.0 41165.0 43515.0 ;
      RECT  40460.0 44860.0 41165.0 46205.0 ;
      RECT  40460.0 47550.0 41165.0 46205.0 ;
      RECT  40460.0 47550.0 41165.0 48895.0 ;
      RECT  40460.0 50240.0 41165.0 48895.0 ;
      RECT  40460.0 50240.0 41165.0 51585.0 ;
      RECT  40460.0 52930.0 41165.0 51585.0 ;
      RECT  40460.0 52930.0 41165.0 54275.0 ;
      RECT  40460.0 55620.0 41165.0 54275.0 ;
      RECT  40460.0 55620.0 41165.0 56965.0 ;
      RECT  40460.0 58310.0 41165.0 56965.0 ;
      RECT  40460.0 58310.0 41165.0 59655.0 ;
      RECT  40460.0 61000.0 41165.0 59655.0 ;
      RECT  40460.0 61000.0 41165.0 62345.0 ;
      RECT  40460.0 63690.0 41165.0 62345.0 ;
      RECT  40460.0 63690.0 41165.0 65035.0 ;
      RECT  40460.0 66380.0 41165.0 65035.0 ;
      RECT  40460.0 66380.0 41165.0 67725.0 ;
      RECT  40460.0 69070.0 41165.0 67725.0 ;
      RECT  40460.0 69070.0 41165.0 70415.0 ;
      RECT  40460.0 71760.0 41165.0 70415.0 ;
      RECT  40460.0 71760.0 41165.0 73105.0 ;
      RECT  40460.0 74450.0 41165.0 73105.0 ;
      RECT  40460.0 74450.0 41165.0 75795.0 ;
      RECT  40460.0 77140.0 41165.0 75795.0 ;
      RECT  40460.0 77140.0 41165.0 78485.0 ;
      RECT  40460.0 79830.0 41165.0 78485.0 ;
      RECT  40460.0 79830.0 41165.0 81175.0 ;
      RECT  40460.0 82520.0 41165.0 81175.0 ;
      RECT  40460.0 82520.0 41165.0 83865.0 ;
      RECT  40460.0 85210.0 41165.0 83865.0 ;
      RECT  40460.0 85210.0 41165.0 86555.0 ;
      RECT  40460.0 87900.0 41165.0 86555.0 ;
      RECT  40460.0 87900.0 41165.0 89245.0 ;
      RECT  40460.0 90590.0 41165.0 89245.0 ;
      RECT  40460.0 90590.0 41165.0 91935.0 ;
      RECT  40460.0 93280.0 41165.0 91935.0 ;
      RECT  40460.0 93280.0 41165.0 94625.0 ;
      RECT  40460.0 95970.0 41165.0 94625.0 ;
      RECT  40460.0 95970.0 41165.0 97315.0 ;
      RECT  40460.0 98660.0 41165.0 97315.0 ;
      RECT  40460.0 98660.0 41165.0 100005.0 ;
      RECT  40460.0 101350.0 41165.0 100005.0 ;
      RECT  40460.0 101350.0 41165.0 102695.0 ;
      RECT  40460.0 104040.0 41165.0 102695.0 ;
      RECT  40460.0 104040.0 41165.0 105385.0 ;
      RECT  40460.0 106730.0 41165.0 105385.0 ;
      RECT  40460.0 106730.0 41165.0 108075.0 ;
      RECT  40460.0 109420.0 41165.0 108075.0 ;
      RECT  40460.0 109420.0 41165.0 110765.0 ;
      RECT  40460.0 112110.0 41165.0 110765.0 ;
      RECT  40460.0 112110.0 41165.0 113455.0 ;
      RECT  40460.0 114800.0 41165.0 113455.0 ;
      RECT  40460.0 114800.0 41165.0 116145.0 ;
      RECT  40460.0 117490.0 41165.0 116145.0 ;
      RECT  40460.0 117490.0 41165.0 118835.0 ;
      RECT  40460.0 120180.0 41165.0 118835.0 ;
      RECT  40460.0 120180.0 41165.0 121525.0 ;
      RECT  40460.0 122870.0 41165.0 121525.0 ;
      RECT  40460.0 122870.0 41165.0 124215.0 ;
      RECT  40460.0 125560.0 41165.0 124215.0 ;
      RECT  40460.0 125560.0 41165.0 126905.0 ;
      RECT  40460.0 128250.0 41165.0 126905.0 ;
      RECT  40460.0 128250.0 41165.0 129595.0 ;
      RECT  40460.0 130940.0 41165.0 129595.0 ;
      RECT  40460.0 130940.0 41165.0 132285.0 ;
      RECT  40460.0 133630.0 41165.0 132285.0 ;
      RECT  40460.0 133630.0 41165.0 134975.0 ;
      RECT  40460.0 136320.0 41165.0 134975.0 ;
      RECT  40460.0 136320.0 41165.0 137665.0 ;
      RECT  40460.0 139010.0 41165.0 137665.0 ;
      RECT  40460.0 139010.0 41165.0 140355.0 ;
      RECT  40460.0 141700.0 41165.0 140355.0 ;
      RECT  40460.0 141700.0 41165.0 143045.0 ;
      RECT  40460.0 144390.0 41165.0 143045.0 ;
      RECT  40460.0 144390.0 41165.0 145735.0 ;
      RECT  40460.0 147080.0 41165.0 145735.0 ;
      RECT  40460.0 147080.0 41165.0 148425.0 ;
      RECT  40460.0 149770.0 41165.0 148425.0 ;
      RECT  40460.0 149770.0 41165.0 151115.0 ;
      RECT  40460.0 152460.0 41165.0 151115.0 ;
      RECT  40460.0 152460.0 41165.0 153805.0 ;
      RECT  40460.0 155150.0 41165.0 153805.0 ;
      RECT  40460.0 155150.0 41165.0 156495.0 ;
      RECT  40460.0 157840.0 41165.0 156495.0 ;
      RECT  40460.0 157840.0 41165.0 159185.0 ;
      RECT  40460.0 160530.0 41165.0 159185.0 ;
      RECT  40460.0 160530.0 41165.0 161875.0 ;
      RECT  40460.0 163220.0 41165.0 161875.0 ;
      RECT  40460.0 163220.0 41165.0 164565.0 ;
      RECT  40460.0 165910.0 41165.0 164565.0 ;
      RECT  40460.0 165910.0 41165.0 167255.0 ;
      RECT  40460.0 168600.0 41165.0 167255.0 ;
      RECT  40460.0 168600.0 41165.0 169945.0 ;
      RECT  40460.0 171290.0 41165.0 169945.0 ;
      RECT  40460.0 171290.0 41165.0 172635.0 ;
      RECT  40460.0 173980.0 41165.0 172635.0 ;
      RECT  40460.0 173980.0 41165.0 175325.0 ;
      RECT  40460.0 176670.0 41165.0 175325.0 ;
      RECT  40460.0 176670.0 41165.0 178015.0 ;
      RECT  40460.0 179360.0 41165.0 178015.0 ;
      RECT  40460.0 179360.0 41165.0 180705.0 ;
      RECT  40460.0 182050.0 41165.0 180705.0 ;
      RECT  40460.0 182050.0 41165.0 183395.0 ;
      RECT  40460.0 184740.0 41165.0 183395.0 ;
      RECT  40460.0 184740.0 41165.0 186085.0 ;
      RECT  40460.0 187430.0 41165.0 186085.0 ;
      RECT  40460.0 187430.0 41165.0 188775.0 ;
      RECT  40460.0 190120.0 41165.0 188775.0 ;
      RECT  40460.0 190120.0 41165.0 191465.0 ;
      RECT  40460.0 192810.0 41165.0 191465.0 ;
      RECT  40460.0 192810.0 41165.0 194155.0 ;
      RECT  40460.0 195500.0 41165.0 194155.0 ;
      RECT  40460.0 195500.0 41165.0 196845.0 ;
      RECT  40460.0 198190.0 41165.0 196845.0 ;
      RECT  40460.0 198190.0 41165.0 199535.0 ;
      RECT  40460.0 200880.0 41165.0 199535.0 ;
      RECT  40460.0 200880.0 41165.0 202225.0 ;
      RECT  40460.0 203570.0 41165.0 202225.0 ;
      RECT  40460.0 203570.0 41165.0 204915.0 ;
      RECT  40460.0 206260.0 41165.0 204915.0 ;
      RECT  41165.0 34100.0 41870.0 35445.0 ;
      RECT  41165.0 36790.0 41870.0 35445.0 ;
      RECT  41165.0 36790.0 41870.0 38135.0 ;
      RECT  41165.0 39480.0 41870.0 38135.0 ;
      RECT  41165.0 39480.0 41870.0 40825.0 ;
      RECT  41165.0 42170.0 41870.0 40825.0 ;
      RECT  41165.0 42170.0 41870.0 43515.0 ;
      RECT  41165.0 44860.0 41870.0 43515.0 ;
      RECT  41165.0 44860.0 41870.0 46205.0 ;
      RECT  41165.0 47550.0 41870.0 46205.0 ;
      RECT  41165.0 47550.0 41870.0 48895.0 ;
      RECT  41165.0 50240.0 41870.0 48895.0 ;
      RECT  41165.0 50240.0 41870.0 51585.0 ;
      RECT  41165.0 52930.0 41870.0 51585.0 ;
      RECT  41165.0 52930.0 41870.0 54275.0 ;
      RECT  41165.0 55620.0 41870.0 54275.0 ;
      RECT  41165.0 55620.0 41870.0 56965.0 ;
      RECT  41165.0 58310.0 41870.0 56965.0 ;
      RECT  41165.0 58310.0 41870.0 59655.0 ;
      RECT  41165.0 61000.0 41870.0 59655.0 ;
      RECT  41165.0 61000.0 41870.0 62345.0 ;
      RECT  41165.0 63690.0 41870.0 62345.0 ;
      RECT  41165.0 63690.0 41870.0 65035.0 ;
      RECT  41165.0 66380.0 41870.0 65035.0 ;
      RECT  41165.0 66380.0 41870.0 67725.0 ;
      RECT  41165.0 69070.0 41870.0 67725.0 ;
      RECT  41165.0 69070.0 41870.0 70415.0 ;
      RECT  41165.0 71760.0 41870.0 70415.0 ;
      RECT  41165.0 71760.0 41870.0 73105.0 ;
      RECT  41165.0 74450.0 41870.0 73105.0 ;
      RECT  41165.0 74450.0 41870.0 75795.0 ;
      RECT  41165.0 77140.0 41870.0 75795.0 ;
      RECT  41165.0 77140.0 41870.0 78485.0 ;
      RECT  41165.0 79830.0 41870.0 78485.0 ;
      RECT  41165.0 79830.0 41870.0 81175.0 ;
      RECT  41165.0 82520.0 41870.0 81175.0 ;
      RECT  41165.0 82520.0 41870.0 83865.0 ;
      RECT  41165.0 85210.0 41870.0 83865.0 ;
      RECT  41165.0 85210.0 41870.0 86555.0 ;
      RECT  41165.0 87900.0 41870.0 86555.0 ;
      RECT  41165.0 87900.0 41870.0 89245.0 ;
      RECT  41165.0 90590.0 41870.0 89245.0 ;
      RECT  41165.0 90590.0 41870.0 91935.0 ;
      RECT  41165.0 93280.0 41870.0 91935.0 ;
      RECT  41165.0 93280.0 41870.0 94625.0 ;
      RECT  41165.0 95970.0 41870.0 94625.0 ;
      RECT  41165.0 95970.0 41870.0 97315.0 ;
      RECT  41165.0 98660.0 41870.0 97315.0 ;
      RECT  41165.0 98660.0 41870.0 100005.0 ;
      RECT  41165.0 101350.0 41870.0 100005.0 ;
      RECT  41165.0 101350.0 41870.0 102695.0 ;
      RECT  41165.0 104040.0 41870.0 102695.0 ;
      RECT  41165.0 104040.0 41870.0 105385.0 ;
      RECT  41165.0 106730.0 41870.0 105385.0 ;
      RECT  41165.0 106730.0 41870.0 108075.0 ;
      RECT  41165.0 109420.0 41870.0 108075.0 ;
      RECT  41165.0 109420.0 41870.0 110765.0 ;
      RECT  41165.0 112110.0 41870.0 110765.0 ;
      RECT  41165.0 112110.0 41870.0 113455.0 ;
      RECT  41165.0 114800.0 41870.0 113455.0 ;
      RECT  41165.0 114800.0 41870.0 116145.0 ;
      RECT  41165.0 117490.0 41870.0 116145.0 ;
      RECT  41165.0 117490.0 41870.0 118835.0 ;
      RECT  41165.0 120180.0 41870.0 118835.0 ;
      RECT  41165.0 120180.0 41870.0 121525.0 ;
      RECT  41165.0 122870.0 41870.0 121525.0 ;
      RECT  41165.0 122870.0 41870.0 124215.0 ;
      RECT  41165.0 125560.0 41870.0 124215.0 ;
      RECT  41165.0 125560.0 41870.0 126905.0 ;
      RECT  41165.0 128250.0 41870.0 126905.0 ;
      RECT  41165.0 128250.0 41870.0 129595.0 ;
      RECT  41165.0 130940.0 41870.0 129595.0 ;
      RECT  41165.0 130940.0 41870.0 132285.0 ;
      RECT  41165.0 133630.0 41870.0 132285.0 ;
      RECT  41165.0 133630.0 41870.0 134975.0 ;
      RECT  41165.0 136320.0 41870.0 134975.0 ;
      RECT  41165.0 136320.0 41870.0 137665.0 ;
      RECT  41165.0 139010.0 41870.0 137665.0 ;
      RECT  41165.0 139010.0 41870.0 140355.0 ;
      RECT  41165.0 141700.0 41870.0 140355.0 ;
      RECT  41165.0 141700.0 41870.0 143045.0 ;
      RECT  41165.0 144390.0 41870.0 143045.0 ;
      RECT  41165.0 144390.0 41870.0 145735.0 ;
      RECT  41165.0 147080.0 41870.0 145735.0 ;
      RECT  41165.0 147080.0 41870.0 148425.0 ;
      RECT  41165.0 149770.0 41870.0 148425.0 ;
      RECT  41165.0 149770.0 41870.0 151115.0 ;
      RECT  41165.0 152460.0 41870.0 151115.0 ;
      RECT  41165.0 152460.0 41870.0 153805.0 ;
      RECT  41165.0 155150.0 41870.0 153805.0 ;
      RECT  41165.0 155150.0 41870.0 156495.0 ;
      RECT  41165.0 157840.0 41870.0 156495.0 ;
      RECT  41165.0 157840.0 41870.0 159185.0 ;
      RECT  41165.0 160530.0 41870.0 159185.0 ;
      RECT  41165.0 160530.0 41870.0 161875.0 ;
      RECT  41165.0 163220.0 41870.0 161875.0 ;
      RECT  41165.0 163220.0 41870.0 164565.0 ;
      RECT  41165.0 165910.0 41870.0 164565.0 ;
      RECT  41165.0 165910.0 41870.0 167255.0 ;
      RECT  41165.0 168600.0 41870.0 167255.0 ;
      RECT  41165.0 168600.0 41870.0 169945.0 ;
      RECT  41165.0 171290.0 41870.0 169945.0 ;
      RECT  41165.0 171290.0 41870.0 172635.0 ;
      RECT  41165.0 173980.0 41870.0 172635.0 ;
      RECT  41165.0 173980.0 41870.0 175325.0 ;
      RECT  41165.0 176670.0 41870.0 175325.0 ;
      RECT  41165.0 176670.0 41870.0 178015.0 ;
      RECT  41165.0 179360.0 41870.0 178015.0 ;
      RECT  41165.0 179360.0 41870.0 180705.0 ;
      RECT  41165.0 182050.0 41870.0 180705.0 ;
      RECT  41165.0 182050.0 41870.0 183395.0 ;
      RECT  41165.0 184740.0 41870.0 183395.0 ;
      RECT  41165.0 184740.0 41870.0 186085.0 ;
      RECT  41165.0 187430.0 41870.0 186085.0 ;
      RECT  41165.0 187430.0 41870.0 188775.0 ;
      RECT  41165.0 190120.0 41870.0 188775.0 ;
      RECT  41165.0 190120.0 41870.0 191465.0 ;
      RECT  41165.0 192810.0 41870.0 191465.0 ;
      RECT  41165.0 192810.0 41870.0 194155.0 ;
      RECT  41165.0 195500.0 41870.0 194155.0 ;
      RECT  41165.0 195500.0 41870.0 196845.0 ;
      RECT  41165.0 198190.0 41870.0 196845.0 ;
      RECT  41165.0 198190.0 41870.0 199535.0 ;
      RECT  41165.0 200880.0 41870.0 199535.0 ;
      RECT  41165.0 200880.0 41870.0 202225.0 ;
      RECT  41165.0 203570.0 41870.0 202225.0 ;
      RECT  41165.0 203570.0 41870.0 204915.0 ;
      RECT  41165.0 206260.0 41870.0 204915.0 ;
      RECT  41870.0 34100.0 42575.0 35445.0 ;
      RECT  41870.0 36790.0 42575.0 35445.0 ;
      RECT  41870.0 36790.0 42575.0 38135.0 ;
      RECT  41870.0 39480.0 42575.0 38135.0 ;
      RECT  41870.0 39480.0 42575.0 40825.0 ;
      RECT  41870.0 42170.0 42575.0 40825.0 ;
      RECT  41870.0 42170.0 42575.0 43515.0 ;
      RECT  41870.0 44860.0 42575.0 43515.0 ;
      RECT  41870.0 44860.0 42575.0 46205.0 ;
      RECT  41870.0 47550.0 42575.0 46205.0 ;
      RECT  41870.0 47550.0 42575.0 48895.0 ;
      RECT  41870.0 50240.0 42575.0 48895.0 ;
      RECT  41870.0 50240.0 42575.0 51585.0 ;
      RECT  41870.0 52930.0 42575.0 51585.0 ;
      RECT  41870.0 52930.0 42575.0 54275.0 ;
      RECT  41870.0 55620.0 42575.0 54275.0 ;
      RECT  41870.0 55620.0 42575.0 56965.0 ;
      RECT  41870.0 58310.0 42575.0 56965.0 ;
      RECT  41870.0 58310.0 42575.0 59655.0 ;
      RECT  41870.0 61000.0 42575.0 59655.0 ;
      RECT  41870.0 61000.0 42575.0 62345.0 ;
      RECT  41870.0 63690.0 42575.0 62345.0 ;
      RECT  41870.0 63690.0 42575.0 65035.0 ;
      RECT  41870.0 66380.0 42575.0 65035.0 ;
      RECT  41870.0 66380.0 42575.0 67725.0 ;
      RECT  41870.0 69070.0 42575.0 67725.0 ;
      RECT  41870.0 69070.0 42575.0 70415.0 ;
      RECT  41870.0 71760.0 42575.0 70415.0 ;
      RECT  41870.0 71760.0 42575.0 73105.0 ;
      RECT  41870.0 74450.0 42575.0 73105.0 ;
      RECT  41870.0 74450.0 42575.0 75795.0 ;
      RECT  41870.0 77140.0 42575.0 75795.0 ;
      RECT  41870.0 77140.0 42575.0 78485.0 ;
      RECT  41870.0 79830.0 42575.0 78485.0 ;
      RECT  41870.0 79830.0 42575.0 81175.0 ;
      RECT  41870.0 82520.0 42575.0 81175.0 ;
      RECT  41870.0 82520.0 42575.0 83865.0 ;
      RECT  41870.0 85210.0 42575.0 83865.0 ;
      RECT  41870.0 85210.0 42575.0 86555.0 ;
      RECT  41870.0 87900.0 42575.0 86555.0 ;
      RECT  41870.0 87900.0 42575.0 89245.0 ;
      RECT  41870.0 90590.0 42575.0 89245.0 ;
      RECT  41870.0 90590.0 42575.0 91935.0 ;
      RECT  41870.0 93280.0 42575.0 91935.0 ;
      RECT  41870.0 93280.0 42575.0 94625.0 ;
      RECT  41870.0 95970.0 42575.0 94625.0 ;
      RECT  41870.0 95970.0 42575.0 97315.0 ;
      RECT  41870.0 98660.0 42575.0 97315.0 ;
      RECT  41870.0 98660.0 42575.0 100005.0 ;
      RECT  41870.0 101350.0 42575.0 100005.0 ;
      RECT  41870.0 101350.0 42575.0 102695.0 ;
      RECT  41870.0 104040.0 42575.0 102695.0 ;
      RECT  41870.0 104040.0 42575.0 105385.0 ;
      RECT  41870.0 106730.0 42575.0 105385.0 ;
      RECT  41870.0 106730.0 42575.0 108075.0 ;
      RECT  41870.0 109420.0 42575.0 108075.0 ;
      RECT  41870.0 109420.0 42575.0 110765.0 ;
      RECT  41870.0 112110.0 42575.0 110765.0 ;
      RECT  41870.0 112110.0 42575.0 113455.0 ;
      RECT  41870.0 114800.0 42575.0 113455.0 ;
      RECT  41870.0 114800.0 42575.0 116145.0 ;
      RECT  41870.0 117490.0 42575.0 116145.0 ;
      RECT  41870.0 117490.0 42575.0 118835.0 ;
      RECT  41870.0 120180.0 42575.0 118835.0 ;
      RECT  41870.0 120180.0 42575.0 121525.0 ;
      RECT  41870.0 122870.0 42575.0 121525.0 ;
      RECT  41870.0 122870.0 42575.0 124215.0 ;
      RECT  41870.0 125560.0 42575.0 124215.0 ;
      RECT  41870.0 125560.0 42575.0 126905.0 ;
      RECT  41870.0 128250.0 42575.0 126905.0 ;
      RECT  41870.0 128250.0 42575.0 129595.0 ;
      RECT  41870.0 130940.0 42575.0 129595.0 ;
      RECT  41870.0 130940.0 42575.0 132285.0 ;
      RECT  41870.0 133630.0 42575.0 132285.0 ;
      RECT  41870.0 133630.0 42575.0 134975.0 ;
      RECT  41870.0 136320.0 42575.0 134975.0 ;
      RECT  41870.0 136320.0 42575.0 137665.0 ;
      RECT  41870.0 139010.0 42575.0 137665.0 ;
      RECT  41870.0 139010.0 42575.0 140355.0 ;
      RECT  41870.0 141700.0 42575.0 140355.0 ;
      RECT  41870.0 141700.0 42575.0 143045.0 ;
      RECT  41870.0 144390.0 42575.0 143045.0 ;
      RECT  41870.0 144390.0 42575.0 145735.0 ;
      RECT  41870.0 147080.0 42575.0 145735.0 ;
      RECT  41870.0 147080.0 42575.0 148425.0 ;
      RECT  41870.0 149770.0 42575.0 148425.0 ;
      RECT  41870.0 149770.0 42575.0 151115.0 ;
      RECT  41870.0 152460.0 42575.0 151115.0 ;
      RECT  41870.0 152460.0 42575.0 153805.0 ;
      RECT  41870.0 155150.0 42575.0 153805.0 ;
      RECT  41870.0 155150.0 42575.0 156495.0 ;
      RECT  41870.0 157840.0 42575.0 156495.0 ;
      RECT  41870.0 157840.0 42575.0 159185.0 ;
      RECT  41870.0 160530.0 42575.0 159185.0 ;
      RECT  41870.0 160530.0 42575.0 161875.0 ;
      RECT  41870.0 163220.0 42575.0 161875.0 ;
      RECT  41870.0 163220.0 42575.0 164565.0 ;
      RECT  41870.0 165910.0 42575.0 164565.0 ;
      RECT  41870.0 165910.0 42575.0 167255.0 ;
      RECT  41870.0 168600.0 42575.0 167255.0 ;
      RECT  41870.0 168600.0 42575.0 169945.0 ;
      RECT  41870.0 171290.0 42575.0 169945.0 ;
      RECT  41870.0 171290.0 42575.0 172635.0 ;
      RECT  41870.0 173980.0 42575.0 172635.0 ;
      RECT  41870.0 173980.0 42575.0 175325.0 ;
      RECT  41870.0 176670.0 42575.0 175325.0 ;
      RECT  41870.0 176670.0 42575.0 178015.0 ;
      RECT  41870.0 179360.0 42575.0 178015.0 ;
      RECT  41870.0 179360.0 42575.0 180705.0 ;
      RECT  41870.0 182050.0 42575.0 180705.0 ;
      RECT  41870.0 182050.0 42575.0 183395.0 ;
      RECT  41870.0 184740.0 42575.0 183395.0 ;
      RECT  41870.0 184740.0 42575.0 186085.0 ;
      RECT  41870.0 187430.0 42575.0 186085.0 ;
      RECT  41870.0 187430.0 42575.0 188775.0 ;
      RECT  41870.0 190120.0 42575.0 188775.0 ;
      RECT  41870.0 190120.0 42575.0 191465.0 ;
      RECT  41870.0 192810.0 42575.0 191465.0 ;
      RECT  41870.0 192810.0 42575.0 194155.0 ;
      RECT  41870.0 195500.0 42575.0 194155.0 ;
      RECT  41870.0 195500.0 42575.0 196845.0 ;
      RECT  41870.0 198190.0 42575.0 196845.0 ;
      RECT  41870.0 198190.0 42575.0 199535.0 ;
      RECT  41870.0 200880.0 42575.0 199535.0 ;
      RECT  41870.0 200880.0 42575.0 202225.0 ;
      RECT  41870.0 203570.0 42575.0 202225.0 ;
      RECT  41870.0 203570.0 42575.0 204915.0 ;
      RECT  41870.0 206260.0 42575.0 204915.0 ;
      RECT  42575.0 34100.0 43280.0 35445.0 ;
      RECT  42575.0 36790.0 43280.0 35445.0 ;
      RECT  42575.0 36790.0 43280.0 38135.0 ;
      RECT  42575.0 39480.0 43280.0 38135.0 ;
      RECT  42575.0 39480.0 43280.0 40825.0 ;
      RECT  42575.0 42170.0 43280.0 40825.0 ;
      RECT  42575.0 42170.0 43280.0 43515.0 ;
      RECT  42575.0 44860.0 43280.0 43515.0 ;
      RECT  42575.0 44860.0 43280.0 46205.0 ;
      RECT  42575.0 47550.0 43280.0 46205.0 ;
      RECT  42575.0 47550.0 43280.0 48895.0 ;
      RECT  42575.0 50240.0 43280.0 48895.0 ;
      RECT  42575.0 50240.0 43280.0 51585.0 ;
      RECT  42575.0 52930.0 43280.0 51585.0 ;
      RECT  42575.0 52930.0 43280.0 54275.0 ;
      RECT  42575.0 55620.0 43280.0 54275.0 ;
      RECT  42575.0 55620.0 43280.0 56965.0 ;
      RECT  42575.0 58310.0 43280.0 56965.0 ;
      RECT  42575.0 58310.0 43280.0 59655.0 ;
      RECT  42575.0 61000.0 43280.0 59655.0 ;
      RECT  42575.0 61000.0 43280.0 62345.0 ;
      RECT  42575.0 63690.0 43280.0 62345.0 ;
      RECT  42575.0 63690.0 43280.0 65035.0 ;
      RECT  42575.0 66380.0 43280.0 65035.0 ;
      RECT  42575.0 66380.0 43280.0 67725.0 ;
      RECT  42575.0 69070.0 43280.0 67725.0 ;
      RECT  42575.0 69070.0 43280.0 70415.0 ;
      RECT  42575.0 71760.0 43280.0 70415.0 ;
      RECT  42575.0 71760.0 43280.0 73105.0 ;
      RECT  42575.0 74450.0 43280.0 73105.0 ;
      RECT  42575.0 74450.0 43280.0 75795.0 ;
      RECT  42575.0 77140.0 43280.0 75795.0 ;
      RECT  42575.0 77140.0 43280.0 78485.0 ;
      RECT  42575.0 79830.0 43280.0 78485.0 ;
      RECT  42575.0 79830.0 43280.0 81175.0 ;
      RECT  42575.0 82520.0 43280.0 81175.0 ;
      RECT  42575.0 82520.0 43280.0 83865.0 ;
      RECT  42575.0 85210.0 43280.0 83865.0 ;
      RECT  42575.0 85210.0 43280.0 86555.0 ;
      RECT  42575.0 87900.0 43280.0 86555.0 ;
      RECT  42575.0 87900.0 43280.0 89245.0 ;
      RECT  42575.0 90590.0 43280.0 89245.0 ;
      RECT  42575.0 90590.0 43280.0 91935.0 ;
      RECT  42575.0 93280.0 43280.0 91935.0 ;
      RECT  42575.0 93280.0 43280.0 94625.0 ;
      RECT  42575.0 95970.0 43280.0 94625.0 ;
      RECT  42575.0 95970.0 43280.0 97315.0 ;
      RECT  42575.0 98660.0 43280.0 97315.0 ;
      RECT  42575.0 98660.0 43280.0 100005.0 ;
      RECT  42575.0 101350.0 43280.0 100005.0 ;
      RECT  42575.0 101350.0 43280.0 102695.0 ;
      RECT  42575.0 104040.0 43280.0 102695.0 ;
      RECT  42575.0 104040.0 43280.0 105385.0 ;
      RECT  42575.0 106730.0 43280.0 105385.0 ;
      RECT  42575.0 106730.0 43280.0 108075.0 ;
      RECT  42575.0 109420.0 43280.0 108075.0 ;
      RECT  42575.0 109420.0 43280.0 110765.0 ;
      RECT  42575.0 112110.0 43280.0 110765.0 ;
      RECT  42575.0 112110.0 43280.0 113455.0 ;
      RECT  42575.0 114800.0 43280.0 113455.0 ;
      RECT  42575.0 114800.0 43280.0 116145.0 ;
      RECT  42575.0 117490.0 43280.0 116145.0 ;
      RECT  42575.0 117490.0 43280.0 118835.0 ;
      RECT  42575.0 120180.0 43280.0 118835.0 ;
      RECT  42575.0 120180.0 43280.0 121525.0 ;
      RECT  42575.0 122870.0 43280.0 121525.0 ;
      RECT  42575.0 122870.0 43280.0 124215.0 ;
      RECT  42575.0 125560.0 43280.0 124215.0 ;
      RECT  42575.0 125560.0 43280.0 126905.0 ;
      RECT  42575.0 128250.0 43280.0 126905.0 ;
      RECT  42575.0 128250.0 43280.0 129595.0 ;
      RECT  42575.0 130940.0 43280.0 129595.0 ;
      RECT  42575.0 130940.0 43280.0 132285.0 ;
      RECT  42575.0 133630.0 43280.0 132285.0 ;
      RECT  42575.0 133630.0 43280.0 134975.0 ;
      RECT  42575.0 136320.0 43280.0 134975.0 ;
      RECT  42575.0 136320.0 43280.0 137665.0 ;
      RECT  42575.0 139010.0 43280.0 137665.0 ;
      RECT  42575.0 139010.0 43280.0 140355.0 ;
      RECT  42575.0 141700.0 43280.0 140355.0 ;
      RECT  42575.0 141700.0 43280.0 143045.0 ;
      RECT  42575.0 144390.0 43280.0 143045.0 ;
      RECT  42575.0 144390.0 43280.0 145735.0 ;
      RECT  42575.0 147080.0 43280.0 145735.0 ;
      RECT  42575.0 147080.0 43280.0 148425.0 ;
      RECT  42575.0 149770.0 43280.0 148425.0 ;
      RECT  42575.0 149770.0 43280.0 151115.0 ;
      RECT  42575.0 152460.0 43280.0 151115.0 ;
      RECT  42575.0 152460.0 43280.0 153805.0 ;
      RECT  42575.0 155150.0 43280.0 153805.0 ;
      RECT  42575.0 155150.0 43280.0 156495.0 ;
      RECT  42575.0 157840.0 43280.0 156495.0 ;
      RECT  42575.0 157840.0 43280.0 159185.0 ;
      RECT  42575.0 160530.0 43280.0 159185.0 ;
      RECT  42575.0 160530.0 43280.0 161875.0 ;
      RECT  42575.0 163220.0 43280.0 161875.0 ;
      RECT  42575.0 163220.0 43280.0 164565.0 ;
      RECT  42575.0 165910.0 43280.0 164565.0 ;
      RECT  42575.0 165910.0 43280.0 167255.0 ;
      RECT  42575.0 168600.0 43280.0 167255.0 ;
      RECT  42575.0 168600.0 43280.0 169945.0 ;
      RECT  42575.0 171290.0 43280.0 169945.0 ;
      RECT  42575.0 171290.0 43280.0 172635.0 ;
      RECT  42575.0 173980.0 43280.0 172635.0 ;
      RECT  42575.0 173980.0 43280.0 175325.0 ;
      RECT  42575.0 176670.0 43280.0 175325.0 ;
      RECT  42575.0 176670.0 43280.0 178015.0 ;
      RECT  42575.0 179360.0 43280.0 178015.0 ;
      RECT  42575.0 179360.0 43280.0 180705.0 ;
      RECT  42575.0 182050.0 43280.0 180705.0 ;
      RECT  42575.0 182050.0 43280.0 183395.0 ;
      RECT  42575.0 184740.0 43280.0 183395.0 ;
      RECT  42575.0 184740.0 43280.0 186085.0 ;
      RECT  42575.0 187430.0 43280.0 186085.0 ;
      RECT  42575.0 187430.0 43280.0 188775.0 ;
      RECT  42575.0 190120.0 43280.0 188775.0 ;
      RECT  42575.0 190120.0 43280.0 191465.0 ;
      RECT  42575.0 192810.0 43280.0 191465.0 ;
      RECT  42575.0 192810.0 43280.0 194155.0 ;
      RECT  42575.0 195500.0 43280.0 194155.0 ;
      RECT  42575.0 195500.0 43280.0 196845.0 ;
      RECT  42575.0 198190.0 43280.0 196845.0 ;
      RECT  42575.0 198190.0 43280.0 199535.0 ;
      RECT  42575.0 200880.0 43280.0 199535.0 ;
      RECT  42575.0 200880.0 43280.0 202225.0 ;
      RECT  42575.0 203570.0 43280.0 202225.0 ;
      RECT  42575.0 203570.0 43280.0 204915.0 ;
      RECT  42575.0 206260.0 43280.0 204915.0 ;
      RECT  43280.0 34100.0 43985.0 35445.0 ;
      RECT  43280.0 36790.0 43985.0 35445.0 ;
      RECT  43280.0 36790.0 43985.0 38135.0 ;
      RECT  43280.0 39480.0 43985.0 38135.0 ;
      RECT  43280.0 39480.0 43985.0 40825.0 ;
      RECT  43280.0 42170.0 43985.0 40825.0 ;
      RECT  43280.0 42170.0 43985.0 43515.0 ;
      RECT  43280.0 44860.0 43985.0 43515.0 ;
      RECT  43280.0 44860.0 43985.0 46205.0 ;
      RECT  43280.0 47550.0 43985.0 46205.0 ;
      RECT  43280.0 47550.0 43985.0 48895.0 ;
      RECT  43280.0 50240.0 43985.0 48895.0 ;
      RECT  43280.0 50240.0 43985.0 51585.0 ;
      RECT  43280.0 52930.0 43985.0 51585.0 ;
      RECT  43280.0 52930.0 43985.0 54275.0 ;
      RECT  43280.0 55620.0 43985.0 54275.0 ;
      RECT  43280.0 55620.0 43985.0 56965.0 ;
      RECT  43280.0 58310.0 43985.0 56965.0 ;
      RECT  43280.0 58310.0 43985.0 59655.0 ;
      RECT  43280.0 61000.0 43985.0 59655.0 ;
      RECT  43280.0 61000.0 43985.0 62345.0 ;
      RECT  43280.0 63690.0 43985.0 62345.0 ;
      RECT  43280.0 63690.0 43985.0 65035.0 ;
      RECT  43280.0 66380.0 43985.0 65035.0 ;
      RECT  43280.0 66380.0 43985.0 67725.0 ;
      RECT  43280.0 69070.0 43985.0 67725.0 ;
      RECT  43280.0 69070.0 43985.0 70415.0 ;
      RECT  43280.0 71760.0 43985.0 70415.0 ;
      RECT  43280.0 71760.0 43985.0 73105.0 ;
      RECT  43280.0 74450.0 43985.0 73105.0 ;
      RECT  43280.0 74450.0 43985.0 75795.0 ;
      RECT  43280.0 77140.0 43985.0 75795.0 ;
      RECT  43280.0 77140.0 43985.0 78485.0 ;
      RECT  43280.0 79830.0 43985.0 78485.0 ;
      RECT  43280.0 79830.0 43985.0 81175.0 ;
      RECT  43280.0 82520.0 43985.0 81175.0 ;
      RECT  43280.0 82520.0 43985.0 83865.0 ;
      RECT  43280.0 85210.0 43985.0 83865.0 ;
      RECT  43280.0 85210.0 43985.0 86555.0 ;
      RECT  43280.0 87900.0 43985.0 86555.0 ;
      RECT  43280.0 87900.0 43985.0 89245.0 ;
      RECT  43280.0 90590.0 43985.0 89245.0 ;
      RECT  43280.0 90590.0 43985.0 91935.0 ;
      RECT  43280.0 93280.0 43985.0 91935.0 ;
      RECT  43280.0 93280.0 43985.0 94625.0 ;
      RECT  43280.0 95970.0 43985.0 94625.0 ;
      RECT  43280.0 95970.0 43985.0 97315.0 ;
      RECT  43280.0 98660.0 43985.0 97315.0 ;
      RECT  43280.0 98660.0 43985.0 100005.0 ;
      RECT  43280.0 101350.0 43985.0 100005.0 ;
      RECT  43280.0 101350.0 43985.0 102695.0 ;
      RECT  43280.0 104040.0 43985.0 102695.0 ;
      RECT  43280.0 104040.0 43985.0 105385.0 ;
      RECT  43280.0 106730.0 43985.0 105385.0 ;
      RECT  43280.0 106730.0 43985.0 108075.0 ;
      RECT  43280.0 109420.0 43985.0 108075.0 ;
      RECT  43280.0 109420.0 43985.0 110765.0 ;
      RECT  43280.0 112110.0 43985.0 110765.0 ;
      RECT  43280.0 112110.0 43985.0 113455.0 ;
      RECT  43280.0 114800.0 43985.0 113455.0 ;
      RECT  43280.0 114800.0 43985.0 116145.0 ;
      RECT  43280.0 117490.0 43985.0 116145.0 ;
      RECT  43280.0 117490.0 43985.0 118835.0 ;
      RECT  43280.0 120180.0 43985.0 118835.0 ;
      RECT  43280.0 120180.0 43985.0 121525.0 ;
      RECT  43280.0 122870.0 43985.0 121525.0 ;
      RECT  43280.0 122870.0 43985.0 124215.0 ;
      RECT  43280.0 125560.0 43985.0 124215.0 ;
      RECT  43280.0 125560.0 43985.0 126905.0 ;
      RECT  43280.0 128250.0 43985.0 126905.0 ;
      RECT  43280.0 128250.0 43985.0 129595.0 ;
      RECT  43280.0 130940.0 43985.0 129595.0 ;
      RECT  43280.0 130940.0 43985.0 132285.0 ;
      RECT  43280.0 133630.0 43985.0 132285.0 ;
      RECT  43280.0 133630.0 43985.0 134975.0 ;
      RECT  43280.0 136320.0 43985.0 134975.0 ;
      RECT  43280.0 136320.0 43985.0 137665.0 ;
      RECT  43280.0 139010.0 43985.0 137665.0 ;
      RECT  43280.0 139010.0 43985.0 140355.0 ;
      RECT  43280.0 141700.0 43985.0 140355.0 ;
      RECT  43280.0 141700.0 43985.0 143045.0 ;
      RECT  43280.0 144390.0 43985.0 143045.0 ;
      RECT  43280.0 144390.0 43985.0 145735.0 ;
      RECT  43280.0 147080.0 43985.0 145735.0 ;
      RECT  43280.0 147080.0 43985.0 148425.0 ;
      RECT  43280.0 149770.0 43985.0 148425.0 ;
      RECT  43280.0 149770.0 43985.0 151115.0 ;
      RECT  43280.0 152460.0 43985.0 151115.0 ;
      RECT  43280.0 152460.0 43985.0 153805.0 ;
      RECT  43280.0 155150.0 43985.0 153805.0 ;
      RECT  43280.0 155150.0 43985.0 156495.0 ;
      RECT  43280.0 157840.0 43985.0 156495.0 ;
      RECT  43280.0 157840.0 43985.0 159185.0 ;
      RECT  43280.0 160530.0 43985.0 159185.0 ;
      RECT  43280.0 160530.0 43985.0 161875.0 ;
      RECT  43280.0 163220.0 43985.0 161875.0 ;
      RECT  43280.0 163220.0 43985.0 164565.0 ;
      RECT  43280.0 165910.0 43985.0 164565.0 ;
      RECT  43280.0 165910.0 43985.0 167255.0 ;
      RECT  43280.0 168600.0 43985.0 167255.0 ;
      RECT  43280.0 168600.0 43985.0 169945.0 ;
      RECT  43280.0 171290.0 43985.0 169945.0 ;
      RECT  43280.0 171290.0 43985.0 172635.0 ;
      RECT  43280.0 173980.0 43985.0 172635.0 ;
      RECT  43280.0 173980.0 43985.0 175325.0 ;
      RECT  43280.0 176670.0 43985.0 175325.0 ;
      RECT  43280.0 176670.0 43985.0 178015.0 ;
      RECT  43280.0 179360.0 43985.0 178015.0 ;
      RECT  43280.0 179360.0 43985.0 180705.0 ;
      RECT  43280.0 182050.0 43985.0 180705.0 ;
      RECT  43280.0 182050.0 43985.0 183395.0 ;
      RECT  43280.0 184740.0 43985.0 183395.0 ;
      RECT  43280.0 184740.0 43985.0 186085.0 ;
      RECT  43280.0 187430.0 43985.0 186085.0 ;
      RECT  43280.0 187430.0 43985.0 188775.0 ;
      RECT  43280.0 190120.0 43985.0 188775.0 ;
      RECT  43280.0 190120.0 43985.0 191465.0 ;
      RECT  43280.0 192810.0 43985.0 191465.0 ;
      RECT  43280.0 192810.0 43985.0 194155.0 ;
      RECT  43280.0 195500.0 43985.0 194155.0 ;
      RECT  43280.0 195500.0 43985.0 196845.0 ;
      RECT  43280.0 198190.0 43985.0 196845.0 ;
      RECT  43280.0 198190.0 43985.0 199535.0 ;
      RECT  43280.0 200880.0 43985.0 199535.0 ;
      RECT  43280.0 200880.0 43985.0 202225.0 ;
      RECT  43280.0 203570.0 43985.0 202225.0 ;
      RECT  43280.0 203570.0 43985.0 204915.0 ;
      RECT  43280.0 206260.0 43985.0 204915.0 ;
      RECT  43985.0 34100.0 44690.0 35445.0 ;
      RECT  43985.0 36790.0 44690.0 35445.0 ;
      RECT  43985.0 36790.0 44690.0 38135.0 ;
      RECT  43985.0 39480.0 44690.0 38135.0 ;
      RECT  43985.0 39480.0 44690.0 40825.0 ;
      RECT  43985.0 42170.0 44690.0 40825.0 ;
      RECT  43985.0 42170.0 44690.0 43515.0 ;
      RECT  43985.0 44860.0 44690.0 43515.0 ;
      RECT  43985.0 44860.0 44690.0 46205.0 ;
      RECT  43985.0 47550.0 44690.0 46205.0 ;
      RECT  43985.0 47550.0 44690.0 48895.0 ;
      RECT  43985.0 50240.0 44690.0 48895.0 ;
      RECT  43985.0 50240.0 44690.0 51585.0 ;
      RECT  43985.0 52930.0 44690.0 51585.0 ;
      RECT  43985.0 52930.0 44690.0 54275.0 ;
      RECT  43985.0 55620.0 44690.0 54275.0 ;
      RECT  43985.0 55620.0 44690.0 56965.0 ;
      RECT  43985.0 58310.0 44690.0 56965.0 ;
      RECT  43985.0 58310.0 44690.0 59655.0 ;
      RECT  43985.0 61000.0 44690.0 59655.0 ;
      RECT  43985.0 61000.0 44690.0 62345.0 ;
      RECT  43985.0 63690.0 44690.0 62345.0 ;
      RECT  43985.0 63690.0 44690.0 65035.0 ;
      RECT  43985.0 66380.0 44690.0 65035.0 ;
      RECT  43985.0 66380.0 44690.0 67725.0 ;
      RECT  43985.0 69070.0 44690.0 67725.0 ;
      RECT  43985.0 69070.0 44690.0 70415.0 ;
      RECT  43985.0 71760.0 44690.0 70415.0 ;
      RECT  43985.0 71760.0 44690.0 73105.0 ;
      RECT  43985.0 74450.0 44690.0 73105.0 ;
      RECT  43985.0 74450.0 44690.0 75795.0 ;
      RECT  43985.0 77140.0 44690.0 75795.0 ;
      RECT  43985.0 77140.0 44690.0 78485.0 ;
      RECT  43985.0 79830.0 44690.0 78485.0 ;
      RECT  43985.0 79830.0 44690.0 81175.0 ;
      RECT  43985.0 82520.0 44690.0 81175.0 ;
      RECT  43985.0 82520.0 44690.0 83865.0 ;
      RECT  43985.0 85210.0 44690.0 83865.0 ;
      RECT  43985.0 85210.0 44690.0 86555.0 ;
      RECT  43985.0 87900.0 44690.0 86555.0 ;
      RECT  43985.0 87900.0 44690.0 89245.0 ;
      RECT  43985.0 90590.0 44690.0 89245.0 ;
      RECT  43985.0 90590.0 44690.0 91935.0 ;
      RECT  43985.0 93280.0 44690.0 91935.0 ;
      RECT  43985.0 93280.0 44690.0 94625.0 ;
      RECT  43985.0 95970.0 44690.0 94625.0 ;
      RECT  43985.0 95970.0 44690.0 97315.0 ;
      RECT  43985.0 98660.0 44690.0 97315.0 ;
      RECT  43985.0 98660.0 44690.0 100005.0 ;
      RECT  43985.0 101350.0 44690.0 100005.0 ;
      RECT  43985.0 101350.0 44690.0 102695.0 ;
      RECT  43985.0 104040.0 44690.0 102695.0 ;
      RECT  43985.0 104040.0 44690.0 105385.0 ;
      RECT  43985.0 106730.0 44690.0 105385.0 ;
      RECT  43985.0 106730.0 44690.0 108075.0 ;
      RECT  43985.0 109420.0 44690.0 108075.0 ;
      RECT  43985.0 109420.0 44690.0 110765.0 ;
      RECT  43985.0 112110.0 44690.0 110765.0 ;
      RECT  43985.0 112110.0 44690.0 113455.0 ;
      RECT  43985.0 114800.0 44690.0 113455.0 ;
      RECT  43985.0 114800.0 44690.0 116145.0 ;
      RECT  43985.0 117490.0 44690.0 116145.0 ;
      RECT  43985.0 117490.0 44690.0 118835.0 ;
      RECT  43985.0 120180.0 44690.0 118835.0 ;
      RECT  43985.0 120180.0 44690.0 121525.0 ;
      RECT  43985.0 122870.0 44690.0 121525.0 ;
      RECT  43985.0 122870.0 44690.0 124215.0 ;
      RECT  43985.0 125560.0 44690.0 124215.0 ;
      RECT  43985.0 125560.0 44690.0 126905.0 ;
      RECT  43985.0 128250.0 44690.0 126905.0 ;
      RECT  43985.0 128250.0 44690.0 129595.0 ;
      RECT  43985.0 130940.0 44690.0 129595.0 ;
      RECT  43985.0 130940.0 44690.0 132285.0 ;
      RECT  43985.0 133630.0 44690.0 132285.0 ;
      RECT  43985.0 133630.0 44690.0 134975.0 ;
      RECT  43985.0 136320.0 44690.0 134975.0 ;
      RECT  43985.0 136320.0 44690.0 137665.0 ;
      RECT  43985.0 139010.0 44690.0 137665.0 ;
      RECT  43985.0 139010.0 44690.0 140355.0 ;
      RECT  43985.0 141700.0 44690.0 140355.0 ;
      RECT  43985.0 141700.0 44690.0 143045.0 ;
      RECT  43985.0 144390.0 44690.0 143045.0 ;
      RECT  43985.0 144390.0 44690.0 145735.0 ;
      RECT  43985.0 147080.0 44690.0 145735.0 ;
      RECT  43985.0 147080.0 44690.0 148425.0 ;
      RECT  43985.0 149770.0 44690.0 148425.0 ;
      RECT  43985.0 149770.0 44690.0 151115.0 ;
      RECT  43985.0 152460.0 44690.0 151115.0 ;
      RECT  43985.0 152460.0 44690.0 153805.0 ;
      RECT  43985.0 155150.0 44690.0 153805.0 ;
      RECT  43985.0 155150.0 44690.0 156495.0 ;
      RECT  43985.0 157840.0 44690.0 156495.0 ;
      RECT  43985.0 157840.0 44690.0 159185.0 ;
      RECT  43985.0 160530.0 44690.0 159185.0 ;
      RECT  43985.0 160530.0 44690.0 161875.0 ;
      RECT  43985.0 163220.0 44690.0 161875.0 ;
      RECT  43985.0 163220.0 44690.0 164565.0 ;
      RECT  43985.0 165910.0 44690.0 164565.0 ;
      RECT  43985.0 165910.0 44690.0 167255.0 ;
      RECT  43985.0 168600.0 44690.0 167255.0 ;
      RECT  43985.0 168600.0 44690.0 169945.0 ;
      RECT  43985.0 171290.0 44690.0 169945.0 ;
      RECT  43985.0 171290.0 44690.0 172635.0 ;
      RECT  43985.0 173980.0 44690.0 172635.0 ;
      RECT  43985.0 173980.0 44690.0 175325.0 ;
      RECT  43985.0 176670.0 44690.0 175325.0 ;
      RECT  43985.0 176670.0 44690.0 178015.0 ;
      RECT  43985.0 179360.0 44690.0 178015.0 ;
      RECT  43985.0 179360.0 44690.0 180705.0 ;
      RECT  43985.0 182050.0 44690.0 180705.0 ;
      RECT  43985.0 182050.0 44690.0 183395.0 ;
      RECT  43985.0 184740.0 44690.0 183395.0 ;
      RECT  43985.0 184740.0 44690.0 186085.0 ;
      RECT  43985.0 187430.0 44690.0 186085.0 ;
      RECT  43985.0 187430.0 44690.0 188775.0 ;
      RECT  43985.0 190120.0 44690.0 188775.0 ;
      RECT  43985.0 190120.0 44690.0 191465.0 ;
      RECT  43985.0 192810.0 44690.0 191465.0 ;
      RECT  43985.0 192810.0 44690.0 194155.0 ;
      RECT  43985.0 195500.0 44690.0 194155.0 ;
      RECT  43985.0 195500.0 44690.0 196845.0 ;
      RECT  43985.0 198190.0 44690.0 196845.0 ;
      RECT  43985.0 198190.0 44690.0 199535.0 ;
      RECT  43985.0 200880.0 44690.0 199535.0 ;
      RECT  43985.0 200880.0 44690.0 202225.0 ;
      RECT  43985.0 203570.0 44690.0 202225.0 ;
      RECT  43985.0 203570.0 44690.0 204915.0 ;
      RECT  43985.0 206260.0 44690.0 204915.0 ;
      RECT  44690.0 34100.0 45395.0 35445.0 ;
      RECT  44690.0 36790.0 45395.0 35445.0 ;
      RECT  44690.0 36790.0 45395.0 38135.0 ;
      RECT  44690.0 39480.0 45395.0 38135.0 ;
      RECT  44690.0 39480.0 45395.0 40825.0 ;
      RECT  44690.0 42170.0 45395.0 40825.0 ;
      RECT  44690.0 42170.0 45395.0 43515.0 ;
      RECT  44690.0 44860.0 45395.0 43515.0 ;
      RECT  44690.0 44860.0 45395.0 46205.0 ;
      RECT  44690.0 47550.0 45395.0 46205.0 ;
      RECT  44690.0 47550.0 45395.0 48895.0 ;
      RECT  44690.0 50240.0 45395.0 48895.0 ;
      RECT  44690.0 50240.0 45395.0 51585.0 ;
      RECT  44690.0 52930.0 45395.0 51585.0 ;
      RECT  44690.0 52930.0 45395.0 54275.0 ;
      RECT  44690.0 55620.0 45395.0 54275.0 ;
      RECT  44690.0 55620.0 45395.0 56965.0 ;
      RECT  44690.0 58310.0 45395.0 56965.0 ;
      RECT  44690.0 58310.0 45395.0 59655.0 ;
      RECT  44690.0 61000.0 45395.0 59655.0 ;
      RECT  44690.0 61000.0 45395.0 62345.0 ;
      RECT  44690.0 63690.0 45395.0 62345.0 ;
      RECT  44690.0 63690.0 45395.0 65035.0 ;
      RECT  44690.0 66380.0 45395.0 65035.0 ;
      RECT  44690.0 66380.0 45395.0 67725.0 ;
      RECT  44690.0 69070.0 45395.0 67725.0 ;
      RECT  44690.0 69070.0 45395.0 70415.0 ;
      RECT  44690.0 71760.0 45395.0 70415.0 ;
      RECT  44690.0 71760.0 45395.0 73105.0 ;
      RECT  44690.0 74450.0 45395.0 73105.0 ;
      RECT  44690.0 74450.0 45395.0 75795.0 ;
      RECT  44690.0 77140.0 45395.0 75795.0 ;
      RECT  44690.0 77140.0 45395.0 78485.0 ;
      RECT  44690.0 79830.0 45395.0 78485.0 ;
      RECT  44690.0 79830.0 45395.0 81175.0 ;
      RECT  44690.0 82520.0 45395.0 81175.0 ;
      RECT  44690.0 82520.0 45395.0 83865.0 ;
      RECT  44690.0 85210.0 45395.0 83865.0 ;
      RECT  44690.0 85210.0 45395.0 86555.0 ;
      RECT  44690.0 87900.0 45395.0 86555.0 ;
      RECT  44690.0 87900.0 45395.0 89245.0 ;
      RECT  44690.0 90590.0 45395.0 89245.0 ;
      RECT  44690.0 90590.0 45395.0 91935.0 ;
      RECT  44690.0 93280.0 45395.0 91935.0 ;
      RECT  44690.0 93280.0 45395.0 94625.0 ;
      RECT  44690.0 95970.0 45395.0 94625.0 ;
      RECT  44690.0 95970.0 45395.0 97315.0 ;
      RECT  44690.0 98660.0 45395.0 97315.0 ;
      RECT  44690.0 98660.0 45395.0 100005.0 ;
      RECT  44690.0 101350.0 45395.0 100005.0 ;
      RECT  44690.0 101350.0 45395.0 102695.0 ;
      RECT  44690.0 104040.0 45395.0 102695.0 ;
      RECT  44690.0 104040.0 45395.0 105385.0 ;
      RECT  44690.0 106730.0 45395.0 105385.0 ;
      RECT  44690.0 106730.0 45395.0 108075.0 ;
      RECT  44690.0 109420.0 45395.0 108075.0 ;
      RECT  44690.0 109420.0 45395.0 110765.0 ;
      RECT  44690.0 112110.0 45395.0 110765.0 ;
      RECT  44690.0 112110.0 45395.0 113455.0 ;
      RECT  44690.0 114800.0 45395.0 113455.0 ;
      RECT  44690.0 114800.0 45395.0 116145.0 ;
      RECT  44690.0 117490.0 45395.0 116145.0 ;
      RECT  44690.0 117490.0 45395.0 118835.0 ;
      RECT  44690.0 120180.0 45395.0 118835.0 ;
      RECT  44690.0 120180.0 45395.0 121525.0 ;
      RECT  44690.0 122870.0 45395.0 121525.0 ;
      RECT  44690.0 122870.0 45395.0 124215.0 ;
      RECT  44690.0 125560.0 45395.0 124215.0 ;
      RECT  44690.0 125560.0 45395.0 126905.0 ;
      RECT  44690.0 128250.0 45395.0 126905.0 ;
      RECT  44690.0 128250.0 45395.0 129595.0 ;
      RECT  44690.0 130940.0 45395.0 129595.0 ;
      RECT  44690.0 130940.0 45395.0 132285.0 ;
      RECT  44690.0 133630.0 45395.0 132285.0 ;
      RECT  44690.0 133630.0 45395.0 134975.0 ;
      RECT  44690.0 136320.0 45395.0 134975.0 ;
      RECT  44690.0 136320.0 45395.0 137665.0 ;
      RECT  44690.0 139010.0 45395.0 137665.0 ;
      RECT  44690.0 139010.0 45395.0 140355.0 ;
      RECT  44690.0 141700.0 45395.0 140355.0 ;
      RECT  44690.0 141700.0 45395.0 143045.0 ;
      RECT  44690.0 144390.0 45395.0 143045.0 ;
      RECT  44690.0 144390.0 45395.0 145735.0 ;
      RECT  44690.0 147080.0 45395.0 145735.0 ;
      RECT  44690.0 147080.0 45395.0 148425.0 ;
      RECT  44690.0 149770.0 45395.0 148425.0 ;
      RECT  44690.0 149770.0 45395.0 151115.0 ;
      RECT  44690.0 152460.0 45395.0 151115.0 ;
      RECT  44690.0 152460.0 45395.0 153805.0 ;
      RECT  44690.0 155150.0 45395.0 153805.0 ;
      RECT  44690.0 155150.0 45395.0 156495.0 ;
      RECT  44690.0 157840.0 45395.0 156495.0 ;
      RECT  44690.0 157840.0 45395.0 159185.0 ;
      RECT  44690.0 160530.0 45395.0 159185.0 ;
      RECT  44690.0 160530.0 45395.0 161875.0 ;
      RECT  44690.0 163220.0 45395.0 161875.0 ;
      RECT  44690.0 163220.0 45395.0 164565.0 ;
      RECT  44690.0 165910.0 45395.0 164565.0 ;
      RECT  44690.0 165910.0 45395.0 167255.0 ;
      RECT  44690.0 168600.0 45395.0 167255.0 ;
      RECT  44690.0 168600.0 45395.0 169945.0 ;
      RECT  44690.0 171290.0 45395.0 169945.0 ;
      RECT  44690.0 171290.0 45395.0 172635.0 ;
      RECT  44690.0 173980.0 45395.0 172635.0 ;
      RECT  44690.0 173980.0 45395.0 175325.0 ;
      RECT  44690.0 176670.0 45395.0 175325.0 ;
      RECT  44690.0 176670.0 45395.0 178015.0 ;
      RECT  44690.0 179360.0 45395.0 178015.0 ;
      RECT  44690.0 179360.0 45395.0 180705.0 ;
      RECT  44690.0 182050.0 45395.0 180705.0 ;
      RECT  44690.0 182050.0 45395.0 183395.0 ;
      RECT  44690.0 184740.0 45395.0 183395.0 ;
      RECT  44690.0 184740.0 45395.0 186085.0 ;
      RECT  44690.0 187430.0 45395.0 186085.0 ;
      RECT  44690.0 187430.0 45395.0 188775.0 ;
      RECT  44690.0 190120.0 45395.0 188775.0 ;
      RECT  44690.0 190120.0 45395.0 191465.0 ;
      RECT  44690.0 192810.0 45395.0 191465.0 ;
      RECT  44690.0 192810.0 45395.0 194155.0 ;
      RECT  44690.0 195500.0 45395.0 194155.0 ;
      RECT  44690.0 195500.0 45395.0 196845.0 ;
      RECT  44690.0 198190.0 45395.0 196845.0 ;
      RECT  44690.0 198190.0 45395.0 199535.0 ;
      RECT  44690.0 200880.0 45395.0 199535.0 ;
      RECT  44690.0 200880.0 45395.0 202225.0 ;
      RECT  44690.0 203570.0 45395.0 202225.0 ;
      RECT  44690.0 203570.0 45395.0 204915.0 ;
      RECT  44690.0 206260.0 45395.0 204915.0 ;
      RECT  45395.0 34100.0 46100.0 35445.0 ;
      RECT  45395.0 36790.0 46100.0 35445.0 ;
      RECT  45395.0 36790.0 46100.0 38135.0 ;
      RECT  45395.0 39480.0 46100.0 38135.0 ;
      RECT  45395.0 39480.0 46100.0 40825.0 ;
      RECT  45395.0 42170.0 46100.0 40825.0 ;
      RECT  45395.0 42170.0 46100.0 43515.0 ;
      RECT  45395.0 44860.0 46100.0 43515.0 ;
      RECT  45395.0 44860.0 46100.0 46205.0 ;
      RECT  45395.0 47550.0 46100.0 46205.0 ;
      RECT  45395.0 47550.0 46100.0 48895.0 ;
      RECT  45395.0 50240.0 46100.0 48895.0 ;
      RECT  45395.0 50240.0 46100.0 51585.0 ;
      RECT  45395.0 52930.0 46100.0 51585.0 ;
      RECT  45395.0 52930.0 46100.0 54275.0 ;
      RECT  45395.0 55620.0 46100.0 54275.0 ;
      RECT  45395.0 55620.0 46100.0 56965.0 ;
      RECT  45395.0 58310.0 46100.0 56965.0 ;
      RECT  45395.0 58310.0 46100.0 59655.0 ;
      RECT  45395.0 61000.0 46100.0 59655.0 ;
      RECT  45395.0 61000.0 46100.0 62345.0 ;
      RECT  45395.0 63690.0 46100.0 62345.0 ;
      RECT  45395.0 63690.0 46100.0 65035.0 ;
      RECT  45395.0 66380.0 46100.0 65035.0 ;
      RECT  45395.0 66380.0 46100.0 67725.0 ;
      RECT  45395.0 69070.0 46100.0 67725.0 ;
      RECT  45395.0 69070.0 46100.0 70415.0 ;
      RECT  45395.0 71760.0 46100.0 70415.0 ;
      RECT  45395.0 71760.0 46100.0 73105.0 ;
      RECT  45395.0 74450.0 46100.0 73105.0 ;
      RECT  45395.0 74450.0 46100.0 75795.0 ;
      RECT  45395.0 77140.0 46100.0 75795.0 ;
      RECT  45395.0 77140.0 46100.0 78485.0 ;
      RECT  45395.0 79830.0 46100.0 78485.0 ;
      RECT  45395.0 79830.0 46100.0 81175.0 ;
      RECT  45395.0 82520.0 46100.0 81175.0 ;
      RECT  45395.0 82520.0 46100.0 83865.0 ;
      RECT  45395.0 85210.0 46100.0 83865.0 ;
      RECT  45395.0 85210.0 46100.0 86555.0 ;
      RECT  45395.0 87900.0 46100.0 86555.0 ;
      RECT  45395.0 87900.0 46100.0 89245.0 ;
      RECT  45395.0 90590.0 46100.0 89245.0 ;
      RECT  45395.0 90590.0 46100.0 91935.0 ;
      RECT  45395.0 93280.0 46100.0 91935.0 ;
      RECT  45395.0 93280.0 46100.0 94625.0 ;
      RECT  45395.0 95970.0 46100.0 94625.0 ;
      RECT  45395.0 95970.0 46100.0 97315.0 ;
      RECT  45395.0 98660.0 46100.0 97315.0 ;
      RECT  45395.0 98660.0 46100.0 100005.0 ;
      RECT  45395.0 101350.0 46100.0 100005.0 ;
      RECT  45395.0 101350.0 46100.0 102695.0 ;
      RECT  45395.0 104040.0 46100.0 102695.0 ;
      RECT  45395.0 104040.0 46100.0 105385.0 ;
      RECT  45395.0 106730.0 46100.0 105385.0 ;
      RECT  45395.0 106730.0 46100.0 108075.0 ;
      RECT  45395.0 109420.0 46100.0 108075.0 ;
      RECT  45395.0 109420.0 46100.0 110765.0 ;
      RECT  45395.0 112110.0 46100.0 110765.0 ;
      RECT  45395.0 112110.0 46100.0 113455.0 ;
      RECT  45395.0 114800.0 46100.0 113455.0 ;
      RECT  45395.0 114800.0 46100.0 116145.0 ;
      RECT  45395.0 117490.0 46100.0 116145.0 ;
      RECT  45395.0 117490.0 46100.0 118835.0 ;
      RECT  45395.0 120180.0 46100.0 118835.0 ;
      RECT  45395.0 120180.0 46100.0 121525.0 ;
      RECT  45395.0 122870.0 46100.0 121525.0 ;
      RECT  45395.0 122870.0 46100.0 124215.0 ;
      RECT  45395.0 125560.0 46100.0 124215.0 ;
      RECT  45395.0 125560.0 46100.0 126905.0 ;
      RECT  45395.0 128250.0 46100.0 126905.0 ;
      RECT  45395.0 128250.0 46100.0 129595.0 ;
      RECT  45395.0 130940.0 46100.0 129595.0 ;
      RECT  45395.0 130940.0 46100.0 132285.0 ;
      RECT  45395.0 133630.0 46100.0 132285.0 ;
      RECT  45395.0 133630.0 46100.0 134975.0 ;
      RECT  45395.0 136320.0 46100.0 134975.0 ;
      RECT  45395.0 136320.0 46100.0 137665.0 ;
      RECT  45395.0 139010.0 46100.0 137665.0 ;
      RECT  45395.0 139010.0 46100.0 140355.0 ;
      RECT  45395.0 141700.0 46100.0 140355.0 ;
      RECT  45395.0 141700.0 46100.0 143045.0 ;
      RECT  45395.0 144390.0 46100.0 143045.0 ;
      RECT  45395.0 144390.0 46100.0 145735.0 ;
      RECT  45395.0 147080.0 46100.0 145735.0 ;
      RECT  45395.0 147080.0 46100.0 148425.0 ;
      RECT  45395.0 149770.0 46100.0 148425.0 ;
      RECT  45395.0 149770.0 46100.0 151115.0 ;
      RECT  45395.0 152460.0 46100.0 151115.0 ;
      RECT  45395.0 152460.0 46100.0 153805.0 ;
      RECT  45395.0 155150.0 46100.0 153805.0 ;
      RECT  45395.0 155150.0 46100.0 156495.0 ;
      RECT  45395.0 157840.0 46100.0 156495.0 ;
      RECT  45395.0 157840.0 46100.0 159185.0 ;
      RECT  45395.0 160530.0 46100.0 159185.0 ;
      RECT  45395.0 160530.0 46100.0 161875.0 ;
      RECT  45395.0 163220.0 46100.0 161875.0 ;
      RECT  45395.0 163220.0 46100.0 164565.0 ;
      RECT  45395.0 165910.0 46100.0 164565.0 ;
      RECT  45395.0 165910.0 46100.0 167255.0 ;
      RECT  45395.0 168600.0 46100.0 167255.0 ;
      RECT  45395.0 168600.0 46100.0 169945.0 ;
      RECT  45395.0 171290.0 46100.0 169945.0 ;
      RECT  45395.0 171290.0 46100.0 172635.0 ;
      RECT  45395.0 173980.0 46100.0 172635.0 ;
      RECT  45395.0 173980.0 46100.0 175325.0 ;
      RECT  45395.0 176670.0 46100.0 175325.0 ;
      RECT  45395.0 176670.0 46100.0 178015.0 ;
      RECT  45395.0 179360.0 46100.0 178015.0 ;
      RECT  45395.0 179360.0 46100.0 180705.0 ;
      RECT  45395.0 182050.0 46100.0 180705.0 ;
      RECT  45395.0 182050.0 46100.0 183395.0 ;
      RECT  45395.0 184740.0 46100.0 183395.0 ;
      RECT  45395.0 184740.0 46100.0 186085.0 ;
      RECT  45395.0 187430.0 46100.0 186085.0 ;
      RECT  45395.0 187430.0 46100.0 188775.0 ;
      RECT  45395.0 190120.0 46100.0 188775.0 ;
      RECT  45395.0 190120.0 46100.0 191465.0 ;
      RECT  45395.0 192810.0 46100.0 191465.0 ;
      RECT  45395.0 192810.0 46100.0 194155.0 ;
      RECT  45395.0 195500.0 46100.0 194155.0 ;
      RECT  45395.0 195500.0 46100.0 196845.0 ;
      RECT  45395.0 198190.0 46100.0 196845.0 ;
      RECT  45395.0 198190.0 46100.0 199535.0 ;
      RECT  45395.0 200880.0 46100.0 199535.0 ;
      RECT  45395.0 200880.0 46100.0 202225.0 ;
      RECT  45395.0 203570.0 46100.0 202225.0 ;
      RECT  45395.0 203570.0 46100.0 204915.0 ;
      RECT  45395.0 206260.0 46100.0 204915.0 ;
      RECT  46100.0 34100.0 46805.0 35445.0 ;
      RECT  46100.0 36790.0 46805.0 35445.0 ;
      RECT  46100.0 36790.0 46805.0 38135.0 ;
      RECT  46100.0 39480.0 46805.0 38135.0 ;
      RECT  46100.0 39480.0 46805.0 40825.0 ;
      RECT  46100.0 42170.0 46805.0 40825.0 ;
      RECT  46100.0 42170.0 46805.0 43515.0 ;
      RECT  46100.0 44860.0 46805.0 43515.0 ;
      RECT  46100.0 44860.0 46805.0 46205.0 ;
      RECT  46100.0 47550.0 46805.0 46205.0 ;
      RECT  46100.0 47550.0 46805.0 48895.0 ;
      RECT  46100.0 50240.0 46805.0 48895.0 ;
      RECT  46100.0 50240.0 46805.0 51585.0 ;
      RECT  46100.0 52930.0 46805.0 51585.0 ;
      RECT  46100.0 52930.0 46805.0 54275.0 ;
      RECT  46100.0 55620.0 46805.0 54275.0 ;
      RECT  46100.0 55620.0 46805.0 56965.0 ;
      RECT  46100.0 58310.0 46805.0 56965.0 ;
      RECT  46100.0 58310.0 46805.0 59655.0 ;
      RECT  46100.0 61000.0 46805.0 59655.0 ;
      RECT  46100.0 61000.0 46805.0 62345.0 ;
      RECT  46100.0 63690.0 46805.0 62345.0 ;
      RECT  46100.0 63690.0 46805.0 65035.0 ;
      RECT  46100.0 66380.0 46805.0 65035.0 ;
      RECT  46100.0 66380.0 46805.0 67725.0 ;
      RECT  46100.0 69070.0 46805.0 67725.0 ;
      RECT  46100.0 69070.0 46805.0 70415.0 ;
      RECT  46100.0 71760.0 46805.0 70415.0 ;
      RECT  46100.0 71760.0 46805.0 73105.0 ;
      RECT  46100.0 74450.0 46805.0 73105.0 ;
      RECT  46100.0 74450.0 46805.0 75795.0 ;
      RECT  46100.0 77140.0 46805.0 75795.0 ;
      RECT  46100.0 77140.0 46805.0 78485.0 ;
      RECT  46100.0 79830.0 46805.0 78485.0 ;
      RECT  46100.0 79830.0 46805.0 81175.0 ;
      RECT  46100.0 82520.0 46805.0 81175.0 ;
      RECT  46100.0 82520.0 46805.0 83865.0 ;
      RECT  46100.0 85210.0 46805.0 83865.0 ;
      RECT  46100.0 85210.0 46805.0 86555.0 ;
      RECT  46100.0 87900.0 46805.0 86555.0 ;
      RECT  46100.0 87900.0 46805.0 89245.0 ;
      RECT  46100.0 90590.0 46805.0 89245.0 ;
      RECT  46100.0 90590.0 46805.0 91935.0 ;
      RECT  46100.0 93280.0 46805.0 91935.0 ;
      RECT  46100.0 93280.0 46805.0 94625.0 ;
      RECT  46100.0 95970.0 46805.0 94625.0 ;
      RECT  46100.0 95970.0 46805.0 97315.0 ;
      RECT  46100.0 98660.0 46805.0 97315.0 ;
      RECT  46100.0 98660.0 46805.0 100005.0 ;
      RECT  46100.0 101350.0 46805.0 100005.0 ;
      RECT  46100.0 101350.0 46805.0 102695.0 ;
      RECT  46100.0 104040.0 46805.0 102695.0 ;
      RECT  46100.0 104040.0 46805.0 105385.0 ;
      RECT  46100.0 106730.0 46805.0 105385.0 ;
      RECT  46100.0 106730.0 46805.0 108075.0 ;
      RECT  46100.0 109420.0 46805.0 108075.0 ;
      RECT  46100.0 109420.0 46805.0 110765.0 ;
      RECT  46100.0 112110.0 46805.0 110765.0 ;
      RECT  46100.0 112110.0 46805.0 113455.0 ;
      RECT  46100.0 114800.0 46805.0 113455.0 ;
      RECT  46100.0 114800.0 46805.0 116145.0 ;
      RECT  46100.0 117490.0 46805.0 116145.0 ;
      RECT  46100.0 117490.0 46805.0 118835.0 ;
      RECT  46100.0 120180.0 46805.0 118835.0 ;
      RECT  46100.0 120180.0 46805.0 121525.0 ;
      RECT  46100.0 122870.0 46805.0 121525.0 ;
      RECT  46100.0 122870.0 46805.0 124215.0 ;
      RECT  46100.0 125560.0 46805.0 124215.0 ;
      RECT  46100.0 125560.0 46805.0 126905.0 ;
      RECT  46100.0 128250.0 46805.0 126905.0 ;
      RECT  46100.0 128250.0 46805.0 129595.0 ;
      RECT  46100.0 130940.0 46805.0 129595.0 ;
      RECT  46100.0 130940.0 46805.0 132285.0 ;
      RECT  46100.0 133630.0 46805.0 132285.0 ;
      RECT  46100.0 133630.0 46805.0 134975.0 ;
      RECT  46100.0 136320.0 46805.0 134975.0 ;
      RECT  46100.0 136320.0 46805.0 137665.0 ;
      RECT  46100.0 139010.0 46805.0 137665.0 ;
      RECT  46100.0 139010.0 46805.0 140355.0 ;
      RECT  46100.0 141700.0 46805.0 140355.0 ;
      RECT  46100.0 141700.0 46805.0 143045.0 ;
      RECT  46100.0 144390.0 46805.0 143045.0 ;
      RECT  46100.0 144390.0 46805.0 145735.0 ;
      RECT  46100.0 147080.0 46805.0 145735.0 ;
      RECT  46100.0 147080.0 46805.0 148425.0 ;
      RECT  46100.0 149770.0 46805.0 148425.0 ;
      RECT  46100.0 149770.0 46805.0 151115.0 ;
      RECT  46100.0 152460.0 46805.0 151115.0 ;
      RECT  46100.0 152460.0 46805.0 153805.0 ;
      RECT  46100.0 155150.0 46805.0 153805.0 ;
      RECT  46100.0 155150.0 46805.0 156495.0 ;
      RECT  46100.0 157840.0 46805.0 156495.0 ;
      RECT  46100.0 157840.0 46805.0 159185.0 ;
      RECT  46100.0 160530.0 46805.0 159185.0 ;
      RECT  46100.0 160530.0 46805.0 161875.0 ;
      RECT  46100.0 163220.0 46805.0 161875.0 ;
      RECT  46100.0 163220.0 46805.0 164565.0 ;
      RECT  46100.0 165910.0 46805.0 164565.0 ;
      RECT  46100.0 165910.0 46805.0 167255.0 ;
      RECT  46100.0 168600.0 46805.0 167255.0 ;
      RECT  46100.0 168600.0 46805.0 169945.0 ;
      RECT  46100.0 171290.0 46805.0 169945.0 ;
      RECT  46100.0 171290.0 46805.0 172635.0 ;
      RECT  46100.0 173980.0 46805.0 172635.0 ;
      RECT  46100.0 173980.0 46805.0 175325.0 ;
      RECT  46100.0 176670.0 46805.0 175325.0 ;
      RECT  46100.0 176670.0 46805.0 178015.0 ;
      RECT  46100.0 179360.0 46805.0 178015.0 ;
      RECT  46100.0 179360.0 46805.0 180705.0 ;
      RECT  46100.0 182050.0 46805.0 180705.0 ;
      RECT  46100.0 182050.0 46805.0 183395.0 ;
      RECT  46100.0 184740.0 46805.0 183395.0 ;
      RECT  46100.0 184740.0 46805.0 186085.0 ;
      RECT  46100.0 187430.0 46805.0 186085.0 ;
      RECT  46100.0 187430.0 46805.0 188775.0 ;
      RECT  46100.0 190120.0 46805.0 188775.0 ;
      RECT  46100.0 190120.0 46805.0 191465.0 ;
      RECT  46100.0 192810.0 46805.0 191465.0 ;
      RECT  46100.0 192810.0 46805.0 194155.0 ;
      RECT  46100.0 195500.0 46805.0 194155.0 ;
      RECT  46100.0 195500.0 46805.0 196845.0 ;
      RECT  46100.0 198190.0 46805.0 196845.0 ;
      RECT  46100.0 198190.0 46805.0 199535.0 ;
      RECT  46100.0 200880.0 46805.0 199535.0 ;
      RECT  46100.0 200880.0 46805.0 202225.0 ;
      RECT  46100.0 203570.0 46805.0 202225.0 ;
      RECT  46100.0 203570.0 46805.0 204915.0 ;
      RECT  46100.0 206260.0 46805.0 204915.0 ;
      RECT  46805.0 34100.0 47510.0 35445.0 ;
      RECT  46805.0 36790.0 47510.0 35445.0 ;
      RECT  46805.0 36790.0 47510.0 38135.0 ;
      RECT  46805.0 39480.0 47510.0 38135.0 ;
      RECT  46805.0 39480.0 47510.0 40825.0 ;
      RECT  46805.0 42170.0 47510.0 40825.0 ;
      RECT  46805.0 42170.0 47510.0 43515.0 ;
      RECT  46805.0 44860.0 47510.0 43515.0 ;
      RECT  46805.0 44860.0 47510.0 46205.0 ;
      RECT  46805.0 47550.0 47510.0 46205.0 ;
      RECT  46805.0 47550.0 47510.0 48895.0 ;
      RECT  46805.0 50240.0 47510.0 48895.0 ;
      RECT  46805.0 50240.0 47510.0 51585.0 ;
      RECT  46805.0 52930.0 47510.0 51585.0 ;
      RECT  46805.0 52930.0 47510.0 54275.0 ;
      RECT  46805.0 55620.0 47510.0 54275.0 ;
      RECT  46805.0 55620.0 47510.0 56965.0 ;
      RECT  46805.0 58310.0 47510.0 56965.0 ;
      RECT  46805.0 58310.0 47510.0 59655.0 ;
      RECT  46805.0 61000.0 47510.0 59655.0 ;
      RECT  46805.0 61000.0 47510.0 62345.0 ;
      RECT  46805.0 63690.0 47510.0 62345.0 ;
      RECT  46805.0 63690.0 47510.0 65035.0 ;
      RECT  46805.0 66380.0 47510.0 65035.0 ;
      RECT  46805.0 66380.0 47510.0 67725.0 ;
      RECT  46805.0 69070.0 47510.0 67725.0 ;
      RECT  46805.0 69070.0 47510.0 70415.0 ;
      RECT  46805.0 71760.0 47510.0 70415.0 ;
      RECT  46805.0 71760.0 47510.0 73105.0 ;
      RECT  46805.0 74450.0 47510.0 73105.0 ;
      RECT  46805.0 74450.0 47510.0 75795.0 ;
      RECT  46805.0 77140.0 47510.0 75795.0 ;
      RECT  46805.0 77140.0 47510.0 78485.0 ;
      RECT  46805.0 79830.0 47510.0 78485.0 ;
      RECT  46805.0 79830.0 47510.0 81175.0 ;
      RECT  46805.0 82520.0 47510.0 81175.0 ;
      RECT  46805.0 82520.0 47510.0 83865.0 ;
      RECT  46805.0 85210.0 47510.0 83865.0 ;
      RECT  46805.0 85210.0 47510.0 86555.0 ;
      RECT  46805.0 87900.0 47510.0 86555.0 ;
      RECT  46805.0 87900.0 47510.0 89245.0 ;
      RECT  46805.0 90590.0 47510.0 89245.0 ;
      RECT  46805.0 90590.0 47510.0 91935.0 ;
      RECT  46805.0 93280.0 47510.0 91935.0 ;
      RECT  46805.0 93280.0 47510.0 94625.0 ;
      RECT  46805.0 95970.0 47510.0 94625.0 ;
      RECT  46805.0 95970.0 47510.0 97315.0 ;
      RECT  46805.0 98660.0 47510.0 97315.0 ;
      RECT  46805.0 98660.0 47510.0 100005.0 ;
      RECT  46805.0 101350.0 47510.0 100005.0 ;
      RECT  46805.0 101350.0 47510.0 102695.0 ;
      RECT  46805.0 104040.0 47510.0 102695.0 ;
      RECT  46805.0 104040.0 47510.0 105385.0 ;
      RECT  46805.0 106730.0 47510.0 105385.0 ;
      RECT  46805.0 106730.0 47510.0 108075.0 ;
      RECT  46805.0 109420.0 47510.0 108075.0 ;
      RECT  46805.0 109420.0 47510.0 110765.0 ;
      RECT  46805.0 112110.0 47510.0 110765.0 ;
      RECT  46805.0 112110.0 47510.0 113455.0 ;
      RECT  46805.0 114800.0 47510.0 113455.0 ;
      RECT  46805.0 114800.0 47510.0 116145.0 ;
      RECT  46805.0 117490.0 47510.0 116145.0 ;
      RECT  46805.0 117490.0 47510.0 118835.0 ;
      RECT  46805.0 120180.0 47510.0 118835.0 ;
      RECT  46805.0 120180.0 47510.0 121525.0 ;
      RECT  46805.0 122870.0 47510.0 121525.0 ;
      RECT  46805.0 122870.0 47510.0 124215.0 ;
      RECT  46805.0 125560.0 47510.0 124215.0 ;
      RECT  46805.0 125560.0 47510.0 126905.0 ;
      RECT  46805.0 128250.0 47510.0 126905.0 ;
      RECT  46805.0 128250.0 47510.0 129595.0 ;
      RECT  46805.0 130940.0 47510.0 129595.0 ;
      RECT  46805.0 130940.0 47510.0 132285.0 ;
      RECT  46805.0 133630.0 47510.0 132285.0 ;
      RECT  46805.0 133630.0 47510.0 134975.0 ;
      RECT  46805.0 136320.0 47510.0 134975.0 ;
      RECT  46805.0 136320.0 47510.0 137665.0 ;
      RECT  46805.0 139010.0 47510.0 137665.0 ;
      RECT  46805.0 139010.0 47510.0 140355.0 ;
      RECT  46805.0 141700.0 47510.0 140355.0 ;
      RECT  46805.0 141700.0 47510.0 143045.0 ;
      RECT  46805.0 144390.0 47510.0 143045.0 ;
      RECT  46805.0 144390.0 47510.0 145735.0 ;
      RECT  46805.0 147080.0 47510.0 145735.0 ;
      RECT  46805.0 147080.0 47510.0 148425.0 ;
      RECT  46805.0 149770.0 47510.0 148425.0 ;
      RECT  46805.0 149770.0 47510.0 151115.0 ;
      RECT  46805.0 152460.0 47510.0 151115.0 ;
      RECT  46805.0 152460.0 47510.0 153805.0 ;
      RECT  46805.0 155150.0 47510.0 153805.0 ;
      RECT  46805.0 155150.0 47510.0 156495.0 ;
      RECT  46805.0 157840.0 47510.0 156495.0 ;
      RECT  46805.0 157840.0 47510.0 159185.0 ;
      RECT  46805.0 160530.0 47510.0 159185.0 ;
      RECT  46805.0 160530.0 47510.0 161875.0 ;
      RECT  46805.0 163220.0 47510.0 161875.0 ;
      RECT  46805.0 163220.0 47510.0 164565.0 ;
      RECT  46805.0 165910.0 47510.0 164565.0 ;
      RECT  46805.0 165910.0 47510.0 167255.0 ;
      RECT  46805.0 168600.0 47510.0 167255.0 ;
      RECT  46805.0 168600.0 47510.0 169945.0 ;
      RECT  46805.0 171290.0 47510.0 169945.0 ;
      RECT  46805.0 171290.0 47510.0 172635.0 ;
      RECT  46805.0 173980.0 47510.0 172635.0 ;
      RECT  46805.0 173980.0 47510.0 175325.0 ;
      RECT  46805.0 176670.0 47510.0 175325.0 ;
      RECT  46805.0 176670.0 47510.0 178015.0 ;
      RECT  46805.0 179360.0 47510.0 178015.0 ;
      RECT  46805.0 179360.0 47510.0 180705.0 ;
      RECT  46805.0 182050.0 47510.0 180705.0 ;
      RECT  46805.0 182050.0 47510.0 183395.0 ;
      RECT  46805.0 184740.0 47510.0 183395.0 ;
      RECT  46805.0 184740.0 47510.0 186085.0 ;
      RECT  46805.0 187430.0 47510.0 186085.0 ;
      RECT  46805.0 187430.0 47510.0 188775.0 ;
      RECT  46805.0 190120.0 47510.0 188775.0 ;
      RECT  46805.0 190120.0 47510.0 191465.0 ;
      RECT  46805.0 192810.0 47510.0 191465.0 ;
      RECT  46805.0 192810.0 47510.0 194155.0 ;
      RECT  46805.0 195500.0 47510.0 194155.0 ;
      RECT  46805.0 195500.0 47510.0 196845.0 ;
      RECT  46805.0 198190.0 47510.0 196845.0 ;
      RECT  46805.0 198190.0 47510.0 199535.0 ;
      RECT  46805.0 200880.0 47510.0 199535.0 ;
      RECT  46805.0 200880.0 47510.0 202225.0 ;
      RECT  46805.0 203570.0 47510.0 202225.0 ;
      RECT  46805.0 203570.0 47510.0 204915.0 ;
      RECT  46805.0 206260.0 47510.0 204915.0 ;
      RECT  47510.0 34100.0 48215.0 35445.0 ;
      RECT  47510.0 36790.0 48215.0 35445.0 ;
      RECT  47510.0 36790.0 48215.0 38135.0 ;
      RECT  47510.0 39480.0 48215.0 38135.0 ;
      RECT  47510.0 39480.0 48215.0 40825.0 ;
      RECT  47510.0 42170.0 48215.0 40825.0 ;
      RECT  47510.0 42170.0 48215.0 43515.0 ;
      RECT  47510.0 44860.0 48215.0 43515.0 ;
      RECT  47510.0 44860.0 48215.0 46205.0 ;
      RECT  47510.0 47550.0 48215.0 46205.0 ;
      RECT  47510.0 47550.0 48215.0 48895.0 ;
      RECT  47510.0 50240.0 48215.0 48895.0 ;
      RECT  47510.0 50240.0 48215.0 51585.0 ;
      RECT  47510.0 52930.0 48215.0 51585.0 ;
      RECT  47510.0 52930.0 48215.0 54275.0 ;
      RECT  47510.0 55620.0 48215.0 54275.0 ;
      RECT  47510.0 55620.0 48215.0 56965.0 ;
      RECT  47510.0 58310.0 48215.0 56965.0 ;
      RECT  47510.0 58310.0 48215.0 59655.0 ;
      RECT  47510.0 61000.0 48215.0 59655.0 ;
      RECT  47510.0 61000.0 48215.0 62345.0 ;
      RECT  47510.0 63690.0 48215.0 62345.0 ;
      RECT  47510.0 63690.0 48215.0 65035.0 ;
      RECT  47510.0 66380.0 48215.0 65035.0 ;
      RECT  47510.0 66380.0 48215.0 67725.0 ;
      RECT  47510.0 69070.0 48215.0 67725.0 ;
      RECT  47510.0 69070.0 48215.0 70415.0 ;
      RECT  47510.0 71760.0 48215.0 70415.0 ;
      RECT  47510.0 71760.0 48215.0 73105.0 ;
      RECT  47510.0 74450.0 48215.0 73105.0 ;
      RECT  47510.0 74450.0 48215.0 75795.0 ;
      RECT  47510.0 77140.0 48215.0 75795.0 ;
      RECT  47510.0 77140.0 48215.0 78485.0 ;
      RECT  47510.0 79830.0 48215.0 78485.0 ;
      RECT  47510.0 79830.0 48215.0 81175.0 ;
      RECT  47510.0 82520.0 48215.0 81175.0 ;
      RECT  47510.0 82520.0 48215.0 83865.0 ;
      RECT  47510.0 85210.0 48215.0 83865.0 ;
      RECT  47510.0 85210.0 48215.0 86555.0 ;
      RECT  47510.0 87900.0 48215.0 86555.0 ;
      RECT  47510.0 87900.0 48215.0 89245.0 ;
      RECT  47510.0 90590.0 48215.0 89245.0 ;
      RECT  47510.0 90590.0 48215.0 91935.0 ;
      RECT  47510.0 93280.0 48215.0 91935.0 ;
      RECT  47510.0 93280.0 48215.0 94625.0 ;
      RECT  47510.0 95970.0 48215.0 94625.0 ;
      RECT  47510.0 95970.0 48215.0 97315.0 ;
      RECT  47510.0 98660.0 48215.0 97315.0 ;
      RECT  47510.0 98660.0 48215.0 100005.0 ;
      RECT  47510.0 101350.0 48215.0 100005.0 ;
      RECT  47510.0 101350.0 48215.0 102695.0 ;
      RECT  47510.0 104040.0 48215.0 102695.0 ;
      RECT  47510.0 104040.0 48215.0 105385.0 ;
      RECT  47510.0 106730.0 48215.0 105385.0 ;
      RECT  47510.0 106730.0 48215.0 108075.0 ;
      RECT  47510.0 109420.0 48215.0 108075.0 ;
      RECT  47510.0 109420.0 48215.0 110765.0 ;
      RECT  47510.0 112110.0 48215.0 110765.0 ;
      RECT  47510.0 112110.0 48215.0 113455.0 ;
      RECT  47510.0 114800.0 48215.0 113455.0 ;
      RECT  47510.0 114800.0 48215.0 116145.0 ;
      RECT  47510.0 117490.0 48215.0 116145.0 ;
      RECT  47510.0 117490.0 48215.0 118835.0 ;
      RECT  47510.0 120180.0 48215.0 118835.0 ;
      RECT  47510.0 120180.0 48215.0 121525.0 ;
      RECT  47510.0 122870.0 48215.0 121525.0 ;
      RECT  47510.0 122870.0 48215.0 124215.0 ;
      RECT  47510.0 125560.0 48215.0 124215.0 ;
      RECT  47510.0 125560.0 48215.0 126905.0 ;
      RECT  47510.0 128250.0 48215.0 126905.0 ;
      RECT  47510.0 128250.0 48215.0 129595.0 ;
      RECT  47510.0 130940.0 48215.0 129595.0 ;
      RECT  47510.0 130940.0 48215.0 132285.0 ;
      RECT  47510.0 133630.0 48215.0 132285.0 ;
      RECT  47510.0 133630.0 48215.0 134975.0 ;
      RECT  47510.0 136320.0 48215.0 134975.0 ;
      RECT  47510.0 136320.0 48215.0 137665.0 ;
      RECT  47510.0 139010.0 48215.0 137665.0 ;
      RECT  47510.0 139010.0 48215.0 140355.0 ;
      RECT  47510.0 141700.0 48215.0 140355.0 ;
      RECT  47510.0 141700.0 48215.0 143045.0 ;
      RECT  47510.0 144390.0 48215.0 143045.0 ;
      RECT  47510.0 144390.0 48215.0 145735.0 ;
      RECT  47510.0 147080.0 48215.0 145735.0 ;
      RECT  47510.0 147080.0 48215.0 148425.0 ;
      RECT  47510.0 149770.0 48215.0 148425.0 ;
      RECT  47510.0 149770.0 48215.0 151115.0 ;
      RECT  47510.0 152460.0 48215.0 151115.0 ;
      RECT  47510.0 152460.0 48215.0 153805.0 ;
      RECT  47510.0 155150.0 48215.0 153805.0 ;
      RECT  47510.0 155150.0 48215.0 156495.0 ;
      RECT  47510.0 157840.0 48215.0 156495.0 ;
      RECT  47510.0 157840.0 48215.0 159185.0 ;
      RECT  47510.0 160530.0 48215.0 159185.0 ;
      RECT  47510.0 160530.0 48215.0 161875.0 ;
      RECT  47510.0 163220.0 48215.0 161875.0 ;
      RECT  47510.0 163220.0 48215.0 164565.0 ;
      RECT  47510.0 165910.0 48215.0 164565.0 ;
      RECT  47510.0 165910.0 48215.0 167255.0 ;
      RECT  47510.0 168600.0 48215.0 167255.0 ;
      RECT  47510.0 168600.0 48215.0 169945.0 ;
      RECT  47510.0 171290.0 48215.0 169945.0 ;
      RECT  47510.0 171290.0 48215.0 172635.0 ;
      RECT  47510.0 173980.0 48215.0 172635.0 ;
      RECT  47510.0 173980.0 48215.0 175325.0 ;
      RECT  47510.0 176670.0 48215.0 175325.0 ;
      RECT  47510.0 176670.0 48215.0 178015.0 ;
      RECT  47510.0 179360.0 48215.0 178015.0 ;
      RECT  47510.0 179360.0 48215.0 180705.0 ;
      RECT  47510.0 182050.0 48215.0 180705.0 ;
      RECT  47510.0 182050.0 48215.0 183395.0 ;
      RECT  47510.0 184740.0 48215.0 183395.0 ;
      RECT  47510.0 184740.0 48215.0 186085.0 ;
      RECT  47510.0 187430.0 48215.0 186085.0 ;
      RECT  47510.0 187430.0 48215.0 188775.0 ;
      RECT  47510.0 190120.0 48215.0 188775.0 ;
      RECT  47510.0 190120.0 48215.0 191465.0 ;
      RECT  47510.0 192810.0 48215.0 191465.0 ;
      RECT  47510.0 192810.0 48215.0 194155.0 ;
      RECT  47510.0 195500.0 48215.0 194155.0 ;
      RECT  47510.0 195500.0 48215.0 196845.0 ;
      RECT  47510.0 198190.0 48215.0 196845.0 ;
      RECT  47510.0 198190.0 48215.0 199535.0 ;
      RECT  47510.0 200880.0 48215.0 199535.0 ;
      RECT  47510.0 200880.0 48215.0 202225.0 ;
      RECT  47510.0 203570.0 48215.0 202225.0 ;
      RECT  47510.0 203570.0 48215.0 204915.0 ;
      RECT  47510.0 206260.0 48215.0 204915.0 ;
      RECT  48215.0 34100.0 48920.0 35445.0 ;
      RECT  48215.0 36790.0 48920.0 35445.0 ;
      RECT  48215.0 36790.0 48920.0 38135.0 ;
      RECT  48215.0 39480.0 48920.0 38135.0 ;
      RECT  48215.0 39480.0 48920.0 40825.0 ;
      RECT  48215.0 42170.0 48920.0 40825.0 ;
      RECT  48215.0 42170.0 48920.0 43515.0 ;
      RECT  48215.0 44860.0 48920.0 43515.0 ;
      RECT  48215.0 44860.0 48920.0 46205.0 ;
      RECT  48215.0 47550.0 48920.0 46205.0 ;
      RECT  48215.0 47550.0 48920.0 48895.0 ;
      RECT  48215.0 50240.0 48920.0 48895.0 ;
      RECT  48215.0 50240.0 48920.0 51585.0 ;
      RECT  48215.0 52930.0 48920.0 51585.0 ;
      RECT  48215.0 52930.0 48920.0 54275.0 ;
      RECT  48215.0 55620.0 48920.0 54275.0 ;
      RECT  48215.0 55620.0 48920.0 56965.0 ;
      RECT  48215.0 58310.0 48920.0 56965.0 ;
      RECT  48215.0 58310.0 48920.0 59655.0 ;
      RECT  48215.0 61000.0 48920.0 59655.0 ;
      RECT  48215.0 61000.0 48920.0 62345.0 ;
      RECT  48215.0 63690.0 48920.0 62345.0 ;
      RECT  48215.0 63690.0 48920.0 65035.0 ;
      RECT  48215.0 66380.0 48920.0 65035.0 ;
      RECT  48215.0 66380.0 48920.0 67725.0 ;
      RECT  48215.0 69070.0 48920.0 67725.0 ;
      RECT  48215.0 69070.0 48920.0 70415.0 ;
      RECT  48215.0 71760.0 48920.0 70415.0 ;
      RECT  48215.0 71760.0 48920.0 73105.0 ;
      RECT  48215.0 74450.0 48920.0 73105.0 ;
      RECT  48215.0 74450.0 48920.0 75795.0 ;
      RECT  48215.0 77140.0 48920.0 75795.0 ;
      RECT  48215.0 77140.0 48920.0 78485.0 ;
      RECT  48215.0 79830.0 48920.0 78485.0 ;
      RECT  48215.0 79830.0 48920.0 81175.0 ;
      RECT  48215.0 82520.0 48920.0 81175.0 ;
      RECT  48215.0 82520.0 48920.0 83865.0 ;
      RECT  48215.0 85210.0 48920.0 83865.0 ;
      RECT  48215.0 85210.0 48920.0 86555.0 ;
      RECT  48215.0 87900.0 48920.0 86555.0 ;
      RECT  48215.0 87900.0 48920.0 89245.0 ;
      RECT  48215.0 90590.0 48920.0 89245.0 ;
      RECT  48215.0 90590.0 48920.0 91935.0 ;
      RECT  48215.0 93280.0 48920.0 91935.0 ;
      RECT  48215.0 93280.0 48920.0 94625.0 ;
      RECT  48215.0 95970.0 48920.0 94625.0 ;
      RECT  48215.0 95970.0 48920.0 97315.0 ;
      RECT  48215.0 98660.0 48920.0 97315.0 ;
      RECT  48215.0 98660.0 48920.0 100005.0 ;
      RECT  48215.0 101350.0 48920.0 100005.0 ;
      RECT  48215.0 101350.0 48920.0 102695.0 ;
      RECT  48215.0 104040.0 48920.0 102695.0 ;
      RECT  48215.0 104040.0 48920.0 105385.0 ;
      RECT  48215.0 106730.0 48920.0 105385.0 ;
      RECT  48215.0 106730.0 48920.0 108075.0 ;
      RECT  48215.0 109420.0 48920.0 108075.0 ;
      RECT  48215.0 109420.0 48920.0 110765.0 ;
      RECT  48215.0 112110.0 48920.0 110765.0 ;
      RECT  48215.0 112110.0 48920.0 113455.0 ;
      RECT  48215.0 114800.0 48920.0 113455.0 ;
      RECT  48215.0 114800.0 48920.0 116145.0 ;
      RECT  48215.0 117490.0 48920.0 116145.0 ;
      RECT  48215.0 117490.0 48920.0 118835.0 ;
      RECT  48215.0 120180.0 48920.0 118835.0 ;
      RECT  48215.0 120180.0 48920.0 121525.0 ;
      RECT  48215.0 122870.0 48920.0 121525.0 ;
      RECT  48215.0 122870.0 48920.0 124215.0 ;
      RECT  48215.0 125560.0 48920.0 124215.0 ;
      RECT  48215.0 125560.0 48920.0 126905.0 ;
      RECT  48215.0 128250.0 48920.0 126905.0 ;
      RECT  48215.0 128250.0 48920.0 129595.0 ;
      RECT  48215.0 130940.0 48920.0 129595.0 ;
      RECT  48215.0 130940.0 48920.0 132285.0 ;
      RECT  48215.0 133630.0 48920.0 132285.0 ;
      RECT  48215.0 133630.0 48920.0 134975.0 ;
      RECT  48215.0 136320.0 48920.0 134975.0 ;
      RECT  48215.0 136320.0 48920.0 137665.0 ;
      RECT  48215.0 139010.0 48920.0 137665.0 ;
      RECT  48215.0 139010.0 48920.0 140355.0 ;
      RECT  48215.0 141700.0 48920.0 140355.0 ;
      RECT  48215.0 141700.0 48920.0 143045.0 ;
      RECT  48215.0 144390.0 48920.0 143045.0 ;
      RECT  48215.0 144390.0 48920.0 145735.0 ;
      RECT  48215.0 147080.0 48920.0 145735.0 ;
      RECT  48215.0 147080.0 48920.0 148425.0 ;
      RECT  48215.0 149770.0 48920.0 148425.0 ;
      RECT  48215.0 149770.0 48920.0 151115.0 ;
      RECT  48215.0 152460.0 48920.0 151115.0 ;
      RECT  48215.0 152460.0 48920.0 153805.0 ;
      RECT  48215.0 155150.0 48920.0 153805.0 ;
      RECT  48215.0 155150.0 48920.0 156495.0 ;
      RECT  48215.0 157840.0 48920.0 156495.0 ;
      RECT  48215.0 157840.0 48920.0 159185.0 ;
      RECT  48215.0 160530.0 48920.0 159185.0 ;
      RECT  48215.0 160530.0 48920.0 161875.0 ;
      RECT  48215.0 163220.0 48920.0 161875.0 ;
      RECT  48215.0 163220.0 48920.0 164565.0 ;
      RECT  48215.0 165910.0 48920.0 164565.0 ;
      RECT  48215.0 165910.0 48920.0 167255.0 ;
      RECT  48215.0 168600.0 48920.0 167255.0 ;
      RECT  48215.0 168600.0 48920.0 169945.0 ;
      RECT  48215.0 171290.0 48920.0 169945.0 ;
      RECT  48215.0 171290.0 48920.0 172635.0 ;
      RECT  48215.0 173980.0 48920.0 172635.0 ;
      RECT  48215.0 173980.0 48920.0 175325.0 ;
      RECT  48215.0 176670.0 48920.0 175325.0 ;
      RECT  48215.0 176670.0 48920.0 178015.0 ;
      RECT  48215.0 179360.0 48920.0 178015.0 ;
      RECT  48215.0 179360.0 48920.0 180705.0 ;
      RECT  48215.0 182050.0 48920.0 180705.0 ;
      RECT  48215.0 182050.0 48920.0 183395.0 ;
      RECT  48215.0 184740.0 48920.0 183395.0 ;
      RECT  48215.0 184740.0 48920.0 186085.0 ;
      RECT  48215.0 187430.0 48920.0 186085.0 ;
      RECT  48215.0 187430.0 48920.0 188775.0 ;
      RECT  48215.0 190120.0 48920.0 188775.0 ;
      RECT  48215.0 190120.0 48920.0 191465.0 ;
      RECT  48215.0 192810.0 48920.0 191465.0 ;
      RECT  48215.0 192810.0 48920.0 194155.0 ;
      RECT  48215.0 195500.0 48920.0 194155.0 ;
      RECT  48215.0 195500.0 48920.0 196845.0 ;
      RECT  48215.0 198190.0 48920.0 196845.0 ;
      RECT  48215.0 198190.0 48920.0 199535.0 ;
      RECT  48215.0 200880.0 48920.0 199535.0 ;
      RECT  48215.0 200880.0 48920.0 202225.0 ;
      RECT  48215.0 203570.0 48920.0 202225.0 ;
      RECT  48215.0 203570.0 48920.0 204915.0 ;
      RECT  48215.0 206260.0 48920.0 204915.0 ;
      RECT  48920.0 34100.0 49625.0 35445.0 ;
      RECT  48920.0 36790.0 49625.0 35445.0 ;
      RECT  48920.0 36790.0 49625.0 38135.0 ;
      RECT  48920.0 39480.0 49625.0 38135.0 ;
      RECT  48920.0 39480.0 49625.0 40825.0 ;
      RECT  48920.0 42170.0 49625.0 40825.0 ;
      RECT  48920.0 42170.0 49625.0 43515.0 ;
      RECT  48920.0 44860.0 49625.0 43515.0 ;
      RECT  48920.0 44860.0 49625.0 46205.0 ;
      RECT  48920.0 47550.0 49625.0 46205.0 ;
      RECT  48920.0 47550.0 49625.0 48895.0 ;
      RECT  48920.0 50240.0 49625.0 48895.0 ;
      RECT  48920.0 50240.0 49625.0 51585.0 ;
      RECT  48920.0 52930.0 49625.0 51585.0 ;
      RECT  48920.0 52930.0 49625.0 54275.0 ;
      RECT  48920.0 55620.0 49625.0 54275.0 ;
      RECT  48920.0 55620.0 49625.0 56965.0 ;
      RECT  48920.0 58310.0 49625.0 56965.0 ;
      RECT  48920.0 58310.0 49625.0 59655.0 ;
      RECT  48920.0 61000.0 49625.0 59655.0 ;
      RECT  48920.0 61000.0 49625.0 62345.0 ;
      RECT  48920.0 63690.0 49625.0 62345.0 ;
      RECT  48920.0 63690.0 49625.0 65035.0 ;
      RECT  48920.0 66380.0 49625.0 65035.0 ;
      RECT  48920.0 66380.0 49625.0 67725.0 ;
      RECT  48920.0 69070.0 49625.0 67725.0 ;
      RECT  48920.0 69070.0 49625.0 70415.0 ;
      RECT  48920.0 71760.0 49625.0 70415.0 ;
      RECT  48920.0 71760.0 49625.0 73105.0 ;
      RECT  48920.0 74450.0 49625.0 73105.0 ;
      RECT  48920.0 74450.0 49625.0 75795.0 ;
      RECT  48920.0 77140.0 49625.0 75795.0 ;
      RECT  48920.0 77140.0 49625.0 78485.0 ;
      RECT  48920.0 79830.0 49625.0 78485.0 ;
      RECT  48920.0 79830.0 49625.0 81175.0 ;
      RECT  48920.0 82520.0 49625.0 81175.0 ;
      RECT  48920.0 82520.0 49625.0 83865.0 ;
      RECT  48920.0 85210.0 49625.0 83865.0 ;
      RECT  48920.0 85210.0 49625.0 86555.0 ;
      RECT  48920.0 87900.0 49625.0 86555.0 ;
      RECT  48920.0 87900.0 49625.0 89245.0 ;
      RECT  48920.0 90590.0 49625.0 89245.0 ;
      RECT  48920.0 90590.0 49625.0 91935.0 ;
      RECT  48920.0 93280.0 49625.0 91935.0 ;
      RECT  48920.0 93280.0 49625.0 94625.0 ;
      RECT  48920.0 95970.0 49625.0 94625.0 ;
      RECT  48920.0 95970.0 49625.0 97315.0 ;
      RECT  48920.0 98660.0 49625.0 97315.0 ;
      RECT  48920.0 98660.0 49625.0 100005.0 ;
      RECT  48920.0 101350.0 49625.0 100005.0 ;
      RECT  48920.0 101350.0 49625.0 102695.0 ;
      RECT  48920.0 104040.0 49625.0 102695.0 ;
      RECT  48920.0 104040.0 49625.0 105385.0 ;
      RECT  48920.0 106730.0 49625.0 105385.0 ;
      RECT  48920.0 106730.0 49625.0 108075.0 ;
      RECT  48920.0 109420.0 49625.0 108075.0 ;
      RECT  48920.0 109420.0 49625.0 110765.0 ;
      RECT  48920.0 112110.0 49625.0 110765.0 ;
      RECT  48920.0 112110.0 49625.0 113455.0 ;
      RECT  48920.0 114800.0 49625.0 113455.0 ;
      RECT  48920.0 114800.0 49625.0 116145.0 ;
      RECT  48920.0 117490.0 49625.0 116145.0 ;
      RECT  48920.0 117490.0 49625.0 118835.0 ;
      RECT  48920.0 120180.0 49625.0 118835.0 ;
      RECT  48920.0 120180.0 49625.0 121525.0 ;
      RECT  48920.0 122870.0 49625.0 121525.0 ;
      RECT  48920.0 122870.0 49625.0 124215.0 ;
      RECT  48920.0 125560.0 49625.0 124215.0 ;
      RECT  48920.0 125560.0 49625.0 126905.0 ;
      RECT  48920.0 128250.0 49625.0 126905.0 ;
      RECT  48920.0 128250.0 49625.0 129595.0 ;
      RECT  48920.0 130940.0 49625.0 129595.0 ;
      RECT  48920.0 130940.0 49625.0 132285.0 ;
      RECT  48920.0 133630.0 49625.0 132285.0 ;
      RECT  48920.0 133630.0 49625.0 134975.0 ;
      RECT  48920.0 136320.0 49625.0 134975.0 ;
      RECT  48920.0 136320.0 49625.0 137665.0 ;
      RECT  48920.0 139010.0 49625.0 137665.0 ;
      RECT  48920.0 139010.0 49625.0 140355.0 ;
      RECT  48920.0 141700.0 49625.0 140355.0 ;
      RECT  48920.0 141700.0 49625.0 143045.0 ;
      RECT  48920.0 144390.0 49625.0 143045.0 ;
      RECT  48920.0 144390.0 49625.0 145735.0 ;
      RECT  48920.0 147080.0 49625.0 145735.0 ;
      RECT  48920.0 147080.0 49625.0 148425.0 ;
      RECT  48920.0 149770.0 49625.0 148425.0 ;
      RECT  48920.0 149770.0 49625.0 151115.0 ;
      RECT  48920.0 152460.0 49625.0 151115.0 ;
      RECT  48920.0 152460.0 49625.0 153805.0 ;
      RECT  48920.0 155150.0 49625.0 153805.0 ;
      RECT  48920.0 155150.0 49625.0 156495.0 ;
      RECT  48920.0 157840.0 49625.0 156495.0 ;
      RECT  48920.0 157840.0 49625.0 159185.0 ;
      RECT  48920.0 160530.0 49625.0 159185.0 ;
      RECT  48920.0 160530.0 49625.0 161875.0 ;
      RECT  48920.0 163220.0 49625.0 161875.0 ;
      RECT  48920.0 163220.0 49625.0 164565.0 ;
      RECT  48920.0 165910.0 49625.0 164565.0 ;
      RECT  48920.0 165910.0 49625.0 167255.0 ;
      RECT  48920.0 168600.0 49625.0 167255.0 ;
      RECT  48920.0 168600.0 49625.0 169945.0 ;
      RECT  48920.0 171290.0 49625.0 169945.0 ;
      RECT  48920.0 171290.0 49625.0 172635.0 ;
      RECT  48920.0 173980.0 49625.0 172635.0 ;
      RECT  48920.0 173980.0 49625.0 175325.0 ;
      RECT  48920.0 176670.0 49625.0 175325.0 ;
      RECT  48920.0 176670.0 49625.0 178015.0 ;
      RECT  48920.0 179360.0 49625.0 178015.0 ;
      RECT  48920.0 179360.0 49625.0 180705.0 ;
      RECT  48920.0 182050.0 49625.0 180705.0 ;
      RECT  48920.0 182050.0 49625.0 183395.0 ;
      RECT  48920.0 184740.0 49625.0 183395.0 ;
      RECT  48920.0 184740.0 49625.0 186085.0 ;
      RECT  48920.0 187430.0 49625.0 186085.0 ;
      RECT  48920.0 187430.0 49625.0 188775.0 ;
      RECT  48920.0 190120.0 49625.0 188775.0 ;
      RECT  48920.0 190120.0 49625.0 191465.0 ;
      RECT  48920.0 192810.0 49625.0 191465.0 ;
      RECT  48920.0 192810.0 49625.0 194155.0 ;
      RECT  48920.0 195500.0 49625.0 194155.0 ;
      RECT  48920.0 195500.0 49625.0 196845.0 ;
      RECT  48920.0 198190.0 49625.0 196845.0 ;
      RECT  48920.0 198190.0 49625.0 199535.0 ;
      RECT  48920.0 200880.0 49625.0 199535.0 ;
      RECT  48920.0 200880.0 49625.0 202225.0 ;
      RECT  48920.0 203570.0 49625.0 202225.0 ;
      RECT  48920.0 203570.0 49625.0 204915.0 ;
      RECT  48920.0 206260.0 49625.0 204915.0 ;
      RECT  49625.0 34100.0 50330.0 35445.0 ;
      RECT  49625.0 36790.0 50330.0 35445.0 ;
      RECT  49625.0 36790.0 50330.0 38135.0 ;
      RECT  49625.0 39480.0 50330.0 38135.0 ;
      RECT  49625.0 39480.0 50330.0 40825.0 ;
      RECT  49625.0 42170.0 50330.0 40825.0 ;
      RECT  49625.0 42170.0 50330.0 43515.0 ;
      RECT  49625.0 44860.0 50330.0 43515.0 ;
      RECT  49625.0 44860.0 50330.0 46205.0 ;
      RECT  49625.0 47550.0 50330.0 46205.0 ;
      RECT  49625.0 47550.0 50330.0 48895.0 ;
      RECT  49625.0 50240.0 50330.0 48895.0 ;
      RECT  49625.0 50240.0 50330.0 51585.0 ;
      RECT  49625.0 52930.0 50330.0 51585.0 ;
      RECT  49625.0 52930.0 50330.0 54275.0 ;
      RECT  49625.0 55620.0 50330.0 54275.0 ;
      RECT  49625.0 55620.0 50330.0 56965.0 ;
      RECT  49625.0 58310.0 50330.0 56965.0 ;
      RECT  49625.0 58310.0 50330.0 59655.0 ;
      RECT  49625.0 61000.0 50330.0 59655.0 ;
      RECT  49625.0 61000.0 50330.0 62345.0 ;
      RECT  49625.0 63690.0 50330.0 62345.0 ;
      RECT  49625.0 63690.0 50330.0 65035.0 ;
      RECT  49625.0 66380.0 50330.0 65035.0 ;
      RECT  49625.0 66380.0 50330.0 67725.0 ;
      RECT  49625.0 69070.0 50330.0 67725.0 ;
      RECT  49625.0 69070.0 50330.0 70415.0 ;
      RECT  49625.0 71760.0 50330.0 70415.0 ;
      RECT  49625.0 71760.0 50330.0 73105.0 ;
      RECT  49625.0 74450.0 50330.0 73105.0 ;
      RECT  49625.0 74450.0 50330.0 75795.0 ;
      RECT  49625.0 77140.0 50330.0 75795.0 ;
      RECT  49625.0 77140.0 50330.0 78485.0 ;
      RECT  49625.0 79830.0 50330.0 78485.0 ;
      RECT  49625.0 79830.0 50330.0 81175.0 ;
      RECT  49625.0 82520.0 50330.0 81175.0 ;
      RECT  49625.0 82520.0 50330.0 83865.0 ;
      RECT  49625.0 85210.0 50330.0 83865.0 ;
      RECT  49625.0 85210.0 50330.0 86555.0 ;
      RECT  49625.0 87900.0 50330.0 86555.0 ;
      RECT  49625.0 87900.0 50330.0 89245.0 ;
      RECT  49625.0 90590.0 50330.0 89245.0 ;
      RECT  49625.0 90590.0 50330.0 91935.0 ;
      RECT  49625.0 93280.0 50330.0 91935.0 ;
      RECT  49625.0 93280.0 50330.0 94625.0 ;
      RECT  49625.0 95970.0 50330.0 94625.0 ;
      RECT  49625.0 95970.0 50330.0 97315.0 ;
      RECT  49625.0 98660.0 50330.0 97315.0 ;
      RECT  49625.0 98660.0 50330.0 100005.0 ;
      RECT  49625.0 101350.0 50330.0 100005.0 ;
      RECT  49625.0 101350.0 50330.0 102695.0 ;
      RECT  49625.0 104040.0 50330.0 102695.0 ;
      RECT  49625.0 104040.0 50330.0 105385.0 ;
      RECT  49625.0 106730.0 50330.0 105385.0 ;
      RECT  49625.0 106730.0 50330.0 108075.0 ;
      RECT  49625.0 109420.0 50330.0 108075.0 ;
      RECT  49625.0 109420.0 50330.0 110765.0 ;
      RECT  49625.0 112110.0 50330.0 110765.0 ;
      RECT  49625.0 112110.0 50330.0 113455.0 ;
      RECT  49625.0 114800.0 50330.0 113455.0 ;
      RECT  49625.0 114800.0 50330.0 116145.0 ;
      RECT  49625.0 117490.0 50330.0 116145.0 ;
      RECT  49625.0 117490.0 50330.0 118835.0 ;
      RECT  49625.0 120180.0 50330.0 118835.0 ;
      RECT  49625.0 120180.0 50330.0 121525.0 ;
      RECT  49625.0 122870.0 50330.0 121525.0 ;
      RECT  49625.0 122870.0 50330.0 124215.0 ;
      RECT  49625.0 125560.0 50330.0 124215.0 ;
      RECT  49625.0 125560.0 50330.0 126905.0 ;
      RECT  49625.0 128250.0 50330.0 126905.0 ;
      RECT  49625.0 128250.0 50330.0 129595.0 ;
      RECT  49625.0 130940.0 50330.0 129595.0 ;
      RECT  49625.0 130940.0 50330.0 132285.0 ;
      RECT  49625.0 133630.0 50330.0 132285.0 ;
      RECT  49625.0 133630.0 50330.0 134975.0 ;
      RECT  49625.0 136320.0 50330.0 134975.0 ;
      RECT  49625.0 136320.0 50330.0 137665.0 ;
      RECT  49625.0 139010.0 50330.0 137665.0 ;
      RECT  49625.0 139010.0 50330.0 140355.0 ;
      RECT  49625.0 141700.0 50330.0 140355.0 ;
      RECT  49625.0 141700.0 50330.0 143045.0 ;
      RECT  49625.0 144390.0 50330.0 143045.0 ;
      RECT  49625.0 144390.0 50330.0 145735.0 ;
      RECT  49625.0 147080.0 50330.0 145735.0 ;
      RECT  49625.0 147080.0 50330.0 148425.0 ;
      RECT  49625.0 149770.0 50330.0 148425.0 ;
      RECT  49625.0 149770.0 50330.0 151115.0 ;
      RECT  49625.0 152460.0 50330.0 151115.0 ;
      RECT  49625.0 152460.0 50330.0 153805.0 ;
      RECT  49625.0 155150.0 50330.0 153805.0 ;
      RECT  49625.0 155150.0 50330.0 156495.0 ;
      RECT  49625.0 157840.0 50330.0 156495.0 ;
      RECT  49625.0 157840.0 50330.0 159185.0 ;
      RECT  49625.0 160530.0 50330.0 159185.0 ;
      RECT  49625.0 160530.0 50330.0 161875.0 ;
      RECT  49625.0 163220.0 50330.0 161875.0 ;
      RECT  49625.0 163220.0 50330.0 164565.0 ;
      RECT  49625.0 165910.0 50330.0 164565.0 ;
      RECT  49625.0 165910.0 50330.0 167255.0 ;
      RECT  49625.0 168600.0 50330.0 167255.0 ;
      RECT  49625.0 168600.0 50330.0 169945.0 ;
      RECT  49625.0 171290.0 50330.0 169945.0 ;
      RECT  49625.0 171290.0 50330.0 172635.0 ;
      RECT  49625.0 173980.0 50330.0 172635.0 ;
      RECT  49625.0 173980.0 50330.0 175325.0 ;
      RECT  49625.0 176670.0 50330.0 175325.0 ;
      RECT  49625.0 176670.0 50330.0 178015.0 ;
      RECT  49625.0 179360.0 50330.0 178015.0 ;
      RECT  49625.0 179360.0 50330.0 180705.0 ;
      RECT  49625.0 182050.0 50330.0 180705.0 ;
      RECT  49625.0 182050.0 50330.0 183395.0 ;
      RECT  49625.0 184740.0 50330.0 183395.0 ;
      RECT  49625.0 184740.0 50330.0 186085.0 ;
      RECT  49625.0 187430.0 50330.0 186085.0 ;
      RECT  49625.0 187430.0 50330.0 188775.0 ;
      RECT  49625.0 190120.0 50330.0 188775.0 ;
      RECT  49625.0 190120.0 50330.0 191465.0 ;
      RECT  49625.0 192810.0 50330.0 191465.0 ;
      RECT  49625.0 192810.0 50330.0 194155.0 ;
      RECT  49625.0 195500.0 50330.0 194155.0 ;
      RECT  49625.0 195500.0 50330.0 196845.0 ;
      RECT  49625.0 198190.0 50330.0 196845.0 ;
      RECT  49625.0 198190.0 50330.0 199535.0 ;
      RECT  49625.0 200880.0 50330.0 199535.0 ;
      RECT  49625.0 200880.0 50330.0 202225.0 ;
      RECT  49625.0 203570.0 50330.0 202225.0 ;
      RECT  49625.0 203570.0 50330.0 204915.0 ;
      RECT  49625.0 206260.0 50330.0 204915.0 ;
      RECT  50330.0 34100.0 51035.0 35445.0 ;
      RECT  50330.0 36790.0 51035.0 35445.0 ;
      RECT  50330.0 36790.0 51035.0 38135.0 ;
      RECT  50330.0 39480.0 51035.0 38135.0 ;
      RECT  50330.0 39480.0 51035.0 40825.0 ;
      RECT  50330.0 42170.0 51035.0 40825.0 ;
      RECT  50330.0 42170.0 51035.0 43515.0 ;
      RECT  50330.0 44860.0 51035.0 43515.0 ;
      RECT  50330.0 44860.0 51035.0 46205.0 ;
      RECT  50330.0 47550.0 51035.0 46205.0 ;
      RECT  50330.0 47550.0 51035.0 48895.0 ;
      RECT  50330.0 50240.0 51035.0 48895.0 ;
      RECT  50330.0 50240.0 51035.0 51585.0 ;
      RECT  50330.0 52930.0 51035.0 51585.0 ;
      RECT  50330.0 52930.0 51035.0 54275.0 ;
      RECT  50330.0 55620.0 51035.0 54275.0 ;
      RECT  50330.0 55620.0 51035.0 56965.0 ;
      RECT  50330.0 58310.0 51035.0 56965.0 ;
      RECT  50330.0 58310.0 51035.0 59655.0 ;
      RECT  50330.0 61000.0 51035.0 59655.0 ;
      RECT  50330.0 61000.0 51035.0 62345.0 ;
      RECT  50330.0 63690.0 51035.0 62345.0 ;
      RECT  50330.0 63690.0 51035.0 65035.0 ;
      RECT  50330.0 66380.0 51035.0 65035.0 ;
      RECT  50330.0 66380.0 51035.0 67725.0 ;
      RECT  50330.0 69070.0 51035.0 67725.0 ;
      RECT  50330.0 69070.0 51035.0 70415.0 ;
      RECT  50330.0 71760.0 51035.0 70415.0 ;
      RECT  50330.0 71760.0 51035.0 73105.0 ;
      RECT  50330.0 74450.0 51035.0 73105.0 ;
      RECT  50330.0 74450.0 51035.0 75795.0 ;
      RECT  50330.0 77140.0 51035.0 75795.0 ;
      RECT  50330.0 77140.0 51035.0 78485.0 ;
      RECT  50330.0 79830.0 51035.0 78485.0 ;
      RECT  50330.0 79830.0 51035.0 81175.0 ;
      RECT  50330.0 82520.0 51035.0 81175.0 ;
      RECT  50330.0 82520.0 51035.0 83865.0 ;
      RECT  50330.0 85210.0 51035.0 83865.0 ;
      RECT  50330.0 85210.0 51035.0 86555.0 ;
      RECT  50330.0 87900.0 51035.0 86555.0 ;
      RECT  50330.0 87900.0 51035.0 89245.0 ;
      RECT  50330.0 90590.0 51035.0 89245.0 ;
      RECT  50330.0 90590.0 51035.0 91935.0 ;
      RECT  50330.0 93280.0 51035.0 91935.0 ;
      RECT  50330.0 93280.0 51035.0 94625.0 ;
      RECT  50330.0 95970.0 51035.0 94625.0 ;
      RECT  50330.0 95970.0 51035.0 97315.0 ;
      RECT  50330.0 98660.0 51035.0 97315.0 ;
      RECT  50330.0 98660.0 51035.0 100005.0 ;
      RECT  50330.0 101350.0 51035.0 100005.0 ;
      RECT  50330.0 101350.0 51035.0 102695.0 ;
      RECT  50330.0 104040.0 51035.0 102695.0 ;
      RECT  50330.0 104040.0 51035.0 105385.0 ;
      RECT  50330.0 106730.0 51035.0 105385.0 ;
      RECT  50330.0 106730.0 51035.0 108075.0 ;
      RECT  50330.0 109420.0 51035.0 108075.0 ;
      RECT  50330.0 109420.0 51035.0 110765.0 ;
      RECT  50330.0 112110.0 51035.0 110765.0 ;
      RECT  50330.0 112110.0 51035.0 113455.0 ;
      RECT  50330.0 114800.0 51035.0 113455.0 ;
      RECT  50330.0 114800.0 51035.0 116145.0 ;
      RECT  50330.0 117490.0 51035.0 116145.0 ;
      RECT  50330.0 117490.0 51035.0 118835.0 ;
      RECT  50330.0 120180.0 51035.0 118835.0 ;
      RECT  50330.0 120180.0 51035.0 121525.0 ;
      RECT  50330.0 122870.0 51035.0 121525.0 ;
      RECT  50330.0 122870.0 51035.0 124215.0 ;
      RECT  50330.0 125560.0 51035.0 124215.0 ;
      RECT  50330.0 125560.0 51035.0 126905.0 ;
      RECT  50330.0 128250.0 51035.0 126905.0 ;
      RECT  50330.0 128250.0 51035.0 129595.0 ;
      RECT  50330.0 130940.0 51035.0 129595.0 ;
      RECT  50330.0 130940.0 51035.0 132285.0 ;
      RECT  50330.0 133630.0 51035.0 132285.0 ;
      RECT  50330.0 133630.0 51035.0 134975.0 ;
      RECT  50330.0 136320.0 51035.0 134975.0 ;
      RECT  50330.0 136320.0 51035.0 137665.0 ;
      RECT  50330.0 139010.0 51035.0 137665.0 ;
      RECT  50330.0 139010.0 51035.0 140355.0 ;
      RECT  50330.0 141700.0 51035.0 140355.0 ;
      RECT  50330.0 141700.0 51035.0 143045.0 ;
      RECT  50330.0 144390.0 51035.0 143045.0 ;
      RECT  50330.0 144390.0 51035.0 145735.0 ;
      RECT  50330.0 147080.0 51035.0 145735.0 ;
      RECT  50330.0 147080.0 51035.0 148425.0 ;
      RECT  50330.0 149770.0 51035.0 148425.0 ;
      RECT  50330.0 149770.0 51035.0 151115.0 ;
      RECT  50330.0 152460.0 51035.0 151115.0 ;
      RECT  50330.0 152460.0 51035.0 153805.0 ;
      RECT  50330.0 155150.0 51035.0 153805.0 ;
      RECT  50330.0 155150.0 51035.0 156495.0 ;
      RECT  50330.0 157840.0 51035.0 156495.0 ;
      RECT  50330.0 157840.0 51035.0 159185.0 ;
      RECT  50330.0 160530.0 51035.0 159185.0 ;
      RECT  50330.0 160530.0 51035.0 161875.0 ;
      RECT  50330.0 163220.0 51035.0 161875.0 ;
      RECT  50330.0 163220.0 51035.0 164565.0 ;
      RECT  50330.0 165910.0 51035.0 164565.0 ;
      RECT  50330.0 165910.0 51035.0 167255.0 ;
      RECT  50330.0 168600.0 51035.0 167255.0 ;
      RECT  50330.0 168600.0 51035.0 169945.0 ;
      RECT  50330.0 171290.0 51035.0 169945.0 ;
      RECT  50330.0 171290.0 51035.0 172635.0 ;
      RECT  50330.0 173980.0 51035.0 172635.0 ;
      RECT  50330.0 173980.0 51035.0 175325.0 ;
      RECT  50330.0 176670.0 51035.0 175325.0 ;
      RECT  50330.0 176670.0 51035.0 178015.0 ;
      RECT  50330.0 179360.0 51035.0 178015.0 ;
      RECT  50330.0 179360.0 51035.0 180705.0 ;
      RECT  50330.0 182050.0 51035.0 180705.0 ;
      RECT  50330.0 182050.0 51035.0 183395.0 ;
      RECT  50330.0 184740.0 51035.0 183395.0 ;
      RECT  50330.0 184740.0 51035.0 186085.0 ;
      RECT  50330.0 187430.0 51035.0 186085.0 ;
      RECT  50330.0 187430.0 51035.0 188775.0 ;
      RECT  50330.0 190120.0 51035.0 188775.0 ;
      RECT  50330.0 190120.0 51035.0 191465.0 ;
      RECT  50330.0 192810.0 51035.0 191465.0 ;
      RECT  50330.0 192810.0 51035.0 194155.0 ;
      RECT  50330.0 195500.0 51035.0 194155.0 ;
      RECT  50330.0 195500.0 51035.0 196845.0 ;
      RECT  50330.0 198190.0 51035.0 196845.0 ;
      RECT  50330.0 198190.0 51035.0 199535.0 ;
      RECT  50330.0 200880.0 51035.0 199535.0 ;
      RECT  50330.0 200880.0 51035.0 202225.0 ;
      RECT  50330.0 203570.0 51035.0 202225.0 ;
      RECT  50330.0 203570.0 51035.0 204915.0 ;
      RECT  50330.0 206260.0 51035.0 204915.0 ;
      RECT  51035.0 34100.0 51740.0 35445.0 ;
      RECT  51035.0 36790.0 51740.0 35445.0 ;
      RECT  51035.0 36790.0 51740.0 38135.0 ;
      RECT  51035.0 39480.0 51740.0 38135.0 ;
      RECT  51035.0 39480.0 51740.0 40825.0 ;
      RECT  51035.0 42170.0 51740.0 40825.0 ;
      RECT  51035.0 42170.0 51740.0 43515.0 ;
      RECT  51035.0 44860.0 51740.0 43515.0 ;
      RECT  51035.0 44860.0 51740.0 46205.0 ;
      RECT  51035.0 47550.0 51740.0 46205.0 ;
      RECT  51035.0 47550.0 51740.0 48895.0 ;
      RECT  51035.0 50240.0 51740.0 48895.0 ;
      RECT  51035.0 50240.0 51740.0 51585.0 ;
      RECT  51035.0 52930.0 51740.0 51585.0 ;
      RECT  51035.0 52930.0 51740.0 54275.0 ;
      RECT  51035.0 55620.0 51740.0 54275.0 ;
      RECT  51035.0 55620.0 51740.0 56965.0 ;
      RECT  51035.0 58310.0 51740.0 56965.0 ;
      RECT  51035.0 58310.0 51740.0 59655.0 ;
      RECT  51035.0 61000.0 51740.0 59655.0 ;
      RECT  51035.0 61000.0 51740.0 62345.0 ;
      RECT  51035.0 63690.0 51740.0 62345.0 ;
      RECT  51035.0 63690.0 51740.0 65035.0 ;
      RECT  51035.0 66380.0 51740.0 65035.0 ;
      RECT  51035.0 66380.0 51740.0 67725.0 ;
      RECT  51035.0 69070.0 51740.0 67725.0 ;
      RECT  51035.0 69070.0 51740.0 70415.0 ;
      RECT  51035.0 71760.0 51740.0 70415.0 ;
      RECT  51035.0 71760.0 51740.0 73105.0 ;
      RECT  51035.0 74450.0 51740.0 73105.0 ;
      RECT  51035.0 74450.0 51740.0 75795.0 ;
      RECT  51035.0 77140.0 51740.0 75795.0 ;
      RECT  51035.0 77140.0 51740.0 78485.0 ;
      RECT  51035.0 79830.0 51740.0 78485.0 ;
      RECT  51035.0 79830.0 51740.0 81175.0 ;
      RECT  51035.0 82520.0 51740.0 81175.0 ;
      RECT  51035.0 82520.0 51740.0 83865.0 ;
      RECT  51035.0 85210.0 51740.0 83865.0 ;
      RECT  51035.0 85210.0 51740.0 86555.0 ;
      RECT  51035.0 87900.0 51740.0 86555.0 ;
      RECT  51035.0 87900.0 51740.0 89245.0 ;
      RECT  51035.0 90590.0 51740.0 89245.0 ;
      RECT  51035.0 90590.0 51740.0 91935.0 ;
      RECT  51035.0 93280.0 51740.0 91935.0 ;
      RECT  51035.0 93280.0 51740.0 94625.0 ;
      RECT  51035.0 95970.0 51740.0 94625.0 ;
      RECT  51035.0 95970.0 51740.0 97315.0 ;
      RECT  51035.0 98660.0 51740.0 97315.0 ;
      RECT  51035.0 98660.0 51740.0 100005.0 ;
      RECT  51035.0 101350.0 51740.0 100005.0 ;
      RECT  51035.0 101350.0 51740.0 102695.0 ;
      RECT  51035.0 104040.0 51740.0 102695.0 ;
      RECT  51035.0 104040.0 51740.0 105385.0 ;
      RECT  51035.0 106730.0 51740.0 105385.0 ;
      RECT  51035.0 106730.0 51740.0 108075.0 ;
      RECT  51035.0 109420.0 51740.0 108075.0 ;
      RECT  51035.0 109420.0 51740.0 110765.0 ;
      RECT  51035.0 112110.0 51740.0 110765.0 ;
      RECT  51035.0 112110.0 51740.0 113455.0 ;
      RECT  51035.0 114800.0 51740.0 113455.0 ;
      RECT  51035.0 114800.0 51740.0 116145.0 ;
      RECT  51035.0 117490.0 51740.0 116145.0 ;
      RECT  51035.0 117490.0 51740.0 118835.0 ;
      RECT  51035.0 120180.0 51740.0 118835.0 ;
      RECT  51035.0 120180.0 51740.0 121525.0 ;
      RECT  51035.0 122870.0 51740.0 121525.0 ;
      RECT  51035.0 122870.0 51740.0 124215.0 ;
      RECT  51035.0 125560.0 51740.0 124215.0 ;
      RECT  51035.0 125560.0 51740.0 126905.0 ;
      RECT  51035.0 128250.0 51740.0 126905.0 ;
      RECT  51035.0 128250.0 51740.0 129595.0 ;
      RECT  51035.0 130940.0 51740.0 129595.0 ;
      RECT  51035.0 130940.0 51740.0 132285.0 ;
      RECT  51035.0 133630.0 51740.0 132285.0 ;
      RECT  51035.0 133630.0 51740.0 134975.0 ;
      RECT  51035.0 136320.0 51740.0 134975.0 ;
      RECT  51035.0 136320.0 51740.0 137665.0 ;
      RECT  51035.0 139010.0 51740.0 137665.0 ;
      RECT  51035.0 139010.0 51740.0 140355.0 ;
      RECT  51035.0 141700.0 51740.0 140355.0 ;
      RECT  51035.0 141700.0 51740.0 143045.0 ;
      RECT  51035.0 144390.0 51740.0 143045.0 ;
      RECT  51035.0 144390.0 51740.0 145735.0 ;
      RECT  51035.0 147080.0 51740.0 145735.0 ;
      RECT  51035.0 147080.0 51740.0 148425.0 ;
      RECT  51035.0 149770.0 51740.0 148425.0 ;
      RECT  51035.0 149770.0 51740.0 151115.0 ;
      RECT  51035.0 152460.0 51740.0 151115.0 ;
      RECT  51035.0 152460.0 51740.0 153805.0 ;
      RECT  51035.0 155150.0 51740.0 153805.0 ;
      RECT  51035.0 155150.0 51740.0 156495.0 ;
      RECT  51035.0 157840.0 51740.0 156495.0 ;
      RECT  51035.0 157840.0 51740.0 159185.0 ;
      RECT  51035.0 160530.0 51740.0 159185.0 ;
      RECT  51035.0 160530.0 51740.0 161875.0 ;
      RECT  51035.0 163220.0 51740.0 161875.0 ;
      RECT  51035.0 163220.0 51740.0 164565.0 ;
      RECT  51035.0 165910.0 51740.0 164565.0 ;
      RECT  51035.0 165910.0 51740.0 167255.0 ;
      RECT  51035.0 168600.0 51740.0 167255.0 ;
      RECT  51035.0 168600.0 51740.0 169945.0 ;
      RECT  51035.0 171290.0 51740.0 169945.0 ;
      RECT  51035.0 171290.0 51740.0 172635.0 ;
      RECT  51035.0 173980.0 51740.0 172635.0 ;
      RECT  51035.0 173980.0 51740.0 175325.0 ;
      RECT  51035.0 176670.0 51740.0 175325.0 ;
      RECT  51035.0 176670.0 51740.0 178015.0 ;
      RECT  51035.0 179360.0 51740.0 178015.0 ;
      RECT  51035.0 179360.0 51740.0 180705.0 ;
      RECT  51035.0 182050.0 51740.0 180705.0 ;
      RECT  51035.0 182050.0 51740.0 183395.0 ;
      RECT  51035.0 184740.0 51740.0 183395.0 ;
      RECT  51035.0 184740.0 51740.0 186085.0 ;
      RECT  51035.0 187430.0 51740.0 186085.0 ;
      RECT  51035.0 187430.0 51740.0 188775.0 ;
      RECT  51035.0 190120.0 51740.0 188775.0 ;
      RECT  51035.0 190120.0 51740.0 191465.0 ;
      RECT  51035.0 192810.0 51740.0 191465.0 ;
      RECT  51035.0 192810.0 51740.0 194155.0 ;
      RECT  51035.0 195500.0 51740.0 194155.0 ;
      RECT  51035.0 195500.0 51740.0 196845.0 ;
      RECT  51035.0 198190.0 51740.0 196845.0 ;
      RECT  51035.0 198190.0 51740.0 199535.0 ;
      RECT  51035.0 200880.0 51740.0 199535.0 ;
      RECT  51035.0 200880.0 51740.0 202225.0 ;
      RECT  51035.0 203570.0 51740.0 202225.0 ;
      RECT  51035.0 203570.0 51740.0 204915.0 ;
      RECT  51035.0 206260.0 51740.0 204915.0 ;
      RECT  51740.0 34100.0 52445.0 35445.0 ;
      RECT  51740.0 36790.0 52445.0 35445.0 ;
      RECT  51740.0 36790.0 52445.0 38135.0 ;
      RECT  51740.0 39480.0 52445.0 38135.0 ;
      RECT  51740.0 39480.0 52445.0 40825.0 ;
      RECT  51740.0 42170.0 52445.0 40825.0 ;
      RECT  51740.0 42170.0 52445.0 43515.0 ;
      RECT  51740.0 44860.0 52445.0 43515.0 ;
      RECT  51740.0 44860.0 52445.0 46205.0 ;
      RECT  51740.0 47550.0 52445.0 46205.0 ;
      RECT  51740.0 47550.0 52445.0 48895.0 ;
      RECT  51740.0 50240.0 52445.0 48895.0 ;
      RECT  51740.0 50240.0 52445.0 51585.0 ;
      RECT  51740.0 52930.0 52445.0 51585.0 ;
      RECT  51740.0 52930.0 52445.0 54275.0 ;
      RECT  51740.0 55620.0 52445.0 54275.0 ;
      RECT  51740.0 55620.0 52445.0 56965.0 ;
      RECT  51740.0 58310.0 52445.0 56965.0 ;
      RECT  51740.0 58310.0 52445.0 59655.0 ;
      RECT  51740.0 61000.0 52445.0 59655.0 ;
      RECT  51740.0 61000.0 52445.0 62345.0 ;
      RECT  51740.0 63690.0 52445.0 62345.0 ;
      RECT  51740.0 63690.0 52445.0 65035.0 ;
      RECT  51740.0 66380.0 52445.0 65035.0 ;
      RECT  51740.0 66380.0 52445.0 67725.0 ;
      RECT  51740.0 69070.0 52445.0 67725.0 ;
      RECT  51740.0 69070.0 52445.0 70415.0 ;
      RECT  51740.0 71760.0 52445.0 70415.0 ;
      RECT  51740.0 71760.0 52445.0 73105.0 ;
      RECT  51740.0 74450.0 52445.0 73105.0 ;
      RECT  51740.0 74450.0 52445.0 75795.0 ;
      RECT  51740.0 77140.0 52445.0 75795.0 ;
      RECT  51740.0 77140.0 52445.0 78485.0 ;
      RECT  51740.0 79830.0 52445.0 78485.0 ;
      RECT  51740.0 79830.0 52445.0 81175.0 ;
      RECT  51740.0 82520.0 52445.0 81175.0 ;
      RECT  51740.0 82520.0 52445.0 83865.0 ;
      RECT  51740.0 85210.0 52445.0 83865.0 ;
      RECT  51740.0 85210.0 52445.0 86555.0 ;
      RECT  51740.0 87900.0 52445.0 86555.0 ;
      RECT  51740.0 87900.0 52445.0 89245.0 ;
      RECT  51740.0 90590.0 52445.0 89245.0 ;
      RECT  51740.0 90590.0 52445.0 91935.0 ;
      RECT  51740.0 93280.0 52445.0 91935.0 ;
      RECT  51740.0 93280.0 52445.0 94625.0 ;
      RECT  51740.0 95970.0 52445.0 94625.0 ;
      RECT  51740.0 95970.0 52445.0 97315.0 ;
      RECT  51740.0 98660.0 52445.0 97315.0 ;
      RECT  51740.0 98660.0 52445.0 100005.0 ;
      RECT  51740.0 101350.0 52445.0 100005.0 ;
      RECT  51740.0 101350.0 52445.0 102695.0 ;
      RECT  51740.0 104040.0 52445.0 102695.0 ;
      RECT  51740.0 104040.0 52445.0 105385.0 ;
      RECT  51740.0 106730.0 52445.0 105385.0 ;
      RECT  51740.0 106730.0 52445.0 108075.0 ;
      RECT  51740.0 109420.0 52445.0 108075.0 ;
      RECT  51740.0 109420.0 52445.0 110765.0 ;
      RECT  51740.0 112110.0 52445.0 110765.0 ;
      RECT  51740.0 112110.0 52445.0 113455.0 ;
      RECT  51740.0 114800.0 52445.0 113455.0 ;
      RECT  51740.0 114800.0 52445.0 116145.0 ;
      RECT  51740.0 117490.0 52445.0 116145.0 ;
      RECT  51740.0 117490.0 52445.0 118835.0 ;
      RECT  51740.0 120180.0 52445.0 118835.0 ;
      RECT  51740.0 120180.0 52445.0 121525.0 ;
      RECT  51740.0 122870.0 52445.0 121525.0 ;
      RECT  51740.0 122870.0 52445.0 124215.0 ;
      RECT  51740.0 125560.0 52445.0 124215.0 ;
      RECT  51740.0 125560.0 52445.0 126905.0 ;
      RECT  51740.0 128250.0 52445.0 126905.0 ;
      RECT  51740.0 128250.0 52445.0 129595.0 ;
      RECT  51740.0 130940.0 52445.0 129595.0 ;
      RECT  51740.0 130940.0 52445.0 132285.0 ;
      RECT  51740.0 133630.0 52445.0 132285.0 ;
      RECT  51740.0 133630.0 52445.0 134975.0 ;
      RECT  51740.0 136320.0 52445.0 134975.0 ;
      RECT  51740.0 136320.0 52445.0 137665.0 ;
      RECT  51740.0 139010.0 52445.0 137665.0 ;
      RECT  51740.0 139010.0 52445.0 140355.0 ;
      RECT  51740.0 141700.0 52445.0 140355.0 ;
      RECT  51740.0 141700.0 52445.0 143045.0 ;
      RECT  51740.0 144390.0 52445.0 143045.0 ;
      RECT  51740.0 144390.0 52445.0 145735.0 ;
      RECT  51740.0 147080.0 52445.0 145735.0 ;
      RECT  51740.0 147080.0 52445.0 148425.0 ;
      RECT  51740.0 149770.0 52445.0 148425.0 ;
      RECT  51740.0 149770.0 52445.0 151115.0 ;
      RECT  51740.0 152460.0 52445.0 151115.0 ;
      RECT  51740.0 152460.0 52445.0 153805.0 ;
      RECT  51740.0 155150.0 52445.0 153805.0 ;
      RECT  51740.0 155150.0 52445.0 156495.0 ;
      RECT  51740.0 157840.0 52445.0 156495.0 ;
      RECT  51740.0 157840.0 52445.0 159185.0 ;
      RECT  51740.0 160530.0 52445.0 159185.0 ;
      RECT  51740.0 160530.0 52445.0 161875.0 ;
      RECT  51740.0 163220.0 52445.0 161875.0 ;
      RECT  51740.0 163220.0 52445.0 164565.0 ;
      RECT  51740.0 165910.0 52445.0 164565.0 ;
      RECT  51740.0 165910.0 52445.0 167255.0 ;
      RECT  51740.0 168600.0 52445.0 167255.0 ;
      RECT  51740.0 168600.0 52445.0 169945.0 ;
      RECT  51740.0 171290.0 52445.0 169945.0 ;
      RECT  51740.0 171290.0 52445.0 172635.0 ;
      RECT  51740.0 173980.0 52445.0 172635.0 ;
      RECT  51740.0 173980.0 52445.0 175325.0 ;
      RECT  51740.0 176670.0 52445.0 175325.0 ;
      RECT  51740.0 176670.0 52445.0 178015.0 ;
      RECT  51740.0 179360.0 52445.0 178015.0 ;
      RECT  51740.0 179360.0 52445.0 180705.0 ;
      RECT  51740.0 182050.0 52445.0 180705.0 ;
      RECT  51740.0 182050.0 52445.0 183395.0 ;
      RECT  51740.0 184740.0 52445.0 183395.0 ;
      RECT  51740.0 184740.0 52445.0 186085.0 ;
      RECT  51740.0 187430.0 52445.0 186085.0 ;
      RECT  51740.0 187430.0 52445.0 188775.0 ;
      RECT  51740.0 190120.0 52445.0 188775.0 ;
      RECT  51740.0 190120.0 52445.0 191465.0 ;
      RECT  51740.0 192810.0 52445.0 191465.0 ;
      RECT  51740.0 192810.0 52445.0 194155.0 ;
      RECT  51740.0 195500.0 52445.0 194155.0 ;
      RECT  51740.0 195500.0 52445.0 196845.0 ;
      RECT  51740.0 198190.0 52445.0 196845.0 ;
      RECT  51740.0 198190.0 52445.0 199535.0 ;
      RECT  51740.0 200880.0 52445.0 199535.0 ;
      RECT  51740.0 200880.0 52445.0 202225.0 ;
      RECT  51740.0 203570.0 52445.0 202225.0 ;
      RECT  51740.0 203570.0 52445.0 204915.0 ;
      RECT  51740.0 206260.0 52445.0 204915.0 ;
      RECT  52445.0 34100.0 53150.0 35445.0 ;
      RECT  52445.0 36790.0 53150.0 35445.0 ;
      RECT  52445.0 36790.0 53150.0 38135.0 ;
      RECT  52445.0 39480.0 53150.0 38135.0 ;
      RECT  52445.0 39480.0 53150.0 40825.0 ;
      RECT  52445.0 42170.0 53150.0 40825.0 ;
      RECT  52445.0 42170.0 53150.0 43515.0 ;
      RECT  52445.0 44860.0 53150.0 43515.0 ;
      RECT  52445.0 44860.0 53150.0 46205.0 ;
      RECT  52445.0 47550.0 53150.0 46205.0 ;
      RECT  52445.0 47550.0 53150.0 48895.0 ;
      RECT  52445.0 50240.0 53150.0 48895.0 ;
      RECT  52445.0 50240.0 53150.0 51585.0 ;
      RECT  52445.0 52930.0 53150.0 51585.0 ;
      RECT  52445.0 52930.0 53150.0 54275.0 ;
      RECT  52445.0 55620.0 53150.0 54275.0 ;
      RECT  52445.0 55620.0 53150.0 56965.0 ;
      RECT  52445.0 58310.0 53150.0 56965.0 ;
      RECT  52445.0 58310.0 53150.0 59655.0 ;
      RECT  52445.0 61000.0 53150.0 59655.0 ;
      RECT  52445.0 61000.0 53150.0 62345.0 ;
      RECT  52445.0 63690.0 53150.0 62345.0 ;
      RECT  52445.0 63690.0 53150.0 65035.0 ;
      RECT  52445.0 66380.0 53150.0 65035.0 ;
      RECT  52445.0 66380.0 53150.0 67725.0 ;
      RECT  52445.0 69070.0 53150.0 67725.0 ;
      RECT  52445.0 69070.0 53150.0 70415.0 ;
      RECT  52445.0 71760.0 53150.0 70415.0 ;
      RECT  52445.0 71760.0 53150.0 73105.0 ;
      RECT  52445.0 74450.0 53150.0 73105.0 ;
      RECT  52445.0 74450.0 53150.0 75795.0 ;
      RECT  52445.0 77140.0 53150.0 75795.0 ;
      RECT  52445.0 77140.0 53150.0 78485.0 ;
      RECT  52445.0 79830.0 53150.0 78485.0 ;
      RECT  52445.0 79830.0 53150.0 81175.0 ;
      RECT  52445.0 82520.0 53150.0 81175.0 ;
      RECT  52445.0 82520.0 53150.0 83865.0 ;
      RECT  52445.0 85210.0 53150.0 83865.0 ;
      RECT  52445.0 85210.0 53150.0 86555.0 ;
      RECT  52445.0 87900.0 53150.0 86555.0 ;
      RECT  52445.0 87900.0 53150.0 89245.0 ;
      RECT  52445.0 90590.0 53150.0 89245.0 ;
      RECT  52445.0 90590.0 53150.0 91935.0 ;
      RECT  52445.0 93280.0 53150.0 91935.0 ;
      RECT  52445.0 93280.0 53150.0 94625.0 ;
      RECT  52445.0 95970.0 53150.0 94625.0 ;
      RECT  52445.0 95970.0 53150.0 97315.0 ;
      RECT  52445.0 98660.0 53150.0 97315.0 ;
      RECT  52445.0 98660.0 53150.0 100005.0 ;
      RECT  52445.0 101350.0 53150.0 100005.0 ;
      RECT  52445.0 101350.0 53150.0 102695.0 ;
      RECT  52445.0 104040.0 53150.0 102695.0 ;
      RECT  52445.0 104040.0 53150.0 105385.0 ;
      RECT  52445.0 106730.0 53150.0 105385.0 ;
      RECT  52445.0 106730.0 53150.0 108075.0 ;
      RECT  52445.0 109420.0 53150.0 108075.0 ;
      RECT  52445.0 109420.0 53150.0 110765.0 ;
      RECT  52445.0 112110.0 53150.0 110765.0 ;
      RECT  52445.0 112110.0 53150.0 113455.0 ;
      RECT  52445.0 114800.0 53150.0 113455.0 ;
      RECT  52445.0 114800.0 53150.0 116145.0 ;
      RECT  52445.0 117490.0 53150.0 116145.0 ;
      RECT  52445.0 117490.0 53150.0 118835.0 ;
      RECT  52445.0 120180.0 53150.0 118835.0 ;
      RECT  52445.0 120180.0 53150.0 121525.0 ;
      RECT  52445.0 122870.0 53150.0 121525.0 ;
      RECT  52445.0 122870.0 53150.0 124215.0 ;
      RECT  52445.0 125560.0 53150.0 124215.0 ;
      RECT  52445.0 125560.0 53150.0 126905.0 ;
      RECT  52445.0 128250.0 53150.0 126905.0 ;
      RECT  52445.0 128250.0 53150.0 129595.0 ;
      RECT  52445.0 130940.0 53150.0 129595.0 ;
      RECT  52445.0 130940.0 53150.0 132285.0 ;
      RECT  52445.0 133630.0 53150.0 132285.0 ;
      RECT  52445.0 133630.0 53150.0 134975.0 ;
      RECT  52445.0 136320.0 53150.0 134975.0 ;
      RECT  52445.0 136320.0 53150.0 137665.0 ;
      RECT  52445.0 139010.0 53150.0 137665.0 ;
      RECT  52445.0 139010.0 53150.0 140355.0 ;
      RECT  52445.0 141700.0 53150.0 140355.0 ;
      RECT  52445.0 141700.0 53150.0 143045.0 ;
      RECT  52445.0 144390.0 53150.0 143045.0 ;
      RECT  52445.0 144390.0 53150.0 145735.0 ;
      RECT  52445.0 147080.0 53150.0 145735.0 ;
      RECT  52445.0 147080.0 53150.0 148425.0 ;
      RECT  52445.0 149770.0 53150.0 148425.0 ;
      RECT  52445.0 149770.0 53150.0 151115.0 ;
      RECT  52445.0 152460.0 53150.0 151115.0 ;
      RECT  52445.0 152460.0 53150.0 153805.0 ;
      RECT  52445.0 155150.0 53150.0 153805.0 ;
      RECT  52445.0 155150.0 53150.0 156495.0 ;
      RECT  52445.0 157840.0 53150.0 156495.0 ;
      RECT  52445.0 157840.0 53150.0 159185.0 ;
      RECT  52445.0 160530.0 53150.0 159185.0 ;
      RECT  52445.0 160530.0 53150.0 161875.0 ;
      RECT  52445.0 163220.0 53150.0 161875.0 ;
      RECT  52445.0 163220.0 53150.0 164565.0 ;
      RECT  52445.0 165910.0 53150.0 164565.0 ;
      RECT  52445.0 165910.0 53150.0 167255.0 ;
      RECT  52445.0 168600.0 53150.0 167255.0 ;
      RECT  52445.0 168600.0 53150.0 169945.0 ;
      RECT  52445.0 171290.0 53150.0 169945.0 ;
      RECT  52445.0 171290.0 53150.0 172635.0 ;
      RECT  52445.0 173980.0 53150.0 172635.0 ;
      RECT  52445.0 173980.0 53150.0 175325.0 ;
      RECT  52445.0 176670.0 53150.0 175325.0 ;
      RECT  52445.0 176670.0 53150.0 178015.0 ;
      RECT  52445.0 179360.0 53150.0 178015.0 ;
      RECT  52445.0 179360.0 53150.0 180705.0 ;
      RECT  52445.0 182050.0 53150.0 180705.0 ;
      RECT  52445.0 182050.0 53150.0 183395.0 ;
      RECT  52445.0 184740.0 53150.0 183395.0 ;
      RECT  52445.0 184740.0 53150.0 186085.0 ;
      RECT  52445.0 187430.0 53150.0 186085.0 ;
      RECT  52445.0 187430.0 53150.0 188775.0 ;
      RECT  52445.0 190120.0 53150.0 188775.0 ;
      RECT  52445.0 190120.0 53150.0 191465.0 ;
      RECT  52445.0 192810.0 53150.0 191465.0 ;
      RECT  52445.0 192810.0 53150.0 194155.0 ;
      RECT  52445.0 195500.0 53150.0 194155.0 ;
      RECT  52445.0 195500.0 53150.0 196845.0 ;
      RECT  52445.0 198190.0 53150.0 196845.0 ;
      RECT  52445.0 198190.0 53150.0 199535.0 ;
      RECT  52445.0 200880.0 53150.0 199535.0 ;
      RECT  52445.0 200880.0 53150.0 202225.0 ;
      RECT  52445.0 203570.0 53150.0 202225.0 ;
      RECT  52445.0 203570.0 53150.0 204915.0 ;
      RECT  52445.0 206260.0 53150.0 204915.0 ;
      RECT  53150.0 34100.0 53855.0 35445.0 ;
      RECT  53150.0 36790.0 53855.0 35445.0 ;
      RECT  53150.0 36790.0 53855.0 38135.0 ;
      RECT  53150.0 39480.0 53855.0 38135.0 ;
      RECT  53150.0 39480.0 53855.0 40825.0 ;
      RECT  53150.0 42170.0 53855.0 40825.0 ;
      RECT  53150.0 42170.0 53855.0 43515.0 ;
      RECT  53150.0 44860.0 53855.0 43515.0 ;
      RECT  53150.0 44860.0 53855.0 46205.0 ;
      RECT  53150.0 47550.0 53855.0 46205.0 ;
      RECT  53150.0 47550.0 53855.0 48895.0 ;
      RECT  53150.0 50240.0 53855.0 48895.0 ;
      RECT  53150.0 50240.0 53855.0 51585.0 ;
      RECT  53150.0 52930.0 53855.0 51585.0 ;
      RECT  53150.0 52930.0 53855.0 54275.0 ;
      RECT  53150.0 55620.0 53855.0 54275.0 ;
      RECT  53150.0 55620.0 53855.0 56965.0 ;
      RECT  53150.0 58310.0 53855.0 56965.0 ;
      RECT  53150.0 58310.0 53855.0 59655.0 ;
      RECT  53150.0 61000.0 53855.0 59655.0 ;
      RECT  53150.0 61000.0 53855.0 62345.0 ;
      RECT  53150.0 63690.0 53855.0 62345.0 ;
      RECT  53150.0 63690.0 53855.0 65035.0 ;
      RECT  53150.0 66380.0 53855.0 65035.0 ;
      RECT  53150.0 66380.0 53855.0 67725.0 ;
      RECT  53150.0 69070.0 53855.0 67725.0 ;
      RECT  53150.0 69070.0 53855.0 70415.0 ;
      RECT  53150.0 71760.0 53855.0 70415.0 ;
      RECT  53150.0 71760.0 53855.0 73105.0 ;
      RECT  53150.0 74450.0 53855.0 73105.0 ;
      RECT  53150.0 74450.0 53855.0 75795.0 ;
      RECT  53150.0 77140.0 53855.0 75795.0 ;
      RECT  53150.0 77140.0 53855.0 78485.0 ;
      RECT  53150.0 79830.0 53855.0 78485.0 ;
      RECT  53150.0 79830.0 53855.0 81175.0 ;
      RECT  53150.0 82520.0 53855.0 81175.0 ;
      RECT  53150.0 82520.0 53855.0 83865.0 ;
      RECT  53150.0 85210.0 53855.0 83865.0 ;
      RECT  53150.0 85210.0 53855.0 86555.0 ;
      RECT  53150.0 87900.0 53855.0 86555.0 ;
      RECT  53150.0 87900.0 53855.0 89245.0 ;
      RECT  53150.0 90590.0 53855.0 89245.0 ;
      RECT  53150.0 90590.0 53855.0 91935.0 ;
      RECT  53150.0 93280.0 53855.0 91935.0 ;
      RECT  53150.0 93280.0 53855.0 94625.0 ;
      RECT  53150.0 95970.0 53855.0 94625.0 ;
      RECT  53150.0 95970.0 53855.0 97315.0 ;
      RECT  53150.0 98660.0 53855.0 97315.0 ;
      RECT  53150.0 98660.0 53855.0 100005.0 ;
      RECT  53150.0 101350.0 53855.0 100005.0 ;
      RECT  53150.0 101350.0 53855.0 102695.0 ;
      RECT  53150.0 104040.0 53855.0 102695.0 ;
      RECT  53150.0 104040.0 53855.0 105385.0 ;
      RECT  53150.0 106730.0 53855.0 105385.0 ;
      RECT  53150.0 106730.0 53855.0 108075.0 ;
      RECT  53150.0 109420.0 53855.0 108075.0 ;
      RECT  53150.0 109420.0 53855.0 110765.0 ;
      RECT  53150.0 112110.0 53855.0 110765.0 ;
      RECT  53150.0 112110.0 53855.0 113455.0 ;
      RECT  53150.0 114800.0 53855.0 113455.0 ;
      RECT  53150.0 114800.0 53855.0 116145.0 ;
      RECT  53150.0 117490.0 53855.0 116145.0 ;
      RECT  53150.0 117490.0 53855.0 118835.0 ;
      RECT  53150.0 120180.0 53855.0 118835.0 ;
      RECT  53150.0 120180.0 53855.0 121525.0 ;
      RECT  53150.0 122870.0 53855.0 121525.0 ;
      RECT  53150.0 122870.0 53855.0 124215.0 ;
      RECT  53150.0 125560.0 53855.0 124215.0 ;
      RECT  53150.0 125560.0 53855.0 126905.0 ;
      RECT  53150.0 128250.0 53855.0 126905.0 ;
      RECT  53150.0 128250.0 53855.0 129595.0 ;
      RECT  53150.0 130940.0 53855.0 129595.0 ;
      RECT  53150.0 130940.0 53855.0 132285.0 ;
      RECT  53150.0 133630.0 53855.0 132285.0 ;
      RECT  53150.0 133630.0 53855.0 134975.0 ;
      RECT  53150.0 136320.0 53855.0 134975.0 ;
      RECT  53150.0 136320.0 53855.0 137665.0 ;
      RECT  53150.0 139010.0 53855.0 137665.0 ;
      RECT  53150.0 139010.0 53855.0 140355.0 ;
      RECT  53150.0 141700.0 53855.0 140355.0 ;
      RECT  53150.0 141700.0 53855.0 143045.0 ;
      RECT  53150.0 144390.0 53855.0 143045.0 ;
      RECT  53150.0 144390.0 53855.0 145735.0 ;
      RECT  53150.0 147080.0 53855.0 145735.0 ;
      RECT  53150.0 147080.0 53855.0 148425.0 ;
      RECT  53150.0 149770.0 53855.0 148425.0 ;
      RECT  53150.0 149770.0 53855.0 151115.0 ;
      RECT  53150.0 152460.0 53855.0 151115.0 ;
      RECT  53150.0 152460.0 53855.0 153805.0 ;
      RECT  53150.0 155150.0 53855.0 153805.0 ;
      RECT  53150.0 155150.0 53855.0 156495.0 ;
      RECT  53150.0 157840.0 53855.0 156495.0 ;
      RECT  53150.0 157840.0 53855.0 159185.0 ;
      RECT  53150.0 160530.0 53855.0 159185.0 ;
      RECT  53150.0 160530.0 53855.0 161875.0 ;
      RECT  53150.0 163220.0 53855.0 161875.0 ;
      RECT  53150.0 163220.0 53855.0 164565.0 ;
      RECT  53150.0 165910.0 53855.0 164565.0 ;
      RECT  53150.0 165910.0 53855.0 167255.0 ;
      RECT  53150.0 168600.0 53855.0 167255.0 ;
      RECT  53150.0 168600.0 53855.0 169945.0 ;
      RECT  53150.0 171290.0 53855.0 169945.0 ;
      RECT  53150.0 171290.0 53855.0 172635.0 ;
      RECT  53150.0 173980.0 53855.0 172635.0 ;
      RECT  53150.0 173980.0 53855.0 175325.0 ;
      RECT  53150.0 176670.0 53855.0 175325.0 ;
      RECT  53150.0 176670.0 53855.0 178015.0 ;
      RECT  53150.0 179360.0 53855.0 178015.0 ;
      RECT  53150.0 179360.0 53855.0 180705.0 ;
      RECT  53150.0 182050.0 53855.0 180705.0 ;
      RECT  53150.0 182050.0 53855.0 183395.0 ;
      RECT  53150.0 184740.0 53855.0 183395.0 ;
      RECT  53150.0 184740.0 53855.0 186085.0 ;
      RECT  53150.0 187430.0 53855.0 186085.0 ;
      RECT  53150.0 187430.0 53855.0 188775.0 ;
      RECT  53150.0 190120.0 53855.0 188775.0 ;
      RECT  53150.0 190120.0 53855.0 191465.0 ;
      RECT  53150.0 192810.0 53855.0 191465.0 ;
      RECT  53150.0 192810.0 53855.0 194155.0 ;
      RECT  53150.0 195500.0 53855.0 194155.0 ;
      RECT  53150.0 195500.0 53855.0 196845.0 ;
      RECT  53150.0 198190.0 53855.0 196845.0 ;
      RECT  53150.0 198190.0 53855.0 199535.0 ;
      RECT  53150.0 200880.0 53855.0 199535.0 ;
      RECT  53150.0 200880.0 53855.0 202225.0 ;
      RECT  53150.0 203570.0 53855.0 202225.0 ;
      RECT  53150.0 203570.0 53855.0 204915.0 ;
      RECT  53150.0 206260.0 53855.0 204915.0 ;
      RECT  53855.0 34100.0 54560.0 35445.0 ;
      RECT  53855.0 36790.0 54560.0 35445.0 ;
      RECT  53855.0 36790.0 54560.0 38135.0 ;
      RECT  53855.0 39480.0 54560.0 38135.0 ;
      RECT  53855.0 39480.0 54560.0 40825.0 ;
      RECT  53855.0 42170.0 54560.0 40825.0 ;
      RECT  53855.0 42170.0 54560.0 43515.0 ;
      RECT  53855.0 44860.0 54560.0 43515.0 ;
      RECT  53855.0 44860.0 54560.0 46205.0 ;
      RECT  53855.0 47550.0 54560.0 46205.0 ;
      RECT  53855.0 47550.0 54560.0 48895.0 ;
      RECT  53855.0 50240.0 54560.0 48895.0 ;
      RECT  53855.0 50240.0 54560.0 51585.0 ;
      RECT  53855.0 52930.0 54560.0 51585.0 ;
      RECT  53855.0 52930.0 54560.0 54275.0 ;
      RECT  53855.0 55620.0 54560.0 54275.0 ;
      RECT  53855.0 55620.0 54560.0 56965.0 ;
      RECT  53855.0 58310.0 54560.0 56965.0 ;
      RECT  53855.0 58310.0 54560.0 59655.0 ;
      RECT  53855.0 61000.0 54560.0 59655.0 ;
      RECT  53855.0 61000.0 54560.0 62345.0 ;
      RECT  53855.0 63690.0 54560.0 62345.0 ;
      RECT  53855.0 63690.0 54560.0 65035.0 ;
      RECT  53855.0 66380.0 54560.0 65035.0 ;
      RECT  53855.0 66380.0 54560.0 67725.0 ;
      RECT  53855.0 69070.0 54560.0 67725.0 ;
      RECT  53855.0 69070.0 54560.0 70415.0 ;
      RECT  53855.0 71760.0 54560.0 70415.0 ;
      RECT  53855.0 71760.0 54560.0 73105.0 ;
      RECT  53855.0 74450.0 54560.0 73105.0 ;
      RECT  53855.0 74450.0 54560.0 75795.0 ;
      RECT  53855.0 77140.0 54560.0 75795.0 ;
      RECT  53855.0 77140.0 54560.0 78485.0 ;
      RECT  53855.0 79830.0 54560.0 78485.0 ;
      RECT  53855.0 79830.0 54560.0 81175.0 ;
      RECT  53855.0 82520.0 54560.0 81175.0 ;
      RECT  53855.0 82520.0 54560.0 83865.0 ;
      RECT  53855.0 85210.0 54560.0 83865.0 ;
      RECT  53855.0 85210.0 54560.0 86555.0 ;
      RECT  53855.0 87900.0 54560.0 86555.0 ;
      RECT  53855.0 87900.0 54560.0 89245.0 ;
      RECT  53855.0 90590.0 54560.0 89245.0 ;
      RECT  53855.0 90590.0 54560.0 91935.0 ;
      RECT  53855.0 93280.0 54560.0 91935.0 ;
      RECT  53855.0 93280.0 54560.0 94625.0 ;
      RECT  53855.0 95970.0 54560.0 94625.0 ;
      RECT  53855.0 95970.0 54560.0 97315.0 ;
      RECT  53855.0 98660.0 54560.0 97315.0 ;
      RECT  53855.0 98660.0 54560.0 100005.0 ;
      RECT  53855.0 101350.0 54560.0 100005.0 ;
      RECT  53855.0 101350.0 54560.0 102695.0 ;
      RECT  53855.0 104040.0 54560.0 102695.0 ;
      RECT  53855.0 104040.0 54560.0 105385.0 ;
      RECT  53855.0 106730.0 54560.0 105385.0 ;
      RECT  53855.0 106730.0 54560.0 108075.0 ;
      RECT  53855.0 109420.0 54560.0 108075.0 ;
      RECT  53855.0 109420.0 54560.0 110765.0 ;
      RECT  53855.0 112110.0 54560.0 110765.0 ;
      RECT  53855.0 112110.0 54560.0 113455.0 ;
      RECT  53855.0 114800.0 54560.0 113455.0 ;
      RECT  53855.0 114800.0 54560.0 116145.0 ;
      RECT  53855.0 117490.0 54560.0 116145.0 ;
      RECT  53855.0 117490.0 54560.0 118835.0 ;
      RECT  53855.0 120180.0 54560.0 118835.0 ;
      RECT  53855.0 120180.0 54560.0 121525.0 ;
      RECT  53855.0 122870.0 54560.0 121525.0 ;
      RECT  53855.0 122870.0 54560.0 124215.0 ;
      RECT  53855.0 125560.0 54560.0 124215.0 ;
      RECT  53855.0 125560.0 54560.0 126905.0 ;
      RECT  53855.0 128250.0 54560.0 126905.0 ;
      RECT  53855.0 128250.0 54560.0 129595.0 ;
      RECT  53855.0 130940.0 54560.0 129595.0 ;
      RECT  53855.0 130940.0 54560.0 132285.0 ;
      RECT  53855.0 133630.0 54560.0 132285.0 ;
      RECT  53855.0 133630.0 54560.0 134975.0 ;
      RECT  53855.0 136320.0 54560.0 134975.0 ;
      RECT  53855.0 136320.0 54560.0 137665.0 ;
      RECT  53855.0 139010.0 54560.0 137665.0 ;
      RECT  53855.0 139010.0 54560.0 140355.0 ;
      RECT  53855.0 141700.0 54560.0 140355.0 ;
      RECT  53855.0 141700.0 54560.0 143045.0 ;
      RECT  53855.0 144390.0 54560.0 143045.0 ;
      RECT  53855.0 144390.0 54560.0 145735.0 ;
      RECT  53855.0 147080.0 54560.0 145735.0 ;
      RECT  53855.0 147080.0 54560.0 148425.0 ;
      RECT  53855.0 149770.0 54560.0 148425.0 ;
      RECT  53855.0 149770.0 54560.0 151115.0 ;
      RECT  53855.0 152460.0 54560.0 151115.0 ;
      RECT  53855.0 152460.0 54560.0 153805.0 ;
      RECT  53855.0 155150.0 54560.0 153805.0 ;
      RECT  53855.0 155150.0 54560.0 156495.0 ;
      RECT  53855.0 157840.0 54560.0 156495.0 ;
      RECT  53855.0 157840.0 54560.0 159185.0 ;
      RECT  53855.0 160530.0 54560.0 159185.0 ;
      RECT  53855.0 160530.0 54560.0 161875.0 ;
      RECT  53855.0 163220.0 54560.0 161875.0 ;
      RECT  53855.0 163220.0 54560.0 164565.0 ;
      RECT  53855.0 165910.0 54560.0 164565.0 ;
      RECT  53855.0 165910.0 54560.0 167255.0 ;
      RECT  53855.0 168600.0 54560.0 167255.0 ;
      RECT  53855.0 168600.0 54560.0 169945.0 ;
      RECT  53855.0 171290.0 54560.0 169945.0 ;
      RECT  53855.0 171290.0 54560.0 172635.0 ;
      RECT  53855.0 173980.0 54560.0 172635.0 ;
      RECT  53855.0 173980.0 54560.0 175325.0 ;
      RECT  53855.0 176670.0 54560.0 175325.0 ;
      RECT  53855.0 176670.0 54560.0 178015.0 ;
      RECT  53855.0 179360.0 54560.0 178015.0 ;
      RECT  53855.0 179360.0 54560.0 180705.0 ;
      RECT  53855.0 182050.0 54560.0 180705.0 ;
      RECT  53855.0 182050.0 54560.0 183395.0 ;
      RECT  53855.0 184740.0 54560.0 183395.0 ;
      RECT  53855.0 184740.0 54560.0 186085.0 ;
      RECT  53855.0 187430.0 54560.0 186085.0 ;
      RECT  53855.0 187430.0 54560.0 188775.0 ;
      RECT  53855.0 190120.0 54560.0 188775.0 ;
      RECT  53855.0 190120.0 54560.0 191465.0 ;
      RECT  53855.0 192810.0 54560.0 191465.0 ;
      RECT  53855.0 192810.0 54560.0 194155.0 ;
      RECT  53855.0 195500.0 54560.0 194155.0 ;
      RECT  53855.0 195500.0 54560.0 196845.0 ;
      RECT  53855.0 198190.0 54560.0 196845.0 ;
      RECT  53855.0 198190.0 54560.0 199535.0 ;
      RECT  53855.0 200880.0 54560.0 199535.0 ;
      RECT  53855.0 200880.0 54560.0 202225.0 ;
      RECT  53855.0 203570.0 54560.0 202225.0 ;
      RECT  53855.0 203570.0 54560.0 204915.0 ;
      RECT  53855.0 206260.0 54560.0 204915.0 ;
      RECT  54560.0 34100.0 55265.0 35445.0 ;
      RECT  54560.0 36790.0 55265.0 35445.0 ;
      RECT  54560.0 36790.0 55265.0 38135.0 ;
      RECT  54560.0 39480.0 55265.0 38135.0 ;
      RECT  54560.0 39480.0 55265.0 40825.0 ;
      RECT  54560.0 42170.0 55265.0 40825.0 ;
      RECT  54560.0 42170.0 55265.0 43515.0 ;
      RECT  54560.0 44860.0 55265.0 43515.0 ;
      RECT  54560.0 44860.0 55265.0 46205.0 ;
      RECT  54560.0 47550.0 55265.0 46205.0 ;
      RECT  54560.0 47550.0 55265.0 48895.0 ;
      RECT  54560.0 50240.0 55265.0 48895.0 ;
      RECT  54560.0 50240.0 55265.0 51585.0 ;
      RECT  54560.0 52930.0 55265.0 51585.0 ;
      RECT  54560.0 52930.0 55265.0 54275.0 ;
      RECT  54560.0 55620.0 55265.0 54275.0 ;
      RECT  54560.0 55620.0 55265.0 56965.0 ;
      RECT  54560.0 58310.0 55265.0 56965.0 ;
      RECT  54560.0 58310.0 55265.0 59655.0 ;
      RECT  54560.0 61000.0 55265.0 59655.0 ;
      RECT  54560.0 61000.0 55265.0 62345.0 ;
      RECT  54560.0 63690.0 55265.0 62345.0 ;
      RECT  54560.0 63690.0 55265.0 65035.0 ;
      RECT  54560.0 66380.0 55265.0 65035.0 ;
      RECT  54560.0 66380.0 55265.0 67725.0 ;
      RECT  54560.0 69070.0 55265.0 67725.0 ;
      RECT  54560.0 69070.0 55265.0 70415.0 ;
      RECT  54560.0 71760.0 55265.0 70415.0 ;
      RECT  54560.0 71760.0 55265.0 73105.0 ;
      RECT  54560.0 74450.0 55265.0 73105.0 ;
      RECT  54560.0 74450.0 55265.0 75795.0 ;
      RECT  54560.0 77140.0 55265.0 75795.0 ;
      RECT  54560.0 77140.0 55265.0 78485.0 ;
      RECT  54560.0 79830.0 55265.0 78485.0 ;
      RECT  54560.0 79830.0 55265.0 81175.0 ;
      RECT  54560.0 82520.0 55265.0 81175.0 ;
      RECT  54560.0 82520.0 55265.0 83865.0 ;
      RECT  54560.0 85210.0 55265.0 83865.0 ;
      RECT  54560.0 85210.0 55265.0 86555.0 ;
      RECT  54560.0 87900.0 55265.0 86555.0 ;
      RECT  54560.0 87900.0 55265.0 89245.0 ;
      RECT  54560.0 90590.0 55265.0 89245.0 ;
      RECT  54560.0 90590.0 55265.0 91935.0 ;
      RECT  54560.0 93280.0 55265.0 91935.0 ;
      RECT  54560.0 93280.0 55265.0 94625.0 ;
      RECT  54560.0 95970.0 55265.0 94625.0 ;
      RECT  54560.0 95970.0 55265.0 97315.0 ;
      RECT  54560.0 98660.0 55265.0 97315.0 ;
      RECT  54560.0 98660.0 55265.0 100005.0 ;
      RECT  54560.0 101350.0 55265.0 100005.0 ;
      RECT  54560.0 101350.0 55265.0 102695.0 ;
      RECT  54560.0 104040.0 55265.0 102695.0 ;
      RECT  54560.0 104040.0 55265.0 105385.0 ;
      RECT  54560.0 106730.0 55265.0 105385.0 ;
      RECT  54560.0 106730.0 55265.0 108075.0 ;
      RECT  54560.0 109420.0 55265.0 108075.0 ;
      RECT  54560.0 109420.0 55265.0 110765.0 ;
      RECT  54560.0 112110.0 55265.0 110765.0 ;
      RECT  54560.0 112110.0 55265.0 113455.0 ;
      RECT  54560.0 114800.0 55265.0 113455.0 ;
      RECT  54560.0 114800.0 55265.0 116145.0 ;
      RECT  54560.0 117490.0 55265.0 116145.0 ;
      RECT  54560.0 117490.0 55265.0 118835.0 ;
      RECT  54560.0 120180.0 55265.0 118835.0 ;
      RECT  54560.0 120180.0 55265.0 121525.0 ;
      RECT  54560.0 122870.0 55265.0 121525.0 ;
      RECT  54560.0 122870.0 55265.0 124215.0 ;
      RECT  54560.0 125560.0 55265.0 124215.0 ;
      RECT  54560.0 125560.0 55265.0 126905.0 ;
      RECT  54560.0 128250.0 55265.0 126905.0 ;
      RECT  54560.0 128250.0 55265.0 129595.0 ;
      RECT  54560.0 130940.0 55265.0 129595.0 ;
      RECT  54560.0 130940.0 55265.0 132285.0 ;
      RECT  54560.0 133630.0 55265.0 132285.0 ;
      RECT  54560.0 133630.0 55265.0 134975.0 ;
      RECT  54560.0 136320.0 55265.0 134975.0 ;
      RECT  54560.0 136320.0 55265.0 137665.0 ;
      RECT  54560.0 139010.0 55265.0 137665.0 ;
      RECT  54560.0 139010.0 55265.0 140355.0 ;
      RECT  54560.0 141700.0 55265.0 140355.0 ;
      RECT  54560.0 141700.0 55265.0 143045.0 ;
      RECT  54560.0 144390.0 55265.0 143045.0 ;
      RECT  54560.0 144390.0 55265.0 145735.0 ;
      RECT  54560.0 147080.0 55265.0 145735.0 ;
      RECT  54560.0 147080.0 55265.0 148425.0 ;
      RECT  54560.0 149770.0 55265.0 148425.0 ;
      RECT  54560.0 149770.0 55265.0 151115.0 ;
      RECT  54560.0 152460.0 55265.0 151115.0 ;
      RECT  54560.0 152460.0 55265.0 153805.0 ;
      RECT  54560.0 155150.0 55265.0 153805.0 ;
      RECT  54560.0 155150.0 55265.0 156495.0 ;
      RECT  54560.0 157840.0 55265.0 156495.0 ;
      RECT  54560.0 157840.0 55265.0 159185.0 ;
      RECT  54560.0 160530.0 55265.0 159185.0 ;
      RECT  54560.0 160530.0 55265.0 161875.0 ;
      RECT  54560.0 163220.0 55265.0 161875.0 ;
      RECT  54560.0 163220.0 55265.0 164565.0 ;
      RECT  54560.0 165910.0 55265.0 164565.0 ;
      RECT  54560.0 165910.0 55265.0 167255.0 ;
      RECT  54560.0 168600.0 55265.0 167255.0 ;
      RECT  54560.0 168600.0 55265.0 169945.0 ;
      RECT  54560.0 171290.0 55265.0 169945.0 ;
      RECT  54560.0 171290.0 55265.0 172635.0 ;
      RECT  54560.0 173980.0 55265.0 172635.0 ;
      RECT  54560.0 173980.0 55265.0 175325.0 ;
      RECT  54560.0 176670.0 55265.0 175325.0 ;
      RECT  54560.0 176670.0 55265.0 178015.0 ;
      RECT  54560.0 179360.0 55265.0 178015.0 ;
      RECT  54560.0 179360.0 55265.0 180705.0 ;
      RECT  54560.0 182050.0 55265.0 180705.0 ;
      RECT  54560.0 182050.0 55265.0 183395.0 ;
      RECT  54560.0 184740.0 55265.0 183395.0 ;
      RECT  54560.0 184740.0 55265.0 186085.0 ;
      RECT  54560.0 187430.0 55265.0 186085.0 ;
      RECT  54560.0 187430.0 55265.0 188775.0 ;
      RECT  54560.0 190120.0 55265.0 188775.0 ;
      RECT  54560.0 190120.0 55265.0 191465.0 ;
      RECT  54560.0 192810.0 55265.0 191465.0 ;
      RECT  54560.0 192810.0 55265.0 194155.0 ;
      RECT  54560.0 195500.0 55265.0 194155.0 ;
      RECT  54560.0 195500.0 55265.0 196845.0 ;
      RECT  54560.0 198190.0 55265.0 196845.0 ;
      RECT  54560.0 198190.0 55265.0 199535.0 ;
      RECT  54560.0 200880.0 55265.0 199535.0 ;
      RECT  54560.0 200880.0 55265.0 202225.0 ;
      RECT  54560.0 203570.0 55265.0 202225.0 ;
      RECT  54560.0 203570.0 55265.0 204915.0 ;
      RECT  54560.0 206260.0 55265.0 204915.0 ;
      RECT  55265.0 34100.0 55970.0 35445.0 ;
      RECT  55265.0 36790.0 55970.0 35445.0 ;
      RECT  55265.0 36790.0 55970.0 38135.0 ;
      RECT  55265.0 39480.0 55970.0 38135.0 ;
      RECT  55265.0 39480.0 55970.0 40825.0 ;
      RECT  55265.0 42170.0 55970.0 40825.0 ;
      RECT  55265.0 42170.0 55970.0 43515.0 ;
      RECT  55265.0 44860.0 55970.0 43515.0 ;
      RECT  55265.0 44860.0 55970.0 46205.0 ;
      RECT  55265.0 47550.0 55970.0 46205.0 ;
      RECT  55265.0 47550.0 55970.0 48895.0 ;
      RECT  55265.0 50240.0 55970.0 48895.0 ;
      RECT  55265.0 50240.0 55970.0 51585.0 ;
      RECT  55265.0 52930.0 55970.0 51585.0 ;
      RECT  55265.0 52930.0 55970.0 54275.0 ;
      RECT  55265.0 55620.0 55970.0 54275.0 ;
      RECT  55265.0 55620.0 55970.0 56965.0 ;
      RECT  55265.0 58310.0 55970.0 56965.0 ;
      RECT  55265.0 58310.0 55970.0 59655.0 ;
      RECT  55265.0 61000.0 55970.0 59655.0 ;
      RECT  55265.0 61000.0 55970.0 62345.0 ;
      RECT  55265.0 63690.0 55970.0 62345.0 ;
      RECT  55265.0 63690.0 55970.0 65035.0 ;
      RECT  55265.0 66380.0 55970.0 65035.0 ;
      RECT  55265.0 66380.0 55970.0 67725.0 ;
      RECT  55265.0 69070.0 55970.0 67725.0 ;
      RECT  55265.0 69070.0 55970.0 70415.0 ;
      RECT  55265.0 71760.0 55970.0 70415.0 ;
      RECT  55265.0 71760.0 55970.0 73105.0 ;
      RECT  55265.0 74450.0 55970.0 73105.0 ;
      RECT  55265.0 74450.0 55970.0 75795.0 ;
      RECT  55265.0 77140.0 55970.0 75795.0 ;
      RECT  55265.0 77140.0 55970.0 78485.0 ;
      RECT  55265.0 79830.0 55970.0 78485.0 ;
      RECT  55265.0 79830.0 55970.0 81175.0 ;
      RECT  55265.0 82520.0 55970.0 81175.0 ;
      RECT  55265.0 82520.0 55970.0 83865.0 ;
      RECT  55265.0 85210.0 55970.0 83865.0 ;
      RECT  55265.0 85210.0 55970.0 86555.0 ;
      RECT  55265.0 87900.0 55970.0 86555.0 ;
      RECT  55265.0 87900.0 55970.0 89245.0 ;
      RECT  55265.0 90590.0 55970.0 89245.0 ;
      RECT  55265.0 90590.0 55970.0 91935.0 ;
      RECT  55265.0 93280.0 55970.0 91935.0 ;
      RECT  55265.0 93280.0 55970.0 94625.0 ;
      RECT  55265.0 95970.0 55970.0 94625.0 ;
      RECT  55265.0 95970.0 55970.0 97315.0 ;
      RECT  55265.0 98660.0 55970.0 97315.0 ;
      RECT  55265.0 98660.0 55970.0 100005.0 ;
      RECT  55265.0 101350.0 55970.0 100005.0 ;
      RECT  55265.0 101350.0 55970.0 102695.0 ;
      RECT  55265.0 104040.0 55970.0 102695.0 ;
      RECT  55265.0 104040.0 55970.0 105385.0 ;
      RECT  55265.0 106730.0 55970.0 105385.0 ;
      RECT  55265.0 106730.0 55970.0 108075.0 ;
      RECT  55265.0 109420.0 55970.0 108075.0 ;
      RECT  55265.0 109420.0 55970.0 110765.0 ;
      RECT  55265.0 112110.0 55970.0 110765.0 ;
      RECT  55265.0 112110.0 55970.0 113455.0 ;
      RECT  55265.0 114800.0 55970.0 113455.0 ;
      RECT  55265.0 114800.0 55970.0 116145.0 ;
      RECT  55265.0 117490.0 55970.0 116145.0 ;
      RECT  55265.0 117490.0 55970.0 118835.0 ;
      RECT  55265.0 120180.0 55970.0 118835.0 ;
      RECT  55265.0 120180.0 55970.0 121525.0 ;
      RECT  55265.0 122870.0 55970.0 121525.0 ;
      RECT  55265.0 122870.0 55970.0 124215.0 ;
      RECT  55265.0 125560.0 55970.0 124215.0 ;
      RECT  55265.0 125560.0 55970.0 126905.0 ;
      RECT  55265.0 128250.0 55970.0 126905.0 ;
      RECT  55265.0 128250.0 55970.0 129595.0 ;
      RECT  55265.0 130940.0 55970.0 129595.0 ;
      RECT  55265.0 130940.0 55970.0 132285.0 ;
      RECT  55265.0 133630.0 55970.0 132285.0 ;
      RECT  55265.0 133630.0 55970.0 134975.0 ;
      RECT  55265.0 136320.0 55970.0 134975.0 ;
      RECT  55265.0 136320.0 55970.0 137665.0 ;
      RECT  55265.0 139010.0 55970.0 137665.0 ;
      RECT  55265.0 139010.0 55970.0 140355.0 ;
      RECT  55265.0 141700.0 55970.0 140355.0 ;
      RECT  55265.0 141700.0 55970.0 143045.0 ;
      RECT  55265.0 144390.0 55970.0 143045.0 ;
      RECT  55265.0 144390.0 55970.0 145735.0 ;
      RECT  55265.0 147080.0 55970.0 145735.0 ;
      RECT  55265.0 147080.0 55970.0 148425.0 ;
      RECT  55265.0 149770.0 55970.0 148425.0 ;
      RECT  55265.0 149770.0 55970.0 151115.0 ;
      RECT  55265.0 152460.0 55970.0 151115.0 ;
      RECT  55265.0 152460.0 55970.0 153805.0 ;
      RECT  55265.0 155150.0 55970.0 153805.0 ;
      RECT  55265.0 155150.0 55970.0 156495.0 ;
      RECT  55265.0 157840.0 55970.0 156495.0 ;
      RECT  55265.0 157840.0 55970.0 159185.0 ;
      RECT  55265.0 160530.0 55970.0 159185.0 ;
      RECT  55265.0 160530.0 55970.0 161875.0 ;
      RECT  55265.0 163220.0 55970.0 161875.0 ;
      RECT  55265.0 163220.0 55970.0 164565.0 ;
      RECT  55265.0 165910.0 55970.0 164565.0 ;
      RECT  55265.0 165910.0 55970.0 167255.0 ;
      RECT  55265.0 168600.0 55970.0 167255.0 ;
      RECT  55265.0 168600.0 55970.0 169945.0 ;
      RECT  55265.0 171290.0 55970.0 169945.0 ;
      RECT  55265.0 171290.0 55970.0 172635.0 ;
      RECT  55265.0 173980.0 55970.0 172635.0 ;
      RECT  55265.0 173980.0 55970.0 175325.0 ;
      RECT  55265.0 176670.0 55970.0 175325.0 ;
      RECT  55265.0 176670.0 55970.0 178015.0 ;
      RECT  55265.0 179360.0 55970.0 178015.0 ;
      RECT  55265.0 179360.0 55970.0 180705.0 ;
      RECT  55265.0 182050.0 55970.0 180705.0 ;
      RECT  55265.0 182050.0 55970.0 183395.0 ;
      RECT  55265.0 184740.0 55970.0 183395.0 ;
      RECT  55265.0 184740.0 55970.0 186085.0 ;
      RECT  55265.0 187430.0 55970.0 186085.0 ;
      RECT  55265.0 187430.0 55970.0 188775.0 ;
      RECT  55265.0 190120.0 55970.0 188775.0 ;
      RECT  55265.0 190120.0 55970.0 191465.0 ;
      RECT  55265.0 192810.0 55970.0 191465.0 ;
      RECT  55265.0 192810.0 55970.0 194155.0 ;
      RECT  55265.0 195500.0 55970.0 194155.0 ;
      RECT  55265.0 195500.0 55970.0 196845.0 ;
      RECT  55265.0 198190.0 55970.0 196845.0 ;
      RECT  55265.0 198190.0 55970.0 199535.0 ;
      RECT  55265.0 200880.0 55970.0 199535.0 ;
      RECT  55265.0 200880.0 55970.0 202225.0 ;
      RECT  55265.0 203570.0 55970.0 202225.0 ;
      RECT  55265.0 203570.0 55970.0 204915.0 ;
      RECT  55265.0 206260.0 55970.0 204915.0 ;
      RECT  55970.0 34100.0 56675.0 35445.0 ;
      RECT  55970.0 36790.0 56675.0 35445.0 ;
      RECT  55970.0 36790.0 56675.0 38135.0 ;
      RECT  55970.0 39480.0 56675.0 38135.0 ;
      RECT  55970.0 39480.0 56675.0 40825.0 ;
      RECT  55970.0 42170.0 56675.0 40825.0 ;
      RECT  55970.0 42170.0 56675.0 43515.0 ;
      RECT  55970.0 44860.0 56675.0 43515.0 ;
      RECT  55970.0 44860.0 56675.0 46205.0 ;
      RECT  55970.0 47550.0 56675.0 46205.0 ;
      RECT  55970.0 47550.0 56675.0 48895.0 ;
      RECT  55970.0 50240.0 56675.0 48895.0 ;
      RECT  55970.0 50240.0 56675.0 51585.0 ;
      RECT  55970.0 52930.0 56675.0 51585.0 ;
      RECT  55970.0 52930.0 56675.0 54275.0 ;
      RECT  55970.0 55620.0 56675.0 54275.0 ;
      RECT  55970.0 55620.0 56675.0 56965.0 ;
      RECT  55970.0 58310.0 56675.0 56965.0 ;
      RECT  55970.0 58310.0 56675.0 59655.0 ;
      RECT  55970.0 61000.0 56675.0 59655.0 ;
      RECT  55970.0 61000.0 56675.0 62345.0 ;
      RECT  55970.0 63690.0 56675.0 62345.0 ;
      RECT  55970.0 63690.0 56675.0 65035.0 ;
      RECT  55970.0 66380.0 56675.0 65035.0 ;
      RECT  55970.0 66380.0 56675.0 67725.0 ;
      RECT  55970.0 69070.0 56675.0 67725.0 ;
      RECT  55970.0 69070.0 56675.0 70415.0 ;
      RECT  55970.0 71760.0 56675.0 70415.0 ;
      RECT  55970.0 71760.0 56675.0 73105.0 ;
      RECT  55970.0 74450.0 56675.0 73105.0 ;
      RECT  55970.0 74450.0 56675.0 75795.0 ;
      RECT  55970.0 77140.0 56675.0 75795.0 ;
      RECT  55970.0 77140.0 56675.0 78485.0 ;
      RECT  55970.0 79830.0 56675.0 78485.0 ;
      RECT  55970.0 79830.0 56675.0 81175.0 ;
      RECT  55970.0 82520.0 56675.0 81175.0 ;
      RECT  55970.0 82520.0 56675.0 83865.0 ;
      RECT  55970.0 85210.0 56675.0 83865.0 ;
      RECT  55970.0 85210.0 56675.0 86555.0 ;
      RECT  55970.0 87900.0 56675.0 86555.0 ;
      RECT  55970.0 87900.0 56675.0 89245.0 ;
      RECT  55970.0 90590.0 56675.0 89245.0 ;
      RECT  55970.0 90590.0 56675.0 91935.0 ;
      RECT  55970.0 93280.0 56675.0 91935.0 ;
      RECT  55970.0 93280.0 56675.0 94625.0 ;
      RECT  55970.0 95970.0 56675.0 94625.0 ;
      RECT  55970.0 95970.0 56675.0 97315.0 ;
      RECT  55970.0 98660.0 56675.0 97315.0 ;
      RECT  55970.0 98660.0 56675.0 100005.0 ;
      RECT  55970.0 101350.0 56675.0 100005.0 ;
      RECT  55970.0 101350.0 56675.0 102695.0 ;
      RECT  55970.0 104040.0 56675.0 102695.0 ;
      RECT  55970.0 104040.0 56675.0 105385.0 ;
      RECT  55970.0 106730.0 56675.0 105385.0 ;
      RECT  55970.0 106730.0 56675.0 108075.0 ;
      RECT  55970.0 109420.0 56675.0 108075.0 ;
      RECT  55970.0 109420.0 56675.0 110765.0 ;
      RECT  55970.0 112110.0 56675.0 110765.0 ;
      RECT  55970.0 112110.0 56675.0 113455.0 ;
      RECT  55970.0 114800.0 56675.0 113455.0 ;
      RECT  55970.0 114800.0 56675.0 116145.0 ;
      RECT  55970.0 117490.0 56675.0 116145.0 ;
      RECT  55970.0 117490.0 56675.0 118835.0 ;
      RECT  55970.0 120180.0 56675.0 118835.0 ;
      RECT  55970.0 120180.0 56675.0 121525.0 ;
      RECT  55970.0 122870.0 56675.0 121525.0 ;
      RECT  55970.0 122870.0 56675.0 124215.0 ;
      RECT  55970.0 125560.0 56675.0 124215.0 ;
      RECT  55970.0 125560.0 56675.0 126905.0 ;
      RECT  55970.0 128250.0 56675.0 126905.0 ;
      RECT  55970.0 128250.0 56675.0 129595.0 ;
      RECT  55970.0 130940.0 56675.0 129595.0 ;
      RECT  55970.0 130940.0 56675.0 132285.0 ;
      RECT  55970.0 133630.0 56675.0 132285.0 ;
      RECT  55970.0 133630.0 56675.0 134975.0 ;
      RECT  55970.0 136320.0 56675.0 134975.0 ;
      RECT  55970.0 136320.0 56675.0 137665.0 ;
      RECT  55970.0 139010.0 56675.0 137665.0 ;
      RECT  55970.0 139010.0 56675.0 140355.0 ;
      RECT  55970.0 141700.0 56675.0 140355.0 ;
      RECT  55970.0 141700.0 56675.0 143045.0 ;
      RECT  55970.0 144390.0 56675.0 143045.0 ;
      RECT  55970.0 144390.0 56675.0 145735.0 ;
      RECT  55970.0 147080.0 56675.0 145735.0 ;
      RECT  55970.0 147080.0 56675.0 148425.0 ;
      RECT  55970.0 149770.0 56675.0 148425.0 ;
      RECT  55970.0 149770.0 56675.0 151115.0 ;
      RECT  55970.0 152460.0 56675.0 151115.0 ;
      RECT  55970.0 152460.0 56675.0 153805.0 ;
      RECT  55970.0 155150.0 56675.0 153805.0 ;
      RECT  55970.0 155150.0 56675.0 156495.0 ;
      RECT  55970.0 157840.0 56675.0 156495.0 ;
      RECT  55970.0 157840.0 56675.0 159185.0 ;
      RECT  55970.0 160530.0 56675.0 159185.0 ;
      RECT  55970.0 160530.0 56675.0 161875.0 ;
      RECT  55970.0 163220.0 56675.0 161875.0 ;
      RECT  55970.0 163220.0 56675.0 164565.0 ;
      RECT  55970.0 165910.0 56675.0 164565.0 ;
      RECT  55970.0 165910.0 56675.0 167255.0 ;
      RECT  55970.0 168600.0 56675.0 167255.0 ;
      RECT  55970.0 168600.0 56675.0 169945.0 ;
      RECT  55970.0 171290.0 56675.0 169945.0 ;
      RECT  55970.0 171290.0 56675.0 172635.0 ;
      RECT  55970.0 173980.0 56675.0 172635.0 ;
      RECT  55970.0 173980.0 56675.0 175325.0 ;
      RECT  55970.0 176670.0 56675.0 175325.0 ;
      RECT  55970.0 176670.0 56675.0 178015.0 ;
      RECT  55970.0 179360.0 56675.0 178015.0 ;
      RECT  55970.0 179360.0 56675.0 180705.0 ;
      RECT  55970.0 182050.0 56675.0 180705.0 ;
      RECT  55970.0 182050.0 56675.0 183395.0 ;
      RECT  55970.0 184740.0 56675.0 183395.0 ;
      RECT  55970.0 184740.0 56675.0 186085.0 ;
      RECT  55970.0 187430.0 56675.0 186085.0 ;
      RECT  55970.0 187430.0 56675.0 188775.0 ;
      RECT  55970.0 190120.0 56675.0 188775.0 ;
      RECT  55970.0 190120.0 56675.0 191465.0 ;
      RECT  55970.0 192810.0 56675.0 191465.0 ;
      RECT  55970.0 192810.0 56675.0 194155.0 ;
      RECT  55970.0 195500.0 56675.0 194155.0 ;
      RECT  55970.0 195500.0 56675.0 196845.0 ;
      RECT  55970.0 198190.0 56675.0 196845.0 ;
      RECT  55970.0 198190.0 56675.0 199535.0 ;
      RECT  55970.0 200880.0 56675.0 199535.0 ;
      RECT  55970.0 200880.0 56675.0 202225.0 ;
      RECT  55970.0 203570.0 56675.0 202225.0 ;
      RECT  55970.0 203570.0 56675.0 204915.0 ;
      RECT  55970.0 206260.0 56675.0 204915.0 ;
      RECT  56675.0 34100.0 57380.0 35445.0 ;
      RECT  56675.0 36790.0 57380.0 35445.0 ;
      RECT  56675.0 36790.0 57380.0 38135.0 ;
      RECT  56675.0 39480.0 57380.0 38135.0 ;
      RECT  56675.0 39480.0 57380.0 40825.0 ;
      RECT  56675.0 42170.0 57380.0 40825.0 ;
      RECT  56675.0 42170.0 57380.0 43515.0 ;
      RECT  56675.0 44860.0 57380.0 43515.0 ;
      RECT  56675.0 44860.0 57380.0 46205.0 ;
      RECT  56675.0 47550.0 57380.0 46205.0 ;
      RECT  56675.0 47550.0 57380.0 48895.0 ;
      RECT  56675.0 50240.0 57380.0 48895.0 ;
      RECT  56675.0 50240.0 57380.0 51585.0 ;
      RECT  56675.0 52930.0 57380.0 51585.0 ;
      RECT  56675.0 52930.0 57380.0 54275.0 ;
      RECT  56675.0 55620.0 57380.0 54275.0 ;
      RECT  56675.0 55620.0 57380.0 56965.0 ;
      RECT  56675.0 58310.0 57380.0 56965.0 ;
      RECT  56675.0 58310.0 57380.0 59655.0 ;
      RECT  56675.0 61000.0 57380.0 59655.0 ;
      RECT  56675.0 61000.0 57380.0 62345.0 ;
      RECT  56675.0 63690.0 57380.0 62345.0 ;
      RECT  56675.0 63690.0 57380.0 65035.0 ;
      RECT  56675.0 66380.0 57380.0 65035.0 ;
      RECT  56675.0 66380.0 57380.0 67725.0 ;
      RECT  56675.0 69070.0 57380.0 67725.0 ;
      RECT  56675.0 69070.0 57380.0 70415.0 ;
      RECT  56675.0 71760.0 57380.0 70415.0 ;
      RECT  56675.0 71760.0 57380.0 73105.0 ;
      RECT  56675.0 74450.0 57380.0 73105.0 ;
      RECT  56675.0 74450.0 57380.0 75795.0 ;
      RECT  56675.0 77140.0 57380.0 75795.0 ;
      RECT  56675.0 77140.0 57380.0 78485.0 ;
      RECT  56675.0 79830.0 57380.0 78485.0 ;
      RECT  56675.0 79830.0 57380.0 81175.0 ;
      RECT  56675.0 82520.0 57380.0 81175.0 ;
      RECT  56675.0 82520.0 57380.0 83865.0 ;
      RECT  56675.0 85210.0 57380.0 83865.0 ;
      RECT  56675.0 85210.0 57380.0 86555.0 ;
      RECT  56675.0 87900.0 57380.0 86555.0 ;
      RECT  56675.0 87900.0 57380.0 89245.0 ;
      RECT  56675.0 90590.0 57380.0 89245.0 ;
      RECT  56675.0 90590.0 57380.0 91935.0 ;
      RECT  56675.0 93280.0 57380.0 91935.0 ;
      RECT  56675.0 93280.0 57380.0 94625.0 ;
      RECT  56675.0 95970.0 57380.0 94625.0 ;
      RECT  56675.0 95970.0 57380.0 97315.0 ;
      RECT  56675.0 98660.0 57380.0 97315.0 ;
      RECT  56675.0 98660.0 57380.0 100005.0 ;
      RECT  56675.0 101350.0 57380.0 100005.0 ;
      RECT  56675.0 101350.0 57380.0 102695.0 ;
      RECT  56675.0 104040.0 57380.0 102695.0 ;
      RECT  56675.0 104040.0 57380.0 105385.0 ;
      RECT  56675.0 106730.0 57380.0 105385.0 ;
      RECT  56675.0 106730.0 57380.0 108075.0 ;
      RECT  56675.0 109420.0 57380.0 108075.0 ;
      RECT  56675.0 109420.0 57380.0 110765.0 ;
      RECT  56675.0 112110.0 57380.0 110765.0 ;
      RECT  56675.0 112110.0 57380.0 113455.0 ;
      RECT  56675.0 114800.0 57380.0 113455.0 ;
      RECT  56675.0 114800.0 57380.0 116145.0 ;
      RECT  56675.0 117490.0 57380.0 116145.0 ;
      RECT  56675.0 117490.0 57380.0 118835.0 ;
      RECT  56675.0 120180.0 57380.0 118835.0 ;
      RECT  56675.0 120180.0 57380.0 121525.0 ;
      RECT  56675.0 122870.0 57380.0 121525.0 ;
      RECT  56675.0 122870.0 57380.0 124215.0 ;
      RECT  56675.0 125560.0 57380.0 124215.0 ;
      RECT  56675.0 125560.0 57380.0 126905.0 ;
      RECT  56675.0 128250.0 57380.0 126905.0 ;
      RECT  56675.0 128250.0 57380.0 129595.0 ;
      RECT  56675.0 130940.0 57380.0 129595.0 ;
      RECT  56675.0 130940.0 57380.0 132285.0 ;
      RECT  56675.0 133630.0 57380.0 132285.0 ;
      RECT  56675.0 133630.0 57380.0 134975.0 ;
      RECT  56675.0 136320.0 57380.0 134975.0 ;
      RECT  56675.0 136320.0 57380.0 137665.0 ;
      RECT  56675.0 139010.0 57380.0 137665.0 ;
      RECT  56675.0 139010.0 57380.0 140355.0 ;
      RECT  56675.0 141700.0 57380.0 140355.0 ;
      RECT  56675.0 141700.0 57380.0 143045.0 ;
      RECT  56675.0 144390.0 57380.0 143045.0 ;
      RECT  56675.0 144390.0 57380.0 145735.0 ;
      RECT  56675.0 147080.0 57380.0 145735.0 ;
      RECT  56675.0 147080.0 57380.0 148425.0 ;
      RECT  56675.0 149770.0 57380.0 148425.0 ;
      RECT  56675.0 149770.0 57380.0 151115.0 ;
      RECT  56675.0 152460.0 57380.0 151115.0 ;
      RECT  56675.0 152460.0 57380.0 153805.0 ;
      RECT  56675.0 155150.0 57380.0 153805.0 ;
      RECT  56675.0 155150.0 57380.0 156495.0 ;
      RECT  56675.0 157840.0 57380.0 156495.0 ;
      RECT  56675.0 157840.0 57380.0 159185.0 ;
      RECT  56675.0 160530.0 57380.0 159185.0 ;
      RECT  56675.0 160530.0 57380.0 161875.0 ;
      RECT  56675.0 163220.0 57380.0 161875.0 ;
      RECT  56675.0 163220.0 57380.0 164565.0 ;
      RECT  56675.0 165910.0 57380.0 164565.0 ;
      RECT  56675.0 165910.0 57380.0 167255.0 ;
      RECT  56675.0 168600.0 57380.0 167255.0 ;
      RECT  56675.0 168600.0 57380.0 169945.0 ;
      RECT  56675.0 171290.0 57380.0 169945.0 ;
      RECT  56675.0 171290.0 57380.0 172635.0 ;
      RECT  56675.0 173980.0 57380.0 172635.0 ;
      RECT  56675.0 173980.0 57380.0 175325.0 ;
      RECT  56675.0 176670.0 57380.0 175325.0 ;
      RECT  56675.0 176670.0 57380.0 178015.0 ;
      RECT  56675.0 179360.0 57380.0 178015.0 ;
      RECT  56675.0 179360.0 57380.0 180705.0 ;
      RECT  56675.0 182050.0 57380.0 180705.0 ;
      RECT  56675.0 182050.0 57380.0 183395.0 ;
      RECT  56675.0 184740.0 57380.0 183395.0 ;
      RECT  56675.0 184740.0 57380.0 186085.0 ;
      RECT  56675.0 187430.0 57380.0 186085.0 ;
      RECT  56675.0 187430.0 57380.0 188775.0 ;
      RECT  56675.0 190120.0 57380.0 188775.0 ;
      RECT  56675.0 190120.0 57380.0 191465.0 ;
      RECT  56675.0 192810.0 57380.0 191465.0 ;
      RECT  56675.0 192810.0 57380.0 194155.0 ;
      RECT  56675.0 195500.0 57380.0 194155.0 ;
      RECT  56675.0 195500.0 57380.0 196845.0 ;
      RECT  56675.0 198190.0 57380.0 196845.0 ;
      RECT  56675.0 198190.0 57380.0 199535.0 ;
      RECT  56675.0 200880.0 57380.0 199535.0 ;
      RECT  56675.0 200880.0 57380.0 202225.0 ;
      RECT  56675.0 203570.0 57380.0 202225.0 ;
      RECT  56675.0 203570.0 57380.0 204915.0 ;
      RECT  56675.0 206260.0 57380.0 204915.0 ;
      RECT  57380.0 34100.0 58085.0 35445.0 ;
      RECT  57380.0 36790.0 58085.0 35445.0 ;
      RECT  57380.0 36790.0 58085.0 38135.0 ;
      RECT  57380.0 39480.0 58085.0 38135.0 ;
      RECT  57380.0 39480.0 58085.0 40825.0 ;
      RECT  57380.0 42170.0 58085.0 40825.0 ;
      RECT  57380.0 42170.0 58085.0 43515.0 ;
      RECT  57380.0 44860.0 58085.0 43515.0 ;
      RECT  57380.0 44860.0 58085.0 46205.0 ;
      RECT  57380.0 47550.0 58085.0 46205.0 ;
      RECT  57380.0 47550.0 58085.0 48895.0 ;
      RECT  57380.0 50240.0 58085.0 48895.0 ;
      RECT  57380.0 50240.0 58085.0 51585.0 ;
      RECT  57380.0 52930.0 58085.0 51585.0 ;
      RECT  57380.0 52930.0 58085.0 54275.0 ;
      RECT  57380.0 55620.0 58085.0 54275.0 ;
      RECT  57380.0 55620.0 58085.0 56965.0 ;
      RECT  57380.0 58310.0 58085.0 56965.0 ;
      RECT  57380.0 58310.0 58085.0 59655.0 ;
      RECT  57380.0 61000.0 58085.0 59655.0 ;
      RECT  57380.0 61000.0 58085.0 62345.0 ;
      RECT  57380.0 63690.0 58085.0 62345.0 ;
      RECT  57380.0 63690.0 58085.0 65035.0 ;
      RECT  57380.0 66380.0 58085.0 65035.0 ;
      RECT  57380.0 66380.0 58085.0 67725.0 ;
      RECT  57380.0 69070.0 58085.0 67725.0 ;
      RECT  57380.0 69070.0 58085.0 70415.0 ;
      RECT  57380.0 71760.0 58085.0 70415.0 ;
      RECT  57380.0 71760.0 58085.0 73105.0 ;
      RECT  57380.0 74450.0 58085.0 73105.0 ;
      RECT  57380.0 74450.0 58085.0 75795.0 ;
      RECT  57380.0 77140.0 58085.0 75795.0 ;
      RECT  57380.0 77140.0 58085.0 78485.0 ;
      RECT  57380.0 79830.0 58085.0 78485.0 ;
      RECT  57380.0 79830.0 58085.0 81175.0 ;
      RECT  57380.0 82520.0 58085.0 81175.0 ;
      RECT  57380.0 82520.0 58085.0 83865.0 ;
      RECT  57380.0 85210.0 58085.0 83865.0 ;
      RECT  57380.0 85210.0 58085.0 86555.0 ;
      RECT  57380.0 87900.0 58085.0 86555.0 ;
      RECT  57380.0 87900.0 58085.0 89245.0 ;
      RECT  57380.0 90590.0 58085.0 89245.0 ;
      RECT  57380.0 90590.0 58085.0 91935.0 ;
      RECT  57380.0 93280.0 58085.0 91935.0 ;
      RECT  57380.0 93280.0 58085.0 94625.0 ;
      RECT  57380.0 95970.0 58085.0 94625.0 ;
      RECT  57380.0 95970.0 58085.0 97315.0 ;
      RECT  57380.0 98660.0 58085.0 97315.0 ;
      RECT  57380.0 98660.0 58085.0 100005.0 ;
      RECT  57380.0 101350.0 58085.0 100005.0 ;
      RECT  57380.0 101350.0 58085.0 102695.0 ;
      RECT  57380.0 104040.0 58085.0 102695.0 ;
      RECT  57380.0 104040.0 58085.0 105385.0 ;
      RECT  57380.0 106730.0 58085.0 105385.0 ;
      RECT  57380.0 106730.0 58085.0 108075.0 ;
      RECT  57380.0 109420.0 58085.0 108075.0 ;
      RECT  57380.0 109420.0 58085.0 110765.0 ;
      RECT  57380.0 112110.0 58085.0 110765.0 ;
      RECT  57380.0 112110.0 58085.0 113455.0 ;
      RECT  57380.0 114800.0 58085.0 113455.0 ;
      RECT  57380.0 114800.0 58085.0 116145.0 ;
      RECT  57380.0 117490.0 58085.0 116145.0 ;
      RECT  57380.0 117490.0 58085.0 118835.0 ;
      RECT  57380.0 120180.0 58085.0 118835.0 ;
      RECT  57380.0 120180.0 58085.0 121525.0 ;
      RECT  57380.0 122870.0 58085.0 121525.0 ;
      RECT  57380.0 122870.0 58085.0 124215.0 ;
      RECT  57380.0 125560.0 58085.0 124215.0 ;
      RECT  57380.0 125560.0 58085.0 126905.0 ;
      RECT  57380.0 128250.0 58085.0 126905.0 ;
      RECT  57380.0 128250.0 58085.0 129595.0 ;
      RECT  57380.0 130940.0 58085.0 129595.0 ;
      RECT  57380.0 130940.0 58085.0 132285.0 ;
      RECT  57380.0 133630.0 58085.0 132285.0 ;
      RECT  57380.0 133630.0 58085.0 134975.0 ;
      RECT  57380.0 136320.0 58085.0 134975.0 ;
      RECT  57380.0 136320.0 58085.0 137665.0 ;
      RECT  57380.0 139010.0 58085.0 137665.0 ;
      RECT  57380.0 139010.0 58085.0 140355.0 ;
      RECT  57380.0 141700.0 58085.0 140355.0 ;
      RECT  57380.0 141700.0 58085.0 143045.0 ;
      RECT  57380.0 144390.0 58085.0 143045.0 ;
      RECT  57380.0 144390.0 58085.0 145735.0 ;
      RECT  57380.0 147080.0 58085.0 145735.0 ;
      RECT  57380.0 147080.0 58085.0 148425.0 ;
      RECT  57380.0 149770.0 58085.0 148425.0 ;
      RECT  57380.0 149770.0 58085.0 151115.0 ;
      RECT  57380.0 152460.0 58085.0 151115.0 ;
      RECT  57380.0 152460.0 58085.0 153805.0 ;
      RECT  57380.0 155150.0 58085.0 153805.0 ;
      RECT  57380.0 155150.0 58085.0 156495.0 ;
      RECT  57380.0 157840.0 58085.0 156495.0 ;
      RECT  57380.0 157840.0 58085.0 159185.0 ;
      RECT  57380.0 160530.0 58085.0 159185.0 ;
      RECT  57380.0 160530.0 58085.0 161875.0 ;
      RECT  57380.0 163220.0 58085.0 161875.0 ;
      RECT  57380.0 163220.0 58085.0 164565.0 ;
      RECT  57380.0 165910.0 58085.0 164565.0 ;
      RECT  57380.0 165910.0 58085.0 167255.0 ;
      RECT  57380.0 168600.0 58085.0 167255.0 ;
      RECT  57380.0 168600.0 58085.0 169945.0 ;
      RECT  57380.0 171290.0 58085.0 169945.0 ;
      RECT  57380.0 171290.0 58085.0 172635.0 ;
      RECT  57380.0 173980.0 58085.0 172635.0 ;
      RECT  57380.0 173980.0 58085.0 175325.0 ;
      RECT  57380.0 176670.0 58085.0 175325.0 ;
      RECT  57380.0 176670.0 58085.0 178015.0 ;
      RECT  57380.0 179360.0 58085.0 178015.0 ;
      RECT  57380.0 179360.0 58085.0 180705.0 ;
      RECT  57380.0 182050.0 58085.0 180705.0 ;
      RECT  57380.0 182050.0 58085.0 183395.0 ;
      RECT  57380.0 184740.0 58085.0 183395.0 ;
      RECT  57380.0 184740.0 58085.0 186085.0 ;
      RECT  57380.0 187430.0 58085.0 186085.0 ;
      RECT  57380.0 187430.0 58085.0 188775.0 ;
      RECT  57380.0 190120.0 58085.0 188775.0 ;
      RECT  57380.0 190120.0 58085.0 191465.0 ;
      RECT  57380.0 192810.0 58085.0 191465.0 ;
      RECT  57380.0 192810.0 58085.0 194155.0 ;
      RECT  57380.0 195500.0 58085.0 194155.0 ;
      RECT  57380.0 195500.0 58085.0 196845.0 ;
      RECT  57380.0 198190.0 58085.0 196845.0 ;
      RECT  57380.0 198190.0 58085.0 199535.0 ;
      RECT  57380.0 200880.0 58085.0 199535.0 ;
      RECT  57380.0 200880.0 58085.0 202225.0 ;
      RECT  57380.0 203570.0 58085.0 202225.0 ;
      RECT  57380.0 203570.0 58085.0 204915.0 ;
      RECT  57380.0 206260.0 58085.0 204915.0 ;
      RECT  58085.0 34100.0 58790.0 35445.0 ;
      RECT  58085.0 36790.0 58790.0 35445.0 ;
      RECT  58085.0 36790.0 58790.0 38135.0 ;
      RECT  58085.0 39480.0 58790.0 38135.0 ;
      RECT  58085.0 39480.0 58790.0 40825.0 ;
      RECT  58085.0 42170.0 58790.0 40825.0 ;
      RECT  58085.0 42170.0 58790.0 43515.0 ;
      RECT  58085.0 44860.0 58790.0 43515.0 ;
      RECT  58085.0 44860.0 58790.0 46205.0 ;
      RECT  58085.0 47550.0 58790.0 46205.0 ;
      RECT  58085.0 47550.0 58790.0 48895.0 ;
      RECT  58085.0 50240.0 58790.0 48895.0 ;
      RECT  58085.0 50240.0 58790.0 51585.0 ;
      RECT  58085.0 52930.0 58790.0 51585.0 ;
      RECT  58085.0 52930.0 58790.0 54275.0 ;
      RECT  58085.0 55620.0 58790.0 54275.0 ;
      RECT  58085.0 55620.0 58790.0 56965.0 ;
      RECT  58085.0 58310.0 58790.0 56965.0 ;
      RECT  58085.0 58310.0 58790.0 59655.0 ;
      RECT  58085.0 61000.0 58790.0 59655.0 ;
      RECT  58085.0 61000.0 58790.0 62345.0 ;
      RECT  58085.0 63690.0 58790.0 62345.0 ;
      RECT  58085.0 63690.0 58790.0 65035.0 ;
      RECT  58085.0 66380.0 58790.0 65035.0 ;
      RECT  58085.0 66380.0 58790.0 67725.0 ;
      RECT  58085.0 69070.0 58790.0 67725.0 ;
      RECT  58085.0 69070.0 58790.0 70415.0 ;
      RECT  58085.0 71760.0 58790.0 70415.0 ;
      RECT  58085.0 71760.0 58790.0 73105.0 ;
      RECT  58085.0 74450.0 58790.0 73105.0 ;
      RECT  58085.0 74450.0 58790.0 75795.0 ;
      RECT  58085.0 77140.0 58790.0 75795.0 ;
      RECT  58085.0 77140.0 58790.0 78485.0 ;
      RECT  58085.0 79830.0 58790.0 78485.0 ;
      RECT  58085.0 79830.0 58790.0 81175.0 ;
      RECT  58085.0 82520.0 58790.0 81175.0 ;
      RECT  58085.0 82520.0 58790.0 83865.0 ;
      RECT  58085.0 85210.0 58790.0 83865.0 ;
      RECT  58085.0 85210.0 58790.0 86555.0 ;
      RECT  58085.0 87900.0 58790.0 86555.0 ;
      RECT  58085.0 87900.0 58790.0 89245.0 ;
      RECT  58085.0 90590.0 58790.0 89245.0 ;
      RECT  58085.0 90590.0 58790.0 91935.0 ;
      RECT  58085.0 93280.0 58790.0 91935.0 ;
      RECT  58085.0 93280.0 58790.0 94625.0 ;
      RECT  58085.0 95970.0 58790.0 94625.0 ;
      RECT  58085.0 95970.0 58790.0 97315.0 ;
      RECT  58085.0 98660.0 58790.0 97315.0 ;
      RECT  58085.0 98660.0 58790.0 100005.0 ;
      RECT  58085.0 101350.0 58790.0 100005.0 ;
      RECT  58085.0 101350.0 58790.0 102695.0 ;
      RECT  58085.0 104040.0 58790.0 102695.0 ;
      RECT  58085.0 104040.0 58790.0 105385.0 ;
      RECT  58085.0 106730.0 58790.0 105385.0 ;
      RECT  58085.0 106730.0 58790.0 108075.0 ;
      RECT  58085.0 109420.0 58790.0 108075.0 ;
      RECT  58085.0 109420.0 58790.0 110765.0 ;
      RECT  58085.0 112110.0 58790.0 110765.0 ;
      RECT  58085.0 112110.0 58790.0 113455.0 ;
      RECT  58085.0 114800.0 58790.0 113455.0 ;
      RECT  58085.0 114800.0 58790.0 116145.0 ;
      RECT  58085.0 117490.0 58790.0 116145.0 ;
      RECT  58085.0 117490.0 58790.0 118835.0 ;
      RECT  58085.0 120180.0 58790.0 118835.0 ;
      RECT  58085.0 120180.0 58790.0 121525.0 ;
      RECT  58085.0 122870.0 58790.0 121525.0 ;
      RECT  58085.0 122870.0 58790.0 124215.0 ;
      RECT  58085.0 125560.0 58790.0 124215.0 ;
      RECT  58085.0 125560.0 58790.0 126905.0 ;
      RECT  58085.0 128250.0 58790.0 126905.0 ;
      RECT  58085.0 128250.0 58790.0 129595.0 ;
      RECT  58085.0 130940.0 58790.0 129595.0 ;
      RECT  58085.0 130940.0 58790.0 132285.0 ;
      RECT  58085.0 133630.0 58790.0 132285.0 ;
      RECT  58085.0 133630.0 58790.0 134975.0 ;
      RECT  58085.0 136320.0 58790.0 134975.0 ;
      RECT  58085.0 136320.0 58790.0 137665.0 ;
      RECT  58085.0 139010.0 58790.0 137665.0 ;
      RECT  58085.0 139010.0 58790.0 140355.0 ;
      RECT  58085.0 141700.0 58790.0 140355.0 ;
      RECT  58085.0 141700.0 58790.0 143045.0 ;
      RECT  58085.0 144390.0 58790.0 143045.0 ;
      RECT  58085.0 144390.0 58790.0 145735.0 ;
      RECT  58085.0 147080.0 58790.0 145735.0 ;
      RECT  58085.0 147080.0 58790.0 148425.0 ;
      RECT  58085.0 149770.0 58790.0 148425.0 ;
      RECT  58085.0 149770.0 58790.0 151115.0 ;
      RECT  58085.0 152460.0 58790.0 151115.0 ;
      RECT  58085.0 152460.0 58790.0 153805.0 ;
      RECT  58085.0 155150.0 58790.0 153805.0 ;
      RECT  58085.0 155150.0 58790.0 156495.0 ;
      RECT  58085.0 157840.0 58790.0 156495.0 ;
      RECT  58085.0 157840.0 58790.0 159185.0 ;
      RECT  58085.0 160530.0 58790.0 159185.0 ;
      RECT  58085.0 160530.0 58790.0 161875.0 ;
      RECT  58085.0 163220.0 58790.0 161875.0 ;
      RECT  58085.0 163220.0 58790.0 164565.0 ;
      RECT  58085.0 165910.0 58790.0 164565.0 ;
      RECT  58085.0 165910.0 58790.0 167255.0 ;
      RECT  58085.0 168600.0 58790.0 167255.0 ;
      RECT  58085.0 168600.0 58790.0 169945.0 ;
      RECT  58085.0 171290.0 58790.0 169945.0 ;
      RECT  58085.0 171290.0 58790.0 172635.0 ;
      RECT  58085.0 173980.0 58790.0 172635.0 ;
      RECT  58085.0 173980.0 58790.0 175325.0 ;
      RECT  58085.0 176670.0 58790.0 175325.0 ;
      RECT  58085.0 176670.0 58790.0 178015.0 ;
      RECT  58085.0 179360.0 58790.0 178015.0 ;
      RECT  58085.0 179360.0 58790.0 180705.0 ;
      RECT  58085.0 182050.0 58790.0 180705.0 ;
      RECT  58085.0 182050.0 58790.0 183395.0 ;
      RECT  58085.0 184740.0 58790.0 183395.0 ;
      RECT  58085.0 184740.0 58790.0 186085.0 ;
      RECT  58085.0 187430.0 58790.0 186085.0 ;
      RECT  58085.0 187430.0 58790.0 188775.0 ;
      RECT  58085.0 190120.0 58790.0 188775.0 ;
      RECT  58085.0 190120.0 58790.0 191465.0 ;
      RECT  58085.0 192810.0 58790.0 191465.0 ;
      RECT  58085.0 192810.0 58790.0 194155.0 ;
      RECT  58085.0 195500.0 58790.0 194155.0 ;
      RECT  58085.0 195500.0 58790.0 196845.0 ;
      RECT  58085.0 198190.0 58790.0 196845.0 ;
      RECT  58085.0 198190.0 58790.0 199535.0 ;
      RECT  58085.0 200880.0 58790.0 199535.0 ;
      RECT  58085.0 200880.0 58790.0 202225.0 ;
      RECT  58085.0 203570.0 58790.0 202225.0 ;
      RECT  58085.0 203570.0 58790.0 204915.0 ;
      RECT  58085.0 206260.0 58790.0 204915.0 ;
      RECT  58790.0 34100.0 59495.0 35445.0 ;
      RECT  58790.0 36790.0 59495.0 35445.0 ;
      RECT  58790.0 36790.0 59495.0 38135.0 ;
      RECT  58790.0 39480.0 59495.0 38135.0 ;
      RECT  58790.0 39480.0 59495.0 40825.0 ;
      RECT  58790.0 42170.0 59495.0 40825.0 ;
      RECT  58790.0 42170.0 59495.0 43515.0 ;
      RECT  58790.0 44860.0 59495.0 43515.0 ;
      RECT  58790.0 44860.0 59495.0 46205.0 ;
      RECT  58790.0 47550.0 59495.0 46205.0 ;
      RECT  58790.0 47550.0 59495.0 48895.0 ;
      RECT  58790.0 50240.0 59495.0 48895.0 ;
      RECT  58790.0 50240.0 59495.0 51585.0 ;
      RECT  58790.0 52930.0 59495.0 51585.0 ;
      RECT  58790.0 52930.0 59495.0 54275.0 ;
      RECT  58790.0 55620.0 59495.0 54275.0 ;
      RECT  58790.0 55620.0 59495.0 56965.0 ;
      RECT  58790.0 58310.0 59495.0 56965.0 ;
      RECT  58790.0 58310.0 59495.0 59655.0 ;
      RECT  58790.0 61000.0 59495.0 59655.0 ;
      RECT  58790.0 61000.0 59495.0 62345.0 ;
      RECT  58790.0 63690.0 59495.0 62345.0 ;
      RECT  58790.0 63690.0 59495.0 65035.0 ;
      RECT  58790.0 66380.0 59495.0 65035.0 ;
      RECT  58790.0 66380.0 59495.0 67725.0 ;
      RECT  58790.0 69070.0 59495.0 67725.0 ;
      RECT  58790.0 69070.0 59495.0 70415.0 ;
      RECT  58790.0 71760.0 59495.0 70415.0 ;
      RECT  58790.0 71760.0 59495.0 73105.0 ;
      RECT  58790.0 74450.0 59495.0 73105.0 ;
      RECT  58790.0 74450.0 59495.0 75795.0 ;
      RECT  58790.0 77140.0 59495.0 75795.0 ;
      RECT  58790.0 77140.0 59495.0 78485.0 ;
      RECT  58790.0 79830.0 59495.0 78485.0 ;
      RECT  58790.0 79830.0 59495.0 81175.0 ;
      RECT  58790.0 82520.0 59495.0 81175.0 ;
      RECT  58790.0 82520.0 59495.0 83865.0 ;
      RECT  58790.0 85210.0 59495.0 83865.0 ;
      RECT  58790.0 85210.0 59495.0 86555.0 ;
      RECT  58790.0 87900.0 59495.0 86555.0 ;
      RECT  58790.0 87900.0 59495.0 89245.0 ;
      RECT  58790.0 90590.0 59495.0 89245.0 ;
      RECT  58790.0 90590.0 59495.0 91935.0 ;
      RECT  58790.0 93280.0 59495.0 91935.0 ;
      RECT  58790.0 93280.0 59495.0 94625.0 ;
      RECT  58790.0 95970.0 59495.0 94625.0 ;
      RECT  58790.0 95970.0 59495.0 97315.0 ;
      RECT  58790.0 98660.0 59495.0 97315.0 ;
      RECT  58790.0 98660.0 59495.0 100005.0 ;
      RECT  58790.0 101350.0 59495.0 100005.0 ;
      RECT  58790.0 101350.0 59495.0 102695.0 ;
      RECT  58790.0 104040.0 59495.0 102695.0 ;
      RECT  58790.0 104040.0 59495.0 105385.0 ;
      RECT  58790.0 106730.0 59495.0 105385.0 ;
      RECT  58790.0 106730.0 59495.0 108075.0 ;
      RECT  58790.0 109420.0 59495.0 108075.0 ;
      RECT  58790.0 109420.0 59495.0 110765.0 ;
      RECT  58790.0 112110.0 59495.0 110765.0 ;
      RECT  58790.0 112110.0 59495.0 113455.0 ;
      RECT  58790.0 114800.0 59495.0 113455.0 ;
      RECT  58790.0 114800.0 59495.0 116145.0 ;
      RECT  58790.0 117490.0 59495.0 116145.0 ;
      RECT  58790.0 117490.0 59495.0 118835.0 ;
      RECT  58790.0 120180.0 59495.0 118835.0 ;
      RECT  58790.0 120180.0 59495.0 121525.0 ;
      RECT  58790.0 122870.0 59495.0 121525.0 ;
      RECT  58790.0 122870.0 59495.0 124215.0 ;
      RECT  58790.0 125560.0 59495.0 124215.0 ;
      RECT  58790.0 125560.0 59495.0 126905.0 ;
      RECT  58790.0 128250.0 59495.0 126905.0 ;
      RECT  58790.0 128250.0 59495.0 129595.0 ;
      RECT  58790.0 130940.0 59495.0 129595.0 ;
      RECT  58790.0 130940.0 59495.0 132285.0 ;
      RECT  58790.0 133630.0 59495.0 132285.0 ;
      RECT  58790.0 133630.0 59495.0 134975.0 ;
      RECT  58790.0 136320.0 59495.0 134975.0 ;
      RECT  58790.0 136320.0 59495.0 137665.0 ;
      RECT  58790.0 139010.0 59495.0 137665.0 ;
      RECT  58790.0 139010.0 59495.0 140355.0 ;
      RECT  58790.0 141700.0 59495.0 140355.0 ;
      RECT  58790.0 141700.0 59495.0 143045.0 ;
      RECT  58790.0 144390.0 59495.0 143045.0 ;
      RECT  58790.0 144390.0 59495.0 145735.0 ;
      RECT  58790.0 147080.0 59495.0 145735.0 ;
      RECT  58790.0 147080.0 59495.0 148425.0 ;
      RECT  58790.0 149770.0 59495.0 148425.0 ;
      RECT  58790.0 149770.0 59495.0 151115.0 ;
      RECT  58790.0 152460.0 59495.0 151115.0 ;
      RECT  58790.0 152460.0 59495.0 153805.0 ;
      RECT  58790.0 155150.0 59495.0 153805.0 ;
      RECT  58790.0 155150.0 59495.0 156495.0 ;
      RECT  58790.0 157840.0 59495.0 156495.0 ;
      RECT  58790.0 157840.0 59495.0 159185.0 ;
      RECT  58790.0 160530.0 59495.0 159185.0 ;
      RECT  58790.0 160530.0 59495.0 161875.0 ;
      RECT  58790.0 163220.0 59495.0 161875.0 ;
      RECT  58790.0 163220.0 59495.0 164565.0 ;
      RECT  58790.0 165910.0 59495.0 164565.0 ;
      RECT  58790.0 165910.0 59495.0 167255.0 ;
      RECT  58790.0 168600.0 59495.0 167255.0 ;
      RECT  58790.0 168600.0 59495.0 169945.0 ;
      RECT  58790.0 171290.0 59495.0 169945.0 ;
      RECT  58790.0 171290.0 59495.0 172635.0 ;
      RECT  58790.0 173980.0 59495.0 172635.0 ;
      RECT  58790.0 173980.0 59495.0 175325.0 ;
      RECT  58790.0 176670.0 59495.0 175325.0 ;
      RECT  58790.0 176670.0 59495.0 178015.0 ;
      RECT  58790.0 179360.0 59495.0 178015.0 ;
      RECT  58790.0 179360.0 59495.0 180705.0 ;
      RECT  58790.0 182050.0 59495.0 180705.0 ;
      RECT  58790.0 182050.0 59495.0 183395.0 ;
      RECT  58790.0 184740.0 59495.0 183395.0 ;
      RECT  58790.0 184740.0 59495.0 186085.0 ;
      RECT  58790.0 187430.0 59495.0 186085.0 ;
      RECT  58790.0 187430.0 59495.0 188775.0 ;
      RECT  58790.0 190120.0 59495.0 188775.0 ;
      RECT  58790.0 190120.0 59495.0 191465.0 ;
      RECT  58790.0 192810.0 59495.0 191465.0 ;
      RECT  58790.0 192810.0 59495.0 194155.0 ;
      RECT  58790.0 195500.0 59495.0 194155.0 ;
      RECT  58790.0 195500.0 59495.0 196845.0 ;
      RECT  58790.0 198190.0 59495.0 196845.0 ;
      RECT  58790.0 198190.0 59495.0 199535.0 ;
      RECT  58790.0 200880.0 59495.0 199535.0 ;
      RECT  58790.0 200880.0 59495.0 202225.0 ;
      RECT  58790.0 203570.0 59495.0 202225.0 ;
      RECT  58790.0 203570.0 59495.0 204915.0 ;
      RECT  58790.0 206260.0 59495.0 204915.0 ;
      RECT  59495.0 34100.0 60200.0 35445.0 ;
      RECT  59495.0 36790.0 60200.0 35445.0 ;
      RECT  59495.0 36790.0 60200.0 38135.0 ;
      RECT  59495.0 39480.0 60200.0 38135.0 ;
      RECT  59495.0 39480.0 60200.0 40825.0 ;
      RECT  59495.0 42170.0 60200.0 40825.0 ;
      RECT  59495.0 42170.0 60200.0 43515.0 ;
      RECT  59495.0 44860.0 60200.0 43515.0 ;
      RECT  59495.0 44860.0 60200.0 46205.0 ;
      RECT  59495.0 47550.0 60200.0 46205.0 ;
      RECT  59495.0 47550.0 60200.0 48895.0 ;
      RECT  59495.0 50240.0 60200.0 48895.0 ;
      RECT  59495.0 50240.0 60200.0 51585.0 ;
      RECT  59495.0 52930.0 60200.0 51585.0 ;
      RECT  59495.0 52930.0 60200.0 54275.0 ;
      RECT  59495.0 55620.0 60200.0 54275.0 ;
      RECT  59495.0 55620.0 60200.0 56965.0 ;
      RECT  59495.0 58310.0 60200.0 56965.0 ;
      RECT  59495.0 58310.0 60200.0 59655.0 ;
      RECT  59495.0 61000.0 60200.0 59655.0 ;
      RECT  59495.0 61000.0 60200.0 62345.0 ;
      RECT  59495.0 63690.0 60200.0 62345.0 ;
      RECT  59495.0 63690.0 60200.0 65035.0 ;
      RECT  59495.0 66380.0 60200.0 65035.0 ;
      RECT  59495.0 66380.0 60200.0 67725.0 ;
      RECT  59495.0 69070.0 60200.0 67725.0 ;
      RECT  59495.0 69070.0 60200.0 70415.0 ;
      RECT  59495.0 71760.0 60200.0 70415.0 ;
      RECT  59495.0 71760.0 60200.0 73105.0 ;
      RECT  59495.0 74450.0 60200.0 73105.0 ;
      RECT  59495.0 74450.0 60200.0 75795.0 ;
      RECT  59495.0 77140.0 60200.0 75795.0 ;
      RECT  59495.0 77140.0 60200.0 78485.0 ;
      RECT  59495.0 79830.0 60200.0 78485.0 ;
      RECT  59495.0 79830.0 60200.0 81175.0 ;
      RECT  59495.0 82520.0 60200.0 81175.0 ;
      RECT  59495.0 82520.0 60200.0 83865.0 ;
      RECT  59495.0 85210.0 60200.0 83865.0 ;
      RECT  59495.0 85210.0 60200.0 86555.0 ;
      RECT  59495.0 87900.0 60200.0 86555.0 ;
      RECT  59495.0 87900.0 60200.0 89245.0 ;
      RECT  59495.0 90590.0 60200.0 89245.0 ;
      RECT  59495.0 90590.0 60200.0 91935.0 ;
      RECT  59495.0 93280.0 60200.0 91935.0 ;
      RECT  59495.0 93280.0 60200.0 94625.0 ;
      RECT  59495.0 95970.0 60200.0 94625.0 ;
      RECT  59495.0 95970.0 60200.0 97315.0 ;
      RECT  59495.0 98660.0 60200.0 97315.0 ;
      RECT  59495.0 98660.0 60200.0 100005.0 ;
      RECT  59495.0 101350.0 60200.0 100005.0 ;
      RECT  59495.0 101350.0 60200.0 102695.0 ;
      RECT  59495.0 104040.0 60200.0 102695.0 ;
      RECT  59495.0 104040.0 60200.0 105385.0 ;
      RECT  59495.0 106730.0 60200.0 105385.0 ;
      RECT  59495.0 106730.0 60200.0 108075.0 ;
      RECT  59495.0 109420.0 60200.0 108075.0 ;
      RECT  59495.0 109420.0 60200.0 110765.0 ;
      RECT  59495.0 112110.0 60200.0 110765.0 ;
      RECT  59495.0 112110.0 60200.0 113455.0 ;
      RECT  59495.0 114800.0 60200.0 113455.0 ;
      RECT  59495.0 114800.0 60200.0 116145.0 ;
      RECT  59495.0 117490.0 60200.0 116145.0 ;
      RECT  59495.0 117490.0 60200.0 118835.0 ;
      RECT  59495.0 120180.0 60200.0 118835.0 ;
      RECT  59495.0 120180.0 60200.0 121525.0 ;
      RECT  59495.0 122870.0 60200.0 121525.0 ;
      RECT  59495.0 122870.0 60200.0 124215.0 ;
      RECT  59495.0 125560.0 60200.0 124215.0 ;
      RECT  59495.0 125560.0 60200.0 126905.0 ;
      RECT  59495.0 128250.0 60200.0 126905.0 ;
      RECT  59495.0 128250.0 60200.0 129595.0 ;
      RECT  59495.0 130940.0 60200.0 129595.0 ;
      RECT  59495.0 130940.0 60200.0 132285.0 ;
      RECT  59495.0 133630.0 60200.0 132285.0 ;
      RECT  59495.0 133630.0 60200.0 134975.0 ;
      RECT  59495.0 136320.0 60200.0 134975.0 ;
      RECT  59495.0 136320.0 60200.0 137665.0 ;
      RECT  59495.0 139010.0 60200.0 137665.0 ;
      RECT  59495.0 139010.0 60200.0 140355.0 ;
      RECT  59495.0 141700.0 60200.0 140355.0 ;
      RECT  59495.0 141700.0 60200.0 143045.0 ;
      RECT  59495.0 144390.0 60200.0 143045.0 ;
      RECT  59495.0 144390.0 60200.0 145735.0 ;
      RECT  59495.0 147080.0 60200.0 145735.0 ;
      RECT  59495.0 147080.0 60200.0 148425.0 ;
      RECT  59495.0 149770.0 60200.0 148425.0 ;
      RECT  59495.0 149770.0 60200.0 151115.0 ;
      RECT  59495.0 152460.0 60200.0 151115.0 ;
      RECT  59495.0 152460.0 60200.0 153805.0 ;
      RECT  59495.0 155150.0 60200.0 153805.0 ;
      RECT  59495.0 155150.0 60200.0 156495.0 ;
      RECT  59495.0 157840.0 60200.0 156495.0 ;
      RECT  59495.0 157840.0 60200.0 159185.0 ;
      RECT  59495.0 160530.0 60200.0 159185.0 ;
      RECT  59495.0 160530.0 60200.0 161875.0 ;
      RECT  59495.0 163220.0 60200.0 161875.0 ;
      RECT  59495.0 163220.0 60200.0 164565.0 ;
      RECT  59495.0 165910.0 60200.0 164565.0 ;
      RECT  59495.0 165910.0 60200.0 167255.0 ;
      RECT  59495.0 168600.0 60200.0 167255.0 ;
      RECT  59495.0 168600.0 60200.0 169945.0 ;
      RECT  59495.0 171290.0 60200.0 169945.0 ;
      RECT  59495.0 171290.0 60200.0 172635.0 ;
      RECT  59495.0 173980.0 60200.0 172635.0 ;
      RECT  59495.0 173980.0 60200.0 175325.0 ;
      RECT  59495.0 176670.0 60200.0 175325.0 ;
      RECT  59495.0 176670.0 60200.0 178015.0 ;
      RECT  59495.0 179360.0 60200.0 178015.0 ;
      RECT  59495.0 179360.0 60200.0 180705.0 ;
      RECT  59495.0 182050.0 60200.0 180705.0 ;
      RECT  59495.0 182050.0 60200.0 183395.0 ;
      RECT  59495.0 184740.0 60200.0 183395.0 ;
      RECT  59495.0 184740.0 60200.0 186085.0 ;
      RECT  59495.0 187430.0 60200.0 186085.0 ;
      RECT  59495.0 187430.0 60200.0 188775.0 ;
      RECT  59495.0 190120.0 60200.0 188775.0 ;
      RECT  59495.0 190120.0 60200.0 191465.0 ;
      RECT  59495.0 192810.0 60200.0 191465.0 ;
      RECT  59495.0 192810.0 60200.0 194155.0 ;
      RECT  59495.0 195500.0 60200.0 194155.0 ;
      RECT  59495.0 195500.0 60200.0 196845.0 ;
      RECT  59495.0 198190.0 60200.0 196845.0 ;
      RECT  59495.0 198190.0 60200.0 199535.0 ;
      RECT  59495.0 200880.0 60200.0 199535.0 ;
      RECT  59495.0 200880.0 60200.0 202225.0 ;
      RECT  59495.0 203570.0 60200.0 202225.0 ;
      RECT  59495.0 203570.0 60200.0 204915.0 ;
      RECT  59495.0 206260.0 60200.0 204915.0 ;
      RECT  60200.0 34100.0 60905.0 35445.0 ;
      RECT  60200.0 36790.0 60905.0 35445.0 ;
      RECT  60200.0 36790.0 60905.0 38135.0 ;
      RECT  60200.0 39480.0 60905.0 38135.0 ;
      RECT  60200.0 39480.0 60905.0 40825.0 ;
      RECT  60200.0 42170.0 60905.0 40825.0 ;
      RECT  60200.0 42170.0 60905.0 43515.0 ;
      RECT  60200.0 44860.0 60905.0 43515.0 ;
      RECT  60200.0 44860.0 60905.0 46205.0 ;
      RECT  60200.0 47550.0 60905.0 46205.0 ;
      RECT  60200.0 47550.0 60905.0 48895.0 ;
      RECT  60200.0 50240.0 60905.0 48895.0 ;
      RECT  60200.0 50240.0 60905.0 51585.0 ;
      RECT  60200.0 52930.0 60905.0 51585.0 ;
      RECT  60200.0 52930.0 60905.0 54275.0 ;
      RECT  60200.0 55620.0 60905.0 54275.0 ;
      RECT  60200.0 55620.0 60905.0 56965.0 ;
      RECT  60200.0 58310.0 60905.0 56965.0 ;
      RECT  60200.0 58310.0 60905.0 59655.0 ;
      RECT  60200.0 61000.0 60905.0 59655.0 ;
      RECT  60200.0 61000.0 60905.0 62345.0 ;
      RECT  60200.0 63690.0 60905.0 62345.0 ;
      RECT  60200.0 63690.0 60905.0 65035.0 ;
      RECT  60200.0 66380.0 60905.0 65035.0 ;
      RECT  60200.0 66380.0 60905.0 67725.0 ;
      RECT  60200.0 69070.0 60905.0 67725.0 ;
      RECT  60200.0 69070.0 60905.0 70415.0 ;
      RECT  60200.0 71760.0 60905.0 70415.0 ;
      RECT  60200.0 71760.0 60905.0 73105.0 ;
      RECT  60200.0 74450.0 60905.0 73105.0 ;
      RECT  60200.0 74450.0 60905.0 75795.0 ;
      RECT  60200.0 77140.0 60905.0 75795.0 ;
      RECT  60200.0 77140.0 60905.0 78485.0 ;
      RECT  60200.0 79830.0 60905.0 78485.0 ;
      RECT  60200.0 79830.0 60905.0 81175.0 ;
      RECT  60200.0 82520.0 60905.0 81175.0 ;
      RECT  60200.0 82520.0 60905.0 83865.0 ;
      RECT  60200.0 85210.0 60905.0 83865.0 ;
      RECT  60200.0 85210.0 60905.0 86555.0 ;
      RECT  60200.0 87900.0 60905.0 86555.0 ;
      RECT  60200.0 87900.0 60905.0 89245.0 ;
      RECT  60200.0 90590.0 60905.0 89245.0 ;
      RECT  60200.0 90590.0 60905.0 91935.0 ;
      RECT  60200.0 93280.0 60905.0 91935.0 ;
      RECT  60200.0 93280.0 60905.0 94625.0 ;
      RECT  60200.0 95970.0 60905.0 94625.0 ;
      RECT  60200.0 95970.0 60905.0 97315.0 ;
      RECT  60200.0 98660.0 60905.0 97315.0 ;
      RECT  60200.0 98660.0 60905.0 100005.0 ;
      RECT  60200.0 101350.0 60905.0 100005.0 ;
      RECT  60200.0 101350.0 60905.0 102695.0 ;
      RECT  60200.0 104040.0 60905.0 102695.0 ;
      RECT  60200.0 104040.0 60905.0 105385.0 ;
      RECT  60200.0 106730.0 60905.0 105385.0 ;
      RECT  60200.0 106730.0 60905.0 108075.0 ;
      RECT  60200.0 109420.0 60905.0 108075.0 ;
      RECT  60200.0 109420.0 60905.0 110765.0 ;
      RECT  60200.0 112110.0 60905.0 110765.0 ;
      RECT  60200.0 112110.0 60905.0 113455.0 ;
      RECT  60200.0 114800.0 60905.0 113455.0 ;
      RECT  60200.0 114800.0 60905.0 116145.0 ;
      RECT  60200.0 117490.0 60905.0 116145.0 ;
      RECT  60200.0 117490.0 60905.0 118835.0 ;
      RECT  60200.0 120180.0 60905.0 118835.0 ;
      RECT  60200.0 120180.0 60905.0 121525.0 ;
      RECT  60200.0 122870.0 60905.0 121525.0 ;
      RECT  60200.0 122870.0 60905.0 124215.0 ;
      RECT  60200.0 125560.0 60905.0 124215.0 ;
      RECT  60200.0 125560.0 60905.0 126905.0 ;
      RECT  60200.0 128250.0 60905.0 126905.0 ;
      RECT  60200.0 128250.0 60905.0 129595.0 ;
      RECT  60200.0 130940.0 60905.0 129595.0 ;
      RECT  60200.0 130940.0 60905.0 132285.0 ;
      RECT  60200.0 133630.0 60905.0 132285.0 ;
      RECT  60200.0 133630.0 60905.0 134975.0 ;
      RECT  60200.0 136320.0 60905.0 134975.0 ;
      RECT  60200.0 136320.0 60905.0 137665.0 ;
      RECT  60200.0 139010.0 60905.0 137665.0 ;
      RECT  60200.0 139010.0 60905.0 140355.0 ;
      RECT  60200.0 141700.0 60905.0 140355.0 ;
      RECT  60200.0 141700.0 60905.0 143045.0 ;
      RECT  60200.0 144390.0 60905.0 143045.0 ;
      RECT  60200.0 144390.0 60905.0 145735.0 ;
      RECT  60200.0 147080.0 60905.0 145735.0 ;
      RECT  60200.0 147080.0 60905.0 148425.0 ;
      RECT  60200.0 149770.0 60905.0 148425.0 ;
      RECT  60200.0 149770.0 60905.0 151115.0 ;
      RECT  60200.0 152460.0 60905.0 151115.0 ;
      RECT  60200.0 152460.0 60905.0 153805.0 ;
      RECT  60200.0 155150.0 60905.0 153805.0 ;
      RECT  60200.0 155150.0 60905.0 156495.0 ;
      RECT  60200.0 157840.0 60905.0 156495.0 ;
      RECT  60200.0 157840.0 60905.0 159185.0 ;
      RECT  60200.0 160530.0 60905.0 159185.0 ;
      RECT  60200.0 160530.0 60905.0 161875.0 ;
      RECT  60200.0 163220.0 60905.0 161875.0 ;
      RECT  60200.0 163220.0 60905.0 164565.0 ;
      RECT  60200.0 165910.0 60905.0 164565.0 ;
      RECT  60200.0 165910.0 60905.0 167255.0 ;
      RECT  60200.0 168600.0 60905.0 167255.0 ;
      RECT  60200.0 168600.0 60905.0 169945.0 ;
      RECT  60200.0 171290.0 60905.0 169945.0 ;
      RECT  60200.0 171290.0 60905.0 172635.0 ;
      RECT  60200.0 173980.0 60905.0 172635.0 ;
      RECT  60200.0 173980.0 60905.0 175325.0 ;
      RECT  60200.0 176670.0 60905.0 175325.0 ;
      RECT  60200.0 176670.0 60905.0 178015.0 ;
      RECT  60200.0 179360.0 60905.0 178015.0 ;
      RECT  60200.0 179360.0 60905.0 180705.0 ;
      RECT  60200.0 182050.0 60905.0 180705.0 ;
      RECT  60200.0 182050.0 60905.0 183395.0 ;
      RECT  60200.0 184740.0 60905.0 183395.0 ;
      RECT  60200.0 184740.0 60905.0 186085.0 ;
      RECT  60200.0 187430.0 60905.0 186085.0 ;
      RECT  60200.0 187430.0 60905.0 188775.0 ;
      RECT  60200.0 190120.0 60905.0 188775.0 ;
      RECT  60200.0 190120.0 60905.0 191465.0 ;
      RECT  60200.0 192810.0 60905.0 191465.0 ;
      RECT  60200.0 192810.0 60905.0 194155.0 ;
      RECT  60200.0 195500.0 60905.0 194155.0 ;
      RECT  60200.0 195500.0 60905.0 196845.0 ;
      RECT  60200.0 198190.0 60905.0 196845.0 ;
      RECT  60200.0 198190.0 60905.0 199535.0 ;
      RECT  60200.0 200880.0 60905.0 199535.0 ;
      RECT  60200.0 200880.0 60905.0 202225.0 ;
      RECT  60200.0 203570.0 60905.0 202225.0 ;
      RECT  60200.0 203570.0 60905.0 204915.0 ;
      RECT  60200.0 206260.0 60905.0 204915.0 ;
      RECT  60905.0 34100.0 61610.0 35445.0 ;
      RECT  60905.0 36790.0 61610.0 35445.0 ;
      RECT  60905.0 36790.0 61610.0 38135.0 ;
      RECT  60905.0 39480.0 61610.0 38135.0 ;
      RECT  60905.0 39480.0 61610.0 40825.0 ;
      RECT  60905.0 42170.0 61610.0 40825.0 ;
      RECT  60905.0 42170.0 61610.0 43515.0 ;
      RECT  60905.0 44860.0 61610.0 43515.0 ;
      RECT  60905.0 44860.0 61610.0 46205.0 ;
      RECT  60905.0 47550.0 61610.0 46205.0 ;
      RECT  60905.0 47550.0 61610.0 48895.0 ;
      RECT  60905.0 50240.0 61610.0 48895.0 ;
      RECT  60905.0 50240.0 61610.0 51585.0 ;
      RECT  60905.0 52930.0 61610.0 51585.0 ;
      RECT  60905.0 52930.0 61610.0 54275.0 ;
      RECT  60905.0 55620.0 61610.0 54275.0 ;
      RECT  60905.0 55620.0 61610.0 56965.0 ;
      RECT  60905.0 58310.0 61610.0 56965.0 ;
      RECT  60905.0 58310.0 61610.0 59655.0 ;
      RECT  60905.0 61000.0 61610.0 59655.0 ;
      RECT  60905.0 61000.0 61610.0 62345.0 ;
      RECT  60905.0 63690.0 61610.0 62345.0 ;
      RECT  60905.0 63690.0 61610.0 65035.0 ;
      RECT  60905.0 66380.0 61610.0 65035.0 ;
      RECT  60905.0 66380.0 61610.0 67725.0 ;
      RECT  60905.0 69070.0 61610.0 67725.0 ;
      RECT  60905.0 69070.0 61610.0 70415.0 ;
      RECT  60905.0 71760.0 61610.0 70415.0 ;
      RECT  60905.0 71760.0 61610.0 73105.0 ;
      RECT  60905.0 74450.0 61610.0 73105.0 ;
      RECT  60905.0 74450.0 61610.0 75795.0 ;
      RECT  60905.0 77140.0 61610.0 75795.0 ;
      RECT  60905.0 77140.0 61610.0 78485.0 ;
      RECT  60905.0 79830.0 61610.0 78485.0 ;
      RECT  60905.0 79830.0 61610.0 81175.0 ;
      RECT  60905.0 82520.0 61610.0 81175.0 ;
      RECT  60905.0 82520.0 61610.0 83865.0 ;
      RECT  60905.0 85210.0 61610.0 83865.0 ;
      RECT  60905.0 85210.0 61610.0 86555.0 ;
      RECT  60905.0 87900.0 61610.0 86555.0 ;
      RECT  60905.0 87900.0 61610.0 89245.0 ;
      RECT  60905.0 90590.0 61610.0 89245.0 ;
      RECT  60905.0 90590.0 61610.0 91935.0 ;
      RECT  60905.0 93280.0 61610.0 91935.0 ;
      RECT  60905.0 93280.0 61610.0 94625.0 ;
      RECT  60905.0 95970.0 61610.0 94625.0 ;
      RECT  60905.0 95970.0 61610.0 97315.0 ;
      RECT  60905.0 98660.0 61610.0 97315.0 ;
      RECT  60905.0 98660.0 61610.0 100005.0 ;
      RECT  60905.0 101350.0 61610.0 100005.0 ;
      RECT  60905.0 101350.0 61610.0 102695.0 ;
      RECT  60905.0 104040.0 61610.0 102695.0 ;
      RECT  60905.0 104040.0 61610.0 105385.0 ;
      RECT  60905.0 106730.0 61610.0 105385.0 ;
      RECT  60905.0 106730.0 61610.0 108075.0 ;
      RECT  60905.0 109420.0 61610.0 108075.0 ;
      RECT  60905.0 109420.0 61610.0 110765.0 ;
      RECT  60905.0 112110.0 61610.0 110765.0 ;
      RECT  60905.0 112110.0 61610.0 113455.0 ;
      RECT  60905.0 114800.0 61610.0 113455.0 ;
      RECT  60905.0 114800.0 61610.0 116145.0 ;
      RECT  60905.0 117490.0 61610.0 116145.0 ;
      RECT  60905.0 117490.0 61610.0 118835.0 ;
      RECT  60905.0 120180.0 61610.0 118835.0 ;
      RECT  60905.0 120180.0 61610.0 121525.0 ;
      RECT  60905.0 122870.0 61610.0 121525.0 ;
      RECT  60905.0 122870.0 61610.0 124215.0 ;
      RECT  60905.0 125560.0 61610.0 124215.0 ;
      RECT  60905.0 125560.0 61610.0 126905.0 ;
      RECT  60905.0 128250.0 61610.0 126905.0 ;
      RECT  60905.0 128250.0 61610.0 129595.0 ;
      RECT  60905.0 130940.0 61610.0 129595.0 ;
      RECT  60905.0 130940.0 61610.0 132285.0 ;
      RECT  60905.0 133630.0 61610.0 132285.0 ;
      RECT  60905.0 133630.0 61610.0 134975.0 ;
      RECT  60905.0 136320.0 61610.0 134975.0 ;
      RECT  60905.0 136320.0 61610.0 137665.0 ;
      RECT  60905.0 139010.0 61610.0 137665.0 ;
      RECT  60905.0 139010.0 61610.0 140355.0 ;
      RECT  60905.0 141700.0 61610.0 140355.0 ;
      RECT  60905.0 141700.0 61610.0 143045.0 ;
      RECT  60905.0 144390.0 61610.0 143045.0 ;
      RECT  60905.0 144390.0 61610.0 145735.0 ;
      RECT  60905.0 147080.0 61610.0 145735.0 ;
      RECT  60905.0 147080.0 61610.0 148425.0 ;
      RECT  60905.0 149770.0 61610.0 148425.0 ;
      RECT  60905.0 149770.0 61610.0 151115.0 ;
      RECT  60905.0 152460.0 61610.0 151115.0 ;
      RECT  60905.0 152460.0 61610.0 153805.0 ;
      RECT  60905.0 155150.0 61610.0 153805.0 ;
      RECT  60905.0 155150.0 61610.0 156495.0 ;
      RECT  60905.0 157840.0 61610.0 156495.0 ;
      RECT  60905.0 157840.0 61610.0 159185.0 ;
      RECT  60905.0 160530.0 61610.0 159185.0 ;
      RECT  60905.0 160530.0 61610.0 161875.0 ;
      RECT  60905.0 163220.0 61610.0 161875.0 ;
      RECT  60905.0 163220.0 61610.0 164565.0 ;
      RECT  60905.0 165910.0 61610.0 164565.0 ;
      RECT  60905.0 165910.0 61610.0 167255.0 ;
      RECT  60905.0 168600.0 61610.0 167255.0 ;
      RECT  60905.0 168600.0 61610.0 169945.0 ;
      RECT  60905.0 171290.0 61610.0 169945.0 ;
      RECT  60905.0 171290.0 61610.0 172635.0 ;
      RECT  60905.0 173980.0 61610.0 172635.0 ;
      RECT  60905.0 173980.0 61610.0 175325.0 ;
      RECT  60905.0 176670.0 61610.0 175325.0 ;
      RECT  60905.0 176670.0 61610.0 178015.0 ;
      RECT  60905.0 179360.0 61610.0 178015.0 ;
      RECT  60905.0 179360.0 61610.0 180705.0 ;
      RECT  60905.0 182050.0 61610.0 180705.0 ;
      RECT  60905.0 182050.0 61610.0 183395.0 ;
      RECT  60905.0 184740.0 61610.0 183395.0 ;
      RECT  60905.0 184740.0 61610.0 186085.0 ;
      RECT  60905.0 187430.0 61610.0 186085.0 ;
      RECT  60905.0 187430.0 61610.0 188775.0 ;
      RECT  60905.0 190120.0 61610.0 188775.0 ;
      RECT  60905.0 190120.0 61610.0 191465.0 ;
      RECT  60905.0 192810.0 61610.0 191465.0 ;
      RECT  60905.0 192810.0 61610.0 194155.0 ;
      RECT  60905.0 195500.0 61610.0 194155.0 ;
      RECT  60905.0 195500.0 61610.0 196845.0 ;
      RECT  60905.0 198190.0 61610.0 196845.0 ;
      RECT  60905.0 198190.0 61610.0 199535.0 ;
      RECT  60905.0 200880.0 61610.0 199535.0 ;
      RECT  60905.0 200880.0 61610.0 202225.0 ;
      RECT  60905.0 203570.0 61610.0 202225.0 ;
      RECT  60905.0 203570.0 61610.0 204915.0 ;
      RECT  60905.0 206260.0 61610.0 204915.0 ;
      RECT  61610.0 34100.0 62315.0 35445.0 ;
      RECT  61610.0 36790.0 62315.0 35445.0 ;
      RECT  61610.0 36790.0 62315.0 38135.0 ;
      RECT  61610.0 39480.0 62315.0 38135.0 ;
      RECT  61610.0 39480.0 62315.0 40825.0 ;
      RECT  61610.0 42170.0 62315.0 40825.0 ;
      RECT  61610.0 42170.0 62315.0 43515.0 ;
      RECT  61610.0 44860.0 62315.0 43515.0 ;
      RECT  61610.0 44860.0 62315.0 46205.0 ;
      RECT  61610.0 47550.0 62315.0 46205.0 ;
      RECT  61610.0 47550.0 62315.0 48895.0 ;
      RECT  61610.0 50240.0 62315.0 48895.0 ;
      RECT  61610.0 50240.0 62315.0 51585.0 ;
      RECT  61610.0 52930.0 62315.0 51585.0 ;
      RECT  61610.0 52930.0 62315.0 54275.0 ;
      RECT  61610.0 55620.0 62315.0 54275.0 ;
      RECT  61610.0 55620.0 62315.0 56965.0 ;
      RECT  61610.0 58310.0 62315.0 56965.0 ;
      RECT  61610.0 58310.0 62315.0 59655.0 ;
      RECT  61610.0 61000.0 62315.0 59655.0 ;
      RECT  61610.0 61000.0 62315.0 62345.0 ;
      RECT  61610.0 63690.0 62315.0 62345.0 ;
      RECT  61610.0 63690.0 62315.0 65035.0 ;
      RECT  61610.0 66380.0 62315.0 65035.0 ;
      RECT  61610.0 66380.0 62315.0 67725.0 ;
      RECT  61610.0 69070.0 62315.0 67725.0 ;
      RECT  61610.0 69070.0 62315.0 70415.0 ;
      RECT  61610.0 71760.0 62315.0 70415.0 ;
      RECT  61610.0 71760.0 62315.0 73105.0 ;
      RECT  61610.0 74450.0 62315.0 73105.0 ;
      RECT  61610.0 74450.0 62315.0 75795.0 ;
      RECT  61610.0 77140.0 62315.0 75795.0 ;
      RECT  61610.0 77140.0 62315.0 78485.0 ;
      RECT  61610.0 79830.0 62315.0 78485.0 ;
      RECT  61610.0 79830.0 62315.0 81175.0 ;
      RECT  61610.0 82520.0 62315.0 81175.0 ;
      RECT  61610.0 82520.0 62315.0 83865.0 ;
      RECT  61610.0 85210.0 62315.0 83865.0 ;
      RECT  61610.0 85210.0 62315.0 86555.0 ;
      RECT  61610.0 87900.0 62315.0 86555.0 ;
      RECT  61610.0 87900.0 62315.0 89245.0 ;
      RECT  61610.0 90590.0 62315.0 89245.0 ;
      RECT  61610.0 90590.0 62315.0 91935.0 ;
      RECT  61610.0 93280.0 62315.0 91935.0 ;
      RECT  61610.0 93280.0 62315.0 94625.0 ;
      RECT  61610.0 95970.0 62315.0 94625.0 ;
      RECT  61610.0 95970.0 62315.0 97315.0 ;
      RECT  61610.0 98660.0 62315.0 97315.0 ;
      RECT  61610.0 98660.0 62315.0 100005.0 ;
      RECT  61610.0 101350.0 62315.0 100005.0 ;
      RECT  61610.0 101350.0 62315.0 102695.0 ;
      RECT  61610.0 104040.0 62315.0 102695.0 ;
      RECT  61610.0 104040.0 62315.0 105385.0 ;
      RECT  61610.0 106730.0 62315.0 105385.0 ;
      RECT  61610.0 106730.0 62315.0 108075.0 ;
      RECT  61610.0 109420.0 62315.0 108075.0 ;
      RECT  61610.0 109420.0 62315.0 110765.0 ;
      RECT  61610.0 112110.0 62315.0 110765.0 ;
      RECT  61610.0 112110.0 62315.0 113455.0 ;
      RECT  61610.0 114800.0 62315.0 113455.0 ;
      RECT  61610.0 114800.0 62315.0 116145.0 ;
      RECT  61610.0 117490.0 62315.0 116145.0 ;
      RECT  61610.0 117490.0 62315.0 118835.0 ;
      RECT  61610.0 120180.0 62315.0 118835.0 ;
      RECT  61610.0 120180.0 62315.0 121525.0 ;
      RECT  61610.0 122870.0 62315.0 121525.0 ;
      RECT  61610.0 122870.0 62315.0 124215.0 ;
      RECT  61610.0 125560.0 62315.0 124215.0 ;
      RECT  61610.0 125560.0 62315.0 126905.0 ;
      RECT  61610.0 128250.0 62315.0 126905.0 ;
      RECT  61610.0 128250.0 62315.0 129595.0 ;
      RECT  61610.0 130940.0 62315.0 129595.0 ;
      RECT  61610.0 130940.0 62315.0 132285.0 ;
      RECT  61610.0 133630.0 62315.0 132285.0 ;
      RECT  61610.0 133630.0 62315.0 134975.0 ;
      RECT  61610.0 136320.0 62315.0 134975.0 ;
      RECT  61610.0 136320.0 62315.0 137665.0 ;
      RECT  61610.0 139010.0 62315.0 137665.0 ;
      RECT  61610.0 139010.0 62315.0 140355.0 ;
      RECT  61610.0 141700.0 62315.0 140355.0 ;
      RECT  61610.0 141700.0 62315.0 143045.0 ;
      RECT  61610.0 144390.0 62315.0 143045.0 ;
      RECT  61610.0 144390.0 62315.0 145735.0 ;
      RECT  61610.0 147080.0 62315.0 145735.0 ;
      RECT  61610.0 147080.0 62315.0 148425.0 ;
      RECT  61610.0 149770.0 62315.0 148425.0 ;
      RECT  61610.0 149770.0 62315.0 151115.0 ;
      RECT  61610.0 152460.0 62315.0 151115.0 ;
      RECT  61610.0 152460.0 62315.0 153805.0 ;
      RECT  61610.0 155150.0 62315.0 153805.0 ;
      RECT  61610.0 155150.0 62315.0 156495.0 ;
      RECT  61610.0 157840.0 62315.0 156495.0 ;
      RECT  61610.0 157840.0 62315.0 159185.0 ;
      RECT  61610.0 160530.0 62315.0 159185.0 ;
      RECT  61610.0 160530.0 62315.0 161875.0 ;
      RECT  61610.0 163220.0 62315.0 161875.0 ;
      RECT  61610.0 163220.0 62315.0 164565.0 ;
      RECT  61610.0 165910.0 62315.0 164565.0 ;
      RECT  61610.0 165910.0 62315.0 167255.0 ;
      RECT  61610.0 168600.0 62315.0 167255.0 ;
      RECT  61610.0 168600.0 62315.0 169945.0 ;
      RECT  61610.0 171290.0 62315.0 169945.0 ;
      RECT  61610.0 171290.0 62315.0 172635.0 ;
      RECT  61610.0 173980.0 62315.0 172635.0 ;
      RECT  61610.0 173980.0 62315.0 175325.0 ;
      RECT  61610.0 176670.0 62315.0 175325.0 ;
      RECT  61610.0 176670.0 62315.0 178015.0 ;
      RECT  61610.0 179360.0 62315.0 178015.0 ;
      RECT  61610.0 179360.0 62315.0 180705.0 ;
      RECT  61610.0 182050.0 62315.0 180705.0 ;
      RECT  61610.0 182050.0 62315.0 183395.0 ;
      RECT  61610.0 184740.0 62315.0 183395.0 ;
      RECT  61610.0 184740.0 62315.0 186085.0 ;
      RECT  61610.0 187430.0 62315.0 186085.0 ;
      RECT  61610.0 187430.0 62315.0 188775.0 ;
      RECT  61610.0 190120.0 62315.0 188775.0 ;
      RECT  61610.0 190120.0 62315.0 191465.0 ;
      RECT  61610.0 192810.0 62315.0 191465.0 ;
      RECT  61610.0 192810.0 62315.0 194155.0 ;
      RECT  61610.0 195500.0 62315.0 194155.0 ;
      RECT  61610.0 195500.0 62315.0 196845.0 ;
      RECT  61610.0 198190.0 62315.0 196845.0 ;
      RECT  61610.0 198190.0 62315.0 199535.0 ;
      RECT  61610.0 200880.0 62315.0 199535.0 ;
      RECT  61610.0 200880.0 62315.0 202225.0 ;
      RECT  61610.0 203570.0 62315.0 202225.0 ;
      RECT  61610.0 203570.0 62315.0 204915.0 ;
      RECT  61610.0 206260.0 62315.0 204915.0 ;
      RECT  62315.0 34100.0 63020.0 35445.0 ;
      RECT  62315.0 36790.0 63020.0 35445.0 ;
      RECT  62315.0 36790.0 63020.0 38135.0 ;
      RECT  62315.0 39480.0 63020.0 38135.0 ;
      RECT  62315.0 39480.0 63020.0 40825.0 ;
      RECT  62315.0 42170.0 63020.0 40825.0 ;
      RECT  62315.0 42170.0 63020.0 43515.0 ;
      RECT  62315.0 44860.0 63020.0 43515.0 ;
      RECT  62315.0 44860.0 63020.0 46205.0 ;
      RECT  62315.0 47550.0 63020.0 46205.0 ;
      RECT  62315.0 47550.0 63020.0 48895.0 ;
      RECT  62315.0 50240.0 63020.0 48895.0 ;
      RECT  62315.0 50240.0 63020.0 51585.0 ;
      RECT  62315.0 52930.0 63020.0 51585.0 ;
      RECT  62315.0 52930.0 63020.0 54275.0 ;
      RECT  62315.0 55620.0 63020.0 54275.0 ;
      RECT  62315.0 55620.0 63020.0 56965.0 ;
      RECT  62315.0 58310.0 63020.0 56965.0 ;
      RECT  62315.0 58310.0 63020.0 59655.0 ;
      RECT  62315.0 61000.0 63020.0 59655.0 ;
      RECT  62315.0 61000.0 63020.0 62345.0 ;
      RECT  62315.0 63690.0 63020.0 62345.0 ;
      RECT  62315.0 63690.0 63020.0 65035.0 ;
      RECT  62315.0 66380.0 63020.0 65035.0 ;
      RECT  62315.0 66380.0 63020.0 67725.0 ;
      RECT  62315.0 69070.0 63020.0 67725.0 ;
      RECT  62315.0 69070.0 63020.0 70415.0 ;
      RECT  62315.0 71760.0 63020.0 70415.0 ;
      RECT  62315.0 71760.0 63020.0 73105.0 ;
      RECT  62315.0 74450.0 63020.0 73105.0 ;
      RECT  62315.0 74450.0 63020.0 75795.0 ;
      RECT  62315.0 77140.0 63020.0 75795.0 ;
      RECT  62315.0 77140.0 63020.0 78485.0 ;
      RECT  62315.0 79830.0 63020.0 78485.0 ;
      RECT  62315.0 79830.0 63020.0 81175.0 ;
      RECT  62315.0 82520.0 63020.0 81175.0 ;
      RECT  62315.0 82520.0 63020.0 83865.0 ;
      RECT  62315.0 85210.0 63020.0 83865.0 ;
      RECT  62315.0 85210.0 63020.0 86555.0 ;
      RECT  62315.0 87900.0 63020.0 86555.0 ;
      RECT  62315.0 87900.0 63020.0 89245.0 ;
      RECT  62315.0 90590.0 63020.0 89245.0 ;
      RECT  62315.0 90590.0 63020.0 91935.0 ;
      RECT  62315.0 93280.0 63020.0 91935.0 ;
      RECT  62315.0 93280.0 63020.0 94625.0 ;
      RECT  62315.0 95970.0 63020.0 94625.0 ;
      RECT  62315.0 95970.0 63020.0 97315.0 ;
      RECT  62315.0 98660.0 63020.0 97315.0 ;
      RECT  62315.0 98660.0 63020.0 100005.0 ;
      RECT  62315.0 101350.0 63020.0 100005.0 ;
      RECT  62315.0 101350.0 63020.0 102695.0 ;
      RECT  62315.0 104040.0 63020.0 102695.0 ;
      RECT  62315.0 104040.0 63020.0 105385.0 ;
      RECT  62315.0 106730.0 63020.0 105385.0 ;
      RECT  62315.0 106730.0 63020.0 108075.0 ;
      RECT  62315.0 109420.0 63020.0 108075.0 ;
      RECT  62315.0 109420.0 63020.0 110765.0 ;
      RECT  62315.0 112110.0 63020.0 110765.0 ;
      RECT  62315.0 112110.0 63020.0 113455.0 ;
      RECT  62315.0 114800.0 63020.0 113455.0 ;
      RECT  62315.0 114800.0 63020.0 116145.0 ;
      RECT  62315.0 117490.0 63020.0 116145.0 ;
      RECT  62315.0 117490.0 63020.0 118835.0 ;
      RECT  62315.0 120180.0 63020.0 118835.0 ;
      RECT  62315.0 120180.0 63020.0 121525.0 ;
      RECT  62315.0 122870.0 63020.0 121525.0 ;
      RECT  62315.0 122870.0 63020.0 124215.0 ;
      RECT  62315.0 125560.0 63020.0 124215.0 ;
      RECT  62315.0 125560.0 63020.0 126905.0 ;
      RECT  62315.0 128250.0 63020.0 126905.0 ;
      RECT  62315.0 128250.0 63020.0 129595.0 ;
      RECT  62315.0 130940.0 63020.0 129595.0 ;
      RECT  62315.0 130940.0 63020.0 132285.0 ;
      RECT  62315.0 133630.0 63020.0 132285.0 ;
      RECT  62315.0 133630.0 63020.0 134975.0 ;
      RECT  62315.0 136320.0 63020.0 134975.0 ;
      RECT  62315.0 136320.0 63020.0 137665.0 ;
      RECT  62315.0 139010.0 63020.0 137665.0 ;
      RECT  62315.0 139010.0 63020.0 140355.0 ;
      RECT  62315.0 141700.0 63020.0 140355.0 ;
      RECT  62315.0 141700.0 63020.0 143045.0 ;
      RECT  62315.0 144390.0 63020.0 143045.0 ;
      RECT  62315.0 144390.0 63020.0 145735.0 ;
      RECT  62315.0 147080.0 63020.0 145735.0 ;
      RECT  62315.0 147080.0 63020.0 148425.0 ;
      RECT  62315.0 149770.0 63020.0 148425.0 ;
      RECT  62315.0 149770.0 63020.0 151115.0 ;
      RECT  62315.0 152460.0 63020.0 151115.0 ;
      RECT  62315.0 152460.0 63020.0 153805.0 ;
      RECT  62315.0 155150.0 63020.0 153805.0 ;
      RECT  62315.0 155150.0 63020.0 156495.0 ;
      RECT  62315.0 157840.0 63020.0 156495.0 ;
      RECT  62315.0 157840.0 63020.0 159185.0 ;
      RECT  62315.0 160530.0 63020.0 159185.0 ;
      RECT  62315.0 160530.0 63020.0 161875.0 ;
      RECT  62315.0 163220.0 63020.0 161875.0 ;
      RECT  62315.0 163220.0 63020.0 164565.0 ;
      RECT  62315.0 165910.0 63020.0 164565.0 ;
      RECT  62315.0 165910.0 63020.0 167255.0 ;
      RECT  62315.0 168600.0 63020.0 167255.0 ;
      RECT  62315.0 168600.0 63020.0 169945.0 ;
      RECT  62315.0 171290.0 63020.0 169945.0 ;
      RECT  62315.0 171290.0 63020.0 172635.0 ;
      RECT  62315.0 173980.0 63020.0 172635.0 ;
      RECT  62315.0 173980.0 63020.0 175325.0 ;
      RECT  62315.0 176670.0 63020.0 175325.0 ;
      RECT  62315.0 176670.0 63020.0 178015.0 ;
      RECT  62315.0 179360.0 63020.0 178015.0 ;
      RECT  62315.0 179360.0 63020.0 180705.0 ;
      RECT  62315.0 182050.0 63020.0 180705.0 ;
      RECT  62315.0 182050.0 63020.0 183395.0 ;
      RECT  62315.0 184740.0 63020.0 183395.0 ;
      RECT  62315.0 184740.0 63020.0 186085.0 ;
      RECT  62315.0 187430.0 63020.0 186085.0 ;
      RECT  62315.0 187430.0 63020.0 188775.0 ;
      RECT  62315.0 190120.0 63020.0 188775.0 ;
      RECT  62315.0 190120.0 63020.0 191465.0 ;
      RECT  62315.0 192810.0 63020.0 191465.0 ;
      RECT  62315.0 192810.0 63020.0 194155.0 ;
      RECT  62315.0 195500.0 63020.0 194155.0 ;
      RECT  62315.0 195500.0 63020.0 196845.0 ;
      RECT  62315.0 198190.0 63020.0 196845.0 ;
      RECT  62315.0 198190.0 63020.0 199535.0 ;
      RECT  62315.0 200880.0 63020.0 199535.0 ;
      RECT  62315.0 200880.0 63020.0 202225.0 ;
      RECT  62315.0 203570.0 63020.0 202225.0 ;
      RECT  62315.0 203570.0 63020.0 204915.0 ;
      RECT  62315.0 206260.0 63020.0 204915.0 ;
      RECT  63020.0 34100.0 63725.0 35445.0 ;
      RECT  63020.0 36790.0 63725.0 35445.0 ;
      RECT  63020.0 36790.0 63725.0 38135.0 ;
      RECT  63020.0 39480.0 63725.0 38135.0 ;
      RECT  63020.0 39480.0 63725.0 40825.0 ;
      RECT  63020.0 42170.0 63725.0 40825.0 ;
      RECT  63020.0 42170.0 63725.0 43515.0 ;
      RECT  63020.0 44860.0 63725.0 43515.0 ;
      RECT  63020.0 44860.0 63725.0 46205.0 ;
      RECT  63020.0 47550.0 63725.0 46205.0 ;
      RECT  63020.0 47550.0 63725.0 48895.0 ;
      RECT  63020.0 50240.0 63725.0 48895.0 ;
      RECT  63020.0 50240.0 63725.0 51585.0 ;
      RECT  63020.0 52930.0 63725.0 51585.0 ;
      RECT  63020.0 52930.0 63725.0 54275.0 ;
      RECT  63020.0 55620.0 63725.0 54275.0 ;
      RECT  63020.0 55620.0 63725.0 56965.0 ;
      RECT  63020.0 58310.0 63725.0 56965.0 ;
      RECT  63020.0 58310.0 63725.0 59655.0 ;
      RECT  63020.0 61000.0 63725.0 59655.0 ;
      RECT  63020.0 61000.0 63725.0 62345.0 ;
      RECT  63020.0 63690.0 63725.0 62345.0 ;
      RECT  63020.0 63690.0 63725.0 65035.0 ;
      RECT  63020.0 66380.0 63725.0 65035.0 ;
      RECT  63020.0 66380.0 63725.0 67725.0 ;
      RECT  63020.0 69070.0 63725.0 67725.0 ;
      RECT  63020.0 69070.0 63725.0 70415.0 ;
      RECT  63020.0 71760.0 63725.0 70415.0 ;
      RECT  63020.0 71760.0 63725.0 73105.0 ;
      RECT  63020.0 74450.0 63725.0 73105.0 ;
      RECT  63020.0 74450.0 63725.0 75795.0 ;
      RECT  63020.0 77140.0 63725.0 75795.0 ;
      RECT  63020.0 77140.0 63725.0 78485.0 ;
      RECT  63020.0 79830.0 63725.0 78485.0 ;
      RECT  63020.0 79830.0 63725.0 81175.0 ;
      RECT  63020.0 82520.0 63725.0 81175.0 ;
      RECT  63020.0 82520.0 63725.0 83865.0 ;
      RECT  63020.0 85210.0 63725.0 83865.0 ;
      RECT  63020.0 85210.0 63725.0 86555.0 ;
      RECT  63020.0 87900.0 63725.0 86555.0 ;
      RECT  63020.0 87900.0 63725.0 89245.0 ;
      RECT  63020.0 90590.0 63725.0 89245.0 ;
      RECT  63020.0 90590.0 63725.0 91935.0 ;
      RECT  63020.0 93280.0 63725.0 91935.0 ;
      RECT  63020.0 93280.0 63725.0 94625.0 ;
      RECT  63020.0 95970.0 63725.0 94625.0 ;
      RECT  63020.0 95970.0 63725.0 97315.0 ;
      RECT  63020.0 98660.0 63725.0 97315.0 ;
      RECT  63020.0 98660.0 63725.0 100005.0 ;
      RECT  63020.0 101350.0 63725.0 100005.0 ;
      RECT  63020.0 101350.0 63725.0 102695.0 ;
      RECT  63020.0 104040.0 63725.0 102695.0 ;
      RECT  63020.0 104040.0 63725.0 105385.0 ;
      RECT  63020.0 106730.0 63725.0 105385.0 ;
      RECT  63020.0 106730.0 63725.0 108075.0 ;
      RECT  63020.0 109420.0 63725.0 108075.0 ;
      RECT  63020.0 109420.0 63725.0 110765.0 ;
      RECT  63020.0 112110.0 63725.0 110765.0 ;
      RECT  63020.0 112110.0 63725.0 113455.0 ;
      RECT  63020.0 114800.0 63725.0 113455.0 ;
      RECT  63020.0 114800.0 63725.0 116145.0 ;
      RECT  63020.0 117490.0 63725.0 116145.0 ;
      RECT  63020.0 117490.0 63725.0 118835.0 ;
      RECT  63020.0 120180.0 63725.0 118835.0 ;
      RECT  63020.0 120180.0 63725.0 121525.0 ;
      RECT  63020.0 122870.0 63725.0 121525.0 ;
      RECT  63020.0 122870.0 63725.0 124215.0 ;
      RECT  63020.0 125560.0 63725.0 124215.0 ;
      RECT  63020.0 125560.0 63725.0 126905.0 ;
      RECT  63020.0 128250.0 63725.0 126905.0 ;
      RECT  63020.0 128250.0 63725.0 129595.0 ;
      RECT  63020.0 130940.0 63725.0 129595.0 ;
      RECT  63020.0 130940.0 63725.0 132285.0 ;
      RECT  63020.0 133630.0 63725.0 132285.0 ;
      RECT  63020.0 133630.0 63725.0 134975.0 ;
      RECT  63020.0 136320.0 63725.0 134975.0 ;
      RECT  63020.0 136320.0 63725.0 137665.0 ;
      RECT  63020.0 139010.0 63725.0 137665.0 ;
      RECT  63020.0 139010.0 63725.0 140355.0 ;
      RECT  63020.0 141700.0 63725.0 140355.0 ;
      RECT  63020.0 141700.0 63725.0 143045.0 ;
      RECT  63020.0 144390.0 63725.0 143045.0 ;
      RECT  63020.0 144390.0 63725.0 145735.0 ;
      RECT  63020.0 147080.0 63725.0 145735.0 ;
      RECT  63020.0 147080.0 63725.0 148425.0 ;
      RECT  63020.0 149770.0 63725.0 148425.0 ;
      RECT  63020.0 149770.0 63725.0 151115.0 ;
      RECT  63020.0 152460.0 63725.0 151115.0 ;
      RECT  63020.0 152460.0 63725.0 153805.0 ;
      RECT  63020.0 155150.0 63725.0 153805.0 ;
      RECT  63020.0 155150.0 63725.0 156495.0 ;
      RECT  63020.0 157840.0 63725.0 156495.0 ;
      RECT  63020.0 157840.0 63725.0 159185.0 ;
      RECT  63020.0 160530.0 63725.0 159185.0 ;
      RECT  63020.0 160530.0 63725.0 161875.0 ;
      RECT  63020.0 163220.0 63725.0 161875.0 ;
      RECT  63020.0 163220.0 63725.0 164565.0 ;
      RECT  63020.0 165910.0 63725.0 164565.0 ;
      RECT  63020.0 165910.0 63725.0 167255.0 ;
      RECT  63020.0 168600.0 63725.0 167255.0 ;
      RECT  63020.0 168600.0 63725.0 169945.0 ;
      RECT  63020.0 171290.0 63725.0 169945.0 ;
      RECT  63020.0 171290.0 63725.0 172635.0 ;
      RECT  63020.0 173980.0 63725.0 172635.0 ;
      RECT  63020.0 173980.0 63725.0 175325.0 ;
      RECT  63020.0 176670.0 63725.0 175325.0 ;
      RECT  63020.0 176670.0 63725.0 178015.0 ;
      RECT  63020.0 179360.0 63725.0 178015.0 ;
      RECT  63020.0 179360.0 63725.0 180705.0 ;
      RECT  63020.0 182050.0 63725.0 180705.0 ;
      RECT  63020.0 182050.0 63725.0 183395.0 ;
      RECT  63020.0 184740.0 63725.0 183395.0 ;
      RECT  63020.0 184740.0 63725.0 186085.0 ;
      RECT  63020.0 187430.0 63725.0 186085.0 ;
      RECT  63020.0 187430.0 63725.0 188775.0 ;
      RECT  63020.0 190120.0 63725.0 188775.0 ;
      RECT  63020.0 190120.0 63725.0 191465.0 ;
      RECT  63020.0 192810.0 63725.0 191465.0 ;
      RECT  63020.0 192810.0 63725.0 194155.0 ;
      RECT  63020.0 195500.0 63725.0 194155.0 ;
      RECT  63020.0 195500.0 63725.0 196845.0 ;
      RECT  63020.0 198190.0 63725.0 196845.0 ;
      RECT  63020.0 198190.0 63725.0 199535.0 ;
      RECT  63020.0 200880.0 63725.0 199535.0 ;
      RECT  63020.0 200880.0 63725.0 202225.0 ;
      RECT  63020.0 203570.0 63725.0 202225.0 ;
      RECT  63020.0 203570.0 63725.0 204915.0 ;
      RECT  63020.0 206260.0 63725.0 204915.0 ;
      RECT  63725.0 34100.0 64430.0 35445.0 ;
      RECT  63725.0 36790.0 64430.0 35445.0 ;
      RECT  63725.0 36790.0 64430.0 38135.0 ;
      RECT  63725.0 39480.0 64430.0 38135.0 ;
      RECT  63725.0 39480.0 64430.0 40825.0 ;
      RECT  63725.0 42170.0 64430.0 40825.0 ;
      RECT  63725.0 42170.0 64430.0 43515.0 ;
      RECT  63725.0 44860.0 64430.0 43515.0 ;
      RECT  63725.0 44860.0 64430.0 46205.0 ;
      RECT  63725.0 47550.0 64430.0 46205.0 ;
      RECT  63725.0 47550.0 64430.0 48895.0 ;
      RECT  63725.0 50240.0 64430.0 48895.0 ;
      RECT  63725.0 50240.0 64430.0 51585.0 ;
      RECT  63725.0 52930.0 64430.0 51585.0 ;
      RECT  63725.0 52930.0 64430.0 54275.0 ;
      RECT  63725.0 55620.0 64430.0 54275.0 ;
      RECT  63725.0 55620.0 64430.0 56965.0 ;
      RECT  63725.0 58310.0 64430.0 56965.0 ;
      RECT  63725.0 58310.0 64430.0 59655.0 ;
      RECT  63725.0 61000.0 64430.0 59655.0 ;
      RECT  63725.0 61000.0 64430.0 62345.0 ;
      RECT  63725.0 63690.0 64430.0 62345.0 ;
      RECT  63725.0 63690.0 64430.0 65035.0 ;
      RECT  63725.0 66380.0 64430.0 65035.0 ;
      RECT  63725.0 66380.0 64430.0 67725.0 ;
      RECT  63725.0 69070.0 64430.0 67725.0 ;
      RECT  63725.0 69070.0 64430.0 70415.0 ;
      RECT  63725.0 71760.0 64430.0 70415.0 ;
      RECT  63725.0 71760.0 64430.0 73105.0 ;
      RECT  63725.0 74450.0 64430.0 73105.0 ;
      RECT  63725.0 74450.0 64430.0 75795.0 ;
      RECT  63725.0 77140.0 64430.0 75795.0 ;
      RECT  63725.0 77140.0 64430.0 78485.0 ;
      RECT  63725.0 79830.0 64430.0 78485.0 ;
      RECT  63725.0 79830.0 64430.0 81175.0 ;
      RECT  63725.0 82520.0 64430.0 81175.0 ;
      RECT  63725.0 82520.0 64430.0 83865.0 ;
      RECT  63725.0 85210.0 64430.0 83865.0 ;
      RECT  63725.0 85210.0 64430.0 86555.0 ;
      RECT  63725.0 87900.0 64430.0 86555.0 ;
      RECT  63725.0 87900.0 64430.0 89245.0 ;
      RECT  63725.0 90590.0 64430.0 89245.0 ;
      RECT  63725.0 90590.0 64430.0 91935.0 ;
      RECT  63725.0 93280.0 64430.0 91935.0 ;
      RECT  63725.0 93280.0 64430.0 94625.0 ;
      RECT  63725.0 95970.0 64430.0 94625.0 ;
      RECT  63725.0 95970.0 64430.0 97315.0 ;
      RECT  63725.0 98660.0 64430.0 97315.0 ;
      RECT  63725.0 98660.0 64430.0 100005.0 ;
      RECT  63725.0 101350.0 64430.0 100005.0 ;
      RECT  63725.0 101350.0 64430.0 102695.0 ;
      RECT  63725.0 104040.0 64430.0 102695.0 ;
      RECT  63725.0 104040.0 64430.0 105385.0 ;
      RECT  63725.0 106730.0 64430.0 105385.0 ;
      RECT  63725.0 106730.0 64430.0 108075.0 ;
      RECT  63725.0 109420.0 64430.0 108075.0 ;
      RECT  63725.0 109420.0 64430.0 110765.0 ;
      RECT  63725.0 112110.0 64430.0 110765.0 ;
      RECT  63725.0 112110.0 64430.0 113455.0 ;
      RECT  63725.0 114800.0 64430.0 113455.0 ;
      RECT  63725.0 114800.0 64430.0 116145.0 ;
      RECT  63725.0 117490.0 64430.0 116145.0 ;
      RECT  63725.0 117490.0 64430.0 118835.0 ;
      RECT  63725.0 120180.0 64430.0 118835.0 ;
      RECT  63725.0 120180.0 64430.0 121525.0 ;
      RECT  63725.0 122870.0 64430.0 121525.0 ;
      RECT  63725.0 122870.0 64430.0 124215.0 ;
      RECT  63725.0 125560.0 64430.0 124215.0 ;
      RECT  63725.0 125560.0 64430.0 126905.0 ;
      RECT  63725.0 128250.0 64430.0 126905.0 ;
      RECT  63725.0 128250.0 64430.0 129595.0 ;
      RECT  63725.0 130940.0 64430.0 129595.0 ;
      RECT  63725.0 130940.0 64430.0 132285.0 ;
      RECT  63725.0 133630.0 64430.0 132285.0 ;
      RECT  63725.0 133630.0 64430.0 134975.0 ;
      RECT  63725.0 136320.0 64430.0 134975.0 ;
      RECT  63725.0 136320.0 64430.0 137665.0 ;
      RECT  63725.0 139010.0 64430.0 137665.0 ;
      RECT  63725.0 139010.0 64430.0 140355.0 ;
      RECT  63725.0 141700.0 64430.0 140355.0 ;
      RECT  63725.0 141700.0 64430.0 143045.0 ;
      RECT  63725.0 144390.0 64430.0 143045.0 ;
      RECT  63725.0 144390.0 64430.0 145735.0 ;
      RECT  63725.0 147080.0 64430.0 145735.0 ;
      RECT  63725.0 147080.0 64430.0 148425.0 ;
      RECT  63725.0 149770.0 64430.0 148425.0 ;
      RECT  63725.0 149770.0 64430.0 151115.0 ;
      RECT  63725.0 152460.0 64430.0 151115.0 ;
      RECT  63725.0 152460.0 64430.0 153805.0 ;
      RECT  63725.0 155150.0 64430.0 153805.0 ;
      RECT  63725.0 155150.0 64430.0 156495.0 ;
      RECT  63725.0 157840.0 64430.0 156495.0 ;
      RECT  63725.0 157840.0 64430.0 159185.0 ;
      RECT  63725.0 160530.0 64430.0 159185.0 ;
      RECT  63725.0 160530.0 64430.0 161875.0 ;
      RECT  63725.0 163220.0 64430.0 161875.0 ;
      RECT  63725.0 163220.0 64430.0 164565.0 ;
      RECT  63725.0 165910.0 64430.0 164565.0 ;
      RECT  63725.0 165910.0 64430.0 167255.0 ;
      RECT  63725.0 168600.0 64430.0 167255.0 ;
      RECT  63725.0 168600.0 64430.0 169945.0 ;
      RECT  63725.0 171290.0 64430.0 169945.0 ;
      RECT  63725.0 171290.0 64430.0 172635.0 ;
      RECT  63725.0 173980.0 64430.0 172635.0 ;
      RECT  63725.0 173980.0 64430.0 175325.0 ;
      RECT  63725.0 176670.0 64430.0 175325.0 ;
      RECT  63725.0 176670.0 64430.0 178015.0 ;
      RECT  63725.0 179360.0 64430.0 178015.0 ;
      RECT  63725.0 179360.0 64430.0 180705.0 ;
      RECT  63725.0 182050.0 64430.0 180705.0 ;
      RECT  63725.0 182050.0 64430.0 183395.0 ;
      RECT  63725.0 184740.0 64430.0 183395.0 ;
      RECT  63725.0 184740.0 64430.0 186085.0 ;
      RECT  63725.0 187430.0 64430.0 186085.0 ;
      RECT  63725.0 187430.0 64430.0 188775.0 ;
      RECT  63725.0 190120.0 64430.0 188775.0 ;
      RECT  63725.0 190120.0 64430.0 191465.0 ;
      RECT  63725.0 192810.0 64430.0 191465.0 ;
      RECT  63725.0 192810.0 64430.0 194155.0 ;
      RECT  63725.0 195500.0 64430.0 194155.0 ;
      RECT  63725.0 195500.0 64430.0 196845.0 ;
      RECT  63725.0 198190.0 64430.0 196845.0 ;
      RECT  63725.0 198190.0 64430.0 199535.0 ;
      RECT  63725.0 200880.0 64430.0 199535.0 ;
      RECT  63725.0 200880.0 64430.0 202225.0 ;
      RECT  63725.0 203570.0 64430.0 202225.0 ;
      RECT  63725.0 203570.0 64430.0 204915.0 ;
      RECT  63725.0 206260.0 64430.0 204915.0 ;
      RECT  64430.0 34100.0 65135.0 35445.0 ;
      RECT  64430.0 36790.0 65135.0 35445.0 ;
      RECT  64430.0 36790.0 65135.0 38135.0 ;
      RECT  64430.0 39480.0 65135.0 38135.0 ;
      RECT  64430.0 39480.0 65135.0 40825.0 ;
      RECT  64430.0 42170.0 65135.0 40825.0 ;
      RECT  64430.0 42170.0 65135.0 43515.0 ;
      RECT  64430.0 44860.0 65135.0 43515.0 ;
      RECT  64430.0 44860.0 65135.0 46205.0 ;
      RECT  64430.0 47550.0 65135.0 46205.0 ;
      RECT  64430.0 47550.0 65135.0 48895.0 ;
      RECT  64430.0 50240.0 65135.0 48895.0 ;
      RECT  64430.0 50240.0 65135.0 51585.0 ;
      RECT  64430.0 52930.0 65135.0 51585.0 ;
      RECT  64430.0 52930.0 65135.0 54275.0 ;
      RECT  64430.0 55620.0 65135.0 54275.0 ;
      RECT  64430.0 55620.0 65135.0 56965.0 ;
      RECT  64430.0 58310.0 65135.0 56965.0 ;
      RECT  64430.0 58310.0 65135.0 59655.0 ;
      RECT  64430.0 61000.0 65135.0 59655.0 ;
      RECT  64430.0 61000.0 65135.0 62345.0 ;
      RECT  64430.0 63690.0 65135.0 62345.0 ;
      RECT  64430.0 63690.0 65135.0 65035.0 ;
      RECT  64430.0 66380.0 65135.0 65035.0 ;
      RECT  64430.0 66380.0 65135.0 67725.0 ;
      RECT  64430.0 69070.0 65135.0 67725.0 ;
      RECT  64430.0 69070.0 65135.0 70415.0 ;
      RECT  64430.0 71760.0 65135.0 70415.0 ;
      RECT  64430.0 71760.0 65135.0 73105.0 ;
      RECT  64430.0 74450.0 65135.0 73105.0 ;
      RECT  64430.0 74450.0 65135.0 75795.0 ;
      RECT  64430.0 77140.0 65135.0 75795.0 ;
      RECT  64430.0 77140.0 65135.0 78485.0 ;
      RECT  64430.0 79830.0 65135.0 78485.0 ;
      RECT  64430.0 79830.0 65135.0 81175.0 ;
      RECT  64430.0 82520.0 65135.0 81175.0 ;
      RECT  64430.0 82520.0 65135.0 83865.0 ;
      RECT  64430.0 85210.0 65135.0 83865.0 ;
      RECT  64430.0 85210.0 65135.0 86555.0 ;
      RECT  64430.0 87900.0 65135.0 86555.0 ;
      RECT  64430.0 87900.0 65135.0 89245.0 ;
      RECT  64430.0 90590.0 65135.0 89245.0 ;
      RECT  64430.0 90590.0 65135.0 91935.0 ;
      RECT  64430.0 93280.0 65135.0 91935.0 ;
      RECT  64430.0 93280.0 65135.0 94625.0 ;
      RECT  64430.0 95970.0 65135.0 94625.0 ;
      RECT  64430.0 95970.0 65135.0 97315.0 ;
      RECT  64430.0 98660.0 65135.0 97315.0 ;
      RECT  64430.0 98660.0 65135.0 100005.0 ;
      RECT  64430.0 101350.0 65135.0 100005.0 ;
      RECT  64430.0 101350.0 65135.0 102695.0 ;
      RECT  64430.0 104040.0 65135.0 102695.0 ;
      RECT  64430.0 104040.0 65135.0 105385.0 ;
      RECT  64430.0 106730.0 65135.0 105385.0 ;
      RECT  64430.0 106730.0 65135.0 108075.0 ;
      RECT  64430.0 109420.0 65135.0 108075.0 ;
      RECT  64430.0 109420.0 65135.0 110765.0 ;
      RECT  64430.0 112110.0 65135.0 110765.0 ;
      RECT  64430.0 112110.0 65135.0 113455.0 ;
      RECT  64430.0 114800.0 65135.0 113455.0 ;
      RECT  64430.0 114800.0 65135.0 116145.0 ;
      RECT  64430.0 117490.0 65135.0 116145.0 ;
      RECT  64430.0 117490.0 65135.0 118835.0 ;
      RECT  64430.0 120180.0 65135.0 118835.0 ;
      RECT  64430.0 120180.0 65135.0 121525.0 ;
      RECT  64430.0 122870.0 65135.0 121525.0 ;
      RECT  64430.0 122870.0 65135.0 124215.0 ;
      RECT  64430.0 125560.0 65135.0 124215.0 ;
      RECT  64430.0 125560.0 65135.0 126905.0 ;
      RECT  64430.0 128250.0 65135.0 126905.0 ;
      RECT  64430.0 128250.0 65135.0 129595.0 ;
      RECT  64430.0 130940.0 65135.0 129595.0 ;
      RECT  64430.0 130940.0 65135.0 132285.0 ;
      RECT  64430.0 133630.0 65135.0 132285.0 ;
      RECT  64430.0 133630.0 65135.0 134975.0 ;
      RECT  64430.0 136320.0 65135.0 134975.0 ;
      RECT  64430.0 136320.0 65135.0 137665.0 ;
      RECT  64430.0 139010.0 65135.0 137665.0 ;
      RECT  64430.0 139010.0 65135.0 140355.0 ;
      RECT  64430.0 141700.0 65135.0 140355.0 ;
      RECT  64430.0 141700.0 65135.0 143045.0 ;
      RECT  64430.0 144390.0 65135.0 143045.0 ;
      RECT  64430.0 144390.0 65135.0 145735.0 ;
      RECT  64430.0 147080.0 65135.0 145735.0 ;
      RECT  64430.0 147080.0 65135.0 148425.0 ;
      RECT  64430.0 149770.0 65135.0 148425.0 ;
      RECT  64430.0 149770.0 65135.0 151115.0 ;
      RECT  64430.0 152460.0 65135.0 151115.0 ;
      RECT  64430.0 152460.0 65135.0 153805.0 ;
      RECT  64430.0 155150.0 65135.0 153805.0 ;
      RECT  64430.0 155150.0 65135.0 156495.0 ;
      RECT  64430.0 157840.0 65135.0 156495.0 ;
      RECT  64430.0 157840.0 65135.0 159185.0 ;
      RECT  64430.0 160530.0 65135.0 159185.0 ;
      RECT  64430.0 160530.0 65135.0 161875.0 ;
      RECT  64430.0 163220.0 65135.0 161875.0 ;
      RECT  64430.0 163220.0 65135.0 164565.0 ;
      RECT  64430.0 165910.0 65135.0 164565.0 ;
      RECT  64430.0 165910.0 65135.0 167255.0 ;
      RECT  64430.0 168600.0 65135.0 167255.0 ;
      RECT  64430.0 168600.0 65135.0 169945.0 ;
      RECT  64430.0 171290.0 65135.0 169945.0 ;
      RECT  64430.0 171290.0 65135.0 172635.0 ;
      RECT  64430.0 173980.0 65135.0 172635.0 ;
      RECT  64430.0 173980.0 65135.0 175325.0 ;
      RECT  64430.0 176670.0 65135.0 175325.0 ;
      RECT  64430.0 176670.0 65135.0 178015.0 ;
      RECT  64430.0 179360.0 65135.0 178015.0 ;
      RECT  64430.0 179360.0 65135.0 180705.0 ;
      RECT  64430.0 182050.0 65135.0 180705.0 ;
      RECT  64430.0 182050.0 65135.0 183395.0 ;
      RECT  64430.0 184740.0 65135.0 183395.0 ;
      RECT  64430.0 184740.0 65135.0 186085.0 ;
      RECT  64430.0 187430.0 65135.0 186085.0 ;
      RECT  64430.0 187430.0 65135.0 188775.0 ;
      RECT  64430.0 190120.0 65135.0 188775.0 ;
      RECT  64430.0 190120.0 65135.0 191465.0 ;
      RECT  64430.0 192810.0 65135.0 191465.0 ;
      RECT  64430.0 192810.0 65135.0 194155.0 ;
      RECT  64430.0 195500.0 65135.0 194155.0 ;
      RECT  64430.0 195500.0 65135.0 196845.0 ;
      RECT  64430.0 198190.0 65135.0 196845.0 ;
      RECT  64430.0 198190.0 65135.0 199535.0 ;
      RECT  64430.0 200880.0 65135.0 199535.0 ;
      RECT  64430.0 200880.0 65135.0 202225.0 ;
      RECT  64430.0 203570.0 65135.0 202225.0 ;
      RECT  64430.0 203570.0 65135.0 204915.0 ;
      RECT  64430.0 206260.0 65135.0 204915.0 ;
      RECT  65135.0 34100.0 65840.0 35445.0 ;
      RECT  65135.0 36790.0 65840.0 35445.0 ;
      RECT  65135.0 36790.0 65840.0 38135.0 ;
      RECT  65135.0 39480.0 65840.0 38135.0 ;
      RECT  65135.0 39480.0 65840.0 40825.0 ;
      RECT  65135.0 42170.0 65840.0 40825.0 ;
      RECT  65135.0 42170.0 65840.0 43515.0 ;
      RECT  65135.0 44860.0 65840.0 43515.0 ;
      RECT  65135.0 44860.0 65840.0 46205.0 ;
      RECT  65135.0 47550.0 65840.0 46205.0 ;
      RECT  65135.0 47550.0 65840.0 48895.0 ;
      RECT  65135.0 50240.0 65840.0 48895.0 ;
      RECT  65135.0 50240.0 65840.0 51585.0 ;
      RECT  65135.0 52930.0 65840.0 51585.0 ;
      RECT  65135.0 52930.0 65840.0 54275.0 ;
      RECT  65135.0 55620.0 65840.0 54275.0 ;
      RECT  65135.0 55620.0 65840.0 56965.0 ;
      RECT  65135.0 58310.0 65840.0 56965.0 ;
      RECT  65135.0 58310.0 65840.0 59655.0 ;
      RECT  65135.0 61000.0 65840.0 59655.0 ;
      RECT  65135.0 61000.0 65840.0 62345.0 ;
      RECT  65135.0 63690.0 65840.0 62345.0 ;
      RECT  65135.0 63690.0 65840.0 65035.0 ;
      RECT  65135.0 66380.0 65840.0 65035.0 ;
      RECT  65135.0 66380.0 65840.0 67725.0 ;
      RECT  65135.0 69070.0 65840.0 67725.0 ;
      RECT  65135.0 69070.0 65840.0 70415.0 ;
      RECT  65135.0 71760.0 65840.0 70415.0 ;
      RECT  65135.0 71760.0 65840.0 73105.0 ;
      RECT  65135.0 74450.0 65840.0 73105.0 ;
      RECT  65135.0 74450.0 65840.0 75795.0 ;
      RECT  65135.0 77140.0 65840.0 75795.0 ;
      RECT  65135.0 77140.0 65840.0 78485.0 ;
      RECT  65135.0 79830.0 65840.0 78485.0 ;
      RECT  65135.0 79830.0 65840.0 81175.0 ;
      RECT  65135.0 82520.0 65840.0 81175.0 ;
      RECT  65135.0 82520.0 65840.0 83865.0 ;
      RECT  65135.0 85210.0 65840.0 83865.0 ;
      RECT  65135.0 85210.0 65840.0 86555.0 ;
      RECT  65135.0 87900.0 65840.0 86555.0 ;
      RECT  65135.0 87900.0 65840.0 89245.0 ;
      RECT  65135.0 90590.0 65840.0 89245.0 ;
      RECT  65135.0 90590.0 65840.0 91935.0 ;
      RECT  65135.0 93280.0 65840.0 91935.0 ;
      RECT  65135.0 93280.0 65840.0 94625.0 ;
      RECT  65135.0 95970.0 65840.0 94625.0 ;
      RECT  65135.0 95970.0 65840.0 97315.0 ;
      RECT  65135.0 98660.0 65840.0 97315.0 ;
      RECT  65135.0 98660.0 65840.0 100005.0 ;
      RECT  65135.0 101350.0 65840.0 100005.0 ;
      RECT  65135.0 101350.0 65840.0 102695.0 ;
      RECT  65135.0 104040.0 65840.0 102695.0 ;
      RECT  65135.0 104040.0 65840.0 105385.0 ;
      RECT  65135.0 106730.0 65840.0 105385.0 ;
      RECT  65135.0 106730.0 65840.0 108075.0 ;
      RECT  65135.0 109420.0 65840.0 108075.0 ;
      RECT  65135.0 109420.0 65840.0 110765.0 ;
      RECT  65135.0 112110.0 65840.0 110765.0 ;
      RECT  65135.0 112110.0 65840.0 113455.0 ;
      RECT  65135.0 114800.0 65840.0 113455.0 ;
      RECT  65135.0 114800.0 65840.0 116145.0 ;
      RECT  65135.0 117490.0 65840.0 116145.0 ;
      RECT  65135.0 117490.0 65840.0 118835.0 ;
      RECT  65135.0 120180.0 65840.0 118835.0 ;
      RECT  65135.0 120180.0 65840.0 121525.0 ;
      RECT  65135.0 122870.0 65840.0 121525.0 ;
      RECT  65135.0 122870.0 65840.0 124215.0 ;
      RECT  65135.0 125560.0 65840.0 124215.0 ;
      RECT  65135.0 125560.0 65840.0 126905.0 ;
      RECT  65135.0 128250.0 65840.0 126905.0 ;
      RECT  65135.0 128250.0 65840.0 129595.0 ;
      RECT  65135.0 130940.0 65840.0 129595.0 ;
      RECT  65135.0 130940.0 65840.0 132285.0 ;
      RECT  65135.0 133630.0 65840.0 132285.0 ;
      RECT  65135.0 133630.0 65840.0 134975.0 ;
      RECT  65135.0 136320.0 65840.0 134975.0 ;
      RECT  65135.0 136320.0 65840.0 137665.0 ;
      RECT  65135.0 139010.0 65840.0 137665.0 ;
      RECT  65135.0 139010.0 65840.0 140355.0 ;
      RECT  65135.0 141700.0 65840.0 140355.0 ;
      RECT  65135.0 141700.0 65840.0 143045.0 ;
      RECT  65135.0 144390.0 65840.0 143045.0 ;
      RECT  65135.0 144390.0 65840.0 145735.0 ;
      RECT  65135.0 147080.0 65840.0 145735.0 ;
      RECT  65135.0 147080.0 65840.0 148425.0 ;
      RECT  65135.0 149770.0 65840.0 148425.0 ;
      RECT  65135.0 149770.0 65840.0 151115.0 ;
      RECT  65135.0 152460.0 65840.0 151115.0 ;
      RECT  65135.0 152460.0 65840.0 153805.0 ;
      RECT  65135.0 155150.0 65840.0 153805.0 ;
      RECT  65135.0 155150.0 65840.0 156495.0 ;
      RECT  65135.0 157840.0 65840.0 156495.0 ;
      RECT  65135.0 157840.0 65840.0 159185.0 ;
      RECT  65135.0 160530.0 65840.0 159185.0 ;
      RECT  65135.0 160530.0 65840.0 161875.0 ;
      RECT  65135.0 163220.0 65840.0 161875.0 ;
      RECT  65135.0 163220.0 65840.0 164565.0 ;
      RECT  65135.0 165910.0 65840.0 164565.0 ;
      RECT  65135.0 165910.0 65840.0 167255.0 ;
      RECT  65135.0 168600.0 65840.0 167255.0 ;
      RECT  65135.0 168600.0 65840.0 169945.0 ;
      RECT  65135.0 171290.0 65840.0 169945.0 ;
      RECT  65135.0 171290.0 65840.0 172635.0 ;
      RECT  65135.0 173980.0 65840.0 172635.0 ;
      RECT  65135.0 173980.0 65840.0 175325.0 ;
      RECT  65135.0 176670.0 65840.0 175325.0 ;
      RECT  65135.0 176670.0 65840.0 178015.0 ;
      RECT  65135.0 179360.0 65840.0 178015.0 ;
      RECT  65135.0 179360.0 65840.0 180705.0 ;
      RECT  65135.0 182050.0 65840.0 180705.0 ;
      RECT  65135.0 182050.0 65840.0 183395.0 ;
      RECT  65135.0 184740.0 65840.0 183395.0 ;
      RECT  65135.0 184740.0 65840.0 186085.0 ;
      RECT  65135.0 187430.0 65840.0 186085.0 ;
      RECT  65135.0 187430.0 65840.0 188775.0 ;
      RECT  65135.0 190120.0 65840.0 188775.0 ;
      RECT  65135.0 190120.0 65840.0 191465.0 ;
      RECT  65135.0 192810.0 65840.0 191465.0 ;
      RECT  65135.0 192810.0 65840.0 194155.0 ;
      RECT  65135.0 195500.0 65840.0 194155.0 ;
      RECT  65135.0 195500.0 65840.0 196845.0 ;
      RECT  65135.0 198190.0 65840.0 196845.0 ;
      RECT  65135.0 198190.0 65840.0 199535.0 ;
      RECT  65135.0 200880.0 65840.0 199535.0 ;
      RECT  65135.0 200880.0 65840.0 202225.0 ;
      RECT  65135.0 203570.0 65840.0 202225.0 ;
      RECT  65135.0 203570.0 65840.0 204915.0 ;
      RECT  65135.0 206260.0 65840.0 204915.0 ;
      RECT  65840.0 34100.0 66545.0 35445.0 ;
      RECT  65840.0 36790.0 66545.0 35445.0 ;
      RECT  65840.0 36790.0 66545.0 38135.0 ;
      RECT  65840.0 39480.0 66545.0 38135.0 ;
      RECT  65840.0 39480.0 66545.0 40825.0 ;
      RECT  65840.0 42170.0 66545.0 40825.0 ;
      RECT  65840.0 42170.0 66545.0 43515.0 ;
      RECT  65840.0 44860.0 66545.0 43515.0 ;
      RECT  65840.0 44860.0 66545.0 46205.0 ;
      RECT  65840.0 47550.0 66545.0 46205.0 ;
      RECT  65840.0 47550.0 66545.0 48895.0 ;
      RECT  65840.0 50240.0 66545.0 48895.0 ;
      RECT  65840.0 50240.0 66545.0 51585.0 ;
      RECT  65840.0 52930.0 66545.0 51585.0 ;
      RECT  65840.0 52930.0 66545.0 54275.0 ;
      RECT  65840.0 55620.0 66545.0 54275.0 ;
      RECT  65840.0 55620.0 66545.0 56965.0 ;
      RECT  65840.0 58310.0 66545.0 56965.0 ;
      RECT  65840.0 58310.0 66545.0 59655.0 ;
      RECT  65840.0 61000.0 66545.0 59655.0 ;
      RECT  65840.0 61000.0 66545.0 62345.0 ;
      RECT  65840.0 63690.0 66545.0 62345.0 ;
      RECT  65840.0 63690.0 66545.0 65035.0 ;
      RECT  65840.0 66380.0 66545.0 65035.0 ;
      RECT  65840.0 66380.0 66545.0 67725.0 ;
      RECT  65840.0 69070.0 66545.0 67725.0 ;
      RECT  65840.0 69070.0 66545.0 70415.0 ;
      RECT  65840.0 71760.0 66545.0 70415.0 ;
      RECT  65840.0 71760.0 66545.0 73105.0 ;
      RECT  65840.0 74450.0 66545.0 73105.0 ;
      RECT  65840.0 74450.0 66545.0 75795.0 ;
      RECT  65840.0 77140.0 66545.0 75795.0 ;
      RECT  65840.0 77140.0 66545.0 78485.0 ;
      RECT  65840.0 79830.0 66545.0 78485.0 ;
      RECT  65840.0 79830.0 66545.0 81175.0 ;
      RECT  65840.0 82520.0 66545.0 81175.0 ;
      RECT  65840.0 82520.0 66545.0 83865.0 ;
      RECT  65840.0 85210.0 66545.0 83865.0 ;
      RECT  65840.0 85210.0 66545.0 86555.0 ;
      RECT  65840.0 87900.0 66545.0 86555.0 ;
      RECT  65840.0 87900.0 66545.0 89245.0 ;
      RECT  65840.0 90590.0 66545.0 89245.0 ;
      RECT  65840.0 90590.0 66545.0 91935.0 ;
      RECT  65840.0 93280.0 66545.0 91935.0 ;
      RECT  65840.0 93280.0 66545.0 94625.0 ;
      RECT  65840.0 95970.0 66545.0 94625.0 ;
      RECT  65840.0 95970.0 66545.0 97315.0 ;
      RECT  65840.0 98660.0 66545.0 97315.0 ;
      RECT  65840.0 98660.0 66545.0 100005.0 ;
      RECT  65840.0 101350.0 66545.0 100005.0 ;
      RECT  65840.0 101350.0 66545.0 102695.0 ;
      RECT  65840.0 104040.0 66545.0 102695.0 ;
      RECT  65840.0 104040.0 66545.0 105385.0 ;
      RECT  65840.0 106730.0 66545.0 105385.0 ;
      RECT  65840.0 106730.0 66545.0 108075.0 ;
      RECT  65840.0 109420.0 66545.0 108075.0 ;
      RECT  65840.0 109420.0 66545.0 110765.0 ;
      RECT  65840.0 112110.0 66545.0 110765.0 ;
      RECT  65840.0 112110.0 66545.0 113455.0 ;
      RECT  65840.0 114800.0 66545.0 113455.0 ;
      RECT  65840.0 114800.0 66545.0 116145.0 ;
      RECT  65840.0 117490.0 66545.0 116145.0 ;
      RECT  65840.0 117490.0 66545.0 118835.0 ;
      RECT  65840.0 120180.0 66545.0 118835.0 ;
      RECT  65840.0 120180.0 66545.0 121525.0 ;
      RECT  65840.0 122870.0 66545.0 121525.0 ;
      RECT  65840.0 122870.0 66545.0 124215.0 ;
      RECT  65840.0 125560.0 66545.0 124215.0 ;
      RECT  65840.0 125560.0 66545.0 126905.0 ;
      RECT  65840.0 128250.0 66545.0 126905.0 ;
      RECT  65840.0 128250.0 66545.0 129595.0 ;
      RECT  65840.0 130940.0 66545.0 129595.0 ;
      RECT  65840.0 130940.0 66545.0 132285.0 ;
      RECT  65840.0 133630.0 66545.0 132285.0 ;
      RECT  65840.0 133630.0 66545.0 134975.0 ;
      RECT  65840.0 136320.0 66545.0 134975.0 ;
      RECT  65840.0 136320.0 66545.0 137665.0 ;
      RECT  65840.0 139010.0 66545.0 137665.0 ;
      RECT  65840.0 139010.0 66545.0 140355.0 ;
      RECT  65840.0 141700.0 66545.0 140355.0 ;
      RECT  65840.0 141700.0 66545.0 143045.0 ;
      RECT  65840.0 144390.0 66545.0 143045.0 ;
      RECT  65840.0 144390.0 66545.0 145735.0 ;
      RECT  65840.0 147080.0 66545.0 145735.0 ;
      RECT  65840.0 147080.0 66545.0 148425.0 ;
      RECT  65840.0 149770.0 66545.0 148425.0 ;
      RECT  65840.0 149770.0 66545.0 151115.0 ;
      RECT  65840.0 152460.0 66545.0 151115.0 ;
      RECT  65840.0 152460.0 66545.0 153805.0 ;
      RECT  65840.0 155150.0 66545.0 153805.0 ;
      RECT  65840.0 155150.0 66545.0 156495.0 ;
      RECT  65840.0 157840.0 66545.0 156495.0 ;
      RECT  65840.0 157840.0 66545.0 159185.0 ;
      RECT  65840.0 160530.0 66545.0 159185.0 ;
      RECT  65840.0 160530.0 66545.0 161875.0 ;
      RECT  65840.0 163220.0 66545.0 161875.0 ;
      RECT  65840.0 163220.0 66545.0 164565.0 ;
      RECT  65840.0 165910.0 66545.0 164565.0 ;
      RECT  65840.0 165910.0 66545.0 167255.0 ;
      RECT  65840.0 168600.0 66545.0 167255.0 ;
      RECT  65840.0 168600.0 66545.0 169945.0 ;
      RECT  65840.0 171290.0 66545.0 169945.0 ;
      RECT  65840.0 171290.0 66545.0 172635.0 ;
      RECT  65840.0 173980.0 66545.0 172635.0 ;
      RECT  65840.0 173980.0 66545.0 175325.0 ;
      RECT  65840.0 176670.0 66545.0 175325.0 ;
      RECT  65840.0 176670.0 66545.0 178015.0 ;
      RECT  65840.0 179360.0 66545.0 178015.0 ;
      RECT  65840.0 179360.0 66545.0 180705.0 ;
      RECT  65840.0 182050.0 66545.0 180705.0 ;
      RECT  65840.0 182050.0 66545.0 183395.0 ;
      RECT  65840.0 184740.0 66545.0 183395.0 ;
      RECT  65840.0 184740.0 66545.0 186085.0 ;
      RECT  65840.0 187430.0 66545.0 186085.0 ;
      RECT  65840.0 187430.0 66545.0 188775.0 ;
      RECT  65840.0 190120.0 66545.0 188775.0 ;
      RECT  65840.0 190120.0 66545.0 191465.0 ;
      RECT  65840.0 192810.0 66545.0 191465.0 ;
      RECT  65840.0 192810.0 66545.0 194155.0 ;
      RECT  65840.0 195500.0 66545.0 194155.0 ;
      RECT  65840.0 195500.0 66545.0 196845.0 ;
      RECT  65840.0 198190.0 66545.0 196845.0 ;
      RECT  65840.0 198190.0 66545.0 199535.0 ;
      RECT  65840.0 200880.0 66545.0 199535.0 ;
      RECT  65840.0 200880.0 66545.0 202225.0 ;
      RECT  65840.0 203570.0 66545.0 202225.0 ;
      RECT  65840.0 203570.0 66545.0 204915.0 ;
      RECT  65840.0 206260.0 66545.0 204915.0 ;
      RECT  66545.0 34100.0 67250.0 35445.0 ;
      RECT  66545.0 36790.0 67250.0 35445.0 ;
      RECT  66545.0 36790.0 67250.0 38135.0 ;
      RECT  66545.0 39480.0 67250.0 38135.0 ;
      RECT  66545.0 39480.0 67250.0 40825.0 ;
      RECT  66545.0 42170.0 67250.0 40825.0 ;
      RECT  66545.0 42170.0 67250.0 43515.0 ;
      RECT  66545.0 44860.0 67250.0 43515.0 ;
      RECT  66545.0 44860.0 67250.0 46205.0 ;
      RECT  66545.0 47550.0 67250.0 46205.0 ;
      RECT  66545.0 47550.0 67250.0 48895.0 ;
      RECT  66545.0 50240.0 67250.0 48895.0 ;
      RECT  66545.0 50240.0 67250.0 51585.0 ;
      RECT  66545.0 52930.0 67250.0 51585.0 ;
      RECT  66545.0 52930.0 67250.0 54275.0 ;
      RECT  66545.0 55620.0 67250.0 54275.0 ;
      RECT  66545.0 55620.0 67250.0 56965.0 ;
      RECT  66545.0 58310.0 67250.0 56965.0 ;
      RECT  66545.0 58310.0 67250.0 59655.0 ;
      RECT  66545.0 61000.0 67250.0 59655.0 ;
      RECT  66545.0 61000.0 67250.0 62345.0 ;
      RECT  66545.0 63690.0 67250.0 62345.0 ;
      RECT  66545.0 63690.0 67250.0 65035.0 ;
      RECT  66545.0 66380.0 67250.0 65035.0 ;
      RECT  66545.0 66380.0 67250.0 67725.0 ;
      RECT  66545.0 69070.0 67250.0 67725.0 ;
      RECT  66545.0 69070.0 67250.0 70415.0 ;
      RECT  66545.0 71760.0 67250.0 70415.0 ;
      RECT  66545.0 71760.0 67250.0 73105.0 ;
      RECT  66545.0 74450.0 67250.0 73105.0 ;
      RECT  66545.0 74450.0 67250.0 75795.0 ;
      RECT  66545.0 77140.0 67250.0 75795.0 ;
      RECT  66545.0 77140.0 67250.0 78485.0 ;
      RECT  66545.0 79830.0 67250.0 78485.0 ;
      RECT  66545.0 79830.0 67250.0 81175.0 ;
      RECT  66545.0 82520.0 67250.0 81175.0 ;
      RECT  66545.0 82520.0 67250.0 83865.0 ;
      RECT  66545.0 85210.0 67250.0 83865.0 ;
      RECT  66545.0 85210.0 67250.0 86555.0 ;
      RECT  66545.0 87900.0 67250.0 86555.0 ;
      RECT  66545.0 87900.0 67250.0 89245.0 ;
      RECT  66545.0 90590.0 67250.0 89245.0 ;
      RECT  66545.0 90590.0 67250.0 91935.0 ;
      RECT  66545.0 93280.0 67250.0 91935.0 ;
      RECT  66545.0 93280.0 67250.0 94625.0 ;
      RECT  66545.0 95970.0 67250.0 94625.0 ;
      RECT  66545.0 95970.0 67250.0 97315.0 ;
      RECT  66545.0 98660.0 67250.0 97315.0 ;
      RECT  66545.0 98660.0 67250.0 100005.0 ;
      RECT  66545.0 101350.0 67250.0 100005.0 ;
      RECT  66545.0 101350.0 67250.0 102695.0 ;
      RECT  66545.0 104040.0 67250.0 102695.0 ;
      RECT  66545.0 104040.0 67250.0 105385.0 ;
      RECT  66545.0 106730.0 67250.0 105385.0 ;
      RECT  66545.0 106730.0 67250.0 108075.0 ;
      RECT  66545.0 109420.0 67250.0 108075.0 ;
      RECT  66545.0 109420.0 67250.0 110765.0 ;
      RECT  66545.0 112110.0 67250.0 110765.0 ;
      RECT  66545.0 112110.0 67250.0 113455.0 ;
      RECT  66545.0 114800.0 67250.0 113455.0 ;
      RECT  66545.0 114800.0 67250.0 116145.0 ;
      RECT  66545.0 117490.0 67250.0 116145.0 ;
      RECT  66545.0 117490.0 67250.0 118835.0 ;
      RECT  66545.0 120180.0 67250.0 118835.0 ;
      RECT  66545.0 120180.0 67250.0 121525.0 ;
      RECT  66545.0 122870.0 67250.0 121525.0 ;
      RECT  66545.0 122870.0 67250.0 124215.0 ;
      RECT  66545.0 125560.0 67250.0 124215.0 ;
      RECT  66545.0 125560.0 67250.0 126905.0 ;
      RECT  66545.0 128250.0 67250.0 126905.0 ;
      RECT  66545.0 128250.0 67250.0 129595.0 ;
      RECT  66545.0 130940.0 67250.0 129595.0 ;
      RECT  66545.0 130940.0 67250.0 132285.0 ;
      RECT  66545.0 133630.0 67250.0 132285.0 ;
      RECT  66545.0 133630.0 67250.0 134975.0 ;
      RECT  66545.0 136320.0 67250.0 134975.0 ;
      RECT  66545.0 136320.0 67250.0 137665.0 ;
      RECT  66545.0 139010.0 67250.0 137665.0 ;
      RECT  66545.0 139010.0 67250.0 140355.0 ;
      RECT  66545.0 141700.0 67250.0 140355.0 ;
      RECT  66545.0 141700.0 67250.0 143045.0 ;
      RECT  66545.0 144390.0 67250.0 143045.0 ;
      RECT  66545.0 144390.0 67250.0 145735.0 ;
      RECT  66545.0 147080.0 67250.0 145735.0 ;
      RECT  66545.0 147080.0 67250.0 148425.0 ;
      RECT  66545.0 149770.0 67250.0 148425.0 ;
      RECT  66545.0 149770.0 67250.0 151115.0 ;
      RECT  66545.0 152460.0 67250.0 151115.0 ;
      RECT  66545.0 152460.0 67250.0 153805.0 ;
      RECT  66545.0 155150.0 67250.0 153805.0 ;
      RECT  66545.0 155150.0 67250.0 156495.0 ;
      RECT  66545.0 157840.0 67250.0 156495.0 ;
      RECT  66545.0 157840.0 67250.0 159185.0 ;
      RECT  66545.0 160530.0 67250.0 159185.0 ;
      RECT  66545.0 160530.0 67250.0 161875.0 ;
      RECT  66545.0 163220.0 67250.0 161875.0 ;
      RECT  66545.0 163220.0 67250.0 164565.0 ;
      RECT  66545.0 165910.0 67250.0 164565.0 ;
      RECT  66545.0 165910.0 67250.0 167255.0 ;
      RECT  66545.0 168600.0 67250.0 167255.0 ;
      RECT  66545.0 168600.0 67250.0 169945.0 ;
      RECT  66545.0 171290.0 67250.0 169945.0 ;
      RECT  66545.0 171290.0 67250.0 172635.0 ;
      RECT  66545.0 173980.0 67250.0 172635.0 ;
      RECT  66545.0 173980.0 67250.0 175325.0 ;
      RECT  66545.0 176670.0 67250.0 175325.0 ;
      RECT  66545.0 176670.0 67250.0 178015.0 ;
      RECT  66545.0 179360.0 67250.0 178015.0 ;
      RECT  66545.0 179360.0 67250.0 180705.0 ;
      RECT  66545.0 182050.0 67250.0 180705.0 ;
      RECT  66545.0 182050.0 67250.0 183395.0 ;
      RECT  66545.0 184740.0 67250.0 183395.0 ;
      RECT  66545.0 184740.0 67250.0 186085.0 ;
      RECT  66545.0 187430.0 67250.0 186085.0 ;
      RECT  66545.0 187430.0 67250.0 188775.0 ;
      RECT  66545.0 190120.0 67250.0 188775.0 ;
      RECT  66545.0 190120.0 67250.0 191465.0 ;
      RECT  66545.0 192810.0 67250.0 191465.0 ;
      RECT  66545.0 192810.0 67250.0 194155.0 ;
      RECT  66545.0 195500.0 67250.0 194155.0 ;
      RECT  66545.0 195500.0 67250.0 196845.0 ;
      RECT  66545.0 198190.0 67250.0 196845.0 ;
      RECT  66545.0 198190.0 67250.0 199535.0 ;
      RECT  66545.0 200880.0 67250.0 199535.0 ;
      RECT  66545.0 200880.0 67250.0 202225.0 ;
      RECT  66545.0 203570.0 67250.0 202225.0 ;
      RECT  66545.0 203570.0 67250.0 204915.0 ;
      RECT  66545.0 206260.0 67250.0 204915.0 ;
      RECT  67250.0 34100.0 67955.0 35445.0 ;
      RECT  67250.0 36790.0 67955.0 35445.0 ;
      RECT  67250.0 36790.0 67955.0 38135.0 ;
      RECT  67250.0 39480.0 67955.0 38135.0 ;
      RECT  67250.0 39480.0 67955.0 40825.0 ;
      RECT  67250.0 42170.0 67955.0 40825.0 ;
      RECT  67250.0 42170.0 67955.0 43515.0 ;
      RECT  67250.0 44860.0 67955.0 43515.0 ;
      RECT  67250.0 44860.0 67955.0 46205.0 ;
      RECT  67250.0 47550.0 67955.0 46205.0 ;
      RECT  67250.0 47550.0 67955.0 48895.0 ;
      RECT  67250.0 50240.0 67955.0 48895.0 ;
      RECT  67250.0 50240.0 67955.0 51585.0 ;
      RECT  67250.0 52930.0 67955.0 51585.0 ;
      RECT  67250.0 52930.0 67955.0 54275.0 ;
      RECT  67250.0 55620.0 67955.0 54275.0 ;
      RECT  67250.0 55620.0 67955.0 56965.0 ;
      RECT  67250.0 58310.0 67955.0 56965.0 ;
      RECT  67250.0 58310.0 67955.0 59655.0 ;
      RECT  67250.0 61000.0 67955.0 59655.0 ;
      RECT  67250.0 61000.0 67955.0 62345.0 ;
      RECT  67250.0 63690.0 67955.0 62345.0 ;
      RECT  67250.0 63690.0 67955.0 65035.0 ;
      RECT  67250.0 66380.0 67955.0 65035.0 ;
      RECT  67250.0 66380.0 67955.0 67725.0 ;
      RECT  67250.0 69070.0 67955.0 67725.0 ;
      RECT  67250.0 69070.0 67955.0 70415.0 ;
      RECT  67250.0 71760.0 67955.0 70415.0 ;
      RECT  67250.0 71760.0 67955.0 73105.0 ;
      RECT  67250.0 74450.0 67955.0 73105.0 ;
      RECT  67250.0 74450.0 67955.0 75795.0 ;
      RECT  67250.0 77140.0 67955.0 75795.0 ;
      RECT  67250.0 77140.0 67955.0 78485.0 ;
      RECT  67250.0 79830.0 67955.0 78485.0 ;
      RECT  67250.0 79830.0 67955.0 81175.0 ;
      RECT  67250.0 82520.0 67955.0 81175.0 ;
      RECT  67250.0 82520.0 67955.0 83865.0 ;
      RECT  67250.0 85210.0 67955.0 83865.0 ;
      RECT  67250.0 85210.0 67955.0 86555.0 ;
      RECT  67250.0 87900.0 67955.0 86555.0 ;
      RECT  67250.0 87900.0 67955.0 89245.0 ;
      RECT  67250.0 90590.0 67955.0 89245.0 ;
      RECT  67250.0 90590.0 67955.0 91935.0 ;
      RECT  67250.0 93280.0 67955.0 91935.0 ;
      RECT  67250.0 93280.0 67955.0 94625.0 ;
      RECT  67250.0 95970.0 67955.0 94625.0 ;
      RECT  67250.0 95970.0 67955.0 97315.0 ;
      RECT  67250.0 98660.0 67955.0 97315.0 ;
      RECT  67250.0 98660.0 67955.0 100005.0 ;
      RECT  67250.0 101350.0 67955.0 100005.0 ;
      RECT  67250.0 101350.0 67955.0 102695.0 ;
      RECT  67250.0 104040.0 67955.0 102695.0 ;
      RECT  67250.0 104040.0 67955.0 105385.0 ;
      RECT  67250.0 106730.0 67955.0 105385.0 ;
      RECT  67250.0 106730.0 67955.0 108075.0 ;
      RECT  67250.0 109420.0 67955.0 108075.0 ;
      RECT  67250.0 109420.0 67955.0 110765.0 ;
      RECT  67250.0 112110.0 67955.0 110765.0 ;
      RECT  67250.0 112110.0 67955.0 113455.0 ;
      RECT  67250.0 114800.0 67955.0 113455.0 ;
      RECT  67250.0 114800.0 67955.0 116145.0 ;
      RECT  67250.0 117490.0 67955.0 116145.0 ;
      RECT  67250.0 117490.0 67955.0 118835.0 ;
      RECT  67250.0 120180.0 67955.0 118835.0 ;
      RECT  67250.0 120180.0 67955.0 121525.0 ;
      RECT  67250.0 122870.0 67955.0 121525.0 ;
      RECT  67250.0 122870.0 67955.0 124215.0 ;
      RECT  67250.0 125560.0 67955.0 124215.0 ;
      RECT  67250.0 125560.0 67955.0 126905.0 ;
      RECT  67250.0 128250.0 67955.0 126905.0 ;
      RECT  67250.0 128250.0 67955.0 129595.0 ;
      RECT  67250.0 130940.0 67955.0 129595.0 ;
      RECT  67250.0 130940.0 67955.0 132285.0 ;
      RECT  67250.0 133630.0 67955.0 132285.0 ;
      RECT  67250.0 133630.0 67955.0 134975.0 ;
      RECT  67250.0 136320.0 67955.0 134975.0 ;
      RECT  67250.0 136320.0 67955.0 137665.0 ;
      RECT  67250.0 139010.0 67955.0 137665.0 ;
      RECT  67250.0 139010.0 67955.0 140355.0 ;
      RECT  67250.0 141700.0 67955.0 140355.0 ;
      RECT  67250.0 141700.0 67955.0 143045.0 ;
      RECT  67250.0 144390.0 67955.0 143045.0 ;
      RECT  67250.0 144390.0 67955.0 145735.0 ;
      RECT  67250.0 147080.0 67955.0 145735.0 ;
      RECT  67250.0 147080.0 67955.0 148425.0 ;
      RECT  67250.0 149770.0 67955.0 148425.0 ;
      RECT  67250.0 149770.0 67955.0 151115.0 ;
      RECT  67250.0 152460.0 67955.0 151115.0 ;
      RECT  67250.0 152460.0 67955.0 153805.0 ;
      RECT  67250.0 155150.0 67955.0 153805.0 ;
      RECT  67250.0 155150.0 67955.0 156495.0 ;
      RECT  67250.0 157840.0 67955.0 156495.0 ;
      RECT  67250.0 157840.0 67955.0 159185.0 ;
      RECT  67250.0 160530.0 67955.0 159185.0 ;
      RECT  67250.0 160530.0 67955.0 161875.0 ;
      RECT  67250.0 163220.0 67955.0 161875.0 ;
      RECT  67250.0 163220.0 67955.0 164565.0 ;
      RECT  67250.0 165910.0 67955.0 164565.0 ;
      RECT  67250.0 165910.0 67955.0 167255.0 ;
      RECT  67250.0 168600.0 67955.0 167255.0 ;
      RECT  67250.0 168600.0 67955.0 169945.0 ;
      RECT  67250.0 171290.0 67955.0 169945.0 ;
      RECT  67250.0 171290.0 67955.0 172635.0 ;
      RECT  67250.0 173980.0 67955.0 172635.0 ;
      RECT  67250.0 173980.0 67955.0 175325.0 ;
      RECT  67250.0 176670.0 67955.0 175325.0 ;
      RECT  67250.0 176670.0 67955.0 178015.0 ;
      RECT  67250.0 179360.0 67955.0 178015.0 ;
      RECT  67250.0 179360.0 67955.0 180705.0 ;
      RECT  67250.0 182050.0 67955.0 180705.0 ;
      RECT  67250.0 182050.0 67955.0 183395.0 ;
      RECT  67250.0 184740.0 67955.0 183395.0 ;
      RECT  67250.0 184740.0 67955.0 186085.0 ;
      RECT  67250.0 187430.0 67955.0 186085.0 ;
      RECT  67250.0 187430.0 67955.0 188775.0 ;
      RECT  67250.0 190120.0 67955.0 188775.0 ;
      RECT  67250.0 190120.0 67955.0 191465.0 ;
      RECT  67250.0 192810.0 67955.0 191465.0 ;
      RECT  67250.0 192810.0 67955.0 194155.0 ;
      RECT  67250.0 195500.0 67955.0 194155.0 ;
      RECT  67250.0 195500.0 67955.0 196845.0 ;
      RECT  67250.0 198190.0 67955.0 196845.0 ;
      RECT  67250.0 198190.0 67955.0 199535.0 ;
      RECT  67250.0 200880.0 67955.0 199535.0 ;
      RECT  67250.0 200880.0 67955.0 202225.0 ;
      RECT  67250.0 203570.0 67955.0 202225.0 ;
      RECT  67250.0 203570.0 67955.0 204915.0 ;
      RECT  67250.0 206260.0 67955.0 204915.0 ;
      RECT  67955.0 34100.0 68660.0 35445.0 ;
      RECT  67955.0 36790.0 68660.0 35445.0 ;
      RECT  67955.0 36790.0 68660.0 38135.0 ;
      RECT  67955.0 39480.0 68660.0 38135.0 ;
      RECT  67955.0 39480.0 68660.0 40825.0 ;
      RECT  67955.0 42170.0 68660.0 40825.0 ;
      RECT  67955.0 42170.0 68660.0 43515.0 ;
      RECT  67955.0 44860.0 68660.0 43515.0 ;
      RECT  67955.0 44860.0 68660.0 46205.0 ;
      RECT  67955.0 47550.0 68660.0 46205.0 ;
      RECT  67955.0 47550.0 68660.0 48895.0 ;
      RECT  67955.0 50240.0 68660.0 48895.0 ;
      RECT  67955.0 50240.0 68660.0 51585.0 ;
      RECT  67955.0 52930.0 68660.0 51585.0 ;
      RECT  67955.0 52930.0 68660.0 54275.0 ;
      RECT  67955.0 55620.0 68660.0 54275.0 ;
      RECT  67955.0 55620.0 68660.0 56965.0 ;
      RECT  67955.0 58310.0 68660.0 56965.0 ;
      RECT  67955.0 58310.0 68660.0 59655.0 ;
      RECT  67955.0 61000.0 68660.0 59655.0 ;
      RECT  67955.0 61000.0 68660.0 62345.0 ;
      RECT  67955.0 63690.0 68660.0 62345.0 ;
      RECT  67955.0 63690.0 68660.0 65035.0 ;
      RECT  67955.0 66380.0 68660.0 65035.0 ;
      RECT  67955.0 66380.0 68660.0 67725.0 ;
      RECT  67955.0 69070.0 68660.0 67725.0 ;
      RECT  67955.0 69070.0 68660.0 70415.0 ;
      RECT  67955.0 71760.0 68660.0 70415.0 ;
      RECT  67955.0 71760.0 68660.0 73105.0 ;
      RECT  67955.0 74450.0 68660.0 73105.0 ;
      RECT  67955.0 74450.0 68660.0 75795.0 ;
      RECT  67955.0 77140.0 68660.0 75795.0 ;
      RECT  67955.0 77140.0 68660.0 78485.0 ;
      RECT  67955.0 79830.0 68660.0 78485.0 ;
      RECT  67955.0 79830.0 68660.0 81175.0 ;
      RECT  67955.0 82520.0 68660.0 81175.0 ;
      RECT  67955.0 82520.0 68660.0 83865.0 ;
      RECT  67955.0 85210.0 68660.0 83865.0 ;
      RECT  67955.0 85210.0 68660.0 86555.0 ;
      RECT  67955.0 87900.0 68660.0 86555.0 ;
      RECT  67955.0 87900.0 68660.0 89245.0 ;
      RECT  67955.0 90590.0 68660.0 89245.0 ;
      RECT  67955.0 90590.0 68660.0 91935.0 ;
      RECT  67955.0 93280.0 68660.0 91935.0 ;
      RECT  67955.0 93280.0 68660.0 94625.0 ;
      RECT  67955.0 95970.0 68660.0 94625.0 ;
      RECT  67955.0 95970.0 68660.0 97315.0 ;
      RECT  67955.0 98660.0 68660.0 97315.0 ;
      RECT  67955.0 98660.0 68660.0 100005.0 ;
      RECT  67955.0 101350.0 68660.0 100005.0 ;
      RECT  67955.0 101350.0 68660.0 102695.0 ;
      RECT  67955.0 104040.0 68660.0 102695.0 ;
      RECT  67955.0 104040.0 68660.0 105385.0 ;
      RECT  67955.0 106730.0 68660.0 105385.0 ;
      RECT  67955.0 106730.0 68660.0 108075.0 ;
      RECT  67955.0 109420.0 68660.0 108075.0 ;
      RECT  67955.0 109420.0 68660.0 110765.0 ;
      RECT  67955.0 112110.0 68660.0 110765.0 ;
      RECT  67955.0 112110.0 68660.0 113455.0 ;
      RECT  67955.0 114800.0 68660.0 113455.0 ;
      RECT  67955.0 114800.0 68660.0 116145.0 ;
      RECT  67955.0 117490.0 68660.0 116145.0 ;
      RECT  67955.0 117490.0 68660.0 118835.0 ;
      RECT  67955.0 120180.0 68660.0 118835.0 ;
      RECT  67955.0 120180.0 68660.0 121525.0 ;
      RECT  67955.0 122870.0 68660.0 121525.0 ;
      RECT  67955.0 122870.0 68660.0 124215.0 ;
      RECT  67955.0 125560.0 68660.0 124215.0 ;
      RECT  67955.0 125560.0 68660.0 126905.0 ;
      RECT  67955.0 128250.0 68660.0 126905.0 ;
      RECT  67955.0 128250.0 68660.0 129595.0 ;
      RECT  67955.0 130940.0 68660.0 129595.0 ;
      RECT  67955.0 130940.0 68660.0 132285.0 ;
      RECT  67955.0 133630.0 68660.0 132285.0 ;
      RECT  67955.0 133630.0 68660.0 134975.0 ;
      RECT  67955.0 136320.0 68660.0 134975.0 ;
      RECT  67955.0 136320.0 68660.0 137665.0 ;
      RECT  67955.0 139010.0 68660.0 137665.0 ;
      RECT  67955.0 139010.0 68660.0 140355.0 ;
      RECT  67955.0 141700.0 68660.0 140355.0 ;
      RECT  67955.0 141700.0 68660.0 143045.0 ;
      RECT  67955.0 144390.0 68660.0 143045.0 ;
      RECT  67955.0 144390.0 68660.0 145735.0 ;
      RECT  67955.0 147080.0 68660.0 145735.0 ;
      RECT  67955.0 147080.0 68660.0 148425.0 ;
      RECT  67955.0 149770.0 68660.0 148425.0 ;
      RECT  67955.0 149770.0 68660.0 151115.0 ;
      RECT  67955.0 152460.0 68660.0 151115.0 ;
      RECT  67955.0 152460.0 68660.0 153805.0 ;
      RECT  67955.0 155150.0 68660.0 153805.0 ;
      RECT  67955.0 155150.0 68660.0 156495.0 ;
      RECT  67955.0 157840.0 68660.0 156495.0 ;
      RECT  67955.0 157840.0 68660.0 159185.0 ;
      RECT  67955.0 160530.0 68660.0 159185.0 ;
      RECT  67955.0 160530.0 68660.0 161875.0 ;
      RECT  67955.0 163220.0 68660.0 161875.0 ;
      RECT  67955.0 163220.0 68660.0 164565.0 ;
      RECT  67955.0 165910.0 68660.0 164565.0 ;
      RECT  67955.0 165910.0 68660.0 167255.0 ;
      RECT  67955.0 168600.0 68660.0 167255.0 ;
      RECT  67955.0 168600.0 68660.0 169945.0 ;
      RECT  67955.0 171290.0 68660.0 169945.0 ;
      RECT  67955.0 171290.0 68660.0 172635.0 ;
      RECT  67955.0 173980.0 68660.0 172635.0 ;
      RECT  67955.0 173980.0 68660.0 175325.0 ;
      RECT  67955.0 176670.0 68660.0 175325.0 ;
      RECT  67955.0 176670.0 68660.0 178015.0 ;
      RECT  67955.0 179360.0 68660.0 178015.0 ;
      RECT  67955.0 179360.0 68660.0 180705.0 ;
      RECT  67955.0 182050.0 68660.0 180705.0 ;
      RECT  67955.0 182050.0 68660.0 183395.0 ;
      RECT  67955.0 184740.0 68660.0 183395.0 ;
      RECT  67955.0 184740.0 68660.0 186085.0 ;
      RECT  67955.0 187430.0 68660.0 186085.0 ;
      RECT  67955.0 187430.0 68660.0 188775.0 ;
      RECT  67955.0 190120.0 68660.0 188775.0 ;
      RECT  67955.0 190120.0 68660.0 191465.0 ;
      RECT  67955.0 192810.0 68660.0 191465.0 ;
      RECT  67955.0 192810.0 68660.0 194155.0 ;
      RECT  67955.0 195500.0 68660.0 194155.0 ;
      RECT  67955.0 195500.0 68660.0 196845.0 ;
      RECT  67955.0 198190.0 68660.0 196845.0 ;
      RECT  67955.0 198190.0 68660.0 199535.0 ;
      RECT  67955.0 200880.0 68660.0 199535.0 ;
      RECT  67955.0 200880.0 68660.0 202225.0 ;
      RECT  67955.0 203570.0 68660.0 202225.0 ;
      RECT  67955.0 203570.0 68660.0 204915.0 ;
      RECT  67955.0 206260.0 68660.0 204915.0 ;
      RECT  68660.0 34100.0 69365.0 35445.0 ;
      RECT  68660.0 36790.0 69365.0 35445.0 ;
      RECT  68660.0 36790.0 69365.0 38135.0 ;
      RECT  68660.0 39480.0 69365.0 38135.0 ;
      RECT  68660.0 39480.0 69365.0 40825.0 ;
      RECT  68660.0 42170.0 69365.0 40825.0 ;
      RECT  68660.0 42170.0 69365.0 43515.0 ;
      RECT  68660.0 44860.0 69365.0 43515.0 ;
      RECT  68660.0 44860.0 69365.0 46205.0 ;
      RECT  68660.0 47550.0 69365.0 46205.0 ;
      RECT  68660.0 47550.0 69365.0 48895.0 ;
      RECT  68660.0 50240.0 69365.0 48895.0 ;
      RECT  68660.0 50240.0 69365.0 51585.0 ;
      RECT  68660.0 52930.0 69365.0 51585.0 ;
      RECT  68660.0 52930.0 69365.0 54275.0 ;
      RECT  68660.0 55620.0 69365.0 54275.0 ;
      RECT  68660.0 55620.0 69365.0 56965.0 ;
      RECT  68660.0 58310.0 69365.0 56965.0 ;
      RECT  68660.0 58310.0 69365.0 59655.0 ;
      RECT  68660.0 61000.0 69365.0 59655.0 ;
      RECT  68660.0 61000.0 69365.0 62345.0 ;
      RECT  68660.0 63690.0 69365.0 62345.0 ;
      RECT  68660.0 63690.0 69365.0 65035.0 ;
      RECT  68660.0 66380.0 69365.0 65035.0 ;
      RECT  68660.0 66380.0 69365.0 67725.0 ;
      RECT  68660.0 69070.0 69365.0 67725.0 ;
      RECT  68660.0 69070.0 69365.0 70415.0 ;
      RECT  68660.0 71760.0 69365.0 70415.0 ;
      RECT  68660.0 71760.0 69365.0 73105.0 ;
      RECT  68660.0 74450.0 69365.0 73105.0 ;
      RECT  68660.0 74450.0 69365.0 75795.0 ;
      RECT  68660.0 77140.0 69365.0 75795.0 ;
      RECT  68660.0 77140.0 69365.0 78485.0 ;
      RECT  68660.0 79830.0 69365.0 78485.0 ;
      RECT  68660.0 79830.0 69365.0 81175.0 ;
      RECT  68660.0 82520.0 69365.0 81175.0 ;
      RECT  68660.0 82520.0 69365.0 83865.0 ;
      RECT  68660.0 85210.0 69365.0 83865.0 ;
      RECT  68660.0 85210.0 69365.0 86555.0 ;
      RECT  68660.0 87900.0 69365.0 86555.0 ;
      RECT  68660.0 87900.0 69365.0 89245.0 ;
      RECT  68660.0 90590.0 69365.0 89245.0 ;
      RECT  68660.0 90590.0 69365.0 91935.0 ;
      RECT  68660.0 93280.0 69365.0 91935.0 ;
      RECT  68660.0 93280.0 69365.0 94625.0 ;
      RECT  68660.0 95970.0 69365.0 94625.0 ;
      RECT  68660.0 95970.0 69365.0 97315.0 ;
      RECT  68660.0 98660.0 69365.0 97315.0 ;
      RECT  68660.0 98660.0 69365.0 100005.0 ;
      RECT  68660.0 101350.0 69365.0 100005.0 ;
      RECT  68660.0 101350.0 69365.0 102695.0 ;
      RECT  68660.0 104040.0 69365.0 102695.0 ;
      RECT  68660.0 104040.0 69365.0 105385.0 ;
      RECT  68660.0 106730.0 69365.0 105385.0 ;
      RECT  68660.0 106730.0 69365.0 108075.0 ;
      RECT  68660.0 109420.0 69365.0 108075.0 ;
      RECT  68660.0 109420.0 69365.0 110765.0 ;
      RECT  68660.0 112110.0 69365.0 110765.0 ;
      RECT  68660.0 112110.0 69365.0 113455.0 ;
      RECT  68660.0 114800.0 69365.0 113455.0 ;
      RECT  68660.0 114800.0 69365.0 116145.0 ;
      RECT  68660.0 117490.0 69365.0 116145.0 ;
      RECT  68660.0 117490.0 69365.0 118835.0 ;
      RECT  68660.0 120180.0 69365.0 118835.0 ;
      RECT  68660.0 120180.0 69365.0 121525.0 ;
      RECT  68660.0 122870.0 69365.0 121525.0 ;
      RECT  68660.0 122870.0 69365.0 124215.0 ;
      RECT  68660.0 125560.0 69365.0 124215.0 ;
      RECT  68660.0 125560.0 69365.0 126905.0 ;
      RECT  68660.0 128250.0 69365.0 126905.0 ;
      RECT  68660.0 128250.0 69365.0 129595.0 ;
      RECT  68660.0 130940.0 69365.0 129595.0 ;
      RECT  68660.0 130940.0 69365.0 132285.0 ;
      RECT  68660.0 133630.0 69365.0 132285.0 ;
      RECT  68660.0 133630.0 69365.0 134975.0 ;
      RECT  68660.0 136320.0 69365.0 134975.0 ;
      RECT  68660.0 136320.0 69365.0 137665.0 ;
      RECT  68660.0 139010.0 69365.0 137665.0 ;
      RECT  68660.0 139010.0 69365.0 140355.0 ;
      RECT  68660.0 141700.0 69365.0 140355.0 ;
      RECT  68660.0 141700.0 69365.0 143045.0 ;
      RECT  68660.0 144390.0 69365.0 143045.0 ;
      RECT  68660.0 144390.0 69365.0 145735.0 ;
      RECT  68660.0 147080.0 69365.0 145735.0 ;
      RECT  68660.0 147080.0 69365.0 148425.0 ;
      RECT  68660.0 149770.0 69365.0 148425.0 ;
      RECT  68660.0 149770.0 69365.0 151115.0 ;
      RECT  68660.0 152460.0 69365.0 151115.0 ;
      RECT  68660.0 152460.0 69365.0 153805.0 ;
      RECT  68660.0 155150.0 69365.0 153805.0 ;
      RECT  68660.0 155150.0 69365.0 156495.0 ;
      RECT  68660.0 157840.0 69365.0 156495.0 ;
      RECT  68660.0 157840.0 69365.0 159185.0 ;
      RECT  68660.0 160530.0 69365.0 159185.0 ;
      RECT  68660.0 160530.0 69365.0 161875.0 ;
      RECT  68660.0 163220.0 69365.0 161875.0 ;
      RECT  68660.0 163220.0 69365.0 164565.0 ;
      RECT  68660.0 165910.0 69365.0 164565.0 ;
      RECT  68660.0 165910.0 69365.0 167255.0 ;
      RECT  68660.0 168600.0 69365.0 167255.0 ;
      RECT  68660.0 168600.0 69365.0 169945.0 ;
      RECT  68660.0 171290.0 69365.0 169945.0 ;
      RECT  68660.0 171290.0 69365.0 172635.0 ;
      RECT  68660.0 173980.0 69365.0 172635.0 ;
      RECT  68660.0 173980.0 69365.0 175325.0 ;
      RECT  68660.0 176670.0 69365.0 175325.0 ;
      RECT  68660.0 176670.0 69365.0 178015.0 ;
      RECT  68660.0 179360.0 69365.0 178015.0 ;
      RECT  68660.0 179360.0 69365.0 180705.0 ;
      RECT  68660.0 182050.0 69365.0 180705.0 ;
      RECT  68660.0 182050.0 69365.0 183395.0 ;
      RECT  68660.0 184740.0 69365.0 183395.0 ;
      RECT  68660.0 184740.0 69365.0 186085.0 ;
      RECT  68660.0 187430.0 69365.0 186085.0 ;
      RECT  68660.0 187430.0 69365.0 188775.0 ;
      RECT  68660.0 190120.0 69365.0 188775.0 ;
      RECT  68660.0 190120.0 69365.0 191465.0 ;
      RECT  68660.0 192810.0 69365.0 191465.0 ;
      RECT  68660.0 192810.0 69365.0 194155.0 ;
      RECT  68660.0 195500.0 69365.0 194155.0 ;
      RECT  68660.0 195500.0 69365.0 196845.0 ;
      RECT  68660.0 198190.0 69365.0 196845.0 ;
      RECT  68660.0 198190.0 69365.0 199535.0 ;
      RECT  68660.0 200880.0 69365.0 199535.0 ;
      RECT  68660.0 200880.0 69365.0 202225.0 ;
      RECT  68660.0 203570.0 69365.0 202225.0 ;
      RECT  68660.0 203570.0 69365.0 204915.0 ;
      RECT  68660.0 206260.0 69365.0 204915.0 ;
      RECT  69365.0 34100.0 70070.0 35445.0 ;
      RECT  69365.0 36790.0 70070.0 35445.0 ;
      RECT  69365.0 36790.0 70070.0 38135.0 ;
      RECT  69365.0 39480.0 70070.0 38135.0 ;
      RECT  69365.0 39480.0 70070.0 40825.0 ;
      RECT  69365.0 42170.0 70070.0 40825.0 ;
      RECT  69365.0 42170.0 70070.0 43515.0 ;
      RECT  69365.0 44860.0 70070.0 43515.0 ;
      RECT  69365.0 44860.0 70070.0 46205.0 ;
      RECT  69365.0 47550.0 70070.0 46205.0 ;
      RECT  69365.0 47550.0 70070.0 48895.0 ;
      RECT  69365.0 50240.0 70070.0 48895.0 ;
      RECT  69365.0 50240.0 70070.0 51585.0 ;
      RECT  69365.0 52930.0 70070.0 51585.0 ;
      RECT  69365.0 52930.0 70070.0 54275.0 ;
      RECT  69365.0 55620.0 70070.0 54275.0 ;
      RECT  69365.0 55620.0 70070.0 56965.0 ;
      RECT  69365.0 58310.0 70070.0 56965.0 ;
      RECT  69365.0 58310.0 70070.0 59655.0 ;
      RECT  69365.0 61000.0 70070.0 59655.0 ;
      RECT  69365.0 61000.0 70070.0 62345.0 ;
      RECT  69365.0 63690.0 70070.0 62345.0 ;
      RECT  69365.0 63690.0 70070.0 65035.0 ;
      RECT  69365.0 66380.0 70070.0 65035.0 ;
      RECT  69365.0 66380.0 70070.0 67725.0 ;
      RECT  69365.0 69070.0 70070.0 67725.0 ;
      RECT  69365.0 69070.0 70070.0 70415.0 ;
      RECT  69365.0 71760.0 70070.0 70415.0 ;
      RECT  69365.0 71760.0 70070.0 73105.0 ;
      RECT  69365.0 74450.0 70070.0 73105.0 ;
      RECT  69365.0 74450.0 70070.0 75795.0 ;
      RECT  69365.0 77140.0 70070.0 75795.0 ;
      RECT  69365.0 77140.0 70070.0 78485.0 ;
      RECT  69365.0 79830.0 70070.0 78485.0 ;
      RECT  69365.0 79830.0 70070.0 81175.0 ;
      RECT  69365.0 82520.0 70070.0 81175.0 ;
      RECT  69365.0 82520.0 70070.0 83865.0 ;
      RECT  69365.0 85210.0 70070.0 83865.0 ;
      RECT  69365.0 85210.0 70070.0 86555.0 ;
      RECT  69365.0 87900.0 70070.0 86555.0 ;
      RECT  69365.0 87900.0 70070.0 89245.0 ;
      RECT  69365.0 90590.0 70070.0 89245.0 ;
      RECT  69365.0 90590.0 70070.0 91935.0 ;
      RECT  69365.0 93280.0 70070.0 91935.0 ;
      RECT  69365.0 93280.0 70070.0 94625.0 ;
      RECT  69365.0 95970.0 70070.0 94625.0 ;
      RECT  69365.0 95970.0 70070.0 97315.0 ;
      RECT  69365.0 98660.0 70070.0 97315.0 ;
      RECT  69365.0 98660.0 70070.0 100005.0 ;
      RECT  69365.0 101350.0 70070.0 100005.0 ;
      RECT  69365.0 101350.0 70070.0 102695.0 ;
      RECT  69365.0 104040.0 70070.0 102695.0 ;
      RECT  69365.0 104040.0 70070.0 105385.0 ;
      RECT  69365.0 106730.0 70070.0 105385.0 ;
      RECT  69365.0 106730.0 70070.0 108075.0 ;
      RECT  69365.0 109420.0 70070.0 108075.0 ;
      RECT  69365.0 109420.0 70070.0 110765.0 ;
      RECT  69365.0 112110.0 70070.0 110765.0 ;
      RECT  69365.0 112110.0 70070.0 113455.0 ;
      RECT  69365.0 114800.0 70070.0 113455.0 ;
      RECT  69365.0 114800.0 70070.0 116145.0 ;
      RECT  69365.0 117490.0 70070.0 116145.0 ;
      RECT  69365.0 117490.0 70070.0 118835.0 ;
      RECT  69365.0 120180.0 70070.0 118835.0 ;
      RECT  69365.0 120180.0 70070.0 121525.0 ;
      RECT  69365.0 122870.0 70070.0 121525.0 ;
      RECT  69365.0 122870.0 70070.0 124215.0 ;
      RECT  69365.0 125560.0 70070.0 124215.0 ;
      RECT  69365.0 125560.0 70070.0 126905.0 ;
      RECT  69365.0 128250.0 70070.0 126905.0 ;
      RECT  69365.0 128250.0 70070.0 129595.0 ;
      RECT  69365.0 130940.0 70070.0 129595.0 ;
      RECT  69365.0 130940.0 70070.0 132285.0 ;
      RECT  69365.0 133630.0 70070.0 132285.0 ;
      RECT  69365.0 133630.0 70070.0 134975.0 ;
      RECT  69365.0 136320.0 70070.0 134975.0 ;
      RECT  69365.0 136320.0 70070.0 137665.0 ;
      RECT  69365.0 139010.0 70070.0 137665.0 ;
      RECT  69365.0 139010.0 70070.0 140355.0 ;
      RECT  69365.0 141700.0 70070.0 140355.0 ;
      RECT  69365.0 141700.0 70070.0 143045.0 ;
      RECT  69365.0 144390.0 70070.0 143045.0 ;
      RECT  69365.0 144390.0 70070.0 145735.0 ;
      RECT  69365.0 147080.0 70070.0 145735.0 ;
      RECT  69365.0 147080.0 70070.0 148425.0 ;
      RECT  69365.0 149770.0 70070.0 148425.0 ;
      RECT  69365.0 149770.0 70070.0 151115.0 ;
      RECT  69365.0 152460.0 70070.0 151115.0 ;
      RECT  69365.0 152460.0 70070.0 153805.0 ;
      RECT  69365.0 155150.0 70070.0 153805.0 ;
      RECT  69365.0 155150.0 70070.0 156495.0 ;
      RECT  69365.0 157840.0 70070.0 156495.0 ;
      RECT  69365.0 157840.0 70070.0 159185.0 ;
      RECT  69365.0 160530.0 70070.0 159185.0 ;
      RECT  69365.0 160530.0 70070.0 161875.0 ;
      RECT  69365.0 163220.0 70070.0 161875.0 ;
      RECT  69365.0 163220.0 70070.0 164565.0 ;
      RECT  69365.0 165910.0 70070.0 164565.0 ;
      RECT  69365.0 165910.0 70070.0 167255.0 ;
      RECT  69365.0 168600.0 70070.0 167255.0 ;
      RECT  69365.0 168600.0 70070.0 169945.0 ;
      RECT  69365.0 171290.0 70070.0 169945.0 ;
      RECT  69365.0 171290.0 70070.0 172635.0 ;
      RECT  69365.0 173980.0 70070.0 172635.0 ;
      RECT  69365.0 173980.0 70070.0 175325.0 ;
      RECT  69365.0 176670.0 70070.0 175325.0 ;
      RECT  69365.0 176670.0 70070.0 178015.0 ;
      RECT  69365.0 179360.0 70070.0 178015.0 ;
      RECT  69365.0 179360.0 70070.0 180705.0 ;
      RECT  69365.0 182050.0 70070.0 180705.0 ;
      RECT  69365.0 182050.0 70070.0 183395.0 ;
      RECT  69365.0 184740.0 70070.0 183395.0 ;
      RECT  69365.0 184740.0 70070.0 186085.0 ;
      RECT  69365.0 187430.0 70070.0 186085.0 ;
      RECT  69365.0 187430.0 70070.0 188775.0 ;
      RECT  69365.0 190120.0 70070.0 188775.0 ;
      RECT  69365.0 190120.0 70070.0 191465.0 ;
      RECT  69365.0 192810.0 70070.0 191465.0 ;
      RECT  69365.0 192810.0 70070.0 194155.0 ;
      RECT  69365.0 195500.0 70070.0 194155.0 ;
      RECT  69365.0 195500.0 70070.0 196845.0 ;
      RECT  69365.0 198190.0 70070.0 196845.0 ;
      RECT  69365.0 198190.0 70070.0 199535.0 ;
      RECT  69365.0 200880.0 70070.0 199535.0 ;
      RECT  69365.0 200880.0 70070.0 202225.0 ;
      RECT  69365.0 203570.0 70070.0 202225.0 ;
      RECT  69365.0 203570.0 70070.0 204915.0 ;
      RECT  69365.0 206260.0 70070.0 204915.0 ;
      RECT  70070.0 34100.0 70775.0 35445.0 ;
      RECT  70070.0 36790.0 70775.0 35445.0 ;
      RECT  70070.0 36790.0 70775.0 38135.0 ;
      RECT  70070.0 39480.0 70775.0 38135.0 ;
      RECT  70070.0 39480.0 70775.0 40825.0 ;
      RECT  70070.0 42170.0 70775.0 40825.0 ;
      RECT  70070.0 42170.0 70775.0 43515.0 ;
      RECT  70070.0 44860.0 70775.0 43515.0 ;
      RECT  70070.0 44860.0 70775.0 46205.0 ;
      RECT  70070.0 47550.0 70775.0 46205.0 ;
      RECT  70070.0 47550.0 70775.0 48895.0 ;
      RECT  70070.0 50240.0 70775.0 48895.0 ;
      RECT  70070.0 50240.0 70775.0 51585.0 ;
      RECT  70070.0 52930.0 70775.0 51585.0 ;
      RECT  70070.0 52930.0 70775.0 54275.0 ;
      RECT  70070.0 55620.0 70775.0 54275.0 ;
      RECT  70070.0 55620.0 70775.0 56965.0 ;
      RECT  70070.0 58310.0 70775.0 56965.0 ;
      RECT  70070.0 58310.0 70775.0 59655.0 ;
      RECT  70070.0 61000.0 70775.0 59655.0 ;
      RECT  70070.0 61000.0 70775.0 62345.0 ;
      RECT  70070.0 63690.0 70775.0 62345.0 ;
      RECT  70070.0 63690.0 70775.0 65035.0 ;
      RECT  70070.0 66380.0 70775.0 65035.0 ;
      RECT  70070.0 66380.0 70775.0 67725.0 ;
      RECT  70070.0 69070.0 70775.0 67725.0 ;
      RECT  70070.0 69070.0 70775.0 70415.0 ;
      RECT  70070.0 71760.0 70775.0 70415.0 ;
      RECT  70070.0 71760.0 70775.0 73105.0 ;
      RECT  70070.0 74450.0 70775.0 73105.0 ;
      RECT  70070.0 74450.0 70775.0 75795.0 ;
      RECT  70070.0 77140.0 70775.0 75795.0 ;
      RECT  70070.0 77140.0 70775.0 78485.0 ;
      RECT  70070.0 79830.0 70775.0 78485.0 ;
      RECT  70070.0 79830.0 70775.0 81175.0 ;
      RECT  70070.0 82520.0 70775.0 81175.0 ;
      RECT  70070.0 82520.0 70775.0 83865.0 ;
      RECT  70070.0 85210.0 70775.0 83865.0 ;
      RECT  70070.0 85210.0 70775.0 86555.0 ;
      RECT  70070.0 87900.0 70775.0 86555.0 ;
      RECT  70070.0 87900.0 70775.0 89245.0 ;
      RECT  70070.0 90590.0 70775.0 89245.0 ;
      RECT  70070.0 90590.0 70775.0 91935.0 ;
      RECT  70070.0 93280.0 70775.0 91935.0 ;
      RECT  70070.0 93280.0 70775.0 94625.0 ;
      RECT  70070.0 95970.0 70775.0 94625.0 ;
      RECT  70070.0 95970.0 70775.0 97315.0 ;
      RECT  70070.0 98660.0 70775.0 97315.0 ;
      RECT  70070.0 98660.0 70775.0 100005.0 ;
      RECT  70070.0 101350.0 70775.0 100005.0 ;
      RECT  70070.0 101350.0 70775.0 102695.0 ;
      RECT  70070.0 104040.0 70775.0 102695.0 ;
      RECT  70070.0 104040.0 70775.0 105385.0 ;
      RECT  70070.0 106730.0 70775.0 105385.0 ;
      RECT  70070.0 106730.0 70775.0 108075.0 ;
      RECT  70070.0 109420.0 70775.0 108075.0 ;
      RECT  70070.0 109420.0 70775.0 110765.0 ;
      RECT  70070.0 112110.0 70775.0 110765.0 ;
      RECT  70070.0 112110.0 70775.0 113455.0 ;
      RECT  70070.0 114800.0 70775.0 113455.0 ;
      RECT  70070.0 114800.0 70775.0 116145.0 ;
      RECT  70070.0 117490.0 70775.0 116145.0 ;
      RECT  70070.0 117490.0 70775.0 118835.0 ;
      RECT  70070.0 120180.0 70775.0 118835.0 ;
      RECT  70070.0 120180.0 70775.0 121525.0 ;
      RECT  70070.0 122870.0 70775.0 121525.0 ;
      RECT  70070.0 122870.0 70775.0 124215.0 ;
      RECT  70070.0 125560.0 70775.0 124215.0 ;
      RECT  70070.0 125560.0 70775.0 126905.0 ;
      RECT  70070.0 128250.0 70775.0 126905.0 ;
      RECT  70070.0 128250.0 70775.0 129595.0 ;
      RECT  70070.0 130940.0 70775.0 129595.0 ;
      RECT  70070.0 130940.0 70775.0 132285.0 ;
      RECT  70070.0 133630.0 70775.0 132285.0 ;
      RECT  70070.0 133630.0 70775.0 134975.0 ;
      RECT  70070.0 136320.0 70775.0 134975.0 ;
      RECT  70070.0 136320.0 70775.0 137665.0 ;
      RECT  70070.0 139010.0 70775.0 137665.0 ;
      RECT  70070.0 139010.0 70775.0 140355.0 ;
      RECT  70070.0 141700.0 70775.0 140355.0 ;
      RECT  70070.0 141700.0 70775.0 143045.0 ;
      RECT  70070.0 144390.0 70775.0 143045.0 ;
      RECT  70070.0 144390.0 70775.0 145735.0 ;
      RECT  70070.0 147080.0 70775.0 145735.0 ;
      RECT  70070.0 147080.0 70775.0 148425.0 ;
      RECT  70070.0 149770.0 70775.0 148425.0 ;
      RECT  70070.0 149770.0 70775.0 151115.0 ;
      RECT  70070.0 152460.0 70775.0 151115.0 ;
      RECT  70070.0 152460.0 70775.0 153805.0 ;
      RECT  70070.0 155150.0 70775.0 153805.0 ;
      RECT  70070.0 155150.0 70775.0 156495.0 ;
      RECT  70070.0 157840.0 70775.0 156495.0 ;
      RECT  70070.0 157840.0 70775.0 159185.0 ;
      RECT  70070.0 160530.0 70775.0 159185.0 ;
      RECT  70070.0 160530.0 70775.0 161875.0 ;
      RECT  70070.0 163220.0 70775.0 161875.0 ;
      RECT  70070.0 163220.0 70775.0 164565.0 ;
      RECT  70070.0 165910.0 70775.0 164565.0 ;
      RECT  70070.0 165910.0 70775.0 167255.0 ;
      RECT  70070.0 168600.0 70775.0 167255.0 ;
      RECT  70070.0 168600.0 70775.0 169945.0 ;
      RECT  70070.0 171290.0 70775.0 169945.0 ;
      RECT  70070.0 171290.0 70775.0 172635.0 ;
      RECT  70070.0 173980.0 70775.0 172635.0 ;
      RECT  70070.0 173980.0 70775.0 175325.0 ;
      RECT  70070.0 176670.0 70775.0 175325.0 ;
      RECT  70070.0 176670.0 70775.0 178015.0 ;
      RECT  70070.0 179360.0 70775.0 178015.0 ;
      RECT  70070.0 179360.0 70775.0 180705.0 ;
      RECT  70070.0 182050.0 70775.0 180705.0 ;
      RECT  70070.0 182050.0 70775.0 183395.0 ;
      RECT  70070.0 184740.0 70775.0 183395.0 ;
      RECT  70070.0 184740.0 70775.0 186085.0 ;
      RECT  70070.0 187430.0 70775.0 186085.0 ;
      RECT  70070.0 187430.0 70775.0 188775.0 ;
      RECT  70070.0 190120.0 70775.0 188775.0 ;
      RECT  70070.0 190120.0 70775.0 191465.0 ;
      RECT  70070.0 192810.0 70775.0 191465.0 ;
      RECT  70070.0 192810.0 70775.0 194155.0 ;
      RECT  70070.0 195500.0 70775.0 194155.0 ;
      RECT  70070.0 195500.0 70775.0 196845.0 ;
      RECT  70070.0 198190.0 70775.0 196845.0 ;
      RECT  70070.0 198190.0 70775.0 199535.0 ;
      RECT  70070.0 200880.0 70775.0 199535.0 ;
      RECT  70070.0 200880.0 70775.0 202225.0 ;
      RECT  70070.0 203570.0 70775.0 202225.0 ;
      RECT  70070.0 203570.0 70775.0 204915.0 ;
      RECT  70070.0 206260.0 70775.0 204915.0 ;
      RECT  70775.0 34100.0 71480.0 35445.0 ;
      RECT  70775.0 36790.0 71480.0 35445.0 ;
      RECT  70775.0 36790.0 71480.0 38135.0 ;
      RECT  70775.0 39480.0 71480.0 38135.0 ;
      RECT  70775.0 39480.0 71480.0 40825.0 ;
      RECT  70775.0 42170.0 71480.0 40825.0 ;
      RECT  70775.0 42170.0 71480.0 43515.0 ;
      RECT  70775.0 44860.0 71480.0 43515.0 ;
      RECT  70775.0 44860.0 71480.0 46205.0 ;
      RECT  70775.0 47550.0 71480.0 46205.0 ;
      RECT  70775.0 47550.0 71480.0 48895.0 ;
      RECT  70775.0 50240.0 71480.0 48895.0 ;
      RECT  70775.0 50240.0 71480.0 51585.0 ;
      RECT  70775.0 52930.0 71480.0 51585.0 ;
      RECT  70775.0 52930.0 71480.0 54275.0 ;
      RECT  70775.0 55620.0 71480.0 54275.0 ;
      RECT  70775.0 55620.0 71480.0 56965.0 ;
      RECT  70775.0 58310.0 71480.0 56965.0 ;
      RECT  70775.0 58310.0 71480.0 59655.0 ;
      RECT  70775.0 61000.0 71480.0 59655.0 ;
      RECT  70775.0 61000.0 71480.0 62345.0 ;
      RECT  70775.0 63690.0 71480.0 62345.0 ;
      RECT  70775.0 63690.0 71480.0 65035.0 ;
      RECT  70775.0 66380.0 71480.0 65035.0 ;
      RECT  70775.0 66380.0 71480.0 67725.0 ;
      RECT  70775.0 69070.0 71480.0 67725.0 ;
      RECT  70775.0 69070.0 71480.0 70415.0 ;
      RECT  70775.0 71760.0 71480.0 70415.0 ;
      RECT  70775.0 71760.0 71480.0 73105.0 ;
      RECT  70775.0 74450.0 71480.0 73105.0 ;
      RECT  70775.0 74450.0 71480.0 75795.0 ;
      RECT  70775.0 77140.0 71480.0 75795.0 ;
      RECT  70775.0 77140.0 71480.0 78485.0 ;
      RECT  70775.0 79830.0 71480.0 78485.0 ;
      RECT  70775.0 79830.0 71480.0 81175.0 ;
      RECT  70775.0 82520.0 71480.0 81175.0 ;
      RECT  70775.0 82520.0 71480.0 83865.0 ;
      RECT  70775.0 85210.0 71480.0 83865.0 ;
      RECT  70775.0 85210.0 71480.0 86555.0 ;
      RECT  70775.0 87900.0 71480.0 86555.0 ;
      RECT  70775.0 87900.0 71480.0 89245.0 ;
      RECT  70775.0 90590.0 71480.0 89245.0 ;
      RECT  70775.0 90590.0 71480.0 91935.0 ;
      RECT  70775.0 93280.0 71480.0 91935.0 ;
      RECT  70775.0 93280.0 71480.0 94625.0 ;
      RECT  70775.0 95970.0 71480.0 94625.0 ;
      RECT  70775.0 95970.0 71480.0 97315.0 ;
      RECT  70775.0 98660.0 71480.0 97315.0 ;
      RECT  70775.0 98660.0 71480.0 100005.0 ;
      RECT  70775.0 101350.0 71480.0 100005.0 ;
      RECT  70775.0 101350.0 71480.0 102695.0 ;
      RECT  70775.0 104040.0 71480.0 102695.0 ;
      RECT  70775.0 104040.0 71480.0 105385.0 ;
      RECT  70775.0 106730.0 71480.0 105385.0 ;
      RECT  70775.0 106730.0 71480.0 108075.0 ;
      RECT  70775.0 109420.0 71480.0 108075.0 ;
      RECT  70775.0 109420.0 71480.0 110765.0 ;
      RECT  70775.0 112110.0 71480.0 110765.0 ;
      RECT  70775.0 112110.0 71480.0 113455.0 ;
      RECT  70775.0 114800.0 71480.0 113455.0 ;
      RECT  70775.0 114800.0 71480.0 116145.0 ;
      RECT  70775.0 117490.0 71480.0 116145.0 ;
      RECT  70775.0 117490.0 71480.0 118835.0 ;
      RECT  70775.0 120180.0 71480.0 118835.0 ;
      RECT  70775.0 120180.0 71480.0 121525.0 ;
      RECT  70775.0 122870.0 71480.0 121525.0 ;
      RECT  70775.0 122870.0 71480.0 124215.0 ;
      RECT  70775.0 125560.0 71480.0 124215.0 ;
      RECT  70775.0 125560.0 71480.0 126905.0 ;
      RECT  70775.0 128250.0 71480.0 126905.0 ;
      RECT  70775.0 128250.0 71480.0 129595.0 ;
      RECT  70775.0 130940.0 71480.0 129595.0 ;
      RECT  70775.0 130940.0 71480.0 132285.0 ;
      RECT  70775.0 133630.0 71480.0 132285.0 ;
      RECT  70775.0 133630.0 71480.0 134975.0 ;
      RECT  70775.0 136320.0 71480.0 134975.0 ;
      RECT  70775.0 136320.0 71480.0 137665.0 ;
      RECT  70775.0 139010.0 71480.0 137665.0 ;
      RECT  70775.0 139010.0 71480.0 140355.0 ;
      RECT  70775.0 141700.0 71480.0 140355.0 ;
      RECT  70775.0 141700.0 71480.0 143045.0 ;
      RECT  70775.0 144390.0 71480.0 143045.0 ;
      RECT  70775.0 144390.0 71480.0 145735.0 ;
      RECT  70775.0 147080.0 71480.0 145735.0 ;
      RECT  70775.0 147080.0 71480.0 148425.0 ;
      RECT  70775.0 149770.0 71480.0 148425.0 ;
      RECT  70775.0 149770.0 71480.0 151115.0 ;
      RECT  70775.0 152460.0 71480.0 151115.0 ;
      RECT  70775.0 152460.0 71480.0 153805.0 ;
      RECT  70775.0 155150.0 71480.0 153805.0 ;
      RECT  70775.0 155150.0 71480.0 156495.0 ;
      RECT  70775.0 157840.0 71480.0 156495.0 ;
      RECT  70775.0 157840.0 71480.0 159185.0 ;
      RECT  70775.0 160530.0 71480.0 159185.0 ;
      RECT  70775.0 160530.0 71480.0 161875.0 ;
      RECT  70775.0 163220.0 71480.0 161875.0 ;
      RECT  70775.0 163220.0 71480.0 164565.0 ;
      RECT  70775.0 165910.0 71480.0 164565.0 ;
      RECT  70775.0 165910.0 71480.0 167255.0 ;
      RECT  70775.0 168600.0 71480.0 167255.0 ;
      RECT  70775.0 168600.0 71480.0 169945.0 ;
      RECT  70775.0 171290.0 71480.0 169945.0 ;
      RECT  70775.0 171290.0 71480.0 172635.0 ;
      RECT  70775.0 173980.0 71480.0 172635.0 ;
      RECT  70775.0 173980.0 71480.0 175325.0 ;
      RECT  70775.0 176670.0 71480.0 175325.0 ;
      RECT  70775.0 176670.0 71480.0 178015.0 ;
      RECT  70775.0 179360.0 71480.0 178015.0 ;
      RECT  70775.0 179360.0 71480.0 180705.0 ;
      RECT  70775.0 182050.0 71480.0 180705.0 ;
      RECT  70775.0 182050.0 71480.0 183395.0 ;
      RECT  70775.0 184740.0 71480.0 183395.0 ;
      RECT  70775.0 184740.0 71480.0 186085.0 ;
      RECT  70775.0 187430.0 71480.0 186085.0 ;
      RECT  70775.0 187430.0 71480.0 188775.0 ;
      RECT  70775.0 190120.0 71480.0 188775.0 ;
      RECT  70775.0 190120.0 71480.0 191465.0 ;
      RECT  70775.0 192810.0 71480.0 191465.0 ;
      RECT  70775.0 192810.0 71480.0 194155.0 ;
      RECT  70775.0 195500.0 71480.0 194155.0 ;
      RECT  70775.0 195500.0 71480.0 196845.0 ;
      RECT  70775.0 198190.0 71480.0 196845.0 ;
      RECT  70775.0 198190.0 71480.0 199535.0 ;
      RECT  70775.0 200880.0 71480.0 199535.0 ;
      RECT  70775.0 200880.0 71480.0 202225.0 ;
      RECT  70775.0 203570.0 71480.0 202225.0 ;
      RECT  70775.0 203570.0 71480.0 204915.0 ;
      RECT  70775.0 206260.0 71480.0 204915.0 ;
      RECT  71480.0 34100.0 72185.0 35445.0 ;
      RECT  71480.0 36790.0 72185.0 35445.0 ;
      RECT  71480.0 36790.0 72185.0 38135.0 ;
      RECT  71480.0 39480.0 72185.0 38135.0 ;
      RECT  71480.0 39480.0 72185.0 40825.0 ;
      RECT  71480.0 42170.0 72185.0 40825.0 ;
      RECT  71480.0 42170.0 72185.0 43515.0 ;
      RECT  71480.0 44860.0 72185.0 43515.0 ;
      RECT  71480.0 44860.0 72185.0 46205.0 ;
      RECT  71480.0 47550.0 72185.0 46205.0 ;
      RECT  71480.0 47550.0 72185.0 48895.0 ;
      RECT  71480.0 50240.0 72185.0 48895.0 ;
      RECT  71480.0 50240.0 72185.0 51585.0 ;
      RECT  71480.0 52930.0 72185.0 51585.0 ;
      RECT  71480.0 52930.0 72185.0 54275.0 ;
      RECT  71480.0 55620.0 72185.0 54275.0 ;
      RECT  71480.0 55620.0 72185.0 56965.0 ;
      RECT  71480.0 58310.0 72185.0 56965.0 ;
      RECT  71480.0 58310.0 72185.0 59655.0 ;
      RECT  71480.0 61000.0 72185.0 59655.0 ;
      RECT  71480.0 61000.0 72185.0 62345.0 ;
      RECT  71480.0 63690.0 72185.0 62345.0 ;
      RECT  71480.0 63690.0 72185.0 65035.0 ;
      RECT  71480.0 66380.0 72185.0 65035.0 ;
      RECT  71480.0 66380.0 72185.0 67725.0 ;
      RECT  71480.0 69070.0 72185.0 67725.0 ;
      RECT  71480.0 69070.0 72185.0 70415.0 ;
      RECT  71480.0 71760.0 72185.0 70415.0 ;
      RECT  71480.0 71760.0 72185.0 73105.0 ;
      RECT  71480.0 74450.0 72185.0 73105.0 ;
      RECT  71480.0 74450.0 72185.0 75795.0 ;
      RECT  71480.0 77140.0 72185.0 75795.0 ;
      RECT  71480.0 77140.0 72185.0 78485.0 ;
      RECT  71480.0 79830.0 72185.0 78485.0 ;
      RECT  71480.0 79830.0 72185.0 81175.0 ;
      RECT  71480.0 82520.0 72185.0 81175.0 ;
      RECT  71480.0 82520.0 72185.0 83865.0 ;
      RECT  71480.0 85210.0 72185.0 83865.0 ;
      RECT  71480.0 85210.0 72185.0 86555.0 ;
      RECT  71480.0 87900.0 72185.0 86555.0 ;
      RECT  71480.0 87900.0 72185.0 89245.0 ;
      RECT  71480.0 90590.0 72185.0 89245.0 ;
      RECT  71480.0 90590.0 72185.0 91935.0 ;
      RECT  71480.0 93280.0 72185.0 91935.0 ;
      RECT  71480.0 93280.0 72185.0 94625.0 ;
      RECT  71480.0 95970.0 72185.0 94625.0 ;
      RECT  71480.0 95970.0 72185.0 97315.0 ;
      RECT  71480.0 98660.0 72185.0 97315.0 ;
      RECT  71480.0 98660.0 72185.0 100005.0 ;
      RECT  71480.0 101350.0 72185.0 100005.0 ;
      RECT  71480.0 101350.0 72185.0 102695.0 ;
      RECT  71480.0 104040.0 72185.0 102695.0 ;
      RECT  71480.0 104040.0 72185.0 105385.0 ;
      RECT  71480.0 106730.0 72185.0 105385.0 ;
      RECT  71480.0 106730.0 72185.0 108075.0 ;
      RECT  71480.0 109420.0 72185.0 108075.0 ;
      RECT  71480.0 109420.0 72185.0 110765.0 ;
      RECT  71480.0 112110.0 72185.0 110765.0 ;
      RECT  71480.0 112110.0 72185.0 113455.0 ;
      RECT  71480.0 114800.0 72185.0 113455.0 ;
      RECT  71480.0 114800.0 72185.0 116145.0 ;
      RECT  71480.0 117490.0 72185.0 116145.0 ;
      RECT  71480.0 117490.0 72185.0 118835.0 ;
      RECT  71480.0 120180.0 72185.0 118835.0 ;
      RECT  71480.0 120180.0 72185.0 121525.0 ;
      RECT  71480.0 122870.0 72185.0 121525.0 ;
      RECT  71480.0 122870.0 72185.0 124215.0 ;
      RECT  71480.0 125560.0 72185.0 124215.0 ;
      RECT  71480.0 125560.0 72185.0 126905.0 ;
      RECT  71480.0 128250.0 72185.0 126905.0 ;
      RECT  71480.0 128250.0 72185.0 129595.0 ;
      RECT  71480.0 130940.0 72185.0 129595.0 ;
      RECT  71480.0 130940.0 72185.0 132285.0 ;
      RECT  71480.0 133630.0 72185.0 132285.0 ;
      RECT  71480.0 133630.0 72185.0 134975.0 ;
      RECT  71480.0 136320.0 72185.0 134975.0 ;
      RECT  71480.0 136320.0 72185.0 137665.0 ;
      RECT  71480.0 139010.0 72185.0 137665.0 ;
      RECT  71480.0 139010.0 72185.0 140355.0 ;
      RECT  71480.0 141700.0 72185.0 140355.0 ;
      RECT  71480.0 141700.0 72185.0 143045.0 ;
      RECT  71480.0 144390.0 72185.0 143045.0 ;
      RECT  71480.0 144390.0 72185.0 145735.0 ;
      RECT  71480.0 147080.0 72185.0 145735.0 ;
      RECT  71480.0 147080.0 72185.0 148425.0 ;
      RECT  71480.0 149770.0 72185.0 148425.0 ;
      RECT  71480.0 149770.0 72185.0 151115.0 ;
      RECT  71480.0 152460.0 72185.0 151115.0 ;
      RECT  71480.0 152460.0 72185.0 153805.0 ;
      RECT  71480.0 155150.0 72185.0 153805.0 ;
      RECT  71480.0 155150.0 72185.0 156495.0 ;
      RECT  71480.0 157840.0 72185.0 156495.0 ;
      RECT  71480.0 157840.0 72185.0 159185.0 ;
      RECT  71480.0 160530.0 72185.0 159185.0 ;
      RECT  71480.0 160530.0 72185.0 161875.0 ;
      RECT  71480.0 163220.0 72185.0 161875.0 ;
      RECT  71480.0 163220.0 72185.0 164565.0 ;
      RECT  71480.0 165910.0 72185.0 164565.0 ;
      RECT  71480.0 165910.0 72185.0 167255.0 ;
      RECT  71480.0 168600.0 72185.0 167255.0 ;
      RECT  71480.0 168600.0 72185.0 169945.0 ;
      RECT  71480.0 171290.0 72185.0 169945.0 ;
      RECT  71480.0 171290.0 72185.0 172635.0 ;
      RECT  71480.0 173980.0 72185.0 172635.0 ;
      RECT  71480.0 173980.0 72185.0 175325.0 ;
      RECT  71480.0 176670.0 72185.0 175325.0 ;
      RECT  71480.0 176670.0 72185.0 178015.0 ;
      RECT  71480.0 179360.0 72185.0 178015.0 ;
      RECT  71480.0 179360.0 72185.0 180705.0 ;
      RECT  71480.0 182050.0 72185.0 180705.0 ;
      RECT  71480.0 182050.0 72185.0 183395.0 ;
      RECT  71480.0 184740.0 72185.0 183395.0 ;
      RECT  71480.0 184740.0 72185.0 186085.0 ;
      RECT  71480.0 187430.0 72185.0 186085.0 ;
      RECT  71480.0 187430.0 72185.0 188775.0 ;
      RECT  71480.0 190120.0 72185.0 188775.0 ;
      RECT  71480.0 190120.0 72185.0 191465.0 ;
      RECT  71480.0 192810.0 72185.0 191465.0 ;
      RECT  71480.0 192810.0 72185.0 194155.0 ;
      RECT  71480.0 195500.0 72185.0 194155.0 ;
      RECT  71480.0 195500.0 72185.0 196845.0 ;
      RECT  71480.0 198190.0 72185.0 196845.0 ;
      RECT  71480.0 198190.0 72185.0 199535.0 ;
      RECT  71480.0 200880.0 72185.0 199535.0 ;
      RECT  71480.0 200880.0 72185.0 202225.0 ;
      RECT  71480.0 203570.0 72185.0 202225.0 ;
      RECT  71480.0 203570.0 72185.0 204915.0 ;
      RECT  71480.0 206260.0 72185.0 204915.0 ;
      RECT  72185.0 34100.0 72890.0 35445.0 ;
      RECT  72185.0 36790.0 72890.0 35445.0 ;
      RECT  72185.0 36790.0 72890.0 38135.0 ;
      RECT  72185.0 39480.0 72890.0 38135.0 ;
      RECT  72185.0 39480.0 72890.0 40825.0 ;
      RECT  72185.0 42170.0 72890.0 40825.0 ;
      RECT  72185.0 42170.0 72890.0 43515.0 ;
      RECT  72185.0 44860.0 72890.0 43515.0 ;
      RECT  72185.0 44860.0 72890.0 46205.0 ;
      RECT  72185.0 47550.0 72890.0 46205.0 ;
      RECT  72185.0 47550.0 72890.0 48895.0 ;
      RECT  72185.0 50240.0 72890.0 48895.0 ;
      RECT  72185.0 50240.0 72890.0 51585.0 ;
      RECT  72185.0 52930.0 72890.0 51585.0 ;
      RECT  72185.0 52930.0 72890.0 54275.0 ;
      RECT  72185.0 55620.0 72890.0 54275.0 ;
      RECT  72185.0 55620.0 72890.0 56965.0 ;
      RECT  72185.0 58310.0 72890.0 56965.0 ;
      RECT  72185.0 58310.0 72890.0 59655.0 ;
      RECT  72185.0 61000.0 72890.0 59655.0 ;
      RECT  72185.0 61000.0 72890.0 62345.0 ;
      RECT  72185.0 63690.0 72890.0 62345.0 ;
      RECT  72185.0 63690.0 72890.0 65035.0 ;
      RECT  72185.0 66380.0 72890.0 65035.0 ;
      RECT  72185.0 66380.0 72890.0 67725.0 ;
      RECT  72185.0 69070.0 72890.0 67725.0 ;
      RECT  72185.0 69070.0 72890.0 70415.0 ;
      RECT  72185.0 71760.0 72890.0 70415.0 ;
      RECT  72185.0 71760.0 72890.0 73105.0 ;
      RECT  72185.0 74450.0 72890.0 73105.0 ;
      RECT  72185.0 74450.0 72890.0 75795.0 ;
      RECT  72185.0 77140.0 72890.0 75795.0 ;
      RECT  72185.0 77140.0 72890.0 78485.0 ;
      RECT  72185.0 79830.0 72890.0 78485.0 ;
      RECT  72185.0 79830.0 72890.0 81175.0 ;
      RECT  72185.0 82520.0 72890.0 81175.0 ;
      RECT  72185.0 82520.0 72890.0 83865.0 ;
      RECT  72185.0 85210.0 72890.0 83865.0 ;
      RECT  72185.0 85210.0 72890.0 86555.0 ;
      RECT  72185.0 87900.0 72890.0 86555.0 ;
      RECT  72185.0 87900.0 72890.0 89245.0 ;
      RECT  72185.0 90590.0 72890.0 89245.0 ;
      RECT  72185.0 90590.0 72890.0 91935.0 ;
      RECT  72185.0 93280.0 72890.0 91935.0 ;
      RECT  72185.0 93280.0 72890.0 94625.0 ;
      RECT  72185.0 95970.0 72890.0 94625.0 ;
      RECT  72185.0 95970.0 72890.0 97315.0 ;
      RECT  72185.0 98660.0 72890.0 97315.0 ;
      RECT  72185.0 98660.0 72890.0 100005.0 ;
      RECT  72185.0 101350.0 72890.0 100005.0 ;
      RECT  72185.0 101350.0 72890.0 102695.0 ;
      RECT  72185.0 104040.0 72890.0 102695.0 ;
      RECT  72185.0 104040.0 72890.0 105385.0 ;
      RECT  72185.0 106730.0 72890.0 105385.0 ;
      RECT  72185.0 106730.0 72890.0 108075.0 ;
      RECT  72185.0 109420.0 72890.0 108075.0 ;
      RECT  72185.0 109420.0 72890.0 110765.0 ;
      RECT  72185.0 112110.0 72890.0 110765.0 ;
      RECT  72185.0 112110.0 72890.0 113455.0 ;
      RECT  72185.0 114800.0 72890.0 113455.0 ;
      RECT  72185.0 114800.0 72890.0 116145.0 ;
      RECT  72185.0 117490.0 72890.0 116145.0 ;
      RECT  72185.0 117490.0 72890.0 118835.0 ;
      RECT  72185.0 120180.0 72890.0 118835.0 ;
      RECT  72185.0 120180.0 72890.0 121525.0 ;
      RECT  72185.0 122870.0 72890.0 121525.0 ;
      RECT  72185.0 122870.0 72890.0 124215.0 ;
      RECT  72185.0 125560.0 72890.0 124215.0 ;
      RECT  72185.0 125560.0 72890.0 126905.0 ;
      RECT  72185.0 128250.0 72890.0 126905.0 ;
      RECT  72185.0 128250.0 72890.0 129595.0 ;
      RECT  72185.0 130940.0 72890.0 129595.0 ;
      RECT  72185.0 130940.0 72890.0 132285.0 ;
      RECT  72185.0 133630.0 72890.0 132285.0 ;
      RECT  72185.0 133630.0 72890.0 134975.0 ;
      RECT  72185.0 136320.0 72890.0 134975.0 ;
      RECT  72185.0 136320.0 72890.0 137665.0 ;
      RECT  72185.0 139010.0 72890.0 137665.0 ;
      RECT  72185.0 139010.0 72890.0 140355.0 ;
      RECT  72185.0 141700.0 72890.0 140355.0 ;
      RECT  72185.0 141700.0 72890.0 143045.0 ;
      RECT  72185.0 144390.0 72890.0 143045.0 ;
      RECT  72185.0 144390.0 72890.0 145735.0 ;
      RECT  72185.0 147080.0 72890.0 145735.0 ;
      RECT  72185.0 147080.0 72890.0 148425.0 ;
      RECT  72185.0 149770.0 72890.0 148425.0 ;
      RECT  72185.0 149770.0 72890.0 151115.0 ;
      RECT  72185.0 152460.0 72890.0 151115.0 ;
      RECT  72185.0 152460.0 72890.0 153805.0 ;
      RECT  72185.0 155150.0 72890.0 153805.0 ;
      RECT  72185.0 155150.0 72890.0 156495.0 ;
      RECT  72185.0 157840.0 72890.0 156495.0 ;
      RECT  72185.0 157840.0 72890.0 159185.0 ;
      RECT  72185.0 160530.0 72890.0 159185.0 ;
      RECT  72185.0 160530.0 72890.0 161875.0 ;
      RECT  72185.0 163220.0 72890.0 161875.0 ;
      RECT  72185.0 163220.0 72890.0 164565.0 ;
      RECT  72185.0 165910.0 72890.0 164565.0 ;
      RECT  72185.0 165910.0 72890.0 167255.0 ;
      RECT  72185.0 168600.0 72890.0 167255.0 ;
      RECT  72185.0 168600.0 72890.0 169945.0 ;
      RECT  72185.0 171290.0 72890.0 169945.0 ;
      RECT  72185.0 171290.0 72890.0 172635.0 ;
      RECT  72185.0 173980.0 72890.0 172635.0 ;
      RECT  72185.0 173980.0 72890.0 175325.0 ;
      RECT  72185.0 176670.0 72890.0 175325.0 ;
      RECT  72185.0 176670.0 72890.0 178015.0 ;
      RECT  72185.0 179360.0 72890.0 178015.0 ;
      RECT  72185.0 179360.0 72890.0 180705.0 ;
      RECT  72185.0 182050.0 72890.0 180705.0 ;
      RECT  72185.0 182050.0 72890.0 183395.0 ;
      RECT  72185.0 184740.0 72890.0 183395.0 ;
      RECT  72185.0 184740.0 72890.0 186085.0 ;
      RECT  72185.0 187430.0 72890.0 186085.0 ;
      RECT  72185.0 187430.0 72890.0 188775.0 ;
      RECT  72185.0 190120.0 72890.0 188775.0 ;
      RECT  72185.0 190120.0 72890.0 191465.0 ;
      RECT  72185.0 192810.0 72890.0 191465.0 ;
      RECT  72185.0 192810.0 72890.0 194155.0 ;
      RECT  72185.0 195500.0 72890.0 194155.0 ;
      RECT  72185.0 195500.0 72890.0 196845.0 ;
      RECT  72185.0 198190.0 72890.0 196845.0 ;
      RECT  72185.0 198190.0 72890.0 199535.0 ;
      RECT  72185.0 200880.0 72890.0 199535.0 ;
      RECT  72185.0 200880.0 72890.0 202225.0 ;
      RECT  72185.0 203570.0 72890.0 202225.0 ;
      RECT  72185.0 203570.0 72890.0 204915.0 ;
      RECT  72185.0 206260.0 72890.0 204915.0 ;
      RECT  72890.0 34100.0 73595.0 35445.0 ;
      RECT  72890.0 36790.0 73595.0 35445.0 ;
      RECT  72890.0 36790.0 73595.0 38135.0 ;
      RECT  72890.0 39480.0 73595.0 38135.0 ;
      RECT  72890.0 39480.0 73595.0 40825.0 ;
      RECT  72890.0 42170.0 73595.0 40825.0 ;
      RECT  72890.0 42170.0 73595.0 43515.0 ;
      RECT  72890.0 44860.0 73595.0 43515.0 ;
      RECT  72890.0 44860.0 73595.0 46205.0 ;
      RECT  72890.0 47550.0 73595.0 46205.0 ;
      RECT  72890.0 47550.0 73595.0 48895.0 ;
      RECT  72890.0 50240.0 73595.0 48895.0 ;
      RECT  72890.0 50240.0 73595.0 51585.0 ;
      RECT  72890.0 52930.0 73595.0 51585.0 ;
      RECT  72890.0 52930.0 73595.0 54275.0 ;
      RECT  72890.0 55620.0 73595.0 54275.0 ;
      RECT  72890.0 55620.0 73595.0 56965.0 ;
      RECT  72890.0 58310.0 73595.0 56965.0 ;
      RECT  72890.0 58310.0 73595.0 59655.0 ;
      RECT  72890.0 61000.0 73595.0 59655.0 ;
      RECT  72890.0 61000.0 73595.0 62345.0 ;
      RECT  72890.0 63690.0 73595.0 62345.0 ;
      RECT  72890.0 63690.0 73595.0 65035.0 ;
      RECT  72890.0 66380.0 73595.0 65035.0 ;
      RECT  72890.0 66380.0 73595.0 67725.0 ;
      RECT  72890.0 69070.0 73595.0 67725.0 ;
      RECT  72890.0 69070.0 73595.0 70415.0 ;
      RECT  72890.0 71760.0 73595.0 70415.0 ;
      RECT  72890.0 71760.0 73595.0 73105.0 ;
      RECT  72890.0 74450.0 73595.0 73105.0 ;
      RECT  72890.0 74450.0 73595.0 75795.0 ;
      RECT  72890.0 77140.0 73595.0 75795.0 ;
      RECT  72890.0 77140.0 73595.0 78485.0 ;
      RECT  72890.0 79830.0 73595.0 78485.0 ;
      RECT  72890.0 79830.0 73595.0 81175.0 ;
      RECT  72890.0 82520.0 73595.0 81175.0 ;
      RECT  72890.0 82520.0 73595.0 83865.0 ;
      RECT  72890.0 85210.0 73595.0 83865.0 ;
      RECT  72890.0 85210.0 73595.0 86555.0 ;
      RECT  72890.0 87900.0 73595.0 86555.0 ;
      RECT  72890.0 87900.0 73595.0 89245.0 ;
      RECT  72890.0 90590.0 73595.0 89245.0 ;
      RECT  72890.0 90590.0 73595.0 91935.0 ;
      RECT  72890.0 93280.0 73595.0 91935.0 ;
      RECT  72890.0 93280.0 73595.0 94625.0 ;
      RECT  72890.0 95970.0 73595.0 94625.0 ;
      RECT  72890.0 95970.0 73595.0 97315.0 ;
      RECT  72890.0 98660.0 73595.0 97315.0 ;
      RECT  72890.0 98660.0 73595.0 100005.0 ;
      RECT  72890.0 101350.0 73595.0 100005.0 ;
      RECT  72890.0 101350.0 73595.0 102695.0 ;
      RECT  72890.0 104040.0 73595.0 102695.0 ;
      RECT  72890.0 104040.0 73595.0 105385.0 ;
      RECT  72890.0 106730.0 73595.0 105385.0 ;
      RECT  72890.0 106730.0 73595.0 108075.0 ;
      RECT  72890.0 109420.0 73595.0 108075.0 ;
      RECT  72890.0 109420.0 73595.0 110765.0 ;
      RECT  72890.0 112110.0 73595.0 110765.0 ;
      RECT  72890.0 112110.0 73595.0 113455.0 ;
      RECT  72890.0 114800.0 73595.0 113455.0 ;
      RECT  72890.0 114800.0 73595.0 116145.0 ;
      RECT  72890.0 117490.0 73595.0 116145.0 ;
      RECT  72890.0 117490.0 73595.0 118835.0 ;
      RECT  72890.0 120180.0 73595.0 118835.0 ;
      RECT  72890.0 120180.0 73595.0 121525.0 ;
      RECT  72890.0 122870.0 73595.0 121525.0 ;
      RECT  72890.0 122870.0 73595.0 124215.0 ;
      RECT  72890.0 125560.0 73595.0 124215.0 ;
      RECT  72890.0 125560.0 73595.0 126905.0 ;
      RECT  72890.0 128250.0 73595.0 126905.0 ;
      RECT  72890.0 128250.0 73595.0 129595.0 ;
      RECT  72890.0 130940.0 73595.0 129595.0 ;
      RECT  72890.0 130940.0 73595.0 132285.0 ;
      RECT  72890.0 133630.0 73595.0 132285.0 ;
      RECT  72890.0 133630.0 73595.0 134975.0 ;
      RECT  72890.0 136320.0 73595.0 134975.0 ;
      RECT  72890.0 136320.0 73595.0 137665.0 ;
      RECT  72890.0 139010.0 73595.0 137665.0 ;
      RECT  72890.0 139010.0 73595.0 140355.0 ;
      RECT  72890.0 141700.0 73595.0 140355.0 ;
      RECT  72890.0 141700.0 73595.0 143045.0 ;
      RECT  72890.0 144390.0 73595.0 143045.0 ;
      RECT  72890.0 144390.0 73595.0 145735.0 ;
      RECT  72890.0 147080.0 73595.0 145735.0 ;
      RECT  72890.0 147080.0 73595.0 148425.0 ;
      RECT  72890.0 149770.0 73595.0 148425.0 ;
      RECT  72890.0 149770.0 73595.0 151115.0 ;
      RECT  72890.0 152460.0 73595.0 151115.0 ;
      RECT  72890.0 152460.0 73595.0 153805.0 ;
      RECT  72890.0 155150.0 73595.0 153805.0 ;
      RECT  72890.0 155150.0 73595.0 156495.0 ;
      RECT  72890.0 157840.0 73595.0 156495.0 ;
      RECT  72890.0 157840.0 73595.0 159185.0 ;
      RECT  72890.0 160530.0 73595.0 159185.0 ;
      RECT  72890.0 160530.0 73595.0 161875.0 ;
      RECT  72890.0 163220.0 73595.0 161875.0 ;
      RECT  72890.0 163220.0 73595.0 164565.0 ;
      RECT  72890.0 165910.0 73595.0 164565.0 ;
      RECT  72890.0 165910.0 73595.0 167255.0 ;
      RECT  72890.0 168600.0 73595.0 167255.0 ;
      RECT  72890.0 168600.0 73595.0 169945.0 ;
      RECT  72890.0 171290.0 73595.0 169945.0 ;
      RECT  72890.0 171290.0 73595.0 172635.0 ;
      RECT  72890.0 173980.0 73595.0 172635.0 ;
      RECT  72890.0 173980.0 73595.0 175325.0 ;
      RECT  72890.0 176670.0 73595.0 175325.0 ;
      RECT  72890.0 176670.0 73595.0 178015.0 ;
      RECT  72890.0 179360.0 73595.0 178015.0 ;
      RECT  72890.0 179360.0 73595.0 180705.0 ;
      RECT  72890.0 182050.0 73595.0 180705.0 ;
      RECT  72890.0 182050.0 73595.0 183395.0 ;
      RECT  72890.0 184740.0 73595.0 183395.0 ;
      RECT  72890.0 184740.0 73595.0 186085.0 ;
      RECT  72890.0 187430.0 73595.0 186085.0 ;
      RECT  72890.0 187430.0 73595.0 188775.0 ;
      RECT  72890.0 190120.0 73595.0 188775.0 ;
      RECT  72890.0 190120.0 73595.0 191465.0 ;
      RECT  72890.0 192810.0 73595.0 191465.0 ;
      RECT  72890.0 192810.0 73595.0 194155.0 ;
      RECT  72890.0 195500.0 73595.0 194155.0 ;
      RECT  72890.0 195500.0 73595.0 196845.0 ;
      RECT  72890.0 198190.0 73595.0 196845.0 ;
      RECT  72890.0 198190.0 73595.0 199535.0 ;
      RECT  72890.0 200880.0 73595.0 199535.0 ;
      RECT  72890.0 200880.0 73595.0 202225.0 ;
      RECT  72890.0 203570.0 73595.0 202225.0 ;
      RECT  72890.0 203570.0 73595.0 204915.0 ;
      RECT  72890.0 206260.0 73595.0 204915.0 ;
      RECT  73595.0 34100.0 74300.0 35445.0 ;
      RECT  73595.0 36790.0 74300.0 35445.0 ;
      RECT  73595.0 36790.0 74300.0 38135.0 ;
      RECT  73595.0 39480.0 74300.0 38135.0 ;
      RECT  73595.0 39480.0 74300.0 40825.0 ;
      RECT  73595.0 42170.0 74300.0 40825.0 ;
      RECT  73595.0 42170.0 74300.0 43515.0 ;
      RECT  73595.0 44860.0 74300.0 43515.0 ;
      RECT  73595.0 44860.0 74300.0 46205.0 ;
      RECT  73595.0 47550.0 74300.0 46205.0 ;
      RECT  73595.0 47550.0 74300.0 48895.0 ;
      RECT  73595.0 50240.0 74300.0 48895.0 ;
      RECT  73595.0 50240.0 74300.0 51585.0 ;
      RECT  73595.0 52930.0 74300.0 51585.0 ;
      RECT  73595.0 52930.0 74300.0 54275.0 ;
      RECT  73595.0 55620.0 74300.0 54275.0 ;
      RECT  73595.0 55620.0 74300.0 56965.0 ;
      RECT  73595.0 58310.0 74300.0 56965.0 ;
      RECT  73595.0 58310.0 74300.0 59655.0 ;
      RECT  73595.0 61000.0 74300.0 59655.0 ;
      RECT  73595.0 61000.0 74300.0 62345.0 ;
      RECT  73595.0 63690.0 74300.0 62345.0 ;
      RECT  73595.0 63690.0 74300.0 65035.0 ;
      RECT  73595.0 66380.0 74300.0 65035.0 ;
      RECT  73595.0 66380.0 74300.0 67725.0 ;
      RECT  73595.0 69070.0 74300.0 67725.0 ;
      RECT  73595.0 69070.0 74300.0 70415.0 ;
      RECT  73595.0 71760.0 74300.0 70415.0 ;
      RECT  73595.0 71760.0 74300.0 73105.0 ;
      RECT  73595.0 74450.0 74300.0 73105.0 ;
      RECT  73595.0 74450.0 74300.0 75795.0 ;
      RECT  73595.0 77140.0 74300.0 75795.0 ;
      RECT  73595.0 77140.0 74300.0 78485.0 ;
      RECT  73595.0 79830.0 74300.0 78485.0 ;
      RECT  73595.0 79830.0 74300.0 81175.0 ;
      RECT  73595.0 82520.0 74300.0 81175.0 ;
      RECT  73595.0 82520.0 74300.0 83865.0 ;
      RECT  73595.0 85210.0 74300.0 83865.0 ;
      RECT  73595.0 85210.0 74300.0 86555.0 ;
      RECT  73595.0 87900.0 74300.0 86555.0 ;
      RECT  73595.0 87900.0 74300.0 89245.0 ;
      RECT  73595.0 90590.0 74300.0 89245.0 ;
      RECT  73595.0 90590.0 74300.0 91935.0 ;
      RECT  73595.0 93280.0 74300.0 91935.0 ;
      RECT  73595.0 93280.0 74300.0 94625.0 ;
      RECT  73595.0 95970.0 74300.0 94625.0 ;
      RECT  73595.0 95970.0 74300.0 97315.0 ;
      RECT  73595.0 98660.0 74300.0 97315.0 ;
      RECT  73595.0 98660.0 74300.0 100005.0 ;
      RECT  73595.0 101350.0 74300.0 100005.0 ;
      RECT  73595.0 101350.0 74300.0 102695.0 ;
      RECT  73595.0 104040.0 74300.0 102695.0 ;
      RECT  73595.0 104040.0 74300.0 105385.0 ;
      RECT  73595.0 106730.0 74300.0 105385.0 ;
      RECT  73595.0 106730.0 74300.0 108075.0 ;
      RECT  73595.0 109420.0 74300.0 108075.0 ;
      RECT  73595.0 109420.0 74300.0 110765.0 ;
      RECT  73595.0 112110.0 74300.0 110765.0 ;
      RECT  73595.0 112110.0 74300.0 113455.0 ;
      RECT  73595.0 114800.0 74300.0 113455.0 ;
      RECT  73595.0 114800.0 74300.0 116145.0 ;
      RECT  73595.0 117490.0 74300.0 116145.0 ;
      RECT  73595.0 117490.0 74300.0 118835.0 ;
      RECT  73595.0 120180.0 74300.0 118835.0 ;
      RECT  73595.0 120180.0 74300.0 121525.0 ;
      RECT  73595.0 122870.0 74300.0 121525.0 ;
      RECT  73595.0 122870.0 74300.0 124215.0 ;
      RECT  73595.0 125560.0 74300.0 124215.0 ;
      RECT  73595.0 125560.0 74300.0 126905.0 ;
      RECT  73595.0 128250.0 74300.0 126905.0 ;
      RECT  73595.0 128250.0 74300.0 129595.0 ;
      RECT  73595.0 130940.0 74300.0 129595.0 ;
      RECT  73595.0 130940.0 74300.0 132285.0 ;
      RECT  73595.0 133630.0 74300.0 132285.0 ;
      RECT  73595.0 133630.0 74300.0 134975.0 ;
      RECT  73595.0 136320.0 74300.0 134975.0 ;
      RECT  73595.0 136320.0 74300.0 137665.0 ;
      RECT  73595.0 139010.0 74300.0 137665.0 ;
      RECT  73595.0 139010.0 74300.0 140355.0 ;
      RECT  73595.0 141700.0 74300.0 140355.0 ;
      RECT  73595.0 141700.0 74300.0 143045.0 ;
      RECT  73595.0 144390.0 74300.0 143045.0 ;
      RECT  73595.0 144390.0 74300.0 145735.0 ;
      RECT  73595.0 147080.0 74300.0 145735.0 ;
      RECT  73595.0 147080.0 74300.0 148425.0 ;
      RECT  73595.0 149770.0 74300.0 148425.0 ;
      RECT  73595.0 149770.0 74300.0 151115.0 ;
      RECT  73595.0 152460.0 74300.0 151115.0 ;
      RECT  73595.0 152460.0 74300.0 153805.0 ;
      RECT  73595.0 155150.0 74300.0 153805.0 ;
      RECT  73595.0 155150.0 74300.0 156495.0 ;
      RECT  73595.0 157840.0 74300.0 156495.0 ;
      RECT  73595.0 157840.0 74300.0 159185.0 ;
      RECT  73595.0 160530.0 74300.0 159185.0 ;
      RECT  73595.0 160530.0 74300.0 161875.0 ;
      RECT  73595.0 163220.0 74300.0 161875.0 ;
      RECT  73595.0 163220.0 74300.0 164565.0 ;
      RECT  73595.0 165910.0 74300.0 164565.0 ;
      RECT  73595.0 165910.0 74300.0 167255.0 ;
      RECT  73595.0 168600.0 74300.0 167255.0 ;
      RECT  73595.0 168600.0 74300.0 169945.0 ;
      RECT  73595.0 171290.0 74300.0 169945.0 ;
      RECT  73595.0 171290.0 74300.0 172635.0 ;
      RECT  73595.0 173980.0 74300.0 172635.0 ;
      RECT  73595.0 173980.0 74300.0 175325.0 ;
      RECT  73595.0 176670.0 74300.0 175325.0 ;
      RECT  73595.0 176670.0 74300.0 178015.0 ;
      RECT  73595.0 179360.0 74300.0 178015.0 ;
      RECT  73595.0 179360.0 74300.0 180705.0 ;
      RECT  73595.0 182050.0 74300.0 180705.0 ;
      RECT  73595.0 182050.0 74300.0 183395.0 ;
      RECT  73595.0 184740.0 74300.0 183395.0 ;
      RECT  73595.0 184740.0 74300.0 186085.0 ;
      RECT  73595.0 187430.0 74300.0 186085.0 ;
      RECT  73595.0 187430.0 74300.0 188775.0 ;
      RECT  73595.0 190120.0 74300.0 188775.0 ;
      RECT  73595.0 190120.0 74300.0 191465.0 ;
      RECT  73595.0 192810.0 74300.0 191465.0 ;
      RECT  73595.0 192810.0 74300.0 194155.0 ;
      RECT  73595.0 195500.0 74300.0 194155.0 ;
      RECT  73595.0 195500.0 74300.0 196845.0 ;
      RECT  73595.0 198190.0 74300.0 196845.0 ;
      RECT  73595.0 198190.0 74300.0 199535.0 ;
      RECT  73595.0 200880.0 74300.0 199535.0 ;
      RECT  73595.0 200880.0 74300.0 202225.0 ;
      RECT  73595.0 203570.0 74300.0 202225.0 ;
      RECT  73595.0 203570.0 74300.0 204915.0 ;
      RECT  73595.0 206260.0 74300.0 204915.0 ;
      RECT  74300.0 34100.0 75005.0 35445.0 ;
      RECT  74300.0 36790.0 75005.0 35445.0 ;
      RECT  74300.0 36790.0 75005.0 38135.0 ;
      RECT  74300.0 39480.0 75005.0 38135.0 ;
      RECT  74300.0 39480.0 75005.0 40825.0 ;
      RECT  74300.0 42170.0 75005.0 40825.0 ;
      RECT  74300.0 42170.0 75005.0 43515.0 ;
      RECT  74300.0 44860.0 75005.0 43515.0 ;
      RECT  74300.0 44860.0 75005.0 46205.0 ;
      RECT  74300.0 47550.0 75005.0 46205.0 ;
      RECT  74300.0 47550.0 75005.0 48895.0 ;
      RECT  74300.0 50240.0 75005.0 48895.0 ;
      RECT  74300.0 50240.0 75005.0 51585.0 ;
      RECT  74300.0 52930.0 75005.0 51585.0 ;
      RECT  74300.0 52930.0 75005.0 54275.0 ;
      RECT  74300.0 55620.0 75005.0 54275.0 ;
      RECT  74300.0 55620.0 75005.0 56965.0 ;
      RECT  74300.0 58310.0 75005.0 56965.0 ;
      RECT  74300.0 58310.0 75005.0 59655.0 ;
      RECT  74300.0 61000.0 75005.0 59655.0 ;
      RECT  74300.0 61000.0 75005.0 62345.0 ;
      RECT  74300.0 63690.0 75005.0 62345.0 ;
      RECT  74300.0 63690.0 75005.0 65035.0 ;
      RECT  74300.0 66380.0 75005.0 65035.0 ;
      RECT  74300.0 66380.0 75005.0 67725.0 ;
      RECT  74300.0 69070.0 75005.0 67725.0 ;
      RECT  74300.0 69070.0 75005.0 70415.0 ;
      RECT  74300.0 71760.0 75005.0 70415.0 ;
      RECT  74300.0 71760.0 75005.0 73105.0 ;
      RECT  74300.0 74450.0 75005.0 73105.0 ;
      RECT  74300.0 74450.0 75005.0 75795.0 ;
      RECT  74300.0 77140.0 75005.0 75795.0 ;
      RECT  74300.0 77140.0 75005.0 78485.0 ;
      RECT  74300.0 79830.0 75005.0 78485.0 ;
      RECT  74300.0 79830.0 75005.0 81175.0 ;
      RECT  74300.0 82520.0 75005.0 81175.0 ;
      RECT  74300.0 82520.0 75005.0 83865.0 ;
      RECT  74300.0 85210.0 75005.0 83865.0 ;
      RECT  74300.0 85210.0 75005.0 86555.0 ;
      RECT  74300.0 87900.0 75005.0 86555.0 ;
      RECT  74300.0 87900.0 75005.0 89245.0 ;
      RECT  74300.0 90590.0 75005.0 89245.0 ;
      RECT  74300.0 90590.0 75005.0 91935.0 ;
      RECT  74300.0 93280.0 75005.0 91935.0 ;
      RECT  74300.0 93280.0 75005.0 94625.0 ;
      RECT  74300.0 95970.0 75005.0 94625.0 ;
      RECT  74300.0 95970.0 75005.0 97315.0 ;
      RECT  74300.0 98660.0 75005.0 97315.0 ;
      RECT  74300.0 98660.0 75005.0 100005.0 ;
      RECT  74300.0 101350.0 75005.0 100005.0 ;
      RECT  74300.0 101350.0 75005.0 102695.0 ;
      RECT  74300.0 104040.0 75005.0 102695.0 ;
      RECT  74300.0 104040.0 75005.0 105385.0 ;
      RECT  74300.0 106730.0 75005.0 105385.0 ;
      RECT  74300.0 106730.0 75005.0 108075.0 ;
      RECT  74300.0 109420.0 75005.0 108075.0 ;
      RECT  74300.0 109420.0 75005.0 110765.0 ;
      RECT  74300.0 112110.0 75005.0 110765.0 ;
      RECT  74300.0 112110.0 75005.0 113455.0 ;
      RECT  74300.0 114800.0 75005.0 113455.0 ;
      RECT  74300.0 114800.0 75005.0 116145.0 ;
      RECT  74300.0 117490.0 75005.0 116145.0 ;
      RECT  74300.0 117490.0 75005.0 118835.0 ;
      RECT  74300.0 120180.0 75005.0 118835.0 ;
      RECT  74300.0 120180.0 75005.0 121525.0 ;
      RECT  74300.0 122870.0 75005.0 121525.0 ;
      RECT  74300.0 122870.0 75005.0 124215.0 ;
      RECT  74300.0 125560.0 75005.0 124215.0 ;
      RECT  74300.0 125560.0 75005.0 126905.0 ;
      RECT  74300.0 128250.0 75005.0 126905.0 ;
      RECT  74300.0 128250.0 75005.0 129595.0 ;
      RECT  74300.0 130940.0 75005.0 129595.0 ;
      RECT  74300.0 130940.0 75005.0 132285.0 ;
      RECT  74300.0 133630.0 75005.0 132285.0 ;
      RECT  74300.0 133630.0 75005.0 134975.0 ;
      RECT  74300.0 136320.0 75005.0 134975.0 ;
      RECT  74300.0 136320.0 75005.0 137665.0 ;
      RECT  74300.0 139010.0 75005.0 137665.0 ;
      RECT  74300.0 139010.0 75005.0 140355.0 ;
      RECT  74300.0 141700.0 75005.0 140355.0 ;
      RECT  74300.0 141700.0 75005.0 143045.0 ;
      RECT  74300.0 144390.0 75005.0 143045.0 ;
      RECT  74300.0 144390.0 75005.0 145735.0 ;
      RECT  74300.0 147080.0 75005.0 145735.0 ;
      RECT  74300.0 147080.0 75005.0 148425.0 ;
      RECT  74300.0 149770.0 75005.0 148425.0 ;
      RECT  74300.0 149770.0 75005.0 151115.0 ;
      RECT  74300.0 152460.0 75005.0 151115.0 ;
      RECT  74300.0 152460.0 75005.0 153805.0 ;
      RECT  74300.0 155150.0 75005.0 153805.0 ;
      RECT  74300.0 155150.0 75005.0 156495.0 ;
      RECT  74300.0 157840.0 75005.0 156495.0 ;
      RECT  74300.0 157840.0 75005.0 159185.0 ;
      RECT  74300.0 160530.0 75005.0 159185.0 ;
      RECT  74300.0 160530.0 75005.0 161875.0 ;
      RECT  74300.0 163220.0 75005.0 161875.0 ;
      RECT  74300.0 163220.0 75005.0 164565.0 ;
      RECT  74300.0 165910.0 75005.0 164565.0 ;
      RECT  74300.0 165910.0 75005.0 167255.0 ;
      RECT  74300.0 168600.0 75005.0 167255.0 ;
      RECT  74300.0 168600.0 75005.0 169945.0 ;
      RECT  74300.0 171290.0 75005.0 169945.0 ;
      RECT  74300.0 171290.0 75005.0 172635.0 ;
      RECT  74300.0 173980.0 75005.0 172635.0 ;
      RECT  74300.0 173980.0 75005.0 175325.0 ;
      RECT  74300.0 176670.0 75005.0 175325.0 ;
      RECT  74300.0 176670.0 75005.0 178015.0 ;
      RECT  74300.0 179360.0 75005.0 178015.0 ;
      RECT  74300.0 179360.0 75005.0 180705.0 ;
      RECT  74300.0 182050.0 75005.0 180705.0 ;
      RECT  74300.0 182050.0 75005.0 183395.0 ;
      RECT  74300.0 184740.0 75005.0 183395.0 ;
      RECT  74300.0 184740.0 75005.0 186085.0 ;
      RECT  74300.0 187430.0 75005.0 186085.0 ;
      RECT  74300.0 187430.0 75005.0 188775.0 ;
      RECT  74300.0 190120.0 75005.0 188775.0 ;
      RECT  74300.0 190120.0 75005.0 191465.0 ;
      RECT  74300.0 192810.0 75005.0 191465.0 ;
      RECT  74300.0 192810.0 75005.0 194155.0 ;
      RECT  74300.0 195500.0 75005.0 194155.0 ;
      RECT  74300.0 195500.0 75005.0 196845.0 ;
      RECT  74300.0 198190.0 75005.0 196845.0 ;
      RECT  74300.0 198190.0 75005.0 199535.0 ;
      RECT  74300.0 200880.0 75005.0 199535.0 ;
      RECT  74300.0 200880.0 75005.0 202225.0 ;
      RECT  74300.0 203570.0 75005.0 202225.0 ;
      RECT  74300.0 203570.0 75005.0 204915.0 ;
      RECT  74300.0 206260.0 75005.0 204915.0 ;
      RECT  75005.0 34100.0 75710.0 35445.0 ;
      RECT  75005.0 36790.0 75710.0 35445.0 ;
      RECT  75005.0 36790.0 75710.0 38135.0 ;
      RECT  75005.0 39480.0 75710.0 38135.0 ;
      RECT  75005.0 39480.0 75710.0 40825.0 ;
      RECT  75005.0 42170.0 75710.0 40825.0 ;
      RECT  75005.0 42170.0 75710.0 43515.0 ;
      RECT  75005.0 44860.0 75710.0 43515.0 ;
      RECT  75005.0 44860.0 75710.0 46205.0 ;
      RECT  75005.0 47550.0 75710.0 46205.0 ;
      RECT  75005.0 47550.0 75710.0 48895.0 ;
      RECT  75005.0 50240.0 75710.0 48895.0 ;
      RECT  75005.0 50240.0 75710.0 51585.0 ;
      RECT  75005.0 52930.0 75710.0 51585.0 ;
      RECT  75005.0 52930.0 75710.0 54275.0 ;
      RECT  75005.0 55620.0 75710.0 54275.0 ;
      RECT  75005.0 55620.0 75710.0 56965.0 ;
      RECT  75005.0 58310.0 75710.0 56965.0 ;
      RECT  75005.0 58310.0 75710.0 59655.0 ;
      RECT  75005.0 61000.0 75710.0 59655.0 ;
      RECT  75005.0 61000.0 75710.0 62345.0 ;
      RECT  75005.0 63690.0 75710.0 62345.0 ;
      RECT  75005.0 63690.0 75710.0 65035.0 ;
      RECT  75005.0 66380.0 75710.0 65035.0 ;
      RECT  75005.0 66380.0 75710.0 67725.0 ;
      RECT  75005.0 69070.0 75710.0 67725.0 ;
      RECT  75005.0 69070.0 75710.0 70415.0 ;
      RECT  75005.0 71760.0 75710.0 70415.0 ;
      RECT  75005.0 71760.0 75710.0 73105.0 ;
      RECT  75005.0 74450.0 75710.0 73105.0 ;
      RECT  75005.0 74450.0 75710.0 75795.0 ;
      RECT  75005.0 77140.0 75710.0 75795.0 ;
      RECT  75005.0 77140.0 75710.0 78485.0 ;
      RECT  75005.0 79830.0 75710.0 78485.0 ;
      RECT  75005.0 79830.0 75710.0 81175.0 ;
      RECT  75005.0 82520.0 75710.0 81175.0 ;
      RECT  75005.0 82520.0 75710.0 83865.0 ;
      RECT  75005.0 85210.0 75710.0 83865.0 ;
      RECT  75005.0 85210.0 75710.0 86555.0 ;
      RECT  75005.0 87900.0 75710.0 86555.0 ;
      RECT  75005.0 87900.0 75710.0 89245.0 ;
      RECT  75005.0 90590.0 75710.0 89245.0 ;
      RECT  75005.0 90590.0 75710.0 91935.0 ;
      RECT  75005.0 93280.0 75710.0 91935.0 ;
      RECT  75005.0 93280.0 75710.0 94625.0 ;
      RECT  75005.0 95970.0 75710.0 94625.0 ;
      RECT  75005.0 95970.0 75710.0 97315.0 ;
      RECT  75005.0 98660.0 75710.0 97315.0 ;
      RECT  75005.0 98660.0 75710.0 100005.0 ;
      RECT  75005.0 101350.0 75710.0 100005.0 ;
      RECT  75005.0 101350.0 75710.0 102695.0 ;
      RECT  75005.0 104040.0 75710.0 102695.0 ;
      RECT  75005.0 104040.0 75710.0 105385.0 ;
      RECT  75005.0 106730.0 75710.0 105385.0 ;
      RECT  75005.0 106730.0 75710.0 108075.0 ;
      RECT  75005.0 109420.0 75710.0 108075.0 ;
      RECT  75005.0 109420.0 75710.0 110765.0 ;
      RECT  75005.0 112110.0 75710.0 110765.0 ;
      RECT  75005.0 112110.0 75710.0 113455.0 ;
      RECT  75005.0 114800.0 75710.0 113455.0 ;
      RECT  75005.0 114800.0 75710.0 116145.0 ;
      RECT  75005.0 117490.0 75710.0 116145.0 ;
      RECT  75005.0 117490.0 75710.0 118835.0 ;
      RECT  75005.0 120180.0 75710.0 118835.0 ;
      RECT  75005.0 120180.0 75710.0 121525.0 ;
      RECT  75005.0 122870.0 75710.0 121525.0 ;
      RECT  75005.0 122870.0 75710.0 124215.0 ;
      RECT  75005.0 125560.0 75710.0 124215.0 ;
      RECT  75005.0 125560.0 75710.0 126905.0 ;
      RECT  75005.0 128250.0 75710.0 126905.0 ;
      RECT  75005.0 128250.0 75710.0 129595.0 ;
      RECT  75005.0 130940.0 75710.0 129595.0 ;
      RECT  75005.0 130940.0 75710.0 132285.0 ;
      RECT  75005.0 133630.0 75710.0 132285.0 ;
      RECT  75005.0 133630.0 75710.0 134975.0 ;
      RECT  75005.0 136320.0 75710.0 134975.0 ;
      RECT  75005.0 136320.0 75710.0 137665.0 ;
      RECT  75005.0 139010.0 75710.0 137665.0 ;
      RECT  75005.0 139010.0 75710.0 140355.0 ;
      RECT  75005.0 141700.0 75710.0 140355.0 ;
      RECT  75005.0 141700.0 75710.0 143045.0 ;
      RECT  75005.0 144390.0 75710.0 143045.0 ;
      RECT  75005.0 144390.0 75710.0 145735.0 ;
      RECT  75005.0 147080.0 75710.0 145735.0 ;
      RECT  75005.0 147080.0 75710.0 148425.0 ;
      RECT  75005.0 149770.0 75710.0 148425.0 ;
      RECT  75005.0 149770.0 75710.0 151115.0 ;
      RECT  75005.0 152460.0 75710.0 151115.0 ;
      RECT  75005.0 152460.0 75710.0 153805.0 ;
      RECT  75005.0 155150.0 75710.0 153805.0 ;
      RECT  75005.0 155150.0 75710.0 156495.0 ;
      RECT  75005.0 157840.0 75710.0 156495.0 ;
      RECT  75005.0 157840.0 75710.0 159185.0 ;
      RECT  75005.0 160530.0 75710.0 159185.0 ;
      RECT  75005.0 160530.0 75710.0 161875.0 ;
      RECT  75005.0 163220.0 75710.0 161875.0 ;
      RECT  75005.0 163220.0 75710.0 164565.0 ;
      RECT  75005.0 165910.0 75710.0 164565.0 ;
      RECT  75005.0 165910.0 75710.0 167255.0 ;
      RECT  75005.0 168600.0 75710.0 167255.0 ;
      RECT  75005.0 168600.0 75710.0 169945.0 ;
      RECT  75005.0 171290.0 75710.0 169945.0 ;
      RECT  75005.0 171290.0 75710.0 172635.0 ;
      RECT  75005.0 173980.0 75710.0 172635.0 ;
      RECT  75005.0 173980.0 75710.0 175325.0 ;
      RECT  75005.0 176670.0 75710.0 175325.0 ;
      RECT  75005.0 176670.0 75710.0 178015.0 ;
      RECT  75005.0 179360.0 75710.0 178015.0 ;
      RECT  75005.0 179360.0 75710.0 180705.0 ;
      RECT  75005.0 182050.0 75710.0 180705.0 ;
      RECT  75005.0 182050.0 75710.0 183395.0 ;
      RECT  75005.0 184740.0 75710.0 183395.0 ;
      RECT  75005.0 184740.0 75710.0 186085.0 ;
      RECT  75005.0 187430.0 75710.0 186085.0 ;
      RECT  75005.0 187430.0 75710.0 188775.0 ;
      RECT  75005.0 190120.0 75710.0 188775.0 ;
      RECT  75005.0 190120.0 75710.0 191465.0 ;
      RECT  75005.0 192810.0 75710.0 191465.0 ;
      RECT  75005.0 192810.0 75710.0 194155.0 ;
      RECT  75005.0 195500.0 75710.0 194155.0 ;
      RECT  75005.0 195500.0 75710.0 196845.0 ;
      RECT  75005.0 198190.0 75710.0 196845.0 ;
      RECT  75005.0 198190.0 75710.0 199535.0 ;
      RECT  75005.0 200880.0 75710.0 199535.0 ;
      RECT  75005.0 200880.0 75710.0 202225.0 ;
      RECT  75005.0 203570.0 75710.0 202225.0 ;
      RECT  75005.0 203570.0 75710.0 204915.0 ;
      RECT  75005.0 206260.0 75710.0 204915.0 ;
      RECT  75710.0 34100.0 76415.0 35445.0 ;
      RECT  75710.0 36790.0 76415.0 35445.0 ;
      RECT  75710.0 36790.0 76415.0 38135.0 ;
      RECT  75710.0 39480.0 76415.0 38135.0 ;
      RECT  75710.0 39480.0 76415.0 40825.0 ;
      RECT  75710.0 42170.0 76415.0 40825.0 ;
      RECT  75710.0 42170.0 76415.0 43515.0 ;
      RECT  75710.0 44860.0 76415.0 43515.0 ;
      RECT  75710.0 44860.0 76415.0 46205.0 ;
      RECT  75710.0 47550.0 76415.0 46205.0 ;
      RECT  75710.0 47550.0 76415.0 48895.0 ;
      RECT  75710.0 50240.0 76415.0 48895.0 ;
      RECT  75710.0 50240.0 76415.0 51585.0 ;
      RECT  75710.0 52930.0 76415.0 51585.0 ;
      RECT  75710.0 52930.0 76415.0 54275.0 ;
      RECT  75710.0 55620.0 76415.0 54275.0 ;
      RECT  75710.0 55620.0 76415.0 56965.0 ;
      RECT  75710.0 58310.0 76415.0 56965.0 ;
      RECT  75710.0 58310.0 76415.0 59655.0 ;
      RECT  75710.0 61000.0 76415.0 59655.0 ;
      RECT  75710.0 61000.0 76415.0 62345.0 ;
      RECT  75710.0 63690.0 76415.0 62345.0 ;
      RECT  75710.0 63690.0 76415.0 65035.0 ;
      RECT  75710.0 66380.0 76415.0 65035.0 ;
      RECT  75710.0 66380.0 76415.0 67725.0 ;
      RECT  75710.0 69070.0 76415.0 67725.0 ;
      RECT  75710.0 69070.0 76415.0 70415.0 ;
      RECT  75710.0 71760.0 76415.0 70415.0 ;
      RECT  75710.0 71760.0 76415.0 73105.0 ;
      RECT  75710.0 74450.0 76415.0 73105.0 ;
      RECT  75710.0 74450.0 76415.0 75795.0 ;
      RECT  75710.0 77140.0 76415.0 75795.0 ;
      RECT  75710.0 77140.0 76415.0 78485.0 ;
      RECT  75710.0 79830.0 76415.0 78485.0 ;
      RECT  75710.0 79830.0 76415.0 81175.0 ;
      RECT  75710.0 82520.0 76415.0 81175.0 ;
      RECT  75710.0 82520.0 76415.0 83865.0 ;
      RECT  75710.0 85210.0 76415.0 83865.0 ;
      RECT  75710.0 85210.0 76415.0 86555.0 ;
      RECT  75710.0 87900.0 76415.0 86555.0 ;
      RECT  75710.0 87900.0 76415.0 89245.0 ;
      RECT  75710.0 90590.0 76415.0 89245.0 ;
      RECT  75710.0 90590.0 76415.0 91935.0 ;
      RECT  75710.0 93280.0 76415.0 91935.0 ;
      RECT  75710.0 93280.0 76415.0 94625.0 ;
      RECT  75710.0 95970.0 76415.0 94625.0 ;
      RECT  75710.0 95970.0 76415.0 97315.0 ;
      RECT  75710.0 98660.0 76415.0 97315.0 ;
      RECT  75710.0 98660.0 76415.0 100005.0 ;
      RECT  75710.0 101350.0 76415.0 100005.0 ;
      RECT  75710.0 101350.0 76415.0 102695.0 ;
      RECT  75710.0 104040.0 76415.0 102695.0 ;
      RECT  75710.0 104040.0 76415.0 105385.0 ;
      RECT  75710.0 106730.0 76415.0 105385.0 ;
      RECT  75710.0 106730.0 76415.0 108075.0 ;
      RECT  75710.0 109420.0 76415.0 108075.0 ;
      RECT  75710.0 109420.0 76415.0 110765.0 ;
      RECT  75710.0 112110.0 76415.0 110765.0 ;
      RECT  75710.0 112110.0 76415.0 113455.0 ;
      RECT  75710.0 114800.0 76415.0 113455.0 ;
      RECT  75710.0 114800.0 76415.0 116145.0 ;
      RECT  75710.0 117490.0 76415.0 116145.0 ;
      RECT  75710.0 117490.0 76415.0 118835.0 ;
      RECT  75710.0 120180.0 76415.0 118835.0 ;
      RECT  75710.0 120180.0 76415.0 121525.0 ;
      RECT  75710.0 122870.0 76415.0 121525.0 ;
      RECT  75710.0 122870.0 76415.0 124215.0 ;
      RECT  75710.0 125560.0 76415.0 124215.0 ;
      RECT  75710.0 125560.0 76415.0 126905.0 ;
      RECT  75710.0 128250.0 76415.0 126905.0 ;
      RECT  75710.0 128250.0 76415.0 129595.0 ;
      RECT  75710.0 130940.0 76415.0 129595.0 ;
      RECT  75710.0 130940.0 76415.0 132285.0 ;
      RECT  75710.0 133630.0 76415.0 132285.0 ;
      RECT  75710.0 133630.0 76415.0 134975.0 ;
      RECT  75710.0 136320.0 76415.0 134975.0 ;
      RECT  75710.0 136320.0 76415.0 137665.0 ;
      RECT  75710.0 139010.0 76415.0 137665.0 ;
      RECT  75710.0 139010.0 76415.0 140355.0 ;
      RECT  75710.0 141700.0 76415.0 140355.0 ;
      RECT  75710.0 141700.0 76415.0 143045.0 ;
      RECT  75710.0 144390.0 76415.0 143045.0 ;
      RECT  75710.0 144390.0 76415.0 145735.0 ;
      RECT  75710.0 147080.0 76415.0 145735.0 ;
      RECT  75710.0 147080.0 76415.0 148425.0 ;
      RECT  75710.0 149770.0 76415.0 148425.0 ;
      RECT  75710.0 149770.0 76415.0 151115.0 ;
      RECT  75710.0 152460.0 76415.0 151115.0 ;
      RECT  75710.0 152460.0 76415.0 153805.0 ;
      RECT  75710.0 155150.0 76415.0 153805.0 ;
      RECT  75710.0 155150.0 76415.0 156495.0 ;
      RECT  75710.0 157840.0 76415.0 156495.0 ;
      RECT  75710.0 157840.0 76415.0 159185.0 ;
      RECT  75710.0 160530.0 76415.0 159185.0 ;
      RECT  75710.0 160530.0 76415.0 161875.0 ;
      RECT  75710.0 163220.0 76415.0 161875.0 ;
      RECT  75710.0 163220.0 76415.0 164565.0 ;
      RECT  75710.0 165910.0 76415.0 164565.0 ;
      RECT  75710.0 165910.0 76415.0 167255.0 ;
      RECT  75710.0 168600.0 76415.0 167255.0 ;
      RECT  75710.0 168600.0 76415.0 169945.0 ;
      RECT  75710.0 171290.0 76415.0 169945.0 ;
      RECT  75710.0 171290.0 76415.0 172635.0 ;
      RECT  75710.0 173980.0 76415.0 172635.0 ;
      RECT  75710.0 173980.0 76415.0 175325.0 ;
      RECT  75710.0 176670.0 76415.0 175325.0 ;
      RECT  75710.0 176670.0 76415.0 178015.0 ;
      RECT  75710.0 179360.0 76415.0 178015.0 ;
      RECT  75710.0 179360.0 76415.0 180705.0 ;
      RECT  75710.0 182050.0 76415.0 180705.0 ;
      RECT  75710.0 182050.0 76415.0 183395.0 ;
      RECT  75710.0 184740.0 76415.0 183395.0 ;
      RECT  75710.0 184740.0 76415.0 186085.0 ;
      RECT  75710.0 187430.0 76415.0 186085.0 ;
      RECT  75710.0 187430.0 76415.0 188775.0 ;
      RECT  75710.0 190120.0 76415.0 188775.0 ;
      RECT  75710.0 190120.0 76415.0 191465.0 ;
      RECT  75710.0 192810.0 76415.0 191465.0 ;
      RECT  75710.0 192810.0 76415.0 194155.0 ;
      RECT  75710.0 195500.0 76415.0 194155.0 ;
      RECT  75710.0 195500.0 76415.0 196845.0 ;
      RECT  75710.0 198190.0 76415.0 196845.0 ;
      RECT  75710.0 198190.0 76415.0 199535.0 ;
      RECT  75710.0 200880.0 76415.0 199535.0 ;
      RECT  75710.0 200880.0 76415.0 202225.0 ;
      RECT  75710.0 203570.0 76415.0 202225.0 ;
      RECT  75710.0 203570.0 76415.0 204915.0 ;
      RECT  75710.0 206260.0 76415.0 204915.0 ;
      RECT  76415.0 34100.0 77120.0 35445.0 ;
      RECT  76415.0 36790.0 77120.0 35445.0 ;
      RECT  76415.0 36790.0 77120.0 38135.0 ;
      RECT  76415.0 39480.0 77120.0 38135.0 ;
      RECT  76415.0 39480.0 77120.0 40825.0 ;
      RECT  76415.0 42170.0 77120.0 40825.0 ;
      RECT  76415.0 42170.0 77120.0 43515.0 ;
      RECT  76415.0 44860.0 77120.0 43515.0 ;
      RECT  76415.0 44860.0 77120.0 46205.0 ;
      RECT  76415.0 47550.0 77120.0 46205.0 ;
      RECT  76415.0 47550.0 77120.0 48895.0 ;
      RECT  76415.0 50240.0 77120.0 48895.0 ;
      RECT  76415.0 50240.0 77120.0 51585.0 ;
      RECT  76415.0 52930.0 77120.0 51585.0 ;
      RECT  76415.0 52930.0 77120.0 54275.0 ;
      RECT  76415.0 55620.0 77120.0 54275.0 ;
      RECT  76415.0 55620.0 77120.0 56965.0 ;
      RECT  76415.0 58310.0 77120.0 56965.0 ;
      RECT  76415.0 58310.0 77120.0 59655.0 ;
      RECT  76415.0 61000.0 77120.0 59655.0 ;
      RECT  76415.0 61000.0 77120.0 62345.0 ;
      RECT  76415.0 63690.0 77120.0 62345.0 ;
      RECT  76415.0 63690.0 77120.0 65035.0 ;
      RECT  76415.0 66380.0 77120.0 65035.0 ;
      RECT  76415.0 66380.0 77120.0 67725.0 ;
      RECT  76415.0 69070.0 77120.0 67725.0 ;
      RECT  76415.0 69070.0 77120.0 70415.0 ;
      RECT  76415.0 71760.0 77120.0 70415.0 ;
      RECT  76415.0 71760.0 77120.0 73105.0 ;
      RECT  76415.0 74450.0 77120.0 73105.0 ;
      RECT  76415.0 74450.0 77120.0 75795.0 ;
      RECT  76415.0 77140.0 77120.0 75795.0 ;
      RECT  76415.0 77140.0 77120.0 78485.0 ;
      RECT  76415.0 79830.0 77120.0 78485.0 ;
      RECT  76415.0 79830.0 77120.0 81175.0 ;
      RECT  76415.0 82520.0 77120.0 81175.0 ;
      RECT  76415.0 82520.0 77120.0 83865.0 ;
      RECT  76415.0 85210.0 77120.0 83865.0 ;
      RECT  76415.0 85210.0 77120.0 86555.0 ;
      RECT  76415.0 87900.0 77120.0 86555.0 ;
      RECT  76415.0 87900.0 77120.0 89245.0 ;
      RECT  76415.0 90590.0 77120.0 89245.0 ;
      RECT  76415.0 90590.0 77120.0 91935.0 ;
      RECT  76415.0 93280.0 77120.0 91935.0 ;
      RECT  76415.0 93280.0 77120.0 94625.0 ;
      RECT  76415.0 95970.0 77120.0 94625.0 ;
      RECT  76415.0 95970.0 77120.0 97315.0 ;
      RECT  76415.0 98660.0 77120.0 97315.0 ;
      RECT  76415.0 98660.0 77120.0 100005.0 ;
      RECT  76415.0 101350.0 77120.0 100005.0 ;
      RECT  76415.0 101350.0 77120.0 102695.0 ;
      RECT  76415.0 104040.0 77120.0 102695.0 ;
      RECT  76415.0 104040.0 77120.0 105385.0 ;
      RECT  76415.0 106730.0 77120.0 105385.0 ;
      RECT  76415.0 106730.0 77120.0 108075.0 ;
      RECT  76415.0 109420.0 77120.0 108075.0 ;
      RECT  76415.0 109420.0 77120.0 110765.0 ;
      RECT  76415.0 112110.0 77120.0 110765.0 ;
      RECT  76415.0 112110.0 77120.0 113455.0 ;
      RECT  76415.0 114800.0 77120.0 113455.0 ;
      RECT  76415.0 114800.0 77120.0 116145.0 ;
      RECT  76415.0 117490.0 77120.0 116145.0 ;
      RECT  76415.0 117490.0 77120.0 118835.0 ;
      RECT  76415.0 120180.0 77120.0 118835.0 ;
      RECT  76415.0 120180.0 77120.0 121525.0 ;
      RECT  76415.0 122870.0 77120.0 121525.0 ;
      RECT  76415.0 122870.0 77120.0 124215.0 ;
      RECT  76415.0 125560.0 77120.0 124215.0 ;
      RECT  76415.0 125560.0 77120.0 126905.0 ;
      RECT  76415.0 128250.0 77120.0 126905.0 ;
      RECT  76415.0 128250.0 77120.0 129595.0 ;
      RECT  76415.0 130940.0 77120.0 129595.0 ;
      RECT  76415.0 130940.0 77120.0 132285.0 ;
      RECT  76415.0 133630.0 77120.0 132285.0 ;
      RECT  76415.0 133630.0 77120.0 134975.0 ;
      RECT  76415.0 136320.0 77120.0 134975.0 ;
      RECT  76415.0 136320.0 77120.0 137665.0 ;
      RECT  76415.0 139010.0 77120.0 137665.0 ;
      RECT  76415.0 139010.0 77120.0 140355.0 ;
      RECT  76415.0 141700.0 77120.0 140355.0 ;
      RECT  76415.0 141700.0 77120.0 143045.0 ;
      RECT  76415.0 144390.0 77120.0 143045.0 ;
      RECT  76415.0 144390.0 77120.0 145735.0 ;
      RECT  76415.0 147080.0 77120.0 145735.0 ;
      RECT  76415.0 147080.0 77120.0 148425.0 ;
      RECT  76415.0 149770.0 77120.0 148425.0 ;
      RECT  76415.0 149770.0 77120.0 151115.0 ;
      RECT  76415.0 152460.0 77120.0 151115.0 ;
      RECT  76415.0 152460.0 77120.0 153805.0 ;
      RECT  76415.0 155150.0 77120.0 153805.0 ;
      RECT  76415.0 155150.0 77120.0 156495.0 ;
      RECT  76415.0 157840.0 77120.0 156495.0 ;
      RECT  76415.0 157840.0 77120.0 159185.0 ;
      RECT  76415.0 160530.0 77120.0 159185.0 ;
      RECT  76415.0 160530.0 77120.0 161875.0 ;
      RECT  76415.0 163220.0 77120.0 161875.0 ;
      RECT  76415.0 163220.0 77120.0 164565.0 ;
      RECT  76415.0 165910.0 77120.0 164565.0 ;
      RECT  76415.0 165910.0 77120.0 167255.0 ;
      RECT  76415.0 168600.0 77120.0 167255.0 ;
      RECT  76415.0 168600.0 77120.0 169945.0 ;
      RECT  76415.0 171290.0 77120.0 169945.0 ;
      RECT  76415.0 171290.0 77120.0 172635.0 ;
      RECT  76415.0 173980.0 77120.0 172635.0 ;
      RECT  76415.0 173980.0 77120.0 175325.0 ;
      RECT  76415.0 176670.0 77120.0 175325.0 ;
      RECT  76415.0 176670.0 77120.0 178015.0 ;
      RECT  76415.0 179360.0 77120.0 178015.0 ;
      RECT  76415.0 179360.0 77120.0 180705.0 ;
      RECT  76415.0 182050.0 77120.0 180705.0 ;
      RECT  76415.0 182050.0 77120.0 183395.0 ;
      RECT  76415.0 184740.0 77120.0 183395.0 ;
      RECT  76415.0 184740.0 77120.0 186085.0 ;
      RECT  76415.0 187430.0 77120.0 186085.0 ;
      RECT  76415.0 187430.0 77120.0 188775.0 ;
      RECT  76415.0 190120.0 77120.0 188775.0 ;
      RECT  76415.0 190120.0 77120.0 191465.0 ;
      RECT  76415.0 192810.0 77120.0 191465.0 ;
      RECT  76415.0 192810.0 77120.0 194155.0 ;
      RECT  76415.0 195500.0 77120.0 194155.0 ;
      RECT  76415.0 195500.0 77120.0 196845.0 ;
      RECT  76415.0 198190.0 77120.0 196845.0 ;
      RECT  76415.0 198190.0 77120.0 199535.0 ;
      RECT  76415.0 200880.0 77120.0 199535.0 ;
      RECT  76415.0 200880.0 77120.0 202225.0 ;
      RECT  76415.0 203570.0 77120.0 202225.0 ;
      RECT  76415.0 203570.0 77120.0 204915.0 ;
      RECT  76415.0 206260.0 77120.0 204915.0 ;
      RECT  77120.0 34100.0 77825.0 35445.0 ;
      RECT  77120.0 36790.0 77825.0 35445.0 ;
      RECT  77120.0 36790.0 77825.0 38135.0 ;
      RECT  77120.0 39480.0 77825.0 38135.0 ;
      RECT  77120.0 39480.0 77825.0 40825.0 ;
      RECT  77120.0 42170.0 77825.0 40825.0 ;
      RECT  77120.0 42170.0 77825.0 43515.0 ;
      RECT  77120.0 44860.0 77825.0 43515.0 ;
      RECT  77120.0 44860.0 77825.0 46205.0 ;
      RECT  77120.0 47550.0 77825.0 46205.0 ;
      RECT  77120.0 47550.0 77825.0 48895.0 ;
      RECT  77120.0 50240.0 77825.0 48895.0 ;
      RECT  77120.0 50240.0 77825.0 51585.0 ;
      RECT  77120.0 52930.0 77825.0 51585.0 ;
      RECT  77120.0 52930.0 77825.0 54275.0 ;
      RECT  77120.0 55620.0 77825.0 54275.0 ;
      RECT  77120.0 55620.0 77825.0 56965.0 ;
      RECT  77120.0 58310.0 77825.0 56965.0 ;
      RECT  77120.0 58310.0 77825.0 59655.0 ;
      RECT  77120.0 61000.0 77825.0 59655.0 ;
      RECT  77120.0 61000.0 77825.0 62345.0 ;
      RECT  77120.0 63690.0 77825.0 62345.0 ;
      RECT  77120.0 63690.0 77825.0 65035.0 ;
      RECT  77120.0 66380.0 77825.0 65035.0 ;
      RECT  77120.0 66380.0 77825.0 67725.0 ;
      RECT  77120.0 69070.0 77825.0 67725.0 ;
      RECT  77120.0 69070.0 77825.0 70415.0 ;
      RECT  77120.0 71760.0 77825.0 70415.0 ;
      RECT  77120.0 71760.0 77825.0 73105.0 ;
      RECT  77120.0 74450.0 77825.0 73105.0 ;
      RECT  77120.0 74450.0 77825.0 75795.0 ;
      RECT  77120.0 77140.0 77825.0 75795.0 ;
      RECT  77120.0 77140.0 77825.0 78485.0 ;
      RECT  77120.0 79830.0 77825.0 78485.0 ;
      RECT  77120.0 79830.0 77825.0 81175.0 ;
      RECT  77120.0 82520.0 77825.0 81175.0 ;
      RECT  77120.0 82520.0 77825.0 83865.0 ;
      RECT  77120.0 85210.0 77825.0 83865.0 ;
      RECT  77120.0 85210.0 77825.0 86555.0 ;
      RECT  77120.0 87900.0 77825.0 86555.0 ;
      RECT  77120.0 87900.0 77825.0 89245.0 ;
      RECT  77120.0 90590.0 77825.0 89245.0 ;
      RECT  77120.0 90590.0 77825.0 91935.0 ;
      RECT  77120.0 93280.0 77825.0 91935.0 ;
      RECT  77120.0 93280.0 77825.0 94625.0 ;
      RECT  77120.0 95970.0 77825.0 94625.0 ;
      RECT  77120.0 95970.0 77825.0 97315.0 ;
      RECT  77120.0 98660.0 77825.0 97315.0 ;
      RECT  77120.0 98660.0 77825.0 100005.0 ;
      RECT  77120.0 101350.0 77825.0 100005.0 ;
      RECT  77120.0 101350.0 77825.0 102695.0 ;
      RECT  77120.0 104040.0 77825.0 102695.0 ;
      RECT  77120.0 104040.0 77825.0 105385.0 ;
      RECT  77120.0 106730.0 77825.0 105385.0 ;
      RECT  77120.0 106730.0 77825.0 108075.0 ;
      RECT  77120.0 109420.0 77825.0 108075.0 ;
      RECT  77120.0 109420.0 77825.0 110765.0 ;
      RECT  77120.0 112110.0 77825.0 110765.0 ;
      RECT  77120.0 112110.0 77825.0 113455.0 ;
      RECT  77120.0 114800.0 77825.0 113455.0 ;
      RECT  77120.0 114800.0 77825.0 116145.0 ;
      RECT  77120.0 117490.0 77825.0 116145.0 ;
      RECT  77120.0 117490.0 77825.0 118835.0 ;
      RECT  77120.0 120180.0 77825.0 118835.0 ;
      RECT  77120.0 120180.0 77825.0 121525.0 ;
      RECT  77120.0 122870.0 77825.0 121525.0 ;
      RECT  77120.0 122870.0 77825.0 124215.0 ;
      RECT  77120.0 125560.0 77825.0 124215.0 ;
      RECT  77120.0 125560.0 77825.0 126905.0 ;
      RECT  77120.0 128250.0 77825.0 126905.0 ;
      RECT  77120.0 128250.0 77825.0 129595.0 ;
      RECT  77120.0 130940.0 77825.0 129595.0 ;
      RECT  77120.0 130940.0 77825.0 132285.0 ;
      RECT  77120.0 133630.0 77825.0 132285.0 ;
      RECT  77120.0 133630.0 77825.0 134975.0 ;
      RECT  77120.0 136320.0 77825.0 134975.0 ;
      RECT  77120.0 136320.0 77825.0 137665.0 ;
      RECT  77120.0 139010.0 77825.0 137665.0 ;
      RECT  77120.0 139010.0 77825.0 140355.0 ;
      RECT  77120.0 141700.0 77825.0 140355.0 ;
      RECT  77120.0 141700.0 77825.0 143045.0 ;
      RECT  77120.0 144390.0 77825.0 143045.0 ;
      RECT  77120.0 144390.0 77825.0 145735.0 ;
      RECT  77120.0 147080.0 77825.0 145735.0 ;
      RECT  77120.0 147080.0 77825.0 148425.0 ;
      RECT  77120.0 149770.0 77825.0 148425.0 ;
      RECT  77120.0 149770.0 77825.0 151115.0 ;
      RECT  77120.0 152460.0 77825.0 151115.0 ;
      RECT  77120.0 152460.0 77825.0 153805.0 ;
      RECT  77120.0 155150.0 77825.0 153805.0 ;
      RECT  77120.0 155150.0 77825.0 156495.0 ;
      RECT  77120.0 157840.0 77825.0 156495.0 ;
      RECT  77120.0 157840.0 77825.0 159185.0 ;
      RECT  77120.0 160530.0 77825.0 159185.0 ;
      RECT  77120.0 160530.0 77825.0 161875.0 ;
      RECT  77120.0 163220.0 77825.0 161875.0 ;
      RECT  77120.0 163220.0 77825.0 164565.0 ;
      RECT  77120.0 165910.0 77825.0 164565.0 ;
      RECT  77120.0 165910.0 77825.0 167255.0 ;
      RECT  77120.0 168600.0 77825.0 167255.0 ;
      RECT  77120.0 168600.0 77825.0 169945.0 ;
      RECT  77120.0 171290.0 77825.0 169945.0 ;
      RECT  77120.0 171290.0 77825.0 172635.0 ;
      RECT  77120.0 173980.0 77825.0 172635.0 ;
      RECT  77120.0 173980.0 77825.0 175325.0 ;
      RECT  77120.0 176670.0 77825.0 175325.0 ;
      RECT  77120.0 176670.0 77825.0 178015.0 ;
      RECT  77120.0 179360.0 77825.0 178015.0 ;
      RECT  77120.0 179360.0 77825.0 180705.0 ;
      RECT  77120.0 182050.0 77825.0 180705.0 ;
      RECT  77120.0 182050.0 77825.0 183395.0 ;
      RECT  77120.0 184740.0 77825.0 183395.0 ;
      RECT  77120.0 184740.0 77825.0 186085.0 ;
      RECT  77120.0 187430.0 77825.0 186085.0 ;
      RECT  77120.0 187430.0 77825.0 188775.0 ;
      RECT  77120.0 190120.0 77825.0 188775.0 ;
      RECT  77120.0 190120.0 77825.0 191465.0 ;
      RECT  77120.0 192810.0 77825.0 191465.0 ;
      RECT  77120.0 192810.0 77825.0 194155.0 ;
      RECT  77120.0 195500.0 77825.0 194155.0 ;
      RECT  77120.0 195500.0 77825.0 196845.0 ;
      RECT  77120.0 198190.0 77825.0 196845.0 ;
      RECT  77120.0 198190.0 77825.0 199535.0 ;
      RECT  77120.0 200880.0 77825.0 199535.0 ;
      RECT  77120.0 200880.0 77825.0 202225.0 ;
      RECT  77120.0 203570.0 77825.0 202225.0 ;
      RECT  77120.0 203570.0 77825.0 204915.0 ;
      RECT  77120.0 206260.0 77825.0 204915.0 ;
      RECT  77825.0 34100.0 78530.0 35445.0 ;
      RECT  77825.0 36790.0 78530.0 35445.0 ;
      RECT  77825.0 36790.0 78530.0 38135.0 ;
      RECT  77825.0 39480.0 78530.0 38135.0 ;
      RECT  77825.0 39480.0 78530.0 40825.0 ;
      RECT  77825.0 42170.0 78530.0 40825.0 ;
      RECT  77825.0 42170.0 78530.0 43515.0 ;
      RECT  77825.0 44860.0 78530.0 43515.0 ;
      RECT  77825.0 44860.0 78530.0 46205.0 ;
      RECT  77825.0 47550.0 78530.0 46205.0 ;
      RECT  77825.0 47550.0 78530.0 48895.0 ;
      RECT  77825.0 50240.0 78530.0 48895.0 ;
      RECT  77825.0 50240.0 78530.0 51585.0 ;
      RECT  77825.0 52930.0 78530.0 51585.0 ;
      RECT  77825.0 52930.0 78530.0 54275.0 ;
      RECT  77825.0 55620.0 78530.0 54275.0 ;
      RECT  77825.0 55620.0 78530.0 56965.0 ;
      RECT  77825.0 58310.0 78530.0 56965.0 ;
      RECT  77825.0 58310.0 78530.0 59655.0 ;
      RECT  77825.0 61000.0 78530.0 59655.0 ;
      RECT  77825.0 61000.0 78530.0 62345.0 ;
      RECT  77825.0 63690.0 78530.0 62345.0 ;
      RECT  77825.0 63690.0 78530.0 65035.0 ;
      RECT  77825.0 66380.0 78530.0 65035.0 ;
      RECT  77825.0 66380.0 78530.0 67725.0 ;
      RECT  77825.0 69070.0 78530.0 67725.0 ;
      RECT  77825.0 69070.0 78530.0 70415.0 ;
      RECT  77825.0 71760.0 78530.0 70415.0 ;
      RECT  77825.0 71760.0 78530.0 73105.0 ;
      RECT  77825.0 74450.0 78530.0 73105.0 ;
      RECT  77825.0 74450.0 78530.0 75795.0 ;
      RECT  77825.0 77140.0 78530.0 75795.0 ;
      RECT  77825.0 77140.0 78530.0 78485.0 ;
      RECT  77825.0 79830.0 78530.0 78485.0 ;
      RECT  77825.0 79830.0 78530.0 81175.0 ;
      RECT  77825.0 82520.0 78530.0 81175.0 ;
      RECT  77825.0 82520.0 78530.0 83865.0 ;
      RECT  77825.0 85210.0 78530.0 83865.0 ;
      RECT  77825.0 85210.0 78530.0 86555.0 ;
      RECT  77825.0 87900.0 78530.0 86555.0 ;
      RECT  77825.0 87900.0 78530.0 89245.0 ;
      RECT  77825.0 90590.0 78530.0 89245.0 ;
      RECT  77825.0 90590.0 78530.0 91935.0 ;
      RECT  77825.0 93280.0 78530.0 91935.0 ;
      RECT  77825.0 93280.0 78530.0 94625.0 ;
      RECT  77825.0 95970.0 78530.0 94625.0 ;
      RECT  77825.0 95970.0 78530.0 97315.0 ;
      RECT  77825.0 98660.0 78530.0 97315.0 ;
      RECT  77825.0 98660.0 78530.0 100005.0 ;
      RECT  77825.0 101350.0 78530.0 100005.0 ;
      RECT  77825.0 101350.0 78530.0 102695.0 ;
      RECT  77825.0 104040.0 78530.0 102695.0 ;
      RECT  77825.0 104040.0 78530.0 105385.0 ;
      RECT  77825.0 106730.0 78530.0 105385.0 ;
      RECT  77825.0 106730.0 78530.0 108075.0 ;
      RECT  77825.0 109420.0 78530.0 108075.0 ;
      RECT  77825.0 109420.0 78530.0 110765.0 ;
      RECT  77825.0 112110.0 78530.0 110765.0 ;
      RECT  77825.0 112110.0 78530.0 113455.0 ;
      RECT  77825.0 114800.0 78530.0 113455.0 ;
      RECT  77825.0 114800.0 78530.0 116145.0 ;
      RECT  77825.0 117490.0 78530.0 116145.0 ;
      RECT  77825.0 117490.0 78530.0 118835.0 ;
      RECT  77825.0 120180.0 78530.0 118835.0 ;
      RECT  77825.0 120180.0 78530.0 121525.0 ;
      RECT  77825.0 122870.0 78530.0 121525.0 ;
      RECT  77825.0 122870.0 78530.0 124215.0 ;
      RECT  77825.0 125560.0 78530.0 124215.0 ;
      RECT  77825.0 125560.0 78530.0 126905.0 ;
      RECT  77825.0 128250.0 78530.0 126905.0 ;
      RECT  77825.0 128250.0 78530.0 129595.0 ;
      RECT  77825.0 130940.0 78530.0 129595.0 ;
      RECT  77825.0 130940.0 78530.0 132285.0 ;
      RECT  77825.0 133630.0 78530.0 132285.0 ;
      RECT  77825.0 133630.0 78530.0 134975.0 ;
      RECT  77825.0 136320.0 78530.0 134975.0 ;
      RECT  77825.0 136320.0 78530.0 137665.0 ;
      RECT  77825.0 139010.0 78530.0 137665.0 ;
      RECT  77825.0 139010.0 78530.0 140355.0 ;
      RECT  77825.0 141700.0 78530.0 140355.0 ;
      RECT  77825.0 141700.0 78530.0 143045.0 ;
      RECT  77825.0 144390.0 78530.0 143045.0 ;
      RECT  77825.0 144390.0 78530.0 145735.0 ;
      RECT  77825.0 147080.0 78530.0 145735.0 ;
      RECT  77825.0 147080.0 78530.0 148425.0 ;
      RECT  77825.0 149770.0 78530.0 148425.0 ;
      RECT  77825.0 149770.0 78530.0 151115.0 ;
      RECT  77825.0 152460.0 78530.0 151115.0 ;
      RECT  77825.0 152460.0 78530.0 153805.0 ;
      RECT  77825.0 155150.0 78530.0 153805.0 ;
      RECT  77825.0 155150.0 78530.0 156495.0 ;
      RECT  77825.0 157840.0 78530.0 156495.0 ;
      RECT  77825.0 157840.0 78530.0 159185.0 ;
      RECT  77825.0 160530.0 78530.0 159185.0 ;
      RECT  77825.0 160530.0 78530.0 161875.0 ;
      RECT  77825.0 163220.0 78530.0 161875.0 ;
      RECT  77825.0 163220.0 78530.0 164565.0 ;
      RECT  77825.0 165910.0 78530.0 164565.0 ;
      RECT  77825.0 165910.0 78530.0 167255.0 ;
      RECT  77825.0 168600.0 78530.0 167255.0 ;
      RECT  77825.0 168600.0 78530.0 169945.0 ;
      RECT  77825.0 171290.0 78530.0 169945.0 ;
      RECT  77825.0 171290.0 78530.0 172635.0 ;
      RECT  77825.0 173980.0 78530.0 172635.0 ;
      RECT  77825.0 173980.0 78530.0 175325.0 ;
      RECT  77825.0 176670.0 78530.0 175325.0 ;
      RECT  77825.0 176670.0 78530.0 178015.0 ;
      RECT  77825.0 179360.0 78530.0 178015.0 ;
      RECT  77825.0 179360.0 78530.0 180705.0 ;
      RECT  77825.0 182050.0 78530.0 180705.0 ;
      RECT  77825.0 182050.0 78530.0 183395.0 ;
      RECT  77825.0 184740.0 78530.0 183395.0 ;
      RECT  77825.0 184740.0 78530.0 186085.0 ;
      RECT  77825.0 187430.0 78530.0 186085.0 ;
      RECT  77825.0 187430.0 78530.0 188775.0 ;
      RECT  77825.0 190120.0 78530.0 188775.0 ;
      RECT  77825.0 190120.0 78530.0 191465.0 ;
      RECT  77825.0 192810.0 78530.0 191465.0 ;
      RECT  77825.0 192810.0 78530.0 194155.0 ;
      RECT  77825.0 195500.0 78530.0 194155.0 ;
      RECT  77825.0 195500.0 78530.0 196845.0 ;
      RECT  77825.0 198190.0 78530.0 196845.0 ;
      RECT  77825.0 198190.0 78530.0 199535.0 ;
      RECT  77825.0 200880.0 78530.0 199535.0 ;
      RECT  77825.0 200880.0 78530.0 202225.0 ;
      RECT  77825.0 203570.0 78530.0 202225.0 ;
      RECT  77825.0 203570.0 78530.0 204915.0 ;
      RECT  77825.0 206260.0 78530.0 204915.0 ;
      RECT  78530.0 34100.0 79235.0 35445.0 ;
      RECT  78530.0 36790.0 79235.0 35445.0 ;
      RECT  78530.0 36790.0 79235.0 38135.0 ;
      RECT  78530.0 39480.0 79235.0 38135.0 ;
      RECT  78530.0 39480.0 79235.0 40825.0 ;
      RECT  78530.0 42170.0 79235.0 40825.0 ;
      RECT  78530.0 42170.0 79235.0 43515.0 ;
      RECT  78530.0 44860.0 79235.0 43515.0 ;
      RECT  78530.0 44860.0 79235.0 46205.0 ;
      RECT  78530.0 47550.0 79235.0 46205.0 ;
      RECT  78530.0 47550.0 79235.0 48895.0 ;
      RECT  78530.0 50240.0 79235.0 48895.0 ;
      RECT  78530.0 50240.0 79235.0 51585.0 ;
      RECT  78530.0 52930.0 79235.0 51585.0 ;
      RECT  78530.0 52930.0 79235.0 54275.0 ;
      RECT  78530.0 55620.0 79235.0 54275.0 ;
      RECT  78530.0 55620.0 79235.0 56965.0 ;
      RECT  78530.0 58310.0 79235.0 56965.0 ;
      RECT  78530.0 58310.0 79235.0 59655.0 ;
      RECT  78530.0 61000.0 79235.0 59655.0 ;
      RECT  78530.0 61000.0 79235.0 62345.0 ;
      RECT  78530.0 63690.0 79235.0 62345.0 ;
      RECT  78530.0 63690.0 79235.0 65035.0 ;
      RECT  78530.0 66380.0 79235.0 65035.0 ;
      RECT  78530.0 66380.0 79235.0 67725.0 ;
      RECT  78530.0 69070.0 79235.0 67725.0 ;
      RECT  78530.0 69070.0 79235.0 70415.0 ;
      RECT  78530.0 71760.0 79235.0 70415.0 ;
      RECT  78530.0 71760.0 79235.0 73105.0 ;
      RECT  78530.0 74450.0 79235.0 73105.0 ;
      RECT  78530.0 74450.0 79235.0 75795.0 ;
      RECT  78530.0 77140.0 79235.0 75795.0 ;
      RECT  78530.0 77140.0 79235.0 78485.0 ;
      RECT  78530.0 79830.0 79235.0 78485.0 ;
      RECT  78530.0 79830.0 79235.0 81175.0 ;
      RECT  78530.0 82520.0 79235.0 81175.0 ;
      RECT  78530.0 82520.0 79235.0 83865.0 ;
      RECT  78530.0 85210.0 79235.0 83865.0 ;
      RECT  78530.0 85210.0 79235.0 86555.0 ;
      RECT  78530.0 87900.0 79235.0 86555.0 ;
      RECT  78530.0 87900.0 79235.0 89245.0 ;
      RECT  78530.0 90590.0 79235.0 89245.0 ;
      RECT  78530.0 90590.0 79235.0 91935.0 ;
      RECT  78530.0 93280.0 79235.0 91935.0 ;
      RECT  78530.0 93280.0 79235.0 94625.0 ;
      RECT  78530.0 95970.0 79235.0 94625.0 ;
      RECT  78530.0 95970.0 79235.0 97315.0 ;
      RECT  78530.0 98660.0 79235.0 97315.0 ;
      RECT  78530.0 98660.0 79235.0 100005.0 ;
      RECT  78530.0 101350.0 79235.0 100005.0 ;
      RECT  78530.0 101350.0 79235.0 102695.0 ;
      RECT  78530.0 104040.0 79235.0 102695.0 ;
      RECT  78530.0 104040.0 79235.0 105385.0 ;
      RECT  78530.0 106730.0 79235.0 105385.0 ;
      RECT  78530.0 106730.0 79235.0 108075.0 ;
      RECT  78530.0 109420.0 79235.0 108075.0 ;
      RECT  78530.0 109420.0 79235.0 110765.0 ;
      RECT  78530.0 112110.0 79235.0 110765.0 ;
      RECT  78530.0 112110.0 79235.0 113455.0 ;
      RECT  78530.0 114800.0 79235.0 113455.0 ;
      RECT  78530.0 114800.0 79235.0 116145.0 ;
      RECT  78530.0 117490.0 79235.0 116145.0 ;
      RECT  78530.0 117490.0 79235.0 118835.0 ;
      RECT  78530.0 120180.0 79235.0 118835.0 ;
      RECT  78530.0 120180.0 79235.0 121525.0 ;
      RECT  78530.0 122870.0 79235.0 121525.0 ;
      RECT  78530.0 122870.0 79235.0 124215.0 ;
      RECT  78530.0 125560.0 79235.0 124215.0 ;
      RECT  78530.0 125560.0 79235.0 126905.0 ;
      RECT  78530.0 128250.0 79235.0 126905.0 ;
      RECT  78530.0 128250.0 79235.0 129595.0 ;
      RECT  78530.0 130940.0 79235.0 129595.0 ;
      RECT  78530.0 130940.0 79235.0 132285.0 ;
      RECT  78530.0 133630.0 79235.0 132285.0 ;
      RECT  78530.0 133630.0 79235.0 134975.0 ;
      RECT  78530.0 136320.0 79235.0 134975.0 ;
      RECT  78530.0 136320.0 79235.0 137665.0 ;
      RECT  78530.0 139010.0 79235.0 137665.0 ;
      RECT  78530.0 139010.0 79235.0 140355.0 ;
      RECT  78530.0 141700.0 79235.0 140355.0 ;
      RECT  78530.0 141700.0 79235.0 143045.0 ;
      RECT  78530.0 144390.0 79235.0 143045.0 ;
      RECT  78530.0 144390.0 79235.0 145735.0 ;
      RECT  78530.0 147080.0 79235.0 145735.0 ;
      RECT  78530.0 147080.0 79235.0 148425.0 ;
      RECT  78530.0 149770.0 79235.0 148425.0 ;
      RECT  78530.0 149770.0 79235.0 151115.0 ;
      RECT  78530.0 152460.0 79235.0 151115.0 ;
      RECT  78530.0 152460.0 79235.0 153805.0 ;
      RECT  78530.0 155150.0 79235.0 153805.0 ;
      RECT  78530.0 155150.0 79235.0 156495.0 ;
      RECT  78530.0 157840.0 79235.0 156495.0 ;
      RECT  78530.0 157840.0 79235.0 159185.0 ;
      RECT  78530.0 160530.0 79235.0 159185.0 ;
      RECT  78530.0 160530.0 79235.0 161875.0 ;
      RECT  78530.0 163220.0 79235.0 161875.0 ;
      RECT  78530.0 163220.0 79235.0 164565.0 ;
      RECT  78530.0 165910.0 79235.0 164565.0 ;
      RECT  78530.0 165910.0 79235.0 167255.0 ;
      RECT  78530.0 168600.0 79235.0 167255.0 ;
      RECT  78530.0 168600.0 79235.0 169945.0 ;
      RECT  78530.0 171290.0 79235.0 169945.0 ;
      RECT  78530.0 171290.0 79235.0 172635.0 ;
      RECT  78530.0 173980.0 79235.0 172635.0 ;
      RECT  78530.0 173980.0 79235.0 175325.0 ;
      RECT  78530.0 176670.0 79235.0 175325.0 ;
      RECT  78530.0 176670.0 79235.0 178015.0 ;
      RECT  78530.0 179360.0 79235.0 178015.0 ;
      RECT  78530.0 179360.0 79235.0 180705.0 ;
      RECT  78530.0 182050.0 79235.0 180705.0 ;
      RECT  78530.0 182050.0 79235.0 183395.0 ;
      RECT  78530.0 184740.0 79235.0 183395.0 ;
      RECT  78530.0 184740.0 79235.0 186085.0 ;
      RECT  78530.0 187430.0 79235.0 186085.0 ;
      RECT  78530.0 187430.0 79235.0 188775.0 ;
      RECT  78530.0 190120.0 79235.0 188775.0 ;
      RECT  78530.0 190120.0 79235.0 191465.0 ;
      RECT  78530.0 192810.0 79235.0 191465.0 ;
      RECT  78530.0 192810.0 79235.0 194155.0 ;
      RECT  78530.0 195500.0 79235.0 194155.0 ;
      RECT  78530.0 195500.0 79235.0 196845.0 ;
      RECT  78530.0 198190.0 79235.0 196845.0 ;
      RECT  78530.0 198190.0 79235.0 199535.0 ;
      RECT  78530.0 200880.0 79235.0 199535.0 ;
      RECT  78530.0 200880.0 79235.0 202225.0 ;
      RECT  78530.0 203570.0 79235.0 202225.0 ;
      RECT  78530.0 203570.0 79235.0 204915.0 ;
      RECT  78530.0 206260.0 79235.0 204915.0 ;
      RECT  79235.0 34100.0 79940.0 35445.0 ;
      RECT  79235.0 36790.0 79940.0 35445.0 ;
      RECT  79235.0 36790.0 79940.0 38135.0 ;
      RECT  79235.0 39480.0 79940.0 38135.0 ;
      RECT  79235.0 39480.0 79940.0 40825.0 ;
      RECT  79235.0 42170.0 79940.0 40825.0 ;
      RECT  79235.0 42170.0 79940.0 43515.0 ;
      RECT  79235.0 44860.0 79940.0 43515.0 ;
      RECT  79235.0 44860.0 79940.0 46205.0 ;
      RECT  79235.0 47550.0 79940.0 46205.0 ;
      RECT  79235.0 47550.0 79940.0 48895.0 ;
      RECT  79235.0 50240.0 79940.0 48895.0 ;
      RECT  79235.0 50240.0 79940.0 51585.0 ;
      RECT  79235.0 52930.0 79940.0 51585.0 ;
      RECT  79235.0 52930.0 79940.0 54275.0 ;
      RECT  79235.0 55620.0 79940.0 54275.0 ;
      RECT  79235.0 55620.0 79940.0 56965.0 ;
      RECT  79235.0 58310.0 79940.0 56965.0 ;
      RECT  79235.0 58310.0 79940.0 59655.0 ;
      RECT  79235.0 61000.0 79940.0 59655.0 ;
      RECT  79235.0 61000.0 79940.0 62345.0 ;
      RECT  79235.0 63690.0 79940.0 62345.0 ;
      RECT  79235.0 63690.0 79940.0 65035.0 ;
      RECT  79235.0 66380.0 79940.0 65035.0 ;
      RECT  79235.0 66380.0 79940.0 67725.0 ;
      RECT  79235.0 69070.0 79940.0 67725.0 ;
      RECT  79235.0 69070.0 79940.0 70415.0 ;
      RECT  79235.0 71760.0 79940.0 70415.0 ;
      RECT  79235.0 71760.0 79940.0 73105.0 ;
      RECT  79235.0 74450.0 79940.0 73105.0 ;
      RECT  79235.0 74450.0 79940.0 75795.0 ;
      RECT  79235.0 77140.0 79940.0 75795.0 ;
      RECT  79235.0 77140.0 79940.0 78485.0 ;
      RECT  79235.0 79830.0 79940.0 78485.0 ;
      RECT  79235.0 79830.0 79940.0 81175.0 ;
      RECT  79235.0 82520.0 79940.0 81175.0 ;
      RECT  79235.0 82520.0 79940.0 83865.0 ;
      RECT  79235.0 85210.0 79940.0 83865.0 ;
      RECT  79235.0 85210.0 79940.0 86555.0 ;
      RECT  79235.0 87900.0 79940.0 86555.0 ;
      RECT  79235.0 87900.0 79940.0 89245.0 ;
      RECT  79235.0 90590.0 79940.0 89245.0 ;
      RECT  79235.0 90590.0 79940.0 91935.0 ;
      RECT  79235.0 93280.0 79940.0 91935.0 ;
      RECT  79235.0 93280.0 79940.0 94625.0 ;
      RECT  79235.0 95970.0 79940.0 94625.0 ;
      RECT  79235.0 95970.0 79940.0 97315.0 ;
      RECT  79235.0 98660.0 79940.0 97315.0 ;
      RECT  79235.0 98660.0 79940.0 100005.0 ;
      RECT  79235.0 101350.0 79940.0 100005.0 ;
      RECT  79235.0 101350.0 79940.0 102695.0 ;
      RECT  79235.0 104040.0 79940.0 102695.0 ;
      RECT  79235.0 104040.0 79940.0 105385.0 ;
      RECT  79235.0 106730.0 79940.0 105385.0 ;
      RECT  79235.0 106730.0 79940.0 108075.0 ;
      RECT  79235.0 109420.0 79940.0 108075.0 ;
      RECT  79235.0 109420.0 79940.0 110765.0 ;
      RECT  79235.0 112110.0 79940.0 110765.0 ;
      RECT  79235.0 112110.0 79940.0 113455.0 ;
      RECT  79235.0 114800.0 79940.0 113455.0 ;
      RECT  79235.0 114800.0 79940.0 116145.0 ;
      RECT  79235.0 117490.0 79940.0 116145.0 ;
      RECT  79235.0 117490.0 79940.0 118835.0 ;
      RECT  79235.0 120180.0 79940.0 118835.0 ;
      RECT  79235.0 120180.0 79940.0 121525.0 ;
      RECT  79235.0 122870.0 79940.0 121525.0 ;
      RECT  79235.0 122870.0 79940.0 124215.0 ;
      RECT  79235.0 125560.0 79940.0 124215.0 ;
      RECT  79235.0 125560.0 79940.0 126905.0 ;
      RECT  79235.0 128250.0 79940.0 126905.0 ;
      RECT  79235.0 128250.0 79940.0 129595.0 ;
      RECT  79235.0 130940.0 79940.0 129595.0 ;
      RECT  79235.0 130940.0 79940.0 132285.0 ;
      RECT  79235.0 133630.0 79940.0 132285.0 ;
      RECT  79235.0 133630.0 79940.0 134975.0 ;
      RECT  79235.0 136320.0 79940.0 134975.0 ;
      RECT  79235.0 136320.0 79940.0 137665.0 ;
      RECT  79235.0 139010.0 79940.0 137665.0 ;
      RECT  79235.0 139010.0 79940.0 140355.0 ;
      RECT  79235.0 141700.0 79940.0 140355.0 ;
      RECT  79235.0 141700.0 79940.0 143045.0 ;
      RECT  79235.0 144390.0 79940.0 143045.0 ;
      RECT  79235.0 144390.0 79940.0 145735.0 ;
      RECT  79235.0 147080.0 79940.0 145735.0 ;
      RECT  79235.0 147080.0 79940.0 148425.0 ;
      RECT  79235.0 149770.0 79940.0 148425.0 ;
      RECT  79235.0 149770.0 79940.0 151115.0 ;
      RECT  79235.0 152460.0 79940.0 151115.0 ;
      RECT  79235.0 152460.0 79940.0 153805.0 ;
      RECT  79235.0 155150.0 79940.0 153805.0 ;
      RECT  79235.0 155150.0 79940.0 156495.0 ;
      RECT  79235.0 157840.0 79940.0 156495.0 ;
      RECT  79235.0 157840.0 79940.0 159185.0 ;
      RECT  79235.0 160530.0 79940.0 159185.0 ;
      RECT  79235.0 160530.0 79940.0 161875.0 ;
      RECT  79235.0 163220.0 79940.0 161875.0 ;
      RECT  79235.0 163220.0 79940.0 164565.0 ;
      RECT  79235.0 165910.0 79940.0 164565.0 ;
      RECT  79235.0 165910.0 79940.0 167255.0 ;
      RECT  79235.0 168600.0 79940.0 167255.0 ;
      RECT  79235.0 168600.0 79940.0 169945.0 ;
      RECT  79235.0 171290.0 79940.0 169945.0 ;
      RECT  79235.0 171290.0 79940.0 172635.0 ;
      RECT  79235.0 173980.0 79940.0 172635.0 ;
      RECT  79235.0 173980.0 79940.0 175325.0 ;
      RECT  79235.0 176670.0 79940.0 175325.0 ;
      RECT  79235.0 176670.0 79940.0 178015.0 ;
      RECT  79235.0 179360.0 79940.0 178015.0 ;
      RECT  79235.0 179360.0 79940.0 180705.0 ;
      RECT  79235.0 182050.0 79940.0 180705.0 ;
      RECT  79235.0 182050.0 79940.0 183395.0 ;
      RECT  79235.0 184740.0 79940.0 183395.0 ;
      RECT  79235.0 184740.0 79940.0 186085.0 ;
      RECT  79235.0 187430.0 79940.0 186085.0 ;
      RECT  79235.0 187430.0 79940.0 188775.0 ;
      RECT  79235.0 190120.0 79940.0 188775.0 ;
      RECT  79235.0 190120.0 79940.0 191465.0 ;
      RECT  79235.0 192810.0 79940.0 191465.0 ;
      RECT  79235.0 192810.0 79940.0 194155.0 ;
      RECT  79235.0 195500.0 79940.0 194155.0 ;
      RECT  79235.0 195500.0 79940.0 196845.0 ;
      RECT  79235.0 198190.0 79940.0 196845.0 ;
      RECT  79235.0 198190.0 79940.0 199535.0 ;
      RECT  79235.0 200880.0 79940.0 199535.0 ;
      RECT  79235.0 200880.0 79940.0 202225.0 ;
      RECT  79235.0 203570.0 79940.0 202225.0 ;
      RECT  79235.0 203570.0 79940.0 204915.0 ;
      RECT  79235.0 206260.0 79940.0 204915.0 ;
      RECT  79940.0 34100.0 80645.0 35445.0 ;
      RECT  79940.0 36790.0 80645.0 35445.0 ;
      RECT  79940.0 36790.0 80645.0 38135.0 ;
      RECT  79940.0 39480.0 80645.0 38135.0 ;
      RECT  79940.0 39480.0 80645.0 40825.0 ;
      RECT  79940.0 42170.0 80645.0 40825.0 ;
      RECT  79940.0 42170.0 80645.0 43515.0 ;
      RECT  79940.0 44860.0 80645.0 43515.0 ;
      RECT  79940.0 44860.0 80645.0 46205.0 ;
      RECT  79940.0 47550.0 80645.0 46205.0 ;
      RECT  79940.0 47550.0 80645.0 48895.0 ;
      RECT  79940.0 50240.0 80645.0 48895.0 ;
      RECT  79940.0 50240.0 80645.0 51585.0 ;
      RECT  79940.0 52930.0 80645.0 51585.0 ;
      RECT  79940.0 52930.0 80645.0 54275.0 ;
      RECT  79940.0 55620.0 80645.0 54275.0 ;
      RECT  79940.0 55620.0 80645.0 56965.0 ;
      RECT  79940.0 58310.0 80645.0 56965.0 ;
      RECT  79940.0 58310.0 80645.0 59655.0 ;
      RECT  79940.0 61000.0 80645.0 59655.0 ;
      RECT  79940.0 61000.0 80645.0 62345.0 ;
      RECT  79940.0 63690.0 80645.0 62345.0 ;
      RECT  79940.0 63690.0 80645.0 65035.0 ;
      RECT  79940.0 66380.0 80645.0 65035.0 ;
      RECT  79940.0 66380.0 80645.0 67725.0 ;
      RECT  79940.0 69070.0 80645.0 67725.0 ;
      RECT  79940.0 69070.0 80645.0 70415.0 ;
      RECT  79940.0 71760.0 80645.0 70415.0 ;
      RECT  79940.0 71760.0 80645.0 73105.0 ;
      RECT  79940.0 74450.0 80645.0 73105.0 ;
      RECT  79940.0 74450.0 80645.0 75795.0 ;
      RECT  79940.0 77140.0 80645.0 75795.0 ;
      RECT  79940.0 77140.0 80645.0 78485.0 ;
      RECT  79940.0 79830.0 80645.0 78485.0 ;
      RECT  79940.0 79830.0 80645.0 81175.0 ;
      RECT  79940.0 82520.0 80645.0 81175.0 ;
      RECT  79940.0 82520.0 80645.0 83865.0 ;
      RECT  79940.0 85210.0 80645.0 83865.0 ;
      RECT  79940.0 85210.0 80645.0 86555.0 ;
      RECT  79940.0 87900.0 80645.0 86555.0 ;
      RECT  79940.0 87900.0 80645.0 89245.0 ;
      RECT  79940.0 90590.0 80645.0 89245.0 ;
      RECT  79940.0 90590.0 80645.0 91935.0 ;
      RECT  79940.0 93280.0 80645.0 91935.0 ;
      RECT  79940.0 93280.0 80645.0 94625.0 ;
      RECT  79940.0 95970.0 80645.0 94625.0 ;
      RECT  79940.0 95970.0 80645.0 97315.0 ;
      RECT  79940.0 98660.0 80645.0 97315.0 ;
      RECT  79940.0 98660.0 80645.0 100005.0 ;
      RECT  79940.0 101350.0 80645.0 100005.0 ;
      RECT  79940.0 101350.0 80645.0 102695.0 ;
      RECT  79940.0 104040.0 80645.0 102695.0 ;
      RECT  79940.0 104040.0 80645.0 105385.0 ;
      RECT  79940.0 106730.0 80645.0 105385.0 ;
      RECT  79940.0 106730.0 80645.0 108075.0 ;
      RECT  79940.0 109420.0 80645.0 108075.0 ;
      RECT  79940.0 109420.0 80645.0 110765.0 ;
      RECT  79940.0 112110.0 80645.0 110765.0 ;
      RECT  79940.0 112110.0 80645.0 113455.0 ;
      RECT  79940.0 114800.0 80645.0 113455.0 ;
      RECT  79940.0 114800.0 80645.0 116145.0 ;
      RECT  79940.0 117490.0 80645.0 116145.0 ;
      RECT  79940.0 117490.0 80645.0 118835.0 ;
      RECT  79940.0 120180.0 80645.0 118835.0 ;
      RECT  79940.0 120180.0 80645.0 121525.0 ;
      RECT  79940.0 122870.0 80645.0 121525.0 ;
      RECT  79940.0 122870.0 80645.0 124215.0 ;
      RECT  79940.0 125560.0 80645.0 124215.0 ;
      RECT  79940.0 125560.0 80645.0 126905.0 ;
      RECT  79940.0 128250.0 80645.0 126905.0 ;
      RECT  79940.0 128250.0 80645.0 129595.0 ;
      RECT  79940.0 130940.0 80645.0 129595.0 ;
      RECT  79940.0 130940.0 80645.0 132285.0 ;
      RECT  79940.0 133630.0 80645.0 132285.0 ;
      RECT  79940.0 133630.0 80645.0 134975.0 ;
      RECT  79940.0 136320.0 80645.0 134975.0 ;
      RECT  79940.0 136320.0 80645.0 137665.0 ;
      RECT  79940.0 139010.0 80645.0 137665.0 ;
      RECT  79940.0 139010.0 80645.0 140355.0 ;
      RECT  79940.0 141700.0 80645.0 140355.0 ;
      RECT  79940.0 141700.0 80645.0 143045.0 ;
      RECT  79940.0 144390.0 80645.0 143045.0 ;
      RECT  79940.0 144390.0 80645.0 145735.0 ;
      RECT  79940.0 147080.0 80645.0 145735.0 ;
      RECT  79940.0 147080.0 80645.0 148425.0 ;
      RECT  79940.0 149770.0 80645.0 148425.0 ;
      RECT  79940.0 149770.0 80645.0 151115.0 ;
      RECT  79940.0 152460.0 80645.0 151115.0 ;
      RECT  79940.0 152460.0 80645.0 153805.0 ;
      RECT  79940.0 155150.0 80645.0 153805.0 ;
      RECT  79940.0 155150.0 80645.0 156495.0 ;
      RECT  79940.0 157840.0 80645.0 156495.0 ;
      RECT  79940.0 157840.0 80645.0 159185.0 ;
      RECT  79940.0 160530.0 80645.0 159185.0 ;
      RECT  79940.0 160530.0 80645.0 161875.0 ;
      RECT  79940.0 163220.0 80645.0 161875.0 ;
      RECT  79940.0 163220.0 80645.0 164565.0 ;
      RECT  79940.0 165910.0 80645.0 164565.0 ;
      RECT  79940.0 165910.0 80645.0 167255.0 ;
      RECT  79940.0 168600.0 80645.0 167255.0 ;
      RECT  79940.0 168600.0 80645.0 169945.0 ;
      RECT  79940.0 171290.0 80645.0 169945.0 ;
      RECT  79940.0 171290.0 80645.0 172635.0 ;
      RECT  79940.0 173980.0 80645.0 172635.0 ;
      RECT  79940.0 173980.0 80645.0 175325.0 ;
      RECT  79940.0 176670.0 80645.0 175325.0 ;
      RECT  79940.0 176670.0 80645.0 178015.0 ;
      RECT  79940.0 179360.0 80645.0 178015.0 ;
      RECT  79940.0 179360.0 80645.0 180705.0 ;
      RECT  79940.0 182050.0 80645.0 180705.0 ;
      RECT  79940.0 182050.0 80645.0 183395.0 ;
      RECT  79940.0 184740.0 80645.0 183395.0 ;
      RECT  79940.0 184740.0 80645.0 186085.0 ;
      RECT  79940.0 187430.0 80645.0 186085.0 ;
      RECT  79940.0 187430.0 80645.0 188775.0 ;
      RECT  79940.0 190120.0 80645.0 188775.0 ;
      RECT  79940.0 190120.0 80645.0 191465.0 ;
      RECT  79940.0 192810.0 80645.0 191465.0 ;
      RECT  79940.0 192810.0 80645.0 194155.0 ;
      RECT  79940.0 195500.0 80645.0 194155.0 ;
      RECT  79940.0 195500.0 80645.0 196845.0 ;
      RECT  79940.0 198190.0 80645.0 196845.0 ;
      RECT  79940.0 198190.0 80645.0 199535.0 ;
      RECT  79940.0 200880.0 80645.0 199535.0 ;
      RECT  79940.0 200880.0 80645.0 202225.0 ;
      RECT  79940.0 203570.0 80645.0 202225.0 ;
      RECT  79940.0 203570.0 80645.0 204915.0 ;
      RECT  79940.0 206260.0 80645.0 204915.0 ;
      RECT  80645.0 34100.0 81350.0 35445.0 ;
      RECT  80645.0 36790.0 81350.0 35445.0 ;
      RECT  80645.0 36790.0 81350.0 38135.0 ;
      RECT  80645.0 39480.0 81350.0 38135.0 ;
      RECT  80645.0 39480.0 81350.0 40825.0 ;
      RECT  80645.0 42170.0 81350.0 40825.0 ;
      RECT  80645.0 42170.0 81350.0 43515.0 ;
      RECT  80645.0 44860.0 81350.0 43515.0 ;
      RECT  80645.0 44860.0 81350.0 46205.0 ;
      RECT  80645.0 47550.0 81350.0 46205.0 ;
      RECT  80645.0 47550.0 81350.0 48895.0 ;
      RECT  80645.0 50240.0 81350.0 48895.0 ;
      RECT  80645.0 50240.0 81350.0 51585.0 ;
      RECT  80645.0 52930.0 81350.0 51585.0 ;
      RECT  80645.0 52930.0 81350.0 54275.0 ;
      RECT  80645.0 55620.0 81350.0 54275.0 ;
      RECT  80645.0 55620.0 81350.0 56965.0 ;
      RECT  80645.0 58310.0 81350.0 56965.0 ;
      RECT  80645.0 58310.0 81350.0 59655.0 ;
      RECT  80645.0 61000.0 81350.0 59655.0 ;
      RECT  80645.0 61000.0 81350.0 62345.0 ;
      RECT  80645.0 63690.0 81350.0 62345.0 ;
      RECT  80645.0 63690.0 81350.0 65035.0 ;
      RECT  80645.0 66380.0 81350.0 65035.0 ;
      RECT  80645.0 66380.0 81350.0 67725.0 ;
      RECT  80645.0 69070.0 81350.0 67725.0 ;
      RECT  80645.0 69070.0 81350.0 70415.0 ;
      RECT  80645.0 71760.0 81350.0 70415.0 ;
      RECT  80645.0 71760.0 81350.0 73105.0 ;
      RECT  80645.0 74450.0 81350.0 73105.0 ;
      RECT  80645.0 74450.0 81350.0 75795.0 ;
      RECT  80645.0 77140.0 81350.0 75795.0 ;
      RECT  80645.0 77140.0 81350.0 78485.0 ;
      RECT  80645.0 79830.0 81350.0 78485.0 ;
      RECT  80645.0 79830.0 81350.0 81175.0 ;
      RECT  80645.0 82520.0 81350.0 81175.0 ;
      RECT  80645.0 82520.0 81350.0 83865.0 ;
      RECT  80645.0 85210.0 81350.0 83865.0 ;
      RECT  80645.0 85210.0 81350.0 86555.0 ;
      RECT  80645.0 87900.0 81350.0 86555.0 ;
      RECT  80645.0 87900.0 81350.0 89245.0 ;
      RECT  80645.0 90590.0 81350.0 89245.0 ;
      RECT  80645.0 90590.0 81350.0 91935.0 ;
      RECT  80645.0 93280.0 81350.0 91935.0 ;
      RECT  80645.0 93280.0 81350.0 94625.0 ;
      RECT  80645.0 95970.0 81350.0 94625.0 ;
      RECT  80645.0 95970.0 81350.0 97315.0 ;
      RECT  80645.0 98660.0 81350.0 97315.0 ;
      RECT  80645.0 98660.0 81350.0 100005.0 ;
      RECT  80645.0 101350.0 81350.0 100005.0 ;
      RECT  80645.0 101350.0 81350.0 102695.0 ;
      RECT  80645.0 104040.0 81350.0 102695.0 ;
      RECT  80645.0 104040.0 81350.0 105385.0 ;
      RECT  80645.0 106730.0 81350.0 105385.0 ;
      RECT  80645.0 106730.0 81350.0 108075.0 ;
      RECT  80645.0 109420.0 81350.0 108075.0 ;
      RECT  80645.0 109420.0 81350.0 110765.0 ;
      RECT  80645.0 112110.0 81350.0 110765.0 ;
      RECT  80645.0 112110.0 81350.0 113455.0 ;
      RECT  80645.0 114800.0 81350.0 113455.0 ;
      RECT  80645.0 114800.0 81350.0 116145.0 ;
      RECT  80645.0 117490.0 81350.0 116145.0 ;
      RECT  80645.0 117490.0 81350.0 118835.0 ;
      RECT  80645.0 120180.0 81350.0 118835.0 ;
      RECT  80645.0 120180.0 81350.0 121525.0 ;
      RECT  80645.0 122870.0 81350.0 121525.0 ;
      RECT  80645.0 122870.0 81350.0 124215.0 ;
      RECT  80645.0 125560.0 81350.0 124215.0 ;
      RECT  80645.0 125560.0 81350.0 126905.0 ;
      RECT  80645.0 128250.0 81350.0 126905.0 ;
      RECT  80645.0 128250.0 81350.0 129595.0 ;
      RECT  80645.0 130940.0 81350.0 129595.0 ;
      RECT  80645.0 130940.0 81350.0 132285.0 ;
      RECT  80645.0 133630.0 81350.0 132285.0 ;
      RECT  80645.0 133630.0 81350.0 134975.0 ;
      RECT  80645.0 136320.0 81350.0 134975.0 ;
      RECT  80645.0 136320.0 81350.0 137665.0 ;
      RECT  80645.0 139010.0 81350.0 137665.0 ;
      RECT  80645.0 139010.0 81350.0 140355.0 ;
      RECT  80645.0 141700.0 81350.0 140355.0 ;
      RECT  80645.0 141700.0 81350.0 143045.0 ;
      RECT  80645.0 144390.0 81350.0 143045.0 ;
      RECT  80645.0 144390.0 81350.0 145735.0 ;
      RECT  80645.0 147080.0 81350.0 145735.0 ;
      RECT  80645.0 147080.0 81350.0 148425.0 ;
      RECT  80645.0 149770.0 81350.0 148425.0 ;
      RECT  80645.0 149770.0 81350.0 151115.0 ;
      RECT  80645.0 152460.0 81350.0 151115.0 ;
      RECT  80645.0 152460.0 81350.0 153805.0 ;
      RECT  80645.0 155150.0 81350.0 153805.0 ;
      RECT  80645.0 155150.0 81350.0 156495.0 ;
      RECT  80645.0 157840.0 81350.0 156495.0 ;
      RECT  80645.0 157840.0 81350.0 159185.0 ;
      RECT  80645.0 160530.0 81350.0 159185.0 ;
      RECT  80645.0 160530.0 81350.0 161875.0 ;
      RECT  80645.0 163220.0 81350.0 161875.0 ;
      RECT  80645.0 163220.0 81350.0 164565.0 ;
      RECT  80645.0 165910.0 81350.0 164565.0 ;
      RECT  80645.0 165910.0 81350.0 167255.0 ;
      RECT  80645.0 168600.0 81350.0 167255.0 ;
      RECT  80645.0 168600.0 81350.0 169945.0 ;
      RECT  80645.0 171290.0 81350.0 169945.0 ;
      RECT  80645.0 171290.0 81350.0 172635.0 ;
      RECT  80645.0 173980.0 81350.0 172635.0 ;
      RECT  80645.0 173980.0 81350.0 175325.0 ;
      RECT  80645.0 176670.0 81350.0 175325.0 ;
      RECT  80645.0 176670.0 81350.0 178015.0 ;
      RECT  80645.0 179360.0 81350.0 178015.0 ;
      RECT  80645.0 179360.0 81350.0 180705.0 ;
      RECT  80645.0 182050.0 81350.0 180705.0 ;
      RECT  80645.0 182050.0 81350.0 183395.0 ;
      RECT  80645.0 184740.0 81350.0 183395.0 ;
      RECT  80645.0 184740.0 81350.0 186085.0 ;
      RECT  80645.0 187430.0 81350.0 186085.0 ;
      RECT  80645.0 187430.0 81350.0 188775.0 ;
      RECT  80645.0 190120.0 81350.0 188775.0 ;
      RECT  80645.0 190120.0 81350.0 191465.0 ;
      RECT  80645.0 192810.0 81350.0 191465.0 ;
      RECT  80645.0 192810.0 81350.0 194155.0 ;
      RECT  80645.0 195500.0 81350.0 194155.0 ;
      RECT  80645.0 195500.0 81350.0 196845.0 ;
      RECT  80645.0 198190.0 81350.0 196845.0 ;
      RECT  80645.0 198190.0 81350.0 199535.0 ;
      RECT  80645.0 200880.0 81350.0 199535.0 ;
      RECT  80645.0 200880.0 81350.0 202225.0 ;
      RECT  80645.0 203570.0 81350.0 202225.0 ;
      RECT  80645.0 203570.0 81350.0 204915.0 ;
      RECT  80645.0 206260.0 81350.0 204915.0 ;
      RECT  81350.0 34100.0 82055.0 35445.0 ;
      RECT  81350.0 36790.0 82055.0 35445.0 ;
      RECT  81350.0 36790.0 82055.0 38135.0 ;
      RECT  81350.0 39480.0 82055.0 38135.0 ;
      RECT  81350.0 39480.0 82055.0 40825.0 ;
      RECT  81350.0 42170.0 82055.0 40825.0 ;
      RECT  81350.0 42170.0 82055.0 43515.0 ;
      RECT  81350.0 44860.0 82055.0 43515.0 ;
      RECT  81350.0 44860.0 82055.0 46205.0 ;
      RECT  81350.0 47550.0 82055.0 46205.0 ;
      RECT  81350.0 47550.0 82055.0 48895.0 ;
      RECT  81350.0 50240.0 82055.0 48895.0 ;
      RECT  81350.0 50240.0 82055.0 51585.0 ;
      RECT  81350.0 52930.0 82055.0 51585.0 ;
      RECT  81350.0 52930.0 82055.0 54275.0 ;
      RECT  81350.0 55620.0 82055.0 54275.0 ;
      RECT  81350.0 55620.0 82055.0 56965.0 ;
      RECT  81350.0 58310.0 82055.0 56965.0 ;
      RECT  81350.0 58310.0 82055.0 59655.0 ;
      RECT  81350.0 61000.0 82055.0 59655.0 ;
      RECT  81350.0 61000.0 82055.0 62345.0 ;
      RECT  81350.0 63690.0 82055.0 62345.0 ;
      RECT  81350.0 63690.0 82055.0 65035.0 ;
      RECT  81350.0 66380.0 82055.0 65035.0 ;
      RECT  81350.0 66380.0 82055.0 67725.0 ;
      RECT  81350.0 69070.0 82055.0 67725.0 ;
      RECT  81350.0 69070.0 82055.0 70415.0 ;
      RECT  81350.0 71760.0 82055.0 70415.0 ;
      RECT  81350.0 71760.0 82055.0 73105.0 ;
      RECT  81350.0 74450.0 82055.0 73105.0 ;
      RECT  81350.0 74450.0 82055.0 75795.0 ;
      RECT  81350.0 77140.0 82055.0 75795.0 ;
      RECT  81350.0 77140.0 82055.0 78485.0 ;
      RECT  81350.0 79830.0 82055.0 78485.0 ;
      RECT  81350.0 79830.0 82055.0 81175.0 ;
      RECT  81350.0 82520.0 82055.0 81175.0 ;
      RECT  81350.0 82520.0 82055.0 83865.0 ;
      RECT  81350.0 85210.0 82055.0 83865.0 ;
      RECT  81350.0 85210.0 82055.0 86555.0 ;
      RECT  81350.0 87900.0 82055.0 86555.0 ;
      RECT  81350.0 87900.0 82055.0 89245.0 ;
      RECT  81350.0 90590.0 82055.0 89245.0 ;
      RECT  81350.0 90590.0 82055.0 91935.0 ;
      RECT  81350.0 93280.0 82055.0 91935.0 ;
      RECT  81350.0 93280.0 82055.0 94625.0 ;
      RECT  81350.0 95970.0 82055.0 94625.0 ;
      RECT  81350.0 95970.0 82055.0 97315.0 ;
      RECT  81350.0 98660.0 82055.0 97315.0 ;
      RECT  81350.0 98660.0 82055.0 100005.0 ;
      RECT  81350.0 101350.0 82055.0 100005.0 ;
      RECT  81350.0 101350.0 82055.0 102695.0 ;
      RECT  81350.0 104040.0 82055.0 102695.0 ;
      RECT  81350.0 104040.0 82055.0 105385.0 ;
      RECT  81350.0 106730.0 82055.0 105385.0 ;
      RECT  81350.0 106730.0 82055.0 108075.0 ;
      RECT  81350.0 109420.0 82055.0 108075.0 ;
      RECT  81350.0 109420.0 82055.0 110765.0 ;
      RECT  81350.0 112110.0 82055.0 110765.0 ;
      RECT  81350.0 112110.0 82055.0 113455.0 ;
      RECT  81350.0 114800.0 82055.0 113455.0 ;
      RECT  81350.0 114800.0 82055.0 116145.0 ;
      RECT  81350.0 117490.0 82055.0 116145.0 ;
      RECT  81350.0 117490.0 82055.0 118835.0 ;
      RECT  81350.0 120180.0 82055.0 118835.0 ;
      RECT  81350.0 120180.0 82055.0 121525.0 ;
      RECT  81350.0 122870.0 82055.0 121525.0 ;
      RECT  81350.0 122870.0 82055.0 124215.0 ;
      RECT  81350.0 125560.0 82055.0 124215.0 ;
      RECT  81350.0 125560.0 82055.0 126905.0 ;
      RECT  81350.0 128250.0 82055.0 126905.0 ;
      RECT  81350.0 128250.0 82055.0 129595.0 ;
      RECT  81350.0 130940.0 82055.0 129595.0 ;
      RECT  81350.0 130940.0 82055.0 132285.0 ;
      RECT  81350.0 133630.0 82055.0 132285.0 ;
      RECT  81350.0 133630.0 82055.0 134975.0 ;
      RECT  81350.0 136320.0 82055.0 134975.0 ;
      RECT  81350.0 136320.0 82055.0 137665.0 ;
      RECT  81350.0 139010.0 82055.0 137665.0 ;
      RECT  81350.0 139010.0 82055.0 140355.0 ;
      RECT  81350.0 141700.0 82055.0 140355.0 ;
      RECT  81350.0 141700.0 82055.0 143045.0 ;
      RECT  81350.0 144390.0 82055.0 143045.0 ;
      RECT  81350.0 144390.0 82055.0 145735.0 ;
      RECT  81350.0 147080.0 82055.0 145735.0 ;
      RECT  81350.0 147080.0 82055.0 148425.0 ;
      RECT  81350.0 149770.0 82055.0 148425.0 ;
      RECT  81350.0 149770.0 82055.0 151115.0 ;
      RECT  81350.0 152460.0 82055.0 151115.0 ;
      RECT  81350.0 152460.0 82055.0 153805.0 ;
      RECT  81350.0 155150.0 82055.0 153805.0 ;
      RECT  81350.0 155150.0 82055.0 156495.0 ;
      RECT  81350.0 157840.0 82055.0 156495.0 ;
      RECT  81350.0 157840.0 82055.0 159185.0 ;
      RECT  81350.0 160530.0 82055.0 159185.0 ;
      RECT  81350.0 160530.0 82055.0 161875.0 ;
      RECT  81350.0 163220.0 82055.0 161875.0 ;
      RECT  81350.0 163220.0 82055.0 164565.0 ;
      RECT  81350.0 165910.0 82055.0 164565.0 ;
      RECT  81350.0 165910.0 82055.0 167255.0 ;
      RECT  81350.0 168600.0 82055.0 167255.0 ;
      RECT  81350.0 168600.0 82055.0 169945.0 ;
      RECT  81350.0 171290.0 82055.0 169945.0 ;
      RECT  81350.0 171290.0 82055.0 172635.0 ;
      RECT  81350.0 173980.0 82055.0 172635.0 ;
      RECT  81350.0 173980.0 82055.0 175325.0 ;
      RECT  81350.0 176670.0 82055.0 175325.0 ;
      RECT  81350.0 176670.0 82055.0 178015.0 ;
      RECT  81350.0 179360.0 82055.0 178015.0 ;
      RECT  81350.0 179360.0 82055.0 180705.0 ;
      RECT  81350.0 182050.0 82055.0 180705.0 ;
      RECT  81350.0 182050.0 82055.0 183395.0 ;
      RECT  81350.0 184740.0 82055.0 183395.0 ;
      RECT  81350.0 184740.0 82055.0 186085.0 ;
      RECT  81350.0 187430.0 82055.0 186085.0 ;
      RECT  81350.0 187430.0 82055.0 188775.0 ;
      RECT  81350.0 190120.0 82055.0 188775.0 ;
      RECT  81350.0 190120.0 82055.0 191465.0 ;
      RECT  81350.0 192810.0 82055.0 191465.0 ;
      RECT  81350.0 192810.0 82055.0 194155.0 ;
      RECT  81350.0 195500.0 82055.0 194155.0 ;
      RECT  81350.0 195500.0 82055.0 196845.0 ;
      RECT  81350.0 198190.0 82055.0 196845.0 ;
      RECT  81350.0 198190.0 82055.0 199535.0 ;
      RECT  81350.0 200880.0 82055.0 199535.0 ;
      RECT  81350.0 200880.0 82055.0 202225.0 ;
      RECT  81350.0 203570.0 82055.0 202225.0 ;
      RECT  81350.0 203570.0 82055.0 204915.0 ;
      RECT  81350.0 206260.0 82055.0 204915.0 ;
      RECT  82055.0 34100.0 82760.0 35445.0 ;
      RECT  82055.0 36790.0 82760.0 35445.0 ;
      RECT  82055.0 36790.0 82760.0 38135.0 ;
      RECT  82055.0 39480.0 82760.0 38135.0 ;
      RECT  82055.0 39480.0 82760.0 40825.0 ;
      RECT  82055.0 42170.0 82760.0 40825.0 ;
      RECT  82055.0 42170.0 82760.0 43515.0 ;
      RECT  82055.0 44860.0 82760.0 43515.0 ;
      RECT  82055.0 44860.0 82760.0 46205.0 ;
      RECT  82055.0 47550.0 82760.0 46205.0 ;
      RECT  82055.0 47550.0 82760.0 48895.0 ;
      RECT  82055.0 50240.0 82760.0 48895.0 ;
      RECT  82055.0 50240.0 82760.0 51585.0 ;
      RECT  82055.0 52930.0 82760.0 51585.0 ;
      RECT  82055.0 52930.0 82760.0 54275.0 ;
      RECT  82055.0 55620.0 82760.0 54275.0 ;
      RECT  82055.0 55620.0 82760.0 56965.0 ;
      RECT  82055.0 58310.0 82760.0 56965.0 ;
      RECT  82055.0 58310.0 82760.0 59655.0 ;
      RECT  82055.0 61000.0 82760.0 59655.0 ;
      RECT  82055.0 61000.0 82760.0 62345.0 ;
      RECT  82055.0 63690.0 82760.0 62345.0 ;
      RECT  82055.0 63690.0 82760.0 65035.0 ;
      RECT  82055.0 66380.0 82760.0 65035.0 ;
      RECT  82055.0 66380.0 82760.0 67725.0 ;
      RECT  82055.0 69070.0 82760.0 67725.0 ;
      RECT  82055.0 69070.0 82760.0 70415.0 ;
      RECT  82055.0 71760.0 82760.0 70415.0 ;
      RECT  82055.0 71760.0 82760.0 73105.0 ;
      RECT  82055.0 74450.0 82760.0 73105.0 ;
      RECT  82055.0 74450.0 82760.0 75795.0 ;
      RECT  82055.0 77140.0 82760.0 75795.0 ;
      RECT  82055.0 77140.0 82760.0 78485.0 ;
      RECT  82055.0 79830.0 82760.0 78485.0 ;
      RECT  82055.0 79830.0 82760.0 81175.0 ;
      RECT  82055.0 82520.0 82760.0 81175.0 ;
      RECT  82055.0 82520.0 82760.0 83865.0 ;
      RECT  82055.0 85210.0 82760.0 83865.0 ;
      RECT  82055.0 85210.0 82760.0 86555.0 ;
      RECT  82055.0 87900.0 82760.0 86555.0 ;
      RECT  82055.0 87900.0 82760.0 89245.0 ;
      RECT  82055.0 90590.0 82760.0 89245.0 ;
      RECT  82055.0 90590.0 82760.0 91935.0 ;
      RECT  82055.0 93280.0 82760.0 91935.0 ;
      RECT  82055.0 93280.0 82760.0 94625.0 ;
      RECT  82055.0 95970.0 82760.0 94625.0 ;
      RECT  82055.0 95970.0 82760.0 97315.0 ;
      RECT  82055.0 98660.0 82760.0 97315.0 ;
      RECT  82055.0 98660.0 82760.0 100005.0 ;
      RECT  82055.0 101350.0 82760.0 100005.0 ;
      RECT  82055.0 101350.0 82760.0 102695.0 ;
      RECT  82055.0 104040.0 82760.0 102695.0 ;
      RECT  82055.0 104040.0 82760.0 105385.0 ;
      RECT  82055.0 106730.0 82760.0 105385.0 ;
      RECT  82055.0 106730.0 82760.0 108075.0 ;
      RECT  82055.0 109420.0 82760.0 108075.0 ;
      RECT  82055.0 109420.0 82760.0 110765.0 ;
      RECT  82055.0 112110.0 82760.0 110765.0 ;
      RECT  82055.0 112110.0 82760.0 113455.0 ;
      RECT  82055.0 114800.0 82760.0 113455.0 ;
      RECT  82055.0 114800.0 82760.0 116145.0 ;
      RECT  82055.0 117490.0 82760.0 116145.0 ;
      RECT  82055.0 117490.0 82760.0 118835.0 ;
      RECT  82055.0 120180.0 82760.0 118835.0 ;
      RECT  82055.0 120180.0 82760.0 121525.0 ;
      RECT  82055.0 122870.0 82760.0 121525.0 ;
      RECT  82055.0 122870.0 82760.0 124215.0 ;
      RECT  82055.0 125560.0 82760.0 124215.0 ;
      RECT  82055.0 125560.0 82760.0 126905.0 ;
      RECT  82055.0 128250.0 82760.0 126905.0 ;
      RECT  82055.0 128250.0 82760.0 129595.0 ;
      RECT  82055.0 130940.0 82760.0 129595.0 ;
      RECT  82055.0 130940.0 82760.0 132285.0 ;
      RECT  82055.0 133630.0 82760.0 132285.0 ;
      RECT  82055.0 133630.0 82760.0 134975.0 ;
      RECT  82055.0 136320.0 82760.0 134975.0 ;
      RECT  82055.0 136320.0 82760.0 137665.0 ;
      RECT  82055.0 139010.0 82760.0 137665.0 ;
      RECT  82055.0 139010.0 82760.0 140355.0 ;
      RECT  82055.0 141700.0 82760.0 140355.0 ;
      RECT  82055.0 141700.0 82760.0 143045.0 ;
      RECT  82055.0 144390.0 82760.0 143045.0 ;
      RECT  82055.0 144390.0 82760.0 145735.0 ;
      RECT  82055.0 147080.0 82760.0 145735.0 ;
      RECT  82055.0 147080.0 82760.0 148425.0 ;
      RECT  82055.0 149770.0 82760.0 148425.0 ;
      RECT  82055.0 149770.0 82760.0 151115.0 ;
      RECT  82055.0 152460.0 82760.0 151115.0 ;
      RECT  82055.0 152460.0 82760.0 153805.0 ;
      RECT  82055.0 155150.0 82760.0 153805.0 ;
      RECT  82055.0 155150.0 82760.0 156495.0 ;
      RECT  82055.0 157840.0 82760.0 156495.0 ;
      RECT  82055.0 157840.0 82760.0 159185.0 ;
      RECT  82055.0 160530.0 82760.0 159185.0 ;
      RECT  82055.0 160530.0 82760.0 161875.0 ;
      RECT  82055.0 163220.0 82760.0 161875.0 ;
      RECT  82055.0 163220.0 82760.0 164565.0 ;
      RECT  82055.0 165910.0 82760.0 164565.0 ;
      RECT  82055.0 165910.0 82760.0 167255.0 ;
      RECT  82055.0 168600.0 82760.0 167255.0 ;
      RECT  82055.0 168600.0 82760.0 169945.0 ;
      RECT  82055.0 171290.0 82760.0 169945.0 ;
      RECT  82055.0 171290.0 82760.0 172635.0 ;
      RECT  82055.0 173980.0 82760.0 172635.0 ;
      RECT  82055.0 173980.0 82760.0 175325.0 ;
      RECT  82055.0 176670.0 82760.0 175325.0 ;
      RECT  82055.0 176670.0 82760.0 178015.0 ;
      RECT  82055.0 179360.0 82760.0 178015.0 ;
      RECT  82055.0 179360.0 82760.0 180705.0 ;
      RECT  82055.0 182050.0 82760.0 180705.0 ;
      RECT  82055.0 182050.0 82760.0 183395.0 ;
      RECT  82055.0 184740.0 82760.0 183395.0 ;
      RECT  82055.0 184740.0 82760.0 186085.0 ;
      RECT  82055.0 187430.0 82760.0 186085.0 ;
      RECT  82055.0 187430.0 82760.0 188775.0 ;
      RECT  82055.0 190120.0 82760.0 188775.0 ;
      RECT  82055.0 190120.0 82760.0 191465.0 ;
      RECT  82055.0 192810.0 82760.0 191465.0 ;
      RECT  82055.0 192810.0 82760.0 194155.0 ;
      RECT  82055.0 195500.0 82760.0 194155.0 ;
      RECT  82055.0 195500.0 82760.0 196845.0 ;
      RECT  82055.0 198190.0 82760.0 196845.0 ;
      RECT  82055.0 198190.0 82760.0 199535.0 ;
      RECT  82055.0 200880.0 82760.0 199535.0 ;
      RECT  82055.0 200880.0 82760.0 202225.0 ;
      RECT  82055.0 203570.0 82760.0 202225.0 ;
      RECT  82055.0 203570.0 82760.0 204915.0 ;
      RECT  82055.0 206260.0 82760.0 204915.0 ;
      RECT  82760.0 34100.0 83465.0 35445.0 ;
      RECT  82760.0 36790.0 83465.0 35445.0 ;
      RECT  82760.0 36790.0 83465.0 38135.0 ;
      RECT  82760.0 39480.0 83465.0 38135.0 ;
      RECT  82760.0 39480.0 83465.0 40825.0 ;
      RECT  82760.0 42170.0 83465.0 40825.0 ;
      RECT  82760.0 42170.0 83465.0 43515.0 ;
      RECT  82760.0 44860.0 83465.0 43515.0 ;
      RECT  82760.0 44860.0 83465.0 46205.0 ;
      RECT  82760.0 47550.0 83465.0 46205.0 ;
      RECT  82760.0 47550.0 83465.0 48895.0 ;
      RECT  82760.0 50240.0 83465.0 48895.0 ;
      RECT  82760.0 50240.0 83465.0 51585.0 ;
      RECT  82760.0 52930.0 83465.0 51585.0 ;
      RECT  82760.0 52930.0 83465.0 54275.0 ;
      RECT  82760.0 55620.0 83465.0 54275.0 ;
      RECT  82760.0 55620.0 83465.0 56965.0 ;
      RECT  82760.0 58310.0 83465.0 56965.0 ;
      RECT  82760.0 58310.0 83465.0 59655.0 ;
      RECT  82760.0 61000.0 83465.0 59655.0 ;
      RECT  82760.0 61000.0 83465.0 62345.0 ;
      RECT  82760.0 63690.0 83465.0 62345.0 ;
      RECT  82760.0 63690.0 83465.0 65035.0 ;
      RECT  82760.0 66380.0 83465.0 65035.0 ;
      RECT  82760.0 66380.0 83465.0 67725.0 ;
      RECT  82760.0 69070.0 83465.0 67725.0 ;
      RECT  82760.0 69070.0 83465.0 70415.0 ;
      RECT  82760.0 71760.0 83465.0 70415.0 ;
      RECT  82760.0 71760.0 83465.0 73105.0 ;
      RECT  82760.0 74450.0 83465.0 73105.0 ;
      RECT  82760.0 74450.0 83465.0 75795.0 ;
      RECT  82760.0 77140.0 83465.0 75795.0 ;
      RECT  82760.0 77140.0 83465.0 78485.0 ;
      RECT  82760.0 79830.0 83465.0 78485.0 ;
      RECT  82760.0 79830.0 83465.0 81175.0 ;
      RECT  82760.0 82520.0 83465.0 81175.0 ;
      RECT  82760.0 82520.0 83465.0 83865.0 ;
      RECT  82760.0 85210.0 83465.0 83865.0 ;
      RECT  82760.0 85210.0 83465.0 86555.0 ;
      RECT  82760.0 87900.0 83465.0 86555.0 ;
      RECT  82760.0 87900.0 83465.0 89245.0 ;
      RECT  82760.0 90590.0 83465.0 89245.0 ;
      RECT  82760.0 90590.0 83465.0 91935.0 ;
      RECT  82760.0 93280.0 83465.0 91935.0 ;
      RECT  82760.0 93280.0 83465.0 94625.0 ;
      RECT  82760.0 95970.0 83465.0 94625.0 ;
      RECT  82760.0 95970.0 83465.0 97315.0 ;
      RECT  82760.0 98660.0 83465.0 97315.0 ;
      RECT  82760.0 98660.0 83465.0 100005.0 ;
      RECT  82760.0 101350.0 83465.0 100005.0 ;
      RECT  82760.0 101350.0 83465.0 102695.0 ;
      RECT  82760.0 104040.0 83465.0 102695.0 ;
      RECT  82760.0 104040.0 83465.0 105385.0 ;
      RECT  82760.0 106730.0 83465.0 105385.0 ;
      RECT  82760.0 106730.0 83465.0 108075.0 ;
      RECT  82760.0 109420.0 83465.0 108075.0 ;
      RECT  82760.0 109420.0 83465.0 110765.0 ;
      RECT  82760.0 112110.0 83465.0 110765.0 ;
      RECT  82760.0 112110.0 83465.0 113455.0 ;
      RECT  82760.0 114800.0 83465.0 113455.0 ;
      RECT  82760.0 114800.0 83465.0 116145.0 ;
      RECT  82760.0 117490.0 83465.0 116145.0 ;
      RECT  82760.0 117490.0 83465.0 118835.0 ;
      RECT  82760.0 120180.0 83465.0 118835.0 ;
      RECT  82760.0 120180.0 83465.0 121525.0 ;
      RECT  82760.0 122870.0 83465.0 121525.0 ;
      RECT  82760.0 122870.0 83465.0 124215.0 ;
      RECT  82760.0 125560.0 83465.0 124215.0 ;
      RECT  82760.0 125560.0 83465.0 126905.0 ;
      RECT  82760.0 128250.0 83465.0 126905.0 ;
      RECT  82760.0 128250.0 83465.0 129595.0 ;
      RECT  82760.0 130940.0 83465.0 129595.0 ;
      RECT  82760.0 130940.0 83465.0 132285.0 ;
      RECT  82760.0 133630.0 83465.0 132285.0 ;
      RECT  82760.0 133630.0 83465.0 134975.0 ;
      RECT  82760.0 136320.0 83465.0 134975.0 ;
      RECT  82760.0 136320.0 83465.0 137665.0 ;
      RECT  82760.0 139010.0 83465.0 137665.0 ;
      RECT  82760.0 139010.0 83465.0 140355.0 ;
      RECT  82760.0 141700.0 83465.0 140355.0 ;
      RECT  82760.0 141700.0 83465.0 143045.0 ;
      RECT  82760.0 144390.0 83465.0 143045.0 ;
      RECT  82760.0 144390.0 83465.0 145735.0 ;
      RECT  82760.0 147080.0 83465.0 145735.0 ;
      RECT  82760.0 147080.0 83465.0 148425.0 ;
      RECT  82760.0 149770.0 83465.0 148425.0 ;
      RECT  82760.0 149770.0 83465.0 151115.0 ;
      RECT  82760.0 152460.0 83465.0 151115.0 ;
      RECT  82760.0 152460.0 83465.0 153805.0 ;
      RECT  82760.0 155150.0 83465.0 153805.0 ;
      RECT  82760.0 155150.0 83465.0 156495.0 ;
      RECT  82760.0 157840.0 83465.0 156495.0 ;
      RECT  82760.0 157840.0 83465.0 159185.0 ;
      RECT  82760.0 160530.0 83465.0 159185.0 ;
      RECT  82760.0 160530.0 83465.0 161875.0 ;
      RECT  82760.0 163220.0 83465.0 161875.0 ;
      RECT  82760.0 163220.0 83465.0 164565.0 ;
      RECT  82760.0 165910.0 83465.0 164565.0 ;
      RECT  82760.0 165910.0 83465.0 167255.0 ;
      RECT  82760.0 168600.0 83465.0 167255.0 ;
      RECT  82760.0 168600.0 83465.0 169945.0 ;
      RECT  82760.0 171290.0 83465.0 169945.0 ;
      RECT  82760.0 171290.0 83465.0 172635.0 ;
      RECT  82760.0 173980.0 83465.0 172635.0 ;
      RECT  82760.0 173980.0 83465.0 175325.0 ;
      RECT  82760.0 176670.0 83465.0 175325.0 ;
      RECT  82760.0 176670.0 83465.0 178015.0 ;
      RECT  82760.0 179360.0 83465.0 178015.0 ;
      RECT  82760.0 179360.0 83465.0 180705.0 ;
      RECT  82760.0 182050.0 83465.0 180705.0 ;
      RECT  82760.0 182050.0 83465.0 183395.0 ;
      RECT  82760.0 184740.0 83465.0 183395.0 ;
      RECT  82760.0 184740.0 83465.0 186085.0 ;
      RECT  82760.0 187430.0 83465.0 186085.0 ;
      RECT  82760.0 187430.0 83465.0 188775.0 ;
      RECT  82760.0 190120.0 83465.0 188775.0 ;
      RECT  82760.0 190120.0 83465.0 191465.0 ;
      RECT  82760.0 192810.0 83465.0 191465.0 ;
      RECT  82760.0 192810.0 83465.0 194155.0 ;
      RECT  82760.0 195500.0 83465.0 194155.0 ;
      RECT  82760.0 195500.0 83465.0 196845.0 ;
      RECT  82760.0 198190.0 83465.0 196845.0 ;
      RECT  82760.0 198190.0 83465.0 199535.0 ;
      RECT  82760.0 200880.0 83465.0 199535.0 ;
      RECT  82760.0 200880.0 83465.0 202225.0 ;
      RECT  82760.0 203570.0 83465.0 202225.0 ;
      RECT  82760.0 203570.0 83465.0 204915.0 ;
      RECT  82760.0 206260.0 83465.0 204915.0 ;
      RECT  83465.0 34100.0 84170.0 35445.0 ;
      RECT  83465.0 36790.0 84170.0 35445.0 ;
      RECT  83465.0 36790.0 84170.0 38135.0 ;
      RECT  83465.0 39480.0 84170.0 38135.0 ;
      RECT  83465.0 39480.0 84170.0 40825.0 ;
      RECT  83465.0 42170.0 84170.0 40825.0 ;
      RECT  83465.0 42170.0 84170.0 43515.0 ;
      RECT  83465.0 44860.0 84170.0 43515.0 ;
      RECT  83465.0 44860.0 84170.0 46205.0 ;
      RECT  83465.0 47550.0 84170.0 46205.0 ;
      RECT  83465.0 47550.0 84170.0 48895.0 ;
      RECT  83465.0 50240.0 84170.0 48895.0 ;
      RECT  83465.0 50240.0 84170.0 51585.0 ;
      RECT  83465.0 52930.0 84170.0 51585.0 ;
      RECT  83465.0 52930.0 84170.0 54275.0 ;
      RECT  83465.0 55620.0 84170.0 54275.0 ;
      RECT  83465.0 55620.0 84170.0 56965.0 ;
      RECT  83465.0 58310.0 84170.0 56965.0 ;
      RECT  83465.0 58310.0 84170.0 59655.0 ;
      RECT  83465.0 61000.0 84170.0 59655.0 ;
      RECT  83465.0 61000.0 84170.0 62345.0 ;
      RECT  83465.0 63690.0 84170.0 62345.0 ;
      RECT  83465.0 63690.0 84170.0 65035.0 ;
      RECT  83465.0 66380.0 84170.0 65035.0 ;
      RECT  83465.0 66380.0 84170.0 67725.0 ;
      RECT  83465.0 69070.0 84170.0 67725.0 ;
      RECT  83465.0 69070.0 84170.0 70415.0 ;
      RECT  83465.0 71760.0 84170.0 70415.0 ;
      RECT  83465.0 71760.0 84170.0 73105.0 ;
      RECT  83465.0 74450.0 84170.0 73105.0 ;
      RECT  83465.0 74450.0 84170.0 75795.0 ;
      RECT  83465.0 77140.0 84170.0 75795.0 ;
      RECT  83465.0 77140.0 84170.0 78485.0 ;
      RECT  83465.0 79830.0 84170.0 78485.0 ;
      RECT  83465.0 79830.0 84170.0 81175.0 ;
      RECT  83465.0 82520.0 84170.0 81175.0 ;
      RECT  83465.0 82520.0 84170.0 83865.0 ;
      RECT  83465.0 85210.0 84170.0 83865.0 ;
      RECT  83465.0 85210.0 84170.0 86555.0 ;
      RECT  83465.0 87900.0 84170.0 86555.0 ;
      RECT  83465.0 87900.0 84170.0 89245.0 ;
      RECT  83465.0 90590.0 84170.0 89245.0 ;
      RECT  83465.0 90590.0 84170.0 91935.0 ;
      RECT  83465.0 93280.0 84170.0 91935.0 ;
      RECT  83465.0 93280.0 84170.0 94625.0 ;
      RECT  83465.0 95970.0 84170.0 94625.0 ;
      RECT  83465.0 95970.0 84170.0 97315.0 ;
      RECT  83465.0 98660.0 84170.0 97315.0 ;
      RECT  83465.0 98660.0 84170.0 100005.0 ;
      RECT  83465.0 101350.0 84170.0 100005.0 ;
      RECT  83465.0 101350.0 84170.0 102695.0 ;
      RECT  83465.0 104040.0 84170.0 102695.0 ;
      RECT  83465.0 104040.0 84170.0 105385.0 ;
      RECT  83465.0 106730.0 84170.0 105385.0 ;
      RECT  83465.0 106730.0 84170.0 108075.0 ;
      RECT  83465.0 109420.0 84170.0 108075.0 ;
      RECT  83465.0 109420.0 84170.0 110765.0 ;
      RECT  83465.0 112110.0 84170.0 110765.0 ;
      RECT  83465.0 112110.0 84170.0 113455.0 ;
      RECT  83465.0 114800.0 84170.0 113455.0 ;
      RECT  83465.0 114800.0 84170.0 116145.0 ;
      RECT  83465.0 117490.0 84170.0 116145.0 ;
      RECT  83465.0 117490.0 84170.0 118835.0 ;
      RECT  83465.0 120180.0 84170.0 118835.0 ;
      RECT  83465.0 120180.0 84170.0 121525.0 ;
      RECT  83465.0 122870.0 84170.0 121525.0 ;
      RECT  83465.0 122870.0 84170.0 124215.0 ;
      RECT  83465.0 125560.0 84170.0 124215.0 ;
      RECT  83465.0 125560.0 84170.0 126905.0 ;
      RECT  83465.0 128250.0 84170.0 126905.0 ;
      RECT  83465.0 128250.0 84170.0 129595.0 ;
      RECT  83465.0 130940.0 84170.0 129595.0 ;
      RECT  83465.0 130940.0 84170.0 132285.0 ;
      RECT  83465.0 133630.0 84170.0 132285.0 ;
      RECT  83465.0 133630.0 84170.0 134975.0 ;
      RECT  83465.0 136320.0 84170.0 134975.0 ;
      RECT  83465.0 136320.0 84170.0 137665.0 ;
      RECT  83465.0 139010.0 84170.0 137665.0 ;
      RECT  83465.0 139010.0 84170.0 140355.0 ;
      RECT  83465.0 141700.0 84170.0 140355.0 ;
      RECT  83465.0 141700.0 84170.0 143045.0 ;
      RECT  83465.0 144390.0 84170.0 143045.0 ;
      RECT  83465.0 144390.0 84170.0 145735.0 ;
      RECT  83465.0 147080.0 84170.0 145735.0 ;
      RECT  83465.0 147080.0 84170.0 148425.0 ;
      RECT  83465.0 149770.0 84170.0 148425.0 ;
      RECT  83465.0 149770.0 84170.0 151115.0 ;
      RECT  83465.0 152460.0 84170.0 151115.0 ;
      RECT  83465.0 152460.0 84170.0 153805.0 ;
      RECT  83465.0 155150.0 84170.0 153805.0 ;
      RECT  83465.0 155150.0 84170.0 156495.0 ;
      RECT  83465.0 157840.0 84170.0 156495.0 ;
      RECT  83465.0 157840.0 84170.0 159185.0 ;
      RECT  83465.0 160530.0 84170.0 159185.0 ;
      RECT  83465.0 160530.0 84170.0 161875.0 ;
      RECT  83465.0 163220.0 84170.0 161875.0 ;
      RECT  83465.0 163220.0 84170.0 164565.0 ;
      RECT  83465.0 165910.0 84170.0 164565.0 ;
      RECT  83465.0 165910.0 84170.0 167255.0 ;
      RECT  83465.0 168600.0 84170.0 167255.0 ;
      RECT  83465.0 168600.0 84170.0 169945.0 ;
      RECT  83465.0 171290.0 84170.0 169945.0 ;
      RECT  83465.0 171290.0 84170.0 172635.0 ;
      RECT  83465.0 173980.0 84170.0 172635.0 ;
      RECT  83465.0 173980.0 84170.0 175325.0 ;
      RECT  83465.0 176670.0 84170.0 175325.0 ;
      RECT  83465.0 176670.0 84170.0 178015.0 ;
      RECT  83465.0 179360.0 84170.0 178015.0 ;
      RECT  83465.0 179360.0 84170.0 180705.0 ;
      RECT  83465.0 182050.0 84170.0 180705.0 ;
      RECT  83465.0 182050.0 84170.0 183395.0 ;
      RECT  83465.0 184740.0 84170.0 183395.0 ;
      RECT  83465.0 184740.0 84170.0 186085.0 ;
      RECT  83465.0 187430.0 84170.0 186085.0 ;
      RECT  83465.0 187430.0 84170.0 188775.0 ;
      RECT  83465.0 190120.0 84170.0 188775.0 ;
      RECT  83465.0 190120.0 84170.0 191465.0 ;
      RECT  83465.0 192810.0 84170.0 191465.0 ;
      RECT  83465.0 192810.0 84170.0 194155.0 ;
      RECT  83465.0 195500.0 84170.0 194155.0 ;
      RECT  83465.0 195500.0 84170.0 196845.0 ;
      RECT  83465.0 198190.0 84170.0 196845.0 ;
      RECT  83465.0 198190.0 84170.0 199535.0 ;
      RECT  83465.0 200880.0 84170.0 199535.0 ;
      RECT  83465.0 200880.0 84170.0 202225.0 ;
      RECT  83465.0 203570.0 84170.0 202225.0 ;
      RECT  83465.0 203570.0 84170.0 204915.0 ;
      RECT  83465.0 206260.0 84170.0 204915.0 ;
      RECT  84170.0 34100.0 84875.0 35445.0 ;
      RECT  84170.0 36790.0 84875.0 35445.0 ;
      RECT  84170.0 36790.0 84875.0 38135.0 ;
      RECT  84170.0 39480.0 84875.0 38135.0 ;
      RECT  84170.0 39480.0 84875.0 40825.0 ;
      RECT  84170.0 42170.0 84875.0 40825.0 ;
      RECT  84170.0 42170.0 84875.0 43515.0 ;
      RECT  84170.0 44860.0 84875.0 43515.0 ;
      RECT  84170.0 44860.0 84875.0 46205.0 ;
      RECT  84170.0 47550.0 84875.0 46205.0 ;
      RECT  84170.0 47550.0 84875.0 48895.0 ;
      RECT  84170.0 50240.0 84875.0 48895.0 ;
      RECT  84170.0 50240.0 84875.0 51585.0 ;
      RECT  84170.0 52930.0 84875.0 51585.0 ;
      RECT  84170.0 52930.0 84875.0 54275.0 ;
      RECT  84170.0 55620.0 84875.0 54275.0 ;
      RECT  84170.0 55620.0 84875.0 56965.0 ;
      RECT  84170.0 58310.0 84875.0 56965.0 ;
      RECT  84170.0 58310.0 84875.0 59655.0 ;
      RECT  84170.0 61000.0 84875.0 59655.0 ;
      RECT  84170.0 61000.0 84875.0 62345.0 ;
      RECT  84170.0 63690.0 84875.0 62345.0 ;
      RECT  84170.0 63690.0 84875.0 65035.0 ;
      RECT  84170.0 66380.0 84875.0 65035.0 ;
      RECT  84170.0 66380.0 84875.0 67725.0 ;
      RECT  84170.0 69070.0 84875.0 67725.0 ;
      RECT  84170.0 69070.0 84875.0 70415.0 ;
      RECT  84170.0 71760.0 84875.0 70415.0 ;
      RECT  84170.0 71760.0 84875.0 73105.0 ;
      RECT  84170.0 74450.0 84875.0 73105.0 ;
      RECT  84170.0 74450.0 84875.0 75795.0 ;
      RECT  84170.0 77140.0 84875.0 75795.0 ;
      RECT  84170.0 77140.0 84875.0 78485.0 ;
      RECT  84170.0 79830.0 84875.0 78485.0 ;
      RECT  84170.0 79830.0 84875.0 81175.0 ;
      RECT  84170.0 82520.0 84875.0 81175.0 ;
      RECT  84170.0 82520.0 84875.0 83865.0 ;
      RECT  84170.0 85210.0 84875.0 83865.0 ;
      RECT  84170.0 85210.0 84875.0 86555.0 ;
      RECT  84170.0 87900.0 84875.0 86555.0 ;
      RECT  84170.0 87900.0 84875.0 89245.0 ;
      RECT  84170.0 90590.0 84875.0 89245.0 ;
      RECT  84170.0 90590.0 84875.0 91935.0 ;
      RECT  84170.0 93280.0 84875.0 91935.0 ;
      RECT  84170.0 93280.0 84875.0 94625.0 ;
      RECT  84170.0 95970.0 84875.0 94625.0 ;
      RECT  84170.0 95970.0 84875.0 97315.0 ;
      RECT  84170.0 98660.0 84875.0 97315.0 ;
      RECT  84170.0 98660.0 84875.0 100005.0 ;
      RECT  84170.0 101350.0 84875.0 100005.0 ;
      RECT  84170.0 101350.0 84875.0 102695.0 ;
      RECT  84170.0 104040.0 84875.0 102695.0 ;
      RECT  84170.0 104040.0 84875.0 105385.0 ;
      RECT  84170.0 106730.0 84875.0 105385.0 ;
      RECT  84170.0 106730.0 84875.0 108075.0 ;
      RECT  84170.0 109420.0 84875.0 108075.0 ;
      RECT  84170.0 109420.0 84875.0 110765.0 ;
      RECT  84170.0 112110.0 84875.0 110765.0 ;
      RECT  84170.0 112110.0 84875.0 113455.0 ;
      RECT  84170.0 114800.0 84875.0 113455.0 ;
      RECT  84170.0 114800.0 84875.0 116145.0 ;
      RECT  84170.0 117490.0 84875.0 116145.0 ;
      RECT  84170.0 117490.0 84875.0 118835.0 ;
      RECT  84170.0 120180.0 84875.0 118835.0 ;
      RECT  84170.0 120180.0 84875.0 121525.0 ;
      RECT  84170.0 122870.0 84875.0 121525.0 ;
      RECT  84170.0 122870.0 84875.0 124215.0 ;
      RECT  84170.0 125560.0 84875.0 124215.0 ;
      RECT  84170.0 125560.0 84875.0 126905.0 ;
      RECT  84170.0 128250.0 84875.0 126905.0 ;
      RECT  84170.0 128250.0 84875.0 129595.0 ;
      RECT  84170.0 130940.0 84875.0 129595.0 ;
      RECT  84170.0 130940.0 84875.0 132285.0 ;
      RECT  84170.0 133630.0 84875.0 132285.0 ;
      RECT  84170.0 133630.0 84875.0 134975.0 ;
      RECT  84170.0 136320.0 84875.0 134975.0 ;
      RECT  84170.0 136320.0 84875.0 137665.0 ;
      RECT  84170.0 139010.0 84875.0 137665.0 ;
      RECT  84170.0 139010.0 84875.0 140355.0 ;
      RECT  84170.0 141700.0 84875.0 140355.0 ;
      RECT  84170.0 141700.0 84875.0 143045.0 ;
      RECT  84170.0 144390.0 84875.0 143045.0 ;
      RECT  84170.0 144390.0 84875.0 145735.0 ;
      RECT  84170.0 147080.0 84875.0 145735.0 ;
      RECT  84170.0 147080.0 84875.0 148425.0 ;
      RECT  84170.0 149770.0 84875.0 148425.0 ;
      RECT  84170.0 149770.0 84875.0 151115.0 ;
      RECT  84170.0 152460.0 84875.0 151115.0 ;
      RECT  84170.0 152460.0 84875.0 153805.0 ;
      RECT  84170.0 155150.0 84875.0 153805.0 ;
      RECT  84170.0 155150.0 84875.0 156495.0 ;
      RECT  84170.0 157840.0 84875.0 156495.0 ;
      RECT  84170.0 157840.0 84875.0 159185.0 ;
      RECT  84170.0 160530.0 84875.0 159185.0 ;
      RECT  84170.0 160530.0 84875.0 161875.0 ;
      RECT  84170.0 163220.0 84875.0 161875.0 ;
      RECT  84170.0 163220.0 84875.0 164565.0 ;
      RECT  84170.0 165910.0 84875.0 164565.0 ;
      RECT  84170.0 165910.0 84875.0 167255.0 ;
      RECT  84170.0 168600.0 84875.0 167255.0 ;
      RECT  84170.0 168600.0 84875.0 169945.0 ;
      RECT  84170.0 171290.0 84875.0 169945.0 ;
      RECT  84170.0 171290.0 84875.0 172635.0 ;
      RECT  84170.0 173980.0 84875.0 172635.0 ;
      RECT  84170.0 173980.0 84875.0 175325.0 ;
      RECT  84170.0 176670.0 84875.0 175325.0 ;
      RECT  84170.0 176670.0 84875.0 178015.0 ;
      RECT  84170.0 179360.0 84875.0 178015.0 ;
      RECT  84170.0 179360.0 84875.0 180705.0 ;
      RECT  84170.0 182050.0 84875.0 180705.0 ;
      RECT  84170.0 182050.0 84875.0 183395.0 ;
      RECT  84170.0 184740.0 84875.0 183395.0 ;
      RECT  84170.0 184740.0 84875.0 186085.0 ;
      RECT  84170.0 187430.0 84875.0 186085.0 ;
      RECT  84170.0 187430.0 84875.0 188775.0 ;
      RECT  84170.0 190120.0 84875.0 188775.0 ;
      RECT  84170.0 190120.0 84875.0 191465.0 ;
      RECT  84170.0 192810.0 84875.0 191465.0 ;
      RECT  84170.0 192810.0 84875.0 194155.0 ;
      RECT  84170.0 195500.0 84875.0 194155.0 ;
      RECT  84170.0 195500.0 84875.0 196845.0 ;
      RECT  84170.0 198190.0 84875.0 196845.0 ;
      RECT  84170.0 198190.0 84875.0 199535.0 ;
      RECT  84170.0 200880.0 84875.0 199535.0 ;
      RECT  84170.0 200880.0 84875.0 202225.0 ;
      RECT  84170.0 203570.0 84875.0 202225.0 ;
      RECT  84170.0 203570.0 84875.0 204915.0 ;
      RECT  84170.0 206260.0 84875.0 204915.0 ;
      RECT  84875.0 34100.0 85580.0 35445.0 ;
      RECT  84875.0 36790.0 85580.0 35445.0 ;
      RECT  84875.0 36790.0 85580.0 38135.0 ;
      RECT  84875.0 39480.0 85580.0 38135.0 ;
      RECT  84875.0 39480.0 85580.0 40825.0 ;
      RECT  84875.0 42170.0 85580.0 40825.0 ;
      RECT  84875.0 42170.0 85580.0 43515.0 ;
      RECT  84875.0 44860.0 85580.0 43515.0 ;
      RECT  84875.0 44860.0 85580.0 46205.0 ;
      RECT  84875.0 47550.0 85580.0 46205.0 ;
      RECT  84875.0 47550.0 85580.0 48895.0 ;
      RECT  84875.0 50240.0 85580.0 48895.0 ;
      RECT  84875.0 50240.0 85580.0 51585.0 ;
      RECT  84875.0 52930.0 85580.0 51585.0 ;
      RECT  84875.0 52930.0 85580.0 54275.0 ;
      RECT  84875.0 55620.0 85580.0 54275.0 ;
      RECT  84875.0 55620.0 85580.0 56965.0 ;
      RECT  84875.0 58310.0 85580.0 56965.0 ;
      RECT  84875.0 58310.0 85580.0 59655.0 ;
      RECT  84875.0 61000.0 85580.0 59655.0 ;
      RECT  84875.0 61000.0 85580.0 62345.0 ;
      RECT  84875.0 63690.0 85580.0 62345.0 ;
      RECT  84875.0 63690.0 85580.0 65035.0 ;
      RECT  84875.0 66380.0 85580.0 65035.0 ;
      RECT  84875.0 66380.0 85580.0 67725.0 ;
      RECT  84875.0 69070.0 85580.0 67725.0 ;
      RECT  84875.0 69070.0 85580.0 70415.0 ;
      RECT  84875.0 71760.0 85580.0 70415.0 ;
      RECT  84875.0 71760.0 85580.0 73105.0 ;
      RECT  84875.0 74450.0 85580.0 73105.0 ;
      RECT  84875.0 74450.0 85580.0 75795.0 ;
      RECT  84875.0 77140.0 85580.0 75795.0 ;
      RECT  84875.0 77140.0 85580.0 78485.0 ;
      RECT  84875.0 79830.0 85580.0 78485.0 ;
      RECT  84875.0 79830.0 85580.0 81175.0 ;
      RECT  84875.0 82520.0 85580.0 81175.0 ;
      RECT  84875.0 82520.0 85580.0 83865.0 ;
      RECT  84875.0 85210.0 85580.0 83865.0 ;
      RECT  84875.0 85210.0 85580.0 86555.0 ;
      RECT  84875.0 87900.0 85580.0 86555.0 ;
      RECT  84875.0 87900.0 85580.0 89245.0 ;
      RECT  84875.0 90590.0 85580.0 89245.0 ;
      RECT  84875.0 90590.0 85580.0 91935.0 ;
      RECT  84875.0 93280.0 85580.0 91935.0 ;
      RECT  84875.0 93280.0 85580.0 94625.0 ;
      RECT  84875.0 95970.0 85580.0 94625.0 ;
      RECT  84875.0 95970.0 85580.0 97315.0 ;
      RECT  84875.0 98660.0 85580.0 97315.0 ;
      RECT  84875.0 98660.0 85580.0 100005.0 ;
      RECT  84875.0 101350.0 85580.0 100005.0 ;
      RECT  84875.0 101350.0 85580.0 102695.0 ;
      RECT  84875.0 104040.0 85580.0 102695.0 ;
      RECT  84875.0 104040.0 85580.0 105385.0 ;
      RECT  84875.0 106730.0 85580.0 105385.0 ;
      RECT  84875.0 106730.0 85580.0 108075.0 ;
      RECT  84875.0 109420.0 85580.0 108075.0 ;
      RECT  84875.0 109420.0 85580.0 110765.0 ;
      RECT  84875.0 112110.0 85580.0 110765.0 ;
      RECT  84875.0 112110.0 85580.0 113455.0 ;
      RECT  84875.0 114800.0 85580.0 113455.0 ;
      RECT  84875.0 114800.0 85580.0 116145.0 ;
      RECT  84875.0 117490.0 85580.0 116145.0 ;
      RECT  84875.0 117490.0 85580.0 118835.0 ;
      RECT  84875.0 120180.0 85580.0 118835.0 ;
      RECT  84875.0 120180.0 85580.0 121525.0 ;
      RECT  84875.0 122870.0 85580.0 121525.0 ;
      RECT  84875.0 122870.0 85580.0 124215.0 ;
      RECT  84875.0 125560.0 85580.0 124215.0 ;
      RECT  84875.0 125560.0 85580.0 126905.0 ;
      RECT  84875.0 128250.0 85580.0 126905.0 ;
      RECT  84875.0 128250.0 85580.0 129595.0 ;
      RECT  84875.0 130940.0 85580.0 129595.0 ;
      RECT  84875.0 130940.0 85580.0 132285.0 ;
      RECT  84875.0 133630.0 85580.0 132285.0 ;
      RECT  84875.0 133630.0 85580.0 134975.0 ;
      RECT  84875.0 136320.0 85580.0 134975.0 ;
      RECT  84875.0 136320.0 85580.0 137665.0 ;
      RECT  84875.0 139010.0 85580.0 137665.0 ;
      RECT  84875.0 139010.0 85580.0 140355.0 ;
      RECT  84875.0 141700.0 85580.0 140355.0 ;
      RECT  84875.0 141700.0 85580.0 143045.0 ;
      RECT  84875.0 144390.0 85580.0 143045.0 ;
      RECT  84875.0 144390.0 85580.0 145735.0 ;
      RECT  84875.0 147080.0 85580.0 145735.0 ;
      RECT  84875.0 147080.0 85580.0 148425.0 ;
      RECT  84875.0 149770.0 85580.0 148425.0 ;
      RECT  84875.0 149770.0 85580.0 151115.0 ;
      RECT  84875.0 152460.0 85580.0 151115.0 ;
      RECT  84875.0 152460.0 85580.0 153805.0 ;
      RECT  84875.0 155150.0 85580.0 153805.0 ;
      RECT  84875.0 155150.0 85580.0 156495.0 ;
      RECT  84875.0 157840.0 85580.0 156495.0 ;
      RECT  84875.0 157840.0 85580.0 159185.0 ;
      RECT  84875.0 160530.0 85580.0 159185.0 ;
      RECT  84875.0 160530.0 85580.0 161875.0 ;
      RECT  84875.0 163220.0 85580.0 161875.0 ;
      RECT  84875.0 163220.0 85580.0 164565.0 ;
      RECT  84875.0 165910.0 85580.0 164565.0 ;
      RECT  84875.0 165910.0 85580.0 167255.0 ;
      RECT  84875.0 168600.0 85580.0 167255.0 ;
      RECT  84875.0 168600.0 85580.0 169945.0 ;
      RECT  84875.0 171290.0 85580.0 169945.0 ;
      RECT  84875.0 171290.0 85580.0 172635.0 ;
      RECT  84875.0 173980.0 85580.0 172635.0 ;
      RECT  84875.0 173980.0 85580.0 175325.0 ;
      RECT  84875.0 176670.0 85580.0 175325.0 ;
      RECT  84875.0 176670.0 85580.0 178015.0 ;
      RECT  84875.0 179360.0 85580.0 178015.0 ;
      RECT  84875.0 179360.0 85580.0 180705.0 ;
      RECT  84875.0 182050.0 85580.0 180705.0 ;
      RECT  84875.0 182050.0 85580.0 183395.0 ;
      RECT  84875.0 184740.0 85580.0 183395.0 ;
      RECT  84875.0 184740.0 85580.0 186085.0 ;
      RECT  84875.0 187430.0 85580.0 186085.0 ;
      RECT  84875.0 187430.0 85580.0 188775.0 ;
      RECT  84875.0 190120.0 85580.0 188775.0 ;
      RECT  84875.0 190120.0 85580.0 191465.0 ;
      RECT  84875.0 192810.0 85580.0 191465.0 ;
      RECT  84875.0 192810.0 85580.0 194155.0 ;
      RECT  84875.0 195500.0 85580.0 194155.0 ;
      RECT  84875.0 195500.0 85580.0 196845.0 ;
      RECT  84875.0 198190.0 85580.0 196845.0 ;
      RECT  84875.0 198190.0 85580.0 199535.0 ;
      RECT  84875.0 200880.0 85580.0 199535.0 ;
      RECT  84875.0 200880.0 85580.0 202225.0 ;
      RECT  84875.0 203570.0 85580.0 202225.0 ;
      RECT  84875.0 203570.0 85580.0 204915.0 ;
      RECT  84875.0 206260.0 85580.0 204915.0 ;
      RECT  85580.0 34100.0 86285.0 35445.0 ;
      RECT  85580.0 36790.0 86285.0 35445.0 ;
      RECT  85580.0 36790.0 86285.0 38135.0 ;
      RECT  85580.0 39480.0 86285.0 38135.0 ;
      RECT  85580.0 39480.0 86285.0 40825.0 ;
      RECT  85580.0 42170.0 86285.0 40825.0 ;
      RECT  85580.0 42170.0 86285.0 43515.0 ;
      RECT  85580.0 44860.0 86285.0 43515.0 ;
      RECT  85580.0 44860.0 86285.0 46205.0 ;
      RECT  85580.0 47550.0 86285.0 46205.0 ;
      RECT  85580.0 47550.0 86285.0 48895.0 ;
      RECT  85580.0 50240.0 86285.0 48895.0 ;
      RECT  85580.0 50240.0 86285.0 51585.0 ;
      RECT  85580.0 52930.0 86285.0 51585.0 ;
      RECT  85580.0 52930.0 86285.0 54275.0 ;
      RECT  85580.0 55620.0 86285.0 54275.0 ;
      RECT  85580.0 55620.0 86285.0 56965.0 ;
      RECT  85580.0 58310.0 86285.0 56965.0 ;
      RECT  85580.0 58310.0 86285.0 59655.0 ;
      RECT  85580.0 61000.0 86285.0 59655.0 ;
      RECT  85580.0 61000.0 86285.0 62345.0 ;
      RECT  85580.0 63690.0 86285.0 62345.0 ;
      RECT  85580.0 63690.0 86285.0 65035.0 ;
      RECT  85580.0 66380.0 86285.0 65035.0 ;
      RECT  85580.0 66380.0 86285.0 67725.0 ;
      RECT  85580.0 69070.0 86285.0 67725.0 ;
      RECT  85580.0 69070.0 86285.0 70415.0 ;
      RECT  85580.0 71760.0 86285.0 70415.0 ;
      RECT  85580.0 71760.0 86285.0 73105.0 ;
      RECT  85580.0 74450.0 86285.0 73105.0 ;
      RECT  85580.0 74450.0 86285.0 75795.0 ;
      RECT  85580.0 77140.0 86285.0 75795.0 ;
      RECT  85580.0 77140.0 86285.0 78485.0 ;
      RECT  85580.0 79830.0 86285.0 78485.0 ;
      RECT  85580.0 79830.0 86285.0 81175.0 ;
      RECT  85580.0 82520.0 86285.0 81175.0 ;
      RECT  85580.0 82520.0 86285.0 83865.0 ;
      RECT  85580.0 85210.0 86285.0 83865.0 ;
      RECT  85580.0 85210.0 86285.0 86555.0 ;
      RECT  85580.0 87900.0 86285.0 86555.0 ;
      RECT  85580.0 87900.0 86285.0 89245.0 ;
      RECT  85580.0 90590.0 86285.0 89245.0 ;
      RECT  85580.0 90590.0 86285.0 91935.0 ;
      RECT  85580.0 93280.0 86285.0 91935.0 ;
      RECT  85580.0 93280.0 86285.0 94625.0 ;
      RECT  85580.0 95970.0 86285.0 94625.0 ;
      RECT  85580.0 95970.0 86285.0 97315.0 ;
      RECT  85580.0 98660.0 86285.0 97315.0 ;
      RECT  85580.0 98660.0 86285.0 100005.0 ;
      RECT  85580.0 101350.0 86285.0 100005.0 ;
      RECT  85580.0 101350.0 86285.0 102695.0 ;
      RECT  85580.0 104040.0 86285.0 102695.0 ;
      RECT  85580.0 104040.0 86285.0 105385.0 ;
      RECT  85580.0 106730.0 86285.0 105385.0 ;
      RECT  85580.0 106730.0 86285.0 108075.0 ;
      RECT  85580.0 109420.0 86285.0 108075.0 ;
      RECT  85580.0 109420.0 86285.0 110765.0 ;
      RECT  85580.0 112110.0 86285.0 110765.0 ;
      RECT  85580.0 112110.0 86285.0 113455.0 ;
      RECT  85580.0 114800.0 86285.0 113455.0 ;
      RECT  85580.0 114800.0 86285.0 116145.0 ;
      RECT  85580.0 117490.0 86285.0 116145.0 ;
      RECT  85580.0 117490.0 86285.0 118835.0 ;
      RECT  85580.0 120180.0 86285.0 118835.0 ;
      RECT  85580.0 120180.0 86285.0 121525.0 ;
      RECT  85580.0 122870.0 86285.0 121525.0 ;
      RECT  85580.0 122870.0 86285.0 124215.0 ;
      RECT  85580.0 125560.0 86285.0 124215.0 ;
      RECT  85580.0 125560.0 86285.0 126905.0 ;
      RECT  85580.0 128250.0 86285.0 126905.0 ;
      RECT  85580.0 128250.0 86285.0 129595.0 ;
      RECT  85580.0 130940.0 86285.0 129595.0 ;
      RECT  85580.0 130940.0 86285.0 132285.0 ;
      RECT  85580.0 133630.0 86285.0 132285.0 ;
      RECT  85580.0 133630.0 86285.0 134975.0 ;
      RECT  85580.0 136320.0 86285.0 134975.0 ;
      RECT  85580.0 136320.0 86285.0 137665.0 ;
      RECT  85580.0 139010.0 86285.0 137665.0 ;
      RECT  85580.0 139010.0 86285.0 140355.0 ;
      RECT  85580.0 141700.0 86285.0 140355.0 ;
      RECT  85580.0 141700.0 86285.0 143045.0 ;
      RECT  85580.0 144390.0 86285.0 143045.0 ;
      RECT  85580.0 144390.0 86285.0 145735.0 ;
      RECT  85580.0 147080.0 86285.0 145735.0 ;
      RECT  85580.0 147080.0 86285.0 148425.0 ;
      RECT  85580.0 149770.0 86285.0 148425.0 ;
      RECT  85580.0 149770.0 86285.0 151115.0 ;
      RECT  85580.0 152460.0 86285.0 151115.0 ;
      RECT  85580.0 152460.0 86285.0 153805.0 ;
      RECT  85580.0 155150.0 86285.0 153805.0 ;
      RECT  85580.0 155150.0 86285.0 156495.0 ;
      RECT  85580.0 157840.0 86285.0 156495.0 ;
      RECT  85580.0 157840.0 86285.0 159185.0 ;
      RECT  85580.0 160530.0 86285.0 159185.0 ;
      RECT  85580.0 160530.0 86285.0 161875.0 ;
      RECT  85580.0 163220.0 86285.0 161875.0 ;
      RECT  85580.0 163220.0 86285.0 164565.0 ;
      RECT  85580.0 165910.0 86285.0 164565.0 ;
      RECT  85580.0 165910.0 86285.0 167255.0 ;
      RECT  85580.0 168600.0 86285.0 167255.0 ;
      RECT  85580.0 168600.0 86285.0 169945.0 ;
      RECT  85580.0 171290.0 86285.0 169945.0 ;
      RECT  85580.0 171290.0 86285.0 172635.0 ;
      RECT  85580.0 173980.0 86285.0 172635.0 ;
      RECT  85580.0 173980.0 86285.0 175325.0 ;
      RECT  85580.0 176670.0 86285.0 175325.0 ;
      RECT  85580.0 176670.0 86285.0 178015.0 ;
      RECT  85580.0 179360.0 86285.0 178015.0 ;
      RECT  85580.0 179360.0 86285.0 180705.0 ;
      RECT  85580.0 182050.0 86285.0 180705.0 ;
      RECT  85580.0 182050.0 86285.0 183395.0 ;
      RECT  85580.0 184740.0 86285.0 183395.0 ;
      RECT  85580.0 184740.0 86285.0 186085.0 ;
      RECT  85580.0 187430.0 86285.0 186085.0 ;
      RECT  85580.0 187430.0 86285.0 188775.0 ;
      RECT  85580.0 190120.0 86285.0 188775.0 ;
      RECT  85580.0 190120.0 86285.0 191465.0 ;
      RECT  85580.0 192810.0 86285.0 191465.0 ;
      RECT  85580.0 192810.0 86285.0 194155.0 ;
      RECT  85580.0 195500.0 86285.0 194155.0 ;
      RECT  85580.0 195500.0 86285.0 196845.0 ;
      RECT  85580.0 198190.0 86285.0 196845.0 ;
      RECT  85580.0 198190.0 86285.0 199535.0 ;
      RECT  85580.0 200880.0 86285.0 199535.0 ;
      RECT  85580.0 200880.0 86285.0 202225.0 ;
      RECT  85580.0 203570.0 86285.0 202225.0 ;
      RECT  85580.0 203570.0 86285.0 204915.0 ;
      RECT  85580.0 206260.0 86285.0 204915.0 ;
      RECT  86285.0 34100.0 86990.0 35445.0 ;
      RECT  86285.0 36790.0 86990.0 35445.0 ;
      RECT  86285.0 36790.0 86990.0 38135.0 ;
      RECT  86285.0 39480.0 86990.0 38135.0 ;
      RECT  86285.0 39480.0 86990.0 40825.0 ;
      RECT  86285.0 42170.0 86990.0 40825.0 ;
      RECT  86285.0 42170.0 86990.0 43515.0 ;
      RECT  86285.0 44860.0 86990.0 43515.0 ;
      RECT  86285.0 44860.0 86990.0 46205.0 ;
      RECT  86285.0 47550.0 86990.0 46205.0 ;
      RECT  86285.0 47550.0 86990.0 48895.0 ;
      RECT  86285.0 50240.0 86990.0 48895.0 ;
      RECT  86285.0 50240.0 86990.0 51585.0 ;
      RECT  86285.0 52930.0 86990.0 51585.0 ;
      RECT  86285.0 52930.0 86990.0 54275.0 ;
      RECT  86285.0 55620.0 86990.0 54275.0 ;
      RECT  86285.0 55620.0 86990.0 56965.0 ;
      RECT  86285.0 58310.0 86990.0 56965.0 ;
      RECT  86285.0 58310.0 86990.0 59655.0 ;
      RECT  86285.0 61000.0 86990.0 59655.0 ;
      RECT  86285.0 61000.0 86990.0 62345.0 ;
      RECT  86285.0 63690.0 86990.0 62345.0 ;
      RECT  86285.0 63690.0 86990.0 65035.0 ;
      RECT  86285.0 66380.0 86990.0 65035.0 ;
      RECT  86285.0 66380.0 86990.0 67725.0 ;
      RECT  86285.0 69070.0 86990.0 67725.0 ;
      RECT  86285.0 69070.0 86990.0 70415.0 ;
      RECT  86285.0 71760.0 86990.0 70415.0 ;
      RECT  86285.0 71760.0 86990.0 73105.0 ;
      RECT  86285.0 74450.0 86990.0 73105.0 ;
      RECT  86285.0 74450.0 86990.0 75795.0 ;
      RECT  86285.0 77140.0 86990.0 75795.0 ;
      RECT  86285.0 77140.0 86990.0 78485.0 ;
      RECT  86285.0 79830.0 86990.0 78485.0 ;
      RECT  86285.0 79830.0 86990.0 81175.0 ;
      RECT  86285.0 82520.0 86990.0 81175.0 ;
      RECT  86285.0 82520.0 86990.0 83865.0 ;
      RECT  86285.0 85210.0 86990.0 83865.0 ;
      RECT  86285.0 85210.0 86990.0 86555.0 ;
      RECT  86285.0 87900.0 86990.0 86555.0 ;
      RECT  86285.0 87900.0 86990.0 89245.0 ;
      RECT  86285.0 90590.0 86990.0 89245.0 ;
      RECT  86285.0 90590.0 86990.0 91935.0 ;
      RECT  86285.0 93280.0 86990.0 91935.0 ;
      RECT  86285.0 93280.0 86990.0 94625.0 ;
      RECT  86285.0 95970.0 86990.0 94625.0 ;
      RECT  86285.0 95970.0 86990.0 97315.0 ;
      RECT  86285.0 98660.0 86990.0 97315.0 ;
      RECT  86285.0 98660.0 86990.0 100005.0 ;
      RECT  86285.0 101350.0 86990.0 100005.0 ;
      RECT  86285.0 101350.0 86990.0 102695.0 ;
      RECT  86285.0 104040.0 86990.0 102695.0 ;
      RECT  86285.0 104040.0 86990.0 105385.0 ;
      RECT  86285.0 106730.0 86990.0 105385.0 ;
      RECT  86285.0 106730.0 86990.0 108075.0 ;
      RECT  86285.0 109420.0 86990.0 108075.0 ;
      RECT  86285.0 109420.0 86990.0 110765.0 ;
      RECT  86285.0 112110.0 86990.0 110765.0 ;
      RECT  86285.0 112110.0 86990.0 113455.0 ;
      RECT  86285.0 114800.0 86990.0 113455.0 ;
      RECT  86285.0 114800.0 86990.0 116145.0 ;
      RECT  86285.0 117490.0 86990.0 116145.0 ;
      RECT  86285.0 117490.0 86990.0 118835.0 ;
      RECT  86285.0 120180.0 86990.0 118835.0 ;
      RECT  86285.0 120180.0 86990.0 121525.0 ;
      RECT  86285.0 122870.0 86990.0 121525.0 ;
      RECT  86285.0 122870.0 86990.0 124215.0 ;
      RECT  86285.0 125560.0 86990.0 124215.0 ;
      RECT  86285.0 125560.0 86990.0 126905.0 ;
      RECT  86285.0 128250.0 86990.0 126905.0 ;
      RECT  86285.0 128250.0 86990.0 129595.0 ;
      RECT  86285.0 130940.0 86990.0 129595.0 ;
      RECT  86285.0 130940.0 86990.0 132285.0 ;
      RECT  86285.0 133630.0 86990.0 132285.0 ;
      RECT  86285.0 133630.0 86990.0 134975.0 ;
      RECT  86285.0 136320.0 86990.0 134975.0 ;
      RECT  86285.0 136320.0 86990.0 137665.0 ;
      RECT  86285.0 139010.0 86990.0 137665.0 ;
      RECT  86285.0 139010.0 86990.0 140355.0 ;
      RECT  86285.0 141700.0 86990.0 140355.0 ;
      RECT  86285.0 141700.0 86990.0 143045.0 ;
      RECT  86285.0 144390.0 86990.0 143045.0 ;
      RECT  86285.0 144390.0 86990.0 145735.0 ;
      RECT  86285.0 147080.0 86990.0 145735.0 ;
      RECT  86285.0 147080.0 86990.0 148425.0 ;
      RECT  86285.0 149770.0 86990.0 148425.0 ;
      RECT  86285.0 149770.0 86990.0 151115.0 ;
      RECT  86285.0 152460.0 86990.0 151115.0 ;
      RECT  86285.0 152460.0 86990.0 153805.0 ;
      RECT  86285.0 155150.0 86990.0 153805.0 ;
      RECT  86285.0 155150.0 86990.0 156495.0 ;
      RECT  86285.0 157840.0 86990.0 156495.0 ;
      RECT  86285.0 157840.0 86990.0 159185.0 ;
      RECT  86285.0 160530.0 86990.0 159185.0 ;
      RECT  86285.0 160530.0 86990.0 161875.0 ;
      RECT  86285.0 163220.0 86990.0 161875.0 ;
      RECT  86285.0 163220.0 86990.0 164565.0 ;
      RECT  86285.0 165910.0 86990.0 164565.0 ;
      RECT  86285.0 165910.0 86990.0 167255.0 ;
      RECT  86285.0 168600.0 86990.0 167255.0 ;
      RECT  86285.0 168600.0 86990.0 169945.0 ;
      RECT  86285.0 171290.0 86990.0 169945.0 ;
      RECT  86285.0 171290.0 86990.0 172635.0 ;
      RECT  86285.0 173980.0 86990.0 172635.0 ;
      RECT  86285.0 173980.0 86990.0 175325.0 ;
      RECT  86285.0 176670.0 86990.0 175325.0 ;
      RECT  86285.0 176670.0 86990.0 178015.0 ;
      RECT  86285.0 179360.0 86990.0 178015.0 ;
      RECT  86285.0 179360.0 86990.0 180705.0 ;
      RECT  86285.0 182050.0 86990.0 180705.0 ;
      RECT  86285.0 182050.0 86990.0 183395.0 ;
      RECT  86285.0 184740.0 86990.0 183395.0 ;
      RECT  86285.0 184740.0 86990.0 186085.0 ;
      RECT  86285.0 187430.0 86990.0 186085.0 ;
      RECT  86285.0 187430.0 86990.0 188775.0 ;
      RECT  86285.0 190120.0 86990.0 188775.0 ;
      RECT  86285.0 190120.0 86990.0 191465.0 ;
      RECT  86285.0 192810.0 86990.0 191465.0 ;
      RECT  86285.0 192810.0 86990.0 194155.0 ;
      RECT  86285.0 195500.0 86990.0 194155.0 ;
      RECT  86285.0 195500.0 86990.0 196845.0 ;
      RECT  86285.0 198190.0 86990.0 196845.0 ;
      RECT  86285.0 198190.0 86990.0 199535.0 ;
      RECT  86285.0 200880.0 86990.0 199535.0 ;
      RECT  86285.0 200880.0 86990.0 202225.0 ;
      RECT  86285.0 203570.0 86990.0 202225.0 ;
      RECT  86285.0 203570.0 86990.0 204915.0 ;
      RECT  86285.0 206260.0 86990.0 204915.0 ;
      RECT  86990.0 34100.0 87695.0 35445.0 ;
      RECT  86990.0 36790.0 87695.0 35445.0 ;
      RECT  86990.0 36790.0 87695.0 38135.0 ;
      RECT  86990.0 39480.0 87695.0 38135.0 ;
      RECT  86990.0 39480.0 87695.0 40825.0 ;
      RECT  86990.0 42170.0 87695.0 40825.0 ;
      RECT  86990.0 42170.0 87695.0 43515.0 ;
      RECT  86990.0 44860.0 87695.0 43515.0 ;
      RECT  86990.0 44860.0 87695.0 46205.0 ;
      RECT  86990.0 47550.0 87695.0 46205.0 ;
      RECT  86990.0 47550.0 87695.0 48895.0 ;
      RECT  86990.0 50240.0 87695.0 48895.0 ;
      RECT  86990.0 50240.0 87695.0 51585.0 ;
      RECT  86990.0 52930.0 87695.0 51585.0 ;
      RECT  86990.0 52930.0 87695.0 54275.0 ;
      RECT  86990.0 55620.0 87695.0 54275.0 ;
      RECT  86990.0 55620.0 87695.0 56965.0 ;
      RECT  86990.0 58310.0 87695.0 56965.0 ;
      RECT  86990.0 58310.0 87695.0 59655.0 ;
      RECT  86990.0 61000.0 87695.0 59655.0 ;
      RECT  86990.0 61000.0 87695.0 62345.0 ;
      RECT  86990.0 63690.0 87695.0 62345.0 ;
      RECT  86990.0 63690.0 87695.0 65035.0 ;
      RECT  86990.0 66380.0 87695.0 65035.0 ;
      RECT  86990.0 66380.0 87695.0 67725.0 ;
      RECT  86990.0 69070.0 87695.0 67725.0 ;
      RECT  86990.0 69070.0 87695.0 70415.0 ;
      RECT  86990.0 71760.0 87695.0 70415.0 ;
      RECT  86990.0 71760.0 87695.0 73105.0 ;
      RECT  86990.0 74450.0 87695.0 73105.0 ;
      RECT  86990.0 74450.0 87695.0 75795.0 ;
      RECT  86990.0 77140.0 87695.0 75795.0 ;
      RECT  86990.0 77140.0 87695.0 78485.0 ;
      RECT  86990.0 79830.0 87695.0 78485.0 ;
      RECT  86990.0 79830.0 87695.0 81175.0 ;
      RECT  86990.0 82520.0 87695.0 81175.0 ;
      RECT  86990.0 82520.0 87695.0 83865.0 ;
      RECT  86990.0 85210.0 87695.0 83865.0 ;
      RECT  86990.0 85210.0 87695.0 86555.0 ;
      RECT  86990.0 87900.0 87695.0 86555.0 ;
      RECT  86990.0 87900.0 87695.0 89245.0 ;
      RECT  86990.0 90590.0 87695.0 89245.0 ;
      RECT  86990.0 90590.0 87695.0 91935.0 ;
      RECT  86990.0 93280.0 87695.0 91935.0 ;
      RECT  86990.0 93280.0 87695.0 94625.0 ;
      RECT  86990.0 95970.0 87695.0 94625.0 ;
      RECT  86990.0 95970.0 87695.0 97315.0 ;
      RECT  86990.0 98660.0 87695.0 97315.0 ;
      RECT  86990.0 98660.0 87695.0 100005.0 ;
      RECT  86990.0 101350.0 87695.0 100005.0 ;
      RECT  86990.0 101350.0 87695.0 102695.0 ;
      RECT  86990.0 104040.0 87695.0 102695.0 ;
      RECT  86990.0 104040.0 87695.0 105385.0 ;
      RECT  86990.0 106730.0 87695.0 105385.0 ;
      RECT  86990.0 106730.0 87695.0 108075.0 ;
      RECT  86990.0 109420.0 87695.0 108075.0 ;
      RECT  86990.0 109420.0 87695.0 110765.0 ;
      RECT  86990.0 112110.0 87695.0 110765.0 ;
      RECT  86990.0 112110.0 87695.0 113455.0 ;
      RECT  86990.0 114800.0 87695.0 113455.0 ;
      RECT  86990.0 114800.0 87695.0 116145.0 ;
      RECT  86990.0 117490.0 87695.0 116145.0 ;
      RECT  86990.0 117490.0 87695.0 118835.0 ;
      RECT  86990.0 120180.0 87695.0 118835.0 ;
      RECT  86990.0 120180.0 87695.0 121525.0 ;
      RECT  86990.0 122870.0 87695.0 121525.0 ;
      RECT  86990.0 122870.0 87695.0 124215.0 ;
      RECT  86990.0 125560.0 87695.0 124215.0 ;
      RECT  86990.0 125560.0 87695.0 126905.0 ;
      RECT  86990.0 128250.0 87695.0 126905.0 ;
      RECT  86990.0 128250.0 87695.0 129595.0 ;
      RECT  86990.0 130940.0 87695.0 129595.0 ;
      RECT  86990.0 130940.0 87695.0 132285.0 ;
      RECT  86990.0 133630.0 87695.0 132285.0 ;
      RECT  86990.0 133630.0 87695.0 134975.0 ;
      RECT  86990.0 136320.0 87695.0 134975.0 ;
      RECT  86990.0 136320.0 87695.0 137665.0 ;
      RECT  86990.0 139010.0 87695.0 137665.0 ;
      RECT  86990.0 139010.0 87695.0 140355.0 ;
      RECT  86990.0 141700.0 87695.0 140355.0 ;
      RECT  86990.0 141700.0 87695.0 143045.0 ;
      RECT  86990.0 144390.0 87695.0 143045.0 ;
      RECT  86990.0 144390.0 87695.0 145735.0 ;
      RECT  86990.0 147080.0 87695.0 145735.0 ;
      RECT  86990.0 147080.0 87695.0 148425.0 ;
      RECT  86990.0 149770.0 87695.0 148425.0 ;
      RECT  86990.0 149770.0 87695.0 151115.0 ;
      RECT  86990.0 152460.0 87695.0 151115.0 ;
      RECT  86990.0 152460.0 87695.0 153805.0 ;
      RECT  86990.0 155150.0 87695.0 153805.0 ;
      RECT  86990.0 155150.0 87695.0 156495.0 ;
      RECT  86990.0 157840.0 87695.0 156495.0 ;
      RECT  86990.0 157840.0 87695.0 159185.0 ;
      RECT  86990.0 160530.0 87695.0 159185.0 ;
      RECT  86990.0 160530.0 87695.0 161875.0 ;
      RECT  86990.0 163220.0 87695.0 161875.0 ;
      RECT  86990.0 163220.0 87695.0 164565.0 ;
      RECT  86990.0 165910.0 87695.0 164565.0 ;
      RECT  86990.0 165910.0 87695.0 167255.0 ;
      RECT  86990.0 168600.0 87695.0 167255.0 ;
      RECT  86990.0 168600.0 87695.0 169945.0 ;
      RECT  86990.0 171290.0 87695.0 169945.0 ;
      RECT  86990.0 171290.0 87695.0 172635.0 ;
      RECT  86990.0 173980.0 87695.0 172635.0 ;
      RECT  86990.0 173980.0 87695.0 175325.0 ;
      RECT  86990.0 176670.0 87695.0 175325.0 ;
      RECT  86990.0 176670.0 87695.0 178015.0 ;
      RECT  86990.0 179360.0 87695.0 178015.0 ;
      RECT  86990.0 179360.0 87695.0 180705.0 ;
      RECT  86990.0 182050.0 87695.0 180705.0 ;
      RECT  86990.0 182050.0 87695.0 183395.0 ;
      RECT  86990.0 184740.0 87695.0 183395.0 ;
      RECT  86990.0 184740.0 87695.0 186085.0 ;
      RECT  86990.0 187430.0 87695.0 186085.0 ;
      RECT  86990.0 187430.0 87695.0 188775.0 ;
      RECT  86990.0 190120.0 87695.0 188775.0 ;
      RECT  86990.0 190120.0 87695.0 191465.0 ;
      RECT  86990.0 192810.0 87695.0 191465.0 ;
      RECT  86990.0 192810.0 87695.0 194155.0 ;
      RECT  86990.0 195500.0 87695.0 194155.0 ;
      RECT  86990.0 195500.0 87695.0 196845.0 ;
      RECT  86990.0 198190.0 87695.0 196845.0 ;
      RECT  86990.0 198190.0 87695.0 199535.0 ;
      RECT  86990.0 200880.0 87695.0 199535.0 ;
      RECT  86990.0 200880.0 87695.0 202225.0 ;
      RECT  86990.0 203570.0 87695.0 202225.0 ;
      RECT  86990.0 203570.0 87695.0 204915.0 ;
      RECT  86990.0 206260.0 87695.0 204915.0 ;
      RECT  87695.0 34100.0 88400.0 35445.0 ;
      RECT  87695.0 36790.0 88400.0 35445.0 ;
      RECT  87695.0 36790.0 88400.0 38135.0 ;
      RECT  87695.0 39480.0 88400.0 38135.0 ;
      RECT  87695.0 39480.0 88400.0 40825.0 ;
      RECT  87695.0 42170.0 88400.0 40825.0 ;
      RECT  87695.0 42170.0 88400.0 43515.0 ;
      RECT  87695.0 44860.0 88400.0 43515.0 ;
      RECT  87695.0 44860.0 88400.0 46205.0 ;
      RECT  87695.0 47550.0 88400.0 46205.0 ;
      RECT  87695.0 47550.0 88400.0 48895.0 ;
      RECT  87695.0 50240.0 88400.0 48895.0 ;
      RECT  87695.0 50240.0 88400.0 51585.0 ;
      RECT  87695.0 52930.0 88400.0 51585.0 ;
      RECT  87695.0 52930.0 88400.0 54275.0 ;
      RECT  87695.0 55620.0 88400.0 54275.0 ;
      RECT  87695.0 55620.0 88400.0 56965.0 ;
      RECT  87695.0 58310.0 88400.0 56965.0 ;
      RECT  87695.0 58310.0 88400.0 59655.0 ;
      RECT  87695.0 61000.0 88400.0 59655.0 ;
      RECT  87695.0 61000.0 88400.0 62345.0 ;
      RECT  87695.0 63690.0 88400.0 62345.0 ;
      RECT  87695.0 63690.0 88400.0 65035.0 ;
      RECT  87695.0 66380.0 88400.0 65035.0 ;
      RECT  87695.0 66380.0 88400.0 67725.0 ;
      RECT  87695.0 69070.0 88400.0 67725.0 ;
      RECT  87695.0 69070.0 88400.0 70415.0 ;
      RECT  87695.0 71760.0 88400.0 70415.0 ;
      RECT  87695.0 71760.0 88400.0 73105.0 ;
      RECT  87695.0 74450.0 88400.0 73105.0 ;
      RECT  87695.0 74450.0 88400.0 75795.0 ;
      RECT  87695.0 77140.0 88400.0 75795.0 ;
      RECT  87695.0 77140.0 88400.0 78485.0 ;
      RECT  87695.0 79830.0 88400.0 78485.0 ;
      RECT  87695.0 79830.0 88400.0 81175.0 ;
      RECT  87695.0 82520.0 88400.0 81175.0 ;
      RECT  87695.0 82520.0 88400.0 83865.0 ;
      RECT  87695.0 85210.0 88400.0 83865.0 ;
      RECT  87695.0 85210.0 88400.0 86555.0 ;
      RECT  87695.0 87900.0 88400.0 86555.0 ;
      RECT  87695.0 87900.0 88400.0 89245.0 ;
      RECT  87695.0 90590.0 88400.0 89245.0 ;
      RECT  87695.0 90590.0 88400.0 91935.0 ;
      RECT  87695.0 93280.0 88400.0 91935.0 ;
      RECT  87695.0 93280.0 88400.0 94625.0 ;
      RECT  87695.0 95970.0 88400.0 94625.0 ;
      RECT  87695.0 95970.0 88400.0 97315.0 ;
      RECT  87695.0 98660.0 88400.0 97315.0 ;
      RECT  87695.0 98660.0 88400.0 100005.0 ;
      RECT  87695.0 101350.0 88400.0 100005.0 ;
      RECT  87695.0 101350.0 88400.0 102695.0 ;
      RECT  87695.0 104040.0 88400.0 102695.0 ;
      RECT  87695.0 104040.0 88400.0 105385.0 ;
      RECT  87695.0 106730.0 88400.0 105385.0 ;
      RECT  87695.0 106730.0 88400.0 108075.0 ;
      RECT  87695.0 109420.0 88400.0 108075.0 ;
      RECT  87695.0 109420.0 88400.0 110765.0 ;
      RECT  87695.0 112110.0 88400.0 110765.0 ;
      RECT  87695.0 112110.0 88400.0 113455.0 ;
      RECT  87695.0 114800.0 88400.0 113455.0 ;
      RECT  87695.0 114800.0 88400.0 116145.0 ;
      RECT  87695.0 117490.0 88400.0 116145.0 ;
      RECT  87695.0 117490.0 88400.0 118835.0 ;
      RECT  87695.0 120180.0 88400.0 118835.0 ;
      RECT  87695.0 120180.0 88400.0 121525.0 ;
      RECT  87695.0 122870.0 88400.0 121525.0 ;
      RECT  87695.0 122870.0 88400.0 124215.0 ;
      RECT  87695.0 125560.0 88400.0 124215.0 ;
      RECT  87695.0 125560.0 88400.0 126905.0 ;
      RECT  87695.0 128250.0 88400.0 126905.0 ;
      RECT  87695.0 128250.0 88400.0 129595.0 ;
      RECT  87695.0 130940.0 88400.0 129595.0 ;
      RECT  87695.0 130940.0 88400.0 132285.0 ;
      RECT  87695.0 133630.0 88400.0 132285.0 ;
      RECT  87695.0 133630.0 88400.0 134975.0 ;
      RECT  87695.0 136320.0 88400.0 134975.0 ;
      RECT  87695.0 136320.0 88400.0 137665.0 ;
      RECT  87695.0 139010.0 88400.0 137665.0 ;
      RECT  87695.0 139010.0 88400.0 140355.0 ;
      RECT  87695.0 141700.0 88400.0 140355.0 ;
      RECT  87695.0 141700.0 88400.0 143045.0 ;
      RECT  87695.0 144390.0 88400.0 143045.0 ;
      RECT  87695.0 144390.0 88400.0 145735.0 ;
      RECT  87695.0 147080.0 88400.0 145735.0 ;
      RECT  87695.0 147080.0 88400.0 148425.0 ;
      RECT  87695.0 149770.0 88400.0 148425.0 ;
      RECT  87695.0 149770.0 88400.0 151115.0 ;
      RECT  87695.0 152460.0 88400.0 151115.0 ;
      RECT  87695.0 152460.0 88400.0 153805.0 ;
      RECT  87695.0 155150.0 88400.0 153805.0 ;
      RECT  87695.0 155150.0 88400.0 156495.0 ;
      RECT  87695.0 157840.0 88400.0 156495.0 ;
      RECT  87695.0 157840.0 88400.0 159185.0 ;
      RECT  87695.0 160530.0 88400.0 159185.0 ;
      RECT  87695.0 160530.0 88400.0 161875.0 ;
      RECT  87695.0 163220.0 88400.0 161875.0 ;
      RECT  87695.0 163220.0 88400.0 164565.0 ;
      RECT  87695.0 165910.0 88400.0 164565.0 ;
      RECT  87695.0 165910.0 88400.0 167255.0 ;
      RECT  87695.0 168600.0 88400.0 167255.0 ;
      RECT  87695.0 168600.0 88400.0 169945.0 ;
      RECT  87695.0 171290.0 88400.0 169945.0 ;
      RECT  87695.0 171290.0 88400.0 172635.0 ;
      RECT  87695.0 173980.0 88400.0 172635.0 ;
      RECT  87695.0 173980.0 88400.0 175325.0 ;
      RECT  87695.0 176670.0 88400.0 175325.0 ;
      RECT  87695.0 176670.0 88400.0 178015.0 ;
      RECT  87695.0 179360.0 88400.0 178015.0 ;
      RECT  87695.0 179360.0 88400.0 180705.0 ;
      RECT  87695.0 182050.0 88400.0 180705.0 ;
      RECT  87695.0 182050.0 88400.0 183395.0 ;
      RECT  87695.0 184740.0 88400.0 183395.0 ;
      RECT  87695.0 184740.0 88400.0 186085.0 ;
      RECT  87695.0 187430.0 88400.0 186085.0 ;
      RECT  87695.0 187430.0 88400.0 188775.0 ;
      RECT  87695.0 190120.0 88400.0 188775.0 ;
      RECT  87695.0 190120.0 88400.0 191465.0 ;
      RECT  87695.0 192810.0 88400.0 191465.0 ;
      RECT  87695.0 192810.0 88400.0 194155.0 ;
      RECT  87695.0 195500.0 88400.0 194155.0 ;
      RECT  87695.0 195500.0 88400.0 196845.0 ;
      RECT  87695.0 198190.0 88400.0 196845.0 ;
      RECT  87695.0 198190.0 88400.0 199535.0 ;
      RECT  87695.0 200880.0 88400.0 199535.0 ;
      RECT  87695.0 200880.0 88400.0 202225.0 ;
      RECT  87695.0 203570.0 88400.0 202225.0 ;
      RECT  87695.0 203570.0 88400.0 204915.0 ;
      RECT  87695.0 206260.0 88400.0 204915.0 ;
      RECT  88400.0 34100.0 89105.0 35445.0 ;
      RECT  88400.0 36790.0 89105.0 35445.0 ;
      RECT  88400.0 36790.0 89105.0 38135.0 ;
      RECT  88400.0 39480.0 89105.0 38135.0 ;
      RECT  88400.0 39480.0 89105.0 40825.0 ;
      RECT  88400.0 42170.0 89105.0 40825.0 ;
      RECT  88400.0 42170.0 89105.0 43515.0 ;
      RECT  88400.0 44860.0 89105.0 43515.0 ;
      RECT  88400.0 44860.0 89105.0 46205.0 ;
      RECT  88400.0 47550.0 89105.0 46205.0 ;
      RECT  88400.0 47550.0 89105.0 48895.0 ;
      RECT  88400.0 50240.0 89105.0 48895.0 ;
      RECT  88400.0 50240.0 89105.0 51585.0 ;
      RECT  88400.0 52930.0 89105.0 51585.0 ;
      RECT  88400.0 52930.0 89105.0 54275.0 ;
      RECT  88400.0 55620.0 89105.0 54275.0 ;
      RECT  88400.0 55620.0 89105.0 56965.0 ;
      RECT  88400.0 58310.0 89105.0 56965.0 ;
      RECT  88400.0 58310.0 89105.0 59655.0 ;
      RECT  88400.0 61000.0 89105.0 59655.0 ;
      RECT  88400.0 61000.0 89105.0 62345.0 ;
      RECT  88400.0 63690.0 89105.0 62345.0 ;
      RECT  88400.0 63690.0 89105.0 65035.0 ;
      RECT  88400.0 66380.0 89105.0 65035.0 ;
      RECT  88400.0 66380.0 89105.0 67725.0 ;
      RECT  88400.0 69070.0 89105.0 67725.0 ;
      RECT  88400.0 69070.0 89105.0 70415.0 ;
      RECT  88400.0 71760.0 89105.0 70415.0 ;
      RECT  88400.0 71760.0 89105.0 73105.0 ;
      RECT  88400.0 74450.0 89105.0 73105.0 ;
      RECT  88400.0 74450.0 89105.0 75795.0 ;
      RECT  88400.0 77140.0 89105.0 75795.0 ;
      RECT  88400.0 77140.0 89105.0 78485.0 ;
      RECT  88400.0 79830.0 89105.0 78485.0 ;
      RECT  88400.0 79830.0 89105.0 81175.0 ;
      RECT  88400.0 82520.0 89105.0 81175.0 ;
      RECT  88400.0 82520.0 89105.0 83865.0 ;
      RECT  88400.0 85210.0 89105.0 83865.0 ;
      RECT  88400.0 85210.0 89105.0 86555.0 ;
      RECT  88400.0 87900.0 89105.0 86555.0 ;
      RECT  88400.0 87900.0 89105.0 89245.0 ;
      RECT  88400.0 90590.0 89105.0 89245.0 ;
      RECT  88400.0 90590.0 89105.0 91935.0 ;
      RECT  88400.0 93280.0 89105.0 91935.0 ;
      RECT  88400.0 93280.0 89105.0 94625.0 ;
      RECT  88400.0 95970.0 89105.0 94625.0 ;
      RECT  88400.0 95970.0 89105.0 97315.0 ;
      RECT  88400.0 98660.0 89105.0 97315.0 ;
      RECT  88400.0 98660.0 89105.0 100005.0 ;
      RECT  88400.0 101350.0 89105.0 100005.0 ;
      RECT  88400.0 101350.0 89105.0 102695.0 ;
      RECT  88400.0 104040.0 89105.0 102695.0 ;
      RECT  88400.0 104040.0 89105.0 105385.0 ;
      RECT  88400.0 106730.0 89105.0 105385.0 ;
      RECT  88400.0 106730.0 89105.0 108075.0 ;
      RECT  88400.0 109420.0 89105.0 108075.0 ;
      RECT  88400.0 109420.0 89105.0 110765.0 ;
      RECT  88400.0 112110.0 89105.0 110765.0 ;
      RECT  88400.0 112110.0 89105.0 113455.0 ;
      RECT  88400.0 114800.0 89105.0 113455.0 ;
      RECT  88400.0 114800.0 89105.0 116145.0 ;
      RECT  88400.0 117490.0 89105.0 116145.0 ;
      RECT  88400.0 117490.0 89105.0 118835.0 ;
      RECT  88400.0 120180.0 89105.0 118835.0 ;
      RECT  88400.0 120180.0 89105.0 121525.0 ;
      RECT  88400.0 122870.0 89105.0 121525.0 ;
      RECT  88400.0 122870.0 89105.0 124215.0 ;
      RECT  88400.0 125560.0 89105.0 124215.0 ;
      RECT  88400.0 125560.0 89105.0 126905.0 ;
      RECT  88400.0 128250.0 89105.0 126905.0 ;
      RECT  88400.0 128250.0 89105.0 129595.0 ;
      RECT  88400.0 130940.0 89105.0 129595.0 ;
      RECT  88400.0 130940.0 89105.0 132285.0 ;
      RECT  88400.0 133630.0 89105.0 132285.0 ;
      RECT  88400.0 133630.0 89105.0 134975.0 ;
      RECT  88400.0 136320.0 89105.0 134975.0 ;
      RECT  88400.0 136320.0 89105.0 137665.0 ;
      RECT  88400.0 139010.0 89105.0 137665.0 ;
      RECT  88400.0 139010.0 89105.0 140355.0 ;
      RECT  88400.0 141700.0 89105.0 140355.0 ;
      RECT  88400.0 141700.0 89105.0 143045.0 ;
      RECT  88400.0 144390.0 89105.0 143045.0 ;
      RECT  88400.0 144390.0 89105.0 145735.0 ;
      RECT  88400.0 147080.0 89105.0 145735.0 ;
      RECT  88400.0 147080.0 89105.0 148425.0 ;
      RECT  88400.0 149770.0 89105.0 148425.0 ;
      RECT  88400.0 149770.0 89105.0 151115.0 ;
      RECT  88400.0 152460.0 89105.0 151115.0 ;
      RECT  88400.0 152460.0 89105.0 153805.0 ;
      RECT  88400.0 155150.0 89105.0 153805.0 ;
      RECT  88400.0 155150.0 89105.0 156495.0 ;
      RECT  88400.0 157840.0 89105.0 156495.0 ;
      RECT  88400.0 157840.0 89105.0 159185.0 ;
      RECT  88400.0 160530.0 89105.0 159185.0 ;
      RECT  88400.0 160530.0 89105.0 161875.0 ;
      RECT  88400.0 163220.0 89105.0 161875.0 ;
      RECT  88400.0 163220.0 89105.0 164565.0 ;
      RECT  88400.0 165910.0 89105.0 164565.0 ;
      RECT  88400.0 165910.0 89105.0 167255.0 ;
      RECT  88400.0 168600.0 89105.0 167255.0 ;
      RECT  88400.0 168600.0 89105.0 169945.0 ;
      RECT  88400.0 171290.0 89105.0 169945.0 ;
      RECT  88400.0 171290.0 89105.0 172635.0 ;
      RECT  88400.0 173980.0 89105.0 172635.0 ;
      RECT  88400.0 173980.0 89105.0 175325.0 ;
      RECT  88400.0 176670.0 89105.0 175325.0 ;
      RECT  88400.0 176670.0 89105.0 178015.0 ;
      RECT  88400.0 179360.0 89105.0 178015.0 ;
      RECT  88400.0 179360.0 89105.0 180705.0 ;
      RECT  88400.0 182050.0 89105.0 180705.0 ;
      RECT  88400.0 182050.0 89105.0 183395.0 ;
      RECT  88400.0 184740.0 89105.0 183395.0 ;
      RECT  88400.0 184740.0 89105.0 186085.0 ;
      RECT  88400.0 187430.0 89105.0 186085.0 ;
      RECT  88400.0 187430.0 89105.0 188775.0 ;
      RECT  88400.0 190120.0 89105.0 188775.0 ;
      RECT  88400.0 190120.0 89105.0 191465.0 ;
      RECT  88400.0 192810.0 89105.0 191465.0 ;
      RECT  88400.0 192810.0 89105.0 194155.0 ;
      RECT  88400.0 195500.0 89105.0 194155.0 ;
      RECT  88400.0 195500.0 89105.0 196845.0 ;
      RECT  88400.0 198190.0 89105.0 196845.0 ;
      RECT  88400.0 198190.0 89105.0 199535.0 ;
      RECT  88400.0 200880.0 89105.0 199535.0 ;
      RECT  88400.0 200880.0 89105.0 202225.0 ;
      RECT  88400.0 203570.0 89105.0 202225.0 ;
      RECT  88400.0 203570.0 89105.0 204915.0 ;
      RECT  88400.0 206260.0 89105.0 204915.0 ;
      RECT  89105.0 34100.0 89810.0 35445.0 ;
      RECT  89105.0 36790.0 89810.0 35445.0 ;
      RECT  89105.0 36790.0 89810.0 38135.0 ;
      RECT  89105.0 39480.0 89810.0 38135.0 ;
      RECT  89105.0 39480.0 89810.0 40825.0 ;
      RECT  89105.0 42170.0 89810.0 40825.0 ;
      RECT  89105.0 42170.0 89810.0 43515.0 ;
      RECT  89105.0 44860.0 89810.0 43515.0 ;
      RECT  89105.0 44860.0 89810.0 46205.0 ;
      RECT  89105.0 47550.0 89810.0 46205.0 ;
      RECT  89105.0 47550.0 89810.0 48895.0 ;
      RECT  89105.0 50240.0 89810.0 48895.0 ;
      RECT  89105.0 50240.0 89810.0 51585.0 ;
      RECT  89105.0 52930.0 89810.0 51585.0 ;
      RECT  89105.0 52930.0 89810.0 54275.0 ;
      RECT  89105.0 55620.0 89810.0 54275.0 ;
      RECT  89105.0 55620.0 89810.0 56965.0 ;
      RECT  89105.0 58310.0 89810.0 56965.0 ;
      RECT  89105.0 58310.0 89810.0 59655.0 ;
      RECT  89105.0 61000.0 89810.0 59655.0 ;
      RECT  89105.0 61000.0 89810.0 62345.0 ;
      RECT  89105.0 63690.0 89810.0 62345.0 ;
      RECT  89105.0 63690.0 89810.0 65035.0 ;
      RECT  89105.0 66380.0 89810.0 65035.0 ;
      RECT  89105.0 66380.0 89810.0 67725.0 ;
      RECT  89105.0 69070.0 89810.0 67725.0 ;
      RECT  89105.0 69070.0 89810.0 70415.0 ;
      RECT  89105.0 71760.0 89810.0 70415.0 ;
      RECT  89105.0 71760.0 89810.0 73105.0 ;
      RECT  89105.0 74450.0 89810.0 73105.0 ;
      RECT  89105.0 74450.0 89810.0 75795.0 ;
      RECT  89105.0 77140.0 89810.0 75795.0 ;
      RECT  89105.0 77140.0 89810.0 78485.0 ;
      RECT  89105.0 79830.0 89810.0 78485.0 ;
      RECT  89105.0 79830.0 89810.0 81175.0 ;
      RECT  89105.0 82520.0 89810.0 81175.0 ;
      RECT  89105.0 82520.0 89810.0 83865.0 ;
      RECT  89105.0 85210.0 89810.0 83865.0 ;
      RECT  89105.0 85210.0 89810.0 86555.0 ;
      RECT  89105.0 87900.0 89810.0 86555.0 ;
      RECT  89105.0 87900.0 89810.0 89245.0 ;
      RECT  89105.0 90590.0 89810.0 89245.0 ;
      RECT  89105.0 90590.0 89810.0 91935.0 ;
      RECT  89105.0 93280.0 89810.0 91935.0 ;
      RECT  89105.0 93280.0 89810.0 94625.0 ;
      RECT  89105.0 95970.0 89810.0 94625.0 ;
      RECT  89105.0 95970.0 89810.0 97315.0 ;
      RECT  89105.0 98660.0 89810.0 97315.0 ;
      RECT  89105.0 98660.0 89810.0 100005.0 ;
      RECT  89105.0 101350.0 89810.0 100005.0 ;
      RECT  89105.0 101350.0 89810.0 102695.0 ;
      RECT  89105.0 104040.0 89810.0 102695.0 ;
      RECT  89105.0 104040.0 89810.0 105385.0 ;
      RECT  89105.0 106730.0 89810.0 105385.0 ;
      RECT  89105.0 106730.0 89810.0 108075.0 ;
      RECT  89105.0 109420.0 89810.0 108075.0 ;
      RECT  89105.0 109420.0 89810.0 110765.0 ;
      RECT  89105.0 112110.0 89810.0 110765.0 ;
      RECT  89105.0 112110.0 89810.0 113455.0 ;
      RECT  89105.0 114800.0 89810.0 113455.0 ;
      RECT  89105.0 114800.0 89810.0 116145.0 ;
      RECT  89105.0 117490.0 89810.0 116145.0 ;
      RECT  89105.0 117490.0 89810.0 118835.0 ;
      RECT  89105.0 120180.0 89810.0 118835.0 ;
      RECT  89105.0 120180.0 89810.0 121525.0 ;
      RECT  89105.0 122870.0 89810.0 121525.0 ;
      RECT  89105.0 122870.0 89810.0 124215.0 ;
      RECT  89105.0 125560.0 89810.0 124215.0 ;
      RECT  89105.0 125560.0 89810.0 126905.0 ;
      RECT  89105.0 128250.0 89810.0 126905.0 ;
      RECT  89105.0 128250.0 89810.0 129595.0 ;
      RECT  89105.0 130940.0 89810.0 129595.0 ;
      RECT  89105.0 130940.0 89810.0 132285.0 ;
      RECT  89105.0 133630.0 89810.0 132285.0 ;
      RECT  89105.0 133630.0 89810.0 134975.0 ;
      RECT  89105.0 136320.0 89810.0 134975.0 ;
      RECT  89105.0 136320.0 89810.0 137665.0 ;
      RECT  89105.0 139010.0 89810.0 137665.0 ;
      RECT  89105.0 139010.0 89810.0 140355.0 ;
      RECT  89105.0 141700.0 89810.0 140355.0 ;
      RECT  89105.0 141700.0 89810.0 143045.0 ;
      RECT  89105.0 144390.0 89810.0 143045.0 ;
      RECT  89105.0 144390.0 89810.0 145735.0 ;
      RECT  89105.0 147080.0 89810.0 145735.0 ;
      RECT  89105.0 147080.0 89810.0 148425.0 ;
      RECT  89105.0 149770.0 89810.0 148425.0 ;
      RECT  89105.0 149770.0 89810.0 151115.0 ;
      RECT  89105.0 152460.0 89810.0 151115.0 ;
      RECT  89105.0 152460.0 89810.0 153805.0 ;
      RECT  89105.0 155150.0 89810.0 153805.0 ;
      RECT  89105.0 155150.0 89810.0 156495.0 ;
      RECT  89105.0 157840.0 89810.0 156495.0 ;
      RECT  89105.0 157840.0 89810.0 159185.0 ;
      RECT  89105.0 160530.0 89810.0 159185.0 ;
      RECT  89105.0 160530.0 89810.0 161875.0 ;
      RECT  89105.0 163220.0 89810.0 161875.0 ;
      RECT  89105.0 163220.0 89810.0 164565.0 ;
      RECT  89105.0 165910.0 89810.0 164565.0 ;
      RECT  89105.0 165910.0 89810.0 167255.0 ;
      RECT  89105.0 168600.0 89810.0 167255.0 ;
      RECT  89105.0 168600.0 89810.0 169945.0 ;
      RECT  89105.0 171290.0 89810.0 169945.0 ;
      RECT  89105.0 171290.0 89810.0 172635.0 ;
      RECT  89105.0 173980.0 89810.0 172635.0 ;
      RECT  89105.0 173980.0 89810.0 175325.0 ;
      RECT  89105.0 176670.0 89810.0 175325.0 ;
      RECT  89105.0 176670.0 89810.0 178015.0 ;
      RECT  89105.0 179360.0 89810.0 178015.0 ;
      RECT  89105.0 179360.0 89810.0 180705.0 ;
      RECT  89105.0 182050.0 89810.0 180705.0 ;
      RECT  89105.0 182050.0 89810.0 183395.0 ;
      RECT  89105.0 184740.0 89810.0 183395.0 ;
      RECT  89105.0 184740.0 89810.0 186085.0 ;
      RECT  89105.0 187430.0 89810.0 186085.0 ;
      RECT  89105.0 187430.0 89810.0 188775.0 ;
      RECT  89105.0 190120.0 89810.0 188775.0 ;
      RECT  89105.0 190120.0 89810.0 191465.0 ;
      RECT  89105.0 192810.0 89810.0 191465.0 ;
      RECT  89105.0 192810.0 89810.0 194155.0 ;
      RECT  89105.0 195500.0 89810.0 194155.0 ;
      RECT  89105.0 195500.0 89810.0 196845.0 ;
      RECT  89105.0 198190.0 89810.0 196845.0 ;
      RECT  89105.0 198190.0 89810.0 199535.0 ;
      RECT  89105.0 200880.0 89810.0 199535.0 ;
      RECT  89105.0 200880.0 89810.0 202225.0 ;
      RECT  89105.0 203570.0 89810.0 202225.0 ;
      RECT  89105.0 203570.0 89810.0 204915.0 ;
      RECT  89105.0 206260.0 89810.0 204915.0 ;
      RECT  89810.0 34100.0 90515.0 35445.0 ;
      RECT  89810.0 36790.0 90515.0 35445.0 ;
      RECT  89810.0 36790.0 90515.0 38135.0 ;
      RECT  89810.0 39480.0 90515.0 38135.0 ;
      RECT  89810.0 39480.0 90515.0 40825.0 ;
      RECT  89810.0 42170.0 90515.0 40825.0 ;
      RECT  89810.0 42170.0 90515.0 43515.0 ;
      RECT  89810.0 44860.0 90515.0 43515.0 ;
      RECT  89810.0 44860.0 90515.0 46205.0 ;
      RECT  89810.0 47550.0 90515.0 46205.0 ;
      RECT  89810.0 47550.0 90515.0 48895.0 ;
      RECT  89810.0 50240.0 90515.0 48895.0 ;
      RECT  89810.0 50240.0 90515.0 51585.0 ;
      RECT  89810.0 52930.0 90515.0 51585.0 ;
      RECT  89810.0 52930.0 90515.0 54275.0 ;
      RECT  89810.0 55620.0 90515.0 54275.0 ;
      RECT  89810.0 55620.0 90515.0 56965.0 ;
      RECT  89810.0 58310.0 90515.0 56965.0 ;
      RECT  89810.0 58310.0 90515.0 59655.0 ;
      RECT  89810.0 61000.0 90515.0 59655.0 ;
      RECT  89810.0 61000.0 90515.0 62345.0 ;
      RECT  89810.0 63690.0 90515.0 62345.0 ;
      RECT  89810.0 63690.0 90515.0 65035.0 ;
      RECT  89810.0 66380.0 90515.0 65035.0 ;
      RECT  89810.0 66380.0 90515.0 67725.0 ;
      RECT  89810.0 69070.0 90515.0 67725.0 ;
      RECT  89810.0 69070.0 90515.0 70415.0 ;
      RECT  89810.0 71760.0 90515.0 70415.0 ;
      RECT  89810.0 71760.0 90515.0 73105.0 ;
      RECT  89810.0 74450.0 90515.0 73105.0 ;
      RECT  89810.0 74450.0 90515.0 75795.0 ;
      RECT  89810.0 77140.0 90515.0 75795.0 ;
      RECT  89810.0 77140.0 90515.0 78485.0 ;
      RECT  89810.0 79830.0 90515.0 78485.0 ;
      RECT  89810.0 79830.0 90515.0 81175.0 ;
      RECT  89810.0 82520.0 90515.0 81175.0 ;
      RECT  89810.0 82520.0 90515.0 83865.0 ;
      RECT  89810.0 85210.0 90515.0 83865.0 ;
      RECT  89810.0 85210.0 90515.0 86555.0 ;
      RECT  89810.0 87900.0 90515.0 86555.0 ;
      RECT  89810.0 87900.0 90515.0 89245.0 ;
      RECT  89810.0 90590.0 90515.0 89245.0 ;
      RECT  89810.0 90590.0 90515.0 91935.0 ;
      RECT  89810.0 93280.0 90515.0 91935.0 ;
      RECT  89810.0 93280.0 90515.0 94625.0 ;
      RECT  89810.0 95970.0 90515.0 94625.0 ;
      RECT  89810.0 95970.0 90515.0 97315.0 ;
      RECT  89810.0 98660.0 90515.0 97315.0 ;
      RECT  89810.0 98660.0 90515.0 100005.0 ;
      RECT  89810.0 101350.0 90515.0 100005.0 ;
      RECT  89810.0 101350.0 90515.0 102695.0 ;
      RECT  89810.0 104040.0 90515.0 102695.0 ;
      RECT  89810.0 104040.0 90515.0 105385.0 ;
      RECT  89810.0 106730.0 90515.0 105385.0 ;
      RECT  89810.0 106730.0 90515.0 108075.0 ;
      RECT  89810.0 109420.0 90515.0 108075.0 ;
      RECT  89810.0 109420.0 90515.0 110765.0 ;
      RECT  89810.0 112110.0 90515.0 110765.0 ;
      RECT  89810.0 112110.0 90515.0 113455.0 ;
      RECT  89810.0 114800.0 90515.0 113455.0 ;
      RECT  89810.0 114800.0 90515.0 116145.0 ;
      RECT  89810.0 117490.0 90515.0 116145.0 ;
      RECT  89810.0 117490.0 90515.0 118835.0 ;
      RECT  89810.0 120180.0 90515.0 118835.0 ;
      RECT  89810.0 120180.0 90515.0 121525.0 ;
      RECT  89810.0 122870.0 90515.0 121525.0 ;
      RECT  89810.0 122870.0 90515.0 124215.0 ;
      RECT  89810.0 125560.0 90515.0 124215.0 ;
      RECT  89810.0 125560.0 90515.0 126905.0 ;
      RECT  89810.0 128250.0 90515.0 126905.0 ;
      RECT  89810.0 128250.0 90515.0 129595.0 ;
      RECT  89810.0 130940.0 90515.0 129595.0 ;
      RECT  89810.0 130940.0 90515.0 132285.0 ;
      RECT  89810.0 133630.0 90515.0 132285.0 ;
      RECT  89810.0 133630.0 90515.0 134975.0 ;
      RECT  89810.0 136320.0 90515.0 134975.0 ;
      RECT  89810.0 136320.0 90515.0 137665.0 ;
      RECT  89810.0 139010.0 90515.0 137665.0 ;
      RECT  89810.0 139010.0 90515.0 140355.0 ;
      RECT  89810.0 141700.0 90515.0 140355.0 ;
      RECT  89810.0 141700.0 90515.0 143045.0 ;
      RECT  89810.0 144390.0 90515.0 143045.0 ;
      RECT  89810.0 144390.0 90515.0 145735.0 ;
      RECT  89810.0 147080.0 90515.0 145735.0 ;
      RECT  89810.0 147080.0 90515.0 148425.0 ;
      RECT  89810.0 149770.0 90515.0 148425.0 ;
      RECT  89810.0 149770.0 90515.0 151115.0 ;
      RECT  89810.0 152460.0 90515.0 151115.0 ;
      RECT  89810.0 152460.0 90515.0 153805.0 ;
      RECT  89810.0 155150.0 90515.0 153805.0 ;
      RECT  89810.0 155150.0 90515.0 156495.0 ;
      RECT  89810.0 157840.0 90515.0 156495.0 ;
      RECT  89810.0 157840.0 90515.0 159185.0 ;
      RECT  89810.0 160530.0 90515.0 159185.0 ;
      RECT  89810.0 160530.0 90515.0 161875.0 ;
      RECT  89810.0 163220.0 90515.0 161875.0 ;
      RECT  89810.0 163220.0 90515.0 164565.0 ;
      RECT  89810.0 165910.0 90515.0 164565.0 ;
      RECT  89810.0 165910.0 90515.0 167255.0 ;
      RECT  89810.0 168600.0 90515.0 167255.0 ;
      RECT  89810.0 168600.0 90515.0 169945.0 ;
      RECT  89810.0 171290.0 90515.0 169945.0 ;
      RECT  89810.0 171290.0 90515.0 172635.0 ;
      RECT  89810.0 173980.0 90515.0 172635.0 ;
      RECT  89810.0 173980.0 90515.0 175325.0 ;
      RECT  89810.0 176670.0 90515.0 175325.0 ;
      RECT  89810.0 176670.0 90515.0 178015.0 ;
      RECT  89810.0 179360.0 90515.0 178015.0 ;
      RECT  89810.0 179360.0 90515.0 180705.0 ;
      RECT  89810.0 182050.0 90515.0 180705.0 ;
      RECT  89810.0 182050.0 90515.0 183395.0 ;
      RECT  89810.0 184740.0 90515.0 183395.0 ;
      RECT  89810.0 184740.0 90515.0 186085.0 ;
      RECT  89810.0 187430.0 90515.0 186085.0 ;
      RECT  89810.0 187430.0 90515.0 188775.0 ;
      RECT  89810.0 190120.0 90515.0 188775.0 ;
      RECT  89810.0 190120.0 90515.0 191465.0 ;
      RECT  89810.0 192810.0 90515.0 191465.0 ;
      RECT  89810.0 192810.0 90515.0 194155.0 ;
      RECT  89810.0 195500.0 90515.0 194155.0 ;
      RECT  89810.0 195500.0 90515.0 196845.0 ;
      RECT  89810.0 198190.0 90515.0 196845.0 ;
      RECT  89810.0 198190.0 90515.0 199535.0 ;
      RECT  89810.0 200880.0 90515.0 199535.0 ;
      RECT  89810.0 200880.0 90515.0 202225.0 ;
      RECT  89810.0 203570.0 90515.0 202225.0 ;
      RECT  89810.0 203570.0 90515.0 204915.0 ;
      RECT  89810.0 206260.0 90515.0 204915.0 ;
      RECT  90515.0 34100.0 91220.0 35445.0 ;
      RECT  90515.0 36790.0 91220.0 35445.0 ;
      RECT  90515.0 36790.0 91220.0 38135.0 ;
      RECT  90515.0 39480.0 91220.0 38135.0 ;
      RECT  90515.0 39480.0 91220.0 40825.0 ;
      RECT  90515.0 42170.0 91220.0 40825.0 ;
      RECT  90515.0 42170.0 91220.0 43515.0 ;
      RECT  90515.0 44860.0 91220.0 43515.0 ;
      RECT  90515.0 44860.0 91220.0 46205.0 ;
      RECT  90515.0 47550.0 91220.0 46205.0 ;
      RECT  90515.0 47550.0 91220.0 48895.0 ;
      RECT  90515.0 50240.0 91220.0 48895.0 ;
      RECT  90515.0 50240.0 91220.0 51585.0 ;
      RECT  90515.0 52930.0 91220.0 51585.0 ;
      RECT  90515.0 52930.0 91220.0 54275.0 ;
      RECT  90515.0 55620.0 91220.0 54275.0 ;
      RECT  90515.0 55620.0 91220.0 56965.0 ;
      RECT  90515.0 58310.0 91220.0 56965.0 ;
      RECT  90515.0 58310.0 91220.0 59655.0 ;
      RECT  90515.0 61000.0 91220.0 59655.0 ;
      RECT  90515.0 61000.0 91220.0 62345.0 ;
      RECT  90515.0 63690.0 91220.0 62345.0 ;
      RECT  90515.0 63690.0 91220.0 65035.0 ;
      RECT  90515.0 66380.0 91220.0 65035.0 ;
      RECT  90515.0 66380.0 91220.0 67725.0 ;
      RECT  90515.0 69070.0 91220.0 67725.0 ;
      RECT  90515.0 69070.0 91220.0 70415.0 ;
      RECT  90515.0 71760.0 91220.0 70415.0 ;
      RECT  90515.0 71760.0 91220.0 73105.0 ;
      RECT  90515.0 74450.0 91220.0 73105.0 ;
      RECT  90515.0 74450.0 91220.0 75795.0 ;
      RECT  90515.0 77140.0 91220.0 75795.0 ;
      RECT  90515.0 77140.0 91220.0 78485.0 ;
      RECT  90515.0 79830.0 91220.0 78485.0 ;
      RECT  90515.0 79830.0 91220.0 81175.0 ;
      RECT  90515.0 82520.0 91220.0 81175.0 ;
      RECT  90515.0 82520.0 91220.0 83865.0 ;
      RECT  90515.0 85210.0 91220.0 83865.0 ;
      RECT  90515.0 85210.0 91220.0 86555.0 ;
      RECT  90515.0 87900.0 91220.0 86555.0 ;
      RECT  90515.0 87900.0 91220.0 89245.0 ;
      RECT  90515.0 90590.0 91220.0 89245.0 ;
      RECT  90515.0 90590.0 91220.0 91935.0 ;
      RECT  90515.0 93280.0 91220.0 91935.0 ;
      RECT  90515.0 93280.0 91220.0 94625.0 ;
      RECT  90515.0 95970.0 91220.0 94625.0 ;
      RECT  90515.0 95970.0 91220.0 97315.0 ;
      RECT  90515.0 98660.0 91220.0 97315.0 ;
      RECT  90515.0 98660.0 91220.0 100005.0 ;
      RECT  90515.0 101350.0 91220.0 100005.0 ;
      RECT  90515.0 101350.0 91220.0 102695.0 ;
      RECT  90515.0 104040.0 91220.0 102695.0 ;
      RECT  90515.0 104040.0 91220.0 105385.0 ;
      RECT  90515.0 106730.0 91220.0 105385.0 ;
      RECT  90515.0 106730.0 91220.0 108075.0 ;
      RECT  90515.0 109420.0 91220.0 108075.0 ;
      RECT  90515.0 109420.0 91220.0 110765.0 ;
      RECT  90515.0 112110.0 91220.0 110765.0 ;
      RECT  90515.0 112110.0 91220.0 113455.0 ;
      RECT  90515.0 114800.0 91220.0 113455.0 ;
      RECT  90515.0 114800.0 91220.0 116145.0 ;
      RECT  90515.0 117490.0 91220.0 116145.0 ;
      RECT  90515.0 117490.0 91220.0 118835.0 ;
      RECT  90515.0 120180.0 91220.0 118835.0 ;
      RECT  90515.0 120180.0 91220.0 121525.0 ;
      RECT  90515.0 122870.0 91220.0 121525.0 ;
      RECT  90515.0 122870.0 91220.0 124215.0 ;
      RECT  90515.0 125560.0 91220.0 124215.0 ;
      RECT  90515.0 125560.0 91220.0 126905.0 ;
      RECT  90515.0 128250.0 91220.0 126905.0 ;
      RECT  90515.0 128250.0 91220.0 129595.0 ;
      RECT  90515.0 130940.0 91220.0 129595.0 ;
      RECT  90515.0 130940.0 91220.0 132285.0 ;
      RECT  90515.0 133630.0 91220.0 132285.0 ;
      RECT  90515.0 133630.0 91220.0 134975.0 ;
      RECT  90515.0 136320.0 91220.0 134975.0 ;
      RECT  90515.0 136320.0 91220.0 137665.0 ;
      RECT  90515.0 139010.0 91220.0 137665.0 ;
      RECT  90515.0 139010.0 91220.0 140355.0 ;
      RECT  90515.0 141700.0 91220.0 140355.0 ;
      RECT  90515.0 141700.0 91220.0 143045.0 ;
      RECT  90515.0 144390.0 91220.0 143045.0 ;
      RECT  90515.0 144390.0 91220.0 145735.0 ;
      RECT  90515.0 147080.0 91220.0 145735.0 ;
      RECT  90515.0 147080.0 91220.0 148425.0 ;
      RECT  90515.0 149770.0 91220.0 148425.0 ;
      RECT  90515.0 149770.0 91220.0 151115.0 ;
      RECT  90515.0 152460.0 91220.0 151115.0 ;
      RECT  90515.0 152460.0 91220.0 153805.0 ;
      RECT  90515.0 155150.0 91220.0 153805.0 ;
      RECT  90515.0 155150.0 91220.0 156495.0 ;
      RECT  90515.0 157840.0 91220.0 156495.0 ;
      RECT  90515.0 157840.0 91220.0 159185.0 ;
      RECT  90515.0 160530.0 91220.0 159185.0 ;
      RECT  90515.0 160530.0 91220.0 161875.0 ;
      RECT  90515.0 163220.0 91220.0 161875.0 ;
      RECT  90515.0 163220.0 91220.0 164565.0 ;
      RECT  90515.0 165910.0 91220.0 164565.0 ;
      RECT  90515.0 165910.0 91220.0 167255.0 ;
      RECT  90515.0 168600.0 91220.0 167255.0 ;
      RECT  90515.0 168600.0 91220.0 169945.0 ;
      RECT  90515.0 171290.0 91220.0 169945.0 ;
      RECT  90515.0 171290.0 91220.0 172635.0 ;
      RECT  90515.0 173980.0 91220.0 172635.0 ;
      RECT  90515.0 173980.0 91220.0 175325.0 ;
      RECT  90515.0 176670.0 91220.0 175325.0 ;
      RECT  90515.0 176670.0 91220.0 178015.0 ;
      RECT  90515.0 179360.0 91220.0 178015.0 ;
      RECT  90515.0 179360.0 91220.0 180705.0 ;
      RECT  90515.0 182050.0 91220.0 180705.0 ;
      RECT  90515.0 182050.0 91220.0 183395.0 ;
      RECT  90515.0 184740.0 91220.0 183395.0 ;
      RECT  90515.0 184740.0 91220.0 186085.0 ;
      RECT  90515.0 187430.0 91220.0 186085.0 ;
      RECT  90515.0 187430.0 91220.0 188775.0 ;
      RECT  90515.0 190120.0 91220.0 188775.0 ;
      RECT  90515.0 190120.0 91220.0 191465.0 ;
      RECT  90515.0 192810.0 91220.0 191465.0 ;
      RECT  90515.0 192810.0 91220.0 194155.0 ;
      RECT  90515.0 195500.0 91220.0 194155.0 ;
      RECT  90515.0 195500.0 91220.0 196845.0 ;
      RECT  90515.0 198190.0 91220.0 196845.0 ;
      RECT  90515.0 198190.0 91220.0 199535.0 ;
      RECT  90515.0 200880.0 91220.0 199535.0 ;
      RECT  90515.0 200880.0 91220.0 202225.0 ;
      RECT  90515.0 203570.0 91220.0 202225.0 ;
      RECT  90515.0 203570.0 91220.0 204915.0 ;
      RECT  90515.0 206260.0 91220.0 204915.0 ;
      RECT  91220.0 34100.0 91925.0 35445.0 ;
      RECT  91220.0 36790.0 91925.0 35445.0 ;
      RECT  91220.0 36790.0 91925.0 38135.0 ;
      RECT  91220.0 39480.0 91925.0 38135.0 ;
      RECT  91220.0 39480.0 91925.0 40825.0 ;
      RECT  91220.0 42170.0 91925.0 40825.0 ;
      RECT  91220.0 42170.0 91925.0 43515.0 ;
      RECT  91220.0 44860.0 91925.0 43515.0 ;
      RECT  91220.0 44860.0 91925.0 46205.0 ;
      RECT  91220.0 47550.0 91925.0 46205.0 ;
      RECT  91220.0 47550.0 91925.0 48895.0 ;
      RECT  91220.0 50240.0 91925.0 48895.0 ;
      RECT  91220.0 50240.0 91925.0 51585.0 ;
      RECT  91220.0 52930.0 91925.0 51585.0 ;
      RECT  91220.0 52930.0 91925.0 54275.0 ;
      RECT  91220.0 55620.0 91925.0 54275.0 ;
      RECT  91220.0 55620.0 91925.0 56965.0 ;
      RECT  91220.0 58310.0 91925.0 56965.0 ;
      RECT  91220.0 58310.0 91925.0 59655.0 ;
      RECT  91220.0 61000.0 91925.0 59655.0 ;
      RECT  91220.0 61000.0 91925.0 62345.0 ;
      RECT  91220.0 63690.0 91925.0 62345.0 ;
      RECT  91220.0 63690.0 91925.0 65035.0 ;
      RECT  91220.0 66380.0 91925.0 65035.0 ;
      RECT  91220.0 66380.0 91925.0 67725.0 ;
      RECT  91220.0 69070.0 91925.0 67725.0 ;
      RECT  91220.0 69070.0 91925.0 70415.0 ;
      RECT  91220.0 71760.0 91925.0 70415.0 ;
      RECT  91220.0 71760.0 91925.0 73105.0 ;
      RECT  91220.0 74450.0 91925.0 73105.0 ;
      RECT  91220.0 74450.0 91925.0 75795.0 ;
      RECT  91220.0 77140.0 91925.0 75795.0 ;
      RECT  91220.0 77140.0 91925.0 78485.0 ;
      RECT  91220.0 79830.0 91925.0 78485.0 ;
      RECT  91220.0 79830.0 91925.0 81175.0 ;
      RECT  91220.0 82520.0 91925.0 81175.0 ;
      RECT  91220.0 82520.0 91925.0 83865.0 ;
      RECT  91220.0 85210.0 91925.0 83865.0 ;
      RECT  91220.0 85210.0 91925.0 86555.0 ;
      RECT  91220.0 87900.0 91925.0 86555.0 ;
      RECT  91220.0 87900.0 91925.0 89245.0 ;
      RECT  91220.0 90590.0 91925.0 89245.0 ;
      RECT  91220.0 90590.0 91925.0 91935.0 ;
      RECT  91220.0 93280.0 91925.0 91935.0 ;
      RECT  91220.0 93280.0 91925.0 94625.0 ;
      RECT  91220.0 95970.0 91925.0 94625.0 ;
      RECT  91220.0 95970.0 91925.0 97315.0 ;
      RECT  91220.0 98660.0 91925.0 97315.0 ;
      RECT  91220.0 98660.0 91925.0 100005.0 ;
      RECT  91220.0 101350.0 91925.0 100005.0 ;
      RECT  91220.0 101350.0 91925.0 102695.0 ;
      RECT  91220.0 104040.0 91925.0 102695.0 ;
      RECT  91220.0 104040.0 91925.0 105385.0 ;
      RECT  91220.0 106730.0 91925.0 105385.0 ;
      RECT  91220.0 106730.0 91925.0 108075.0 ;
      RECT  91220.0 109420.0 91925.0 108075.0 ;
      RECT  91220.0 109420.0 91925.0 110765.0 ;
      RECT  91220.0 112110.0 91925.0 110765.0 ;
      RECT  91220.0 112110.0 91925.0 113455.0 ;
      RECT  91220.0 114800.0 91925.0 113455.0 ;
      RECT  91220.0 114800.0 91925.0 116145.0 ;
      RECT  91220.0 117490.0 91925.0 116145.0 ;
      RECT  91220.0 117490.0 91925.0 118835.0 ;
      RECT  91220.0 120180.0 91925.0 118835.0 ;
      RECT  91220.0 120180.0 91925.0 121525.0 ;
      RECT  91220.0 122870.0 91925.0 121525.0 ;
      RECT  91220.0 122870.0 91925.0 124215.0 ;
      RECT  91220.0 125560.0 91925.0 124215.0 ;
      RECT  91220.0 125560.0 91925.0 126905.0 ;
      RECT  91220.0 128250.0 91925.0 126905.0 ;
      RECT  91220.0 128250.0 91925.0 129595.0 ;
      RECT  91220.0 130940.0 91925.0 129595.0 ;
      RECT  91220.0 130940.0 91925.0 132285.0 ;
      RECT  91220.0 133630.0 91925.0 132285.0 ;
      RECT  91220.0 133630.0 91925.0 134975.0 ;
      RECT  91220.0 136320.0 91925.0 134975.0 ;
      RECT  91220.0 136320.0 91925.0 137665.0 ;
      RECT  91220.0 139010.0 91925.0 137665.0 ;
      RECT  91220.0 139010.0 91925.0 140355.0 ;
      RECT  91220.0 141700.0 91925.0 140355.0 ;
      RECT  91220.0 141700.0 91925.0 143045.0 ;
      RECT  91220.0 144390.0 91925.0 143045.0 ;
      RECT  91220.0 144390.0 91925.0 145735.0 ;
      RECT  91220.0 147080.0 91925.0 145735.0 ;
      RECT  91220.0 147080.0 91925.0 148425.0 ;
      RECT  91220.0 149770.0 91925.0 148425.0 ;
      RECT  91220.0 149770.0 91925.0 151115.0 ;
      RECT  91220.0 152460.0 91925.0 151115.0 ;
      RECT  91220.0 152460.0 91925.0 153805.0 ;
      RECT  91220.0 155150.0 91925.0 153805.0 ;
      RECT  91220.0 155150.0 91925.0 156495.0 ;
      RECT  91220.0 157840.0 91925.0 156495.0 ;
      RECT  91220.0 157840.0 91925.0 159185.0 ;
      RECT  91220.0 160530.0 91925.0 159185.0 ;
      RECT  91220.0 160530.0 91925.0 161875.0 ;
      RECT  91220.0 163220.0 91925.0 161875.0 ;
      RECT  91220.0 163220.0 91925.0 164565.0 ;
      RECT  91220.0 165910.0 91925.0 164565.0 ;
      RECT  91220.0 165910.0 91925.0 167255.0 ;
      RECT  91220.0 168600.0 91925.0 167255.0 ;
      RECT  91220.0 168600.0 91925.0 169945.0 ;
      RECT  91220.0 171290.0 91925.0 169945.0 ;
      RECT  91220.0 171290.0 91925.0 172635.0 ;
      RECT  91220.0 173980.0 91925.0 172635.0 ;
      RECT  91220.0 173980.0 91925.0 175325.0 ;
      RECT  91220.0 176670.0 91925.0 175325.0 ;
      RECT  91220.0 176670.0 91925.0 178015.0 ;
      RECT  91220.0 179360.0 91925.0 178015.0 ;
      RECT  91220.0 179360.0 91925.0 180705.0 ;
      RECT  91220.0 182050.0 91925.0 180705.0 ;
      RECT  91220.0 182050.0 91925.0 183395.0 ;
      RECT  91220.0 184740.0 91925.0 183395.0 ;
      RECT  91220.0 184740.0 91925.0 186085.0 ;
      RECT  91220.0 187430.0 91925.0 186085.0 ;
      RECT  91220.0 187430.0 91925.0 188775.0 ;
      RECT  91220.0 190120.0 91925.0 188775.0 ;
      RECT  91220.0 190120.0 91925.0 191465.0 ;
      RECT  91220.0 192810.0 91925.0 191465.0 ;
      RECT  91220.0 192810.0 91925.0 194155.0 ;
      RECT  91220.0 195500.0 91925.0 194155.0 ;
      RECT  91220.0 195500.0 91925.0 196845.0 ;
      RECT  91220.0 198190.0 91925.0 196845.0 ;
      RECT  91220.0 198190.0 91925.0 199535.0 ;
      RECT  91220.0 200880.0 91925.0 199535.0 ;
      RECT  91220.0 200880.0 91925.0 202225.0 ;
      RECT  91220.0 203570.0 91925.0 202225.0 ;
      RECT  91220.0 203570.0 91925.0 204915.0 ;
      RECT  91220.0 206260.0 91925.0 204915.0 ;
      RECT  91925.0 34100.0 92630.0 35445.0 ;
      RECT  91925.0 36790.0 92630.0 35445.0 ;
      RECT  91925.0 36790.0 92630.0 38135.0 ;
      RECT  91925.0 39480.0 92630.0 38135.0 ;
      RECT  91925.0 39480.0 92630.0 40825.0 ;
      RECT  91925.0 42170.0 92630.0 40825.0 ;
      RECT  91925.0 42170.0 92630.0 43515.0 ;
      RECT  91925.0 44860.0 92630.0 43515.0 ;
      RECT  91925.0 44860.0 92630.0 46205.0 ;
      RECT  91925.0 47550.0 92630.0 46205.0 ;
      RECT  91925.0 47550.0 92630.0 48895.0 ;
      RECT  91925.0 50240.0 92630.0 48895.0 ;
      RECT  91925.0 50240.0 92630.0 51585.0 ;
      RECT  91925.0 52930.0 92630.0 51585.0 ;
      RECT  91925.0 52930.0 92630.0 54275.0 ;
      RECT  91925.0 55620.0 92630.0 54275.0 ;
      RECT  91925.0 55620.0 92630.0 56965.0 ;
      RECT  91925.0 58310.0 92630.0 56965.0 ;
      RECT  91925.0 58310.0 92630.0 59655.0 ;
      RECT  91925.0 61000.0 92630.0 59655.0 ;
      RECT  91925.0 61000.0 92630.0 62345.0 ;
      RECT  91925.0 63690.0 92630.0 62345.0 ;
      RECT  91925.0 63690.0 92630.0 65035.0 ;
      RECT  91925.0 66380.0 92630.0 65035.0 ;
      RECT  91925.0 66380.0 92630.0 67725.0 ;
      RECT  91925.0 69070.0 92630.0 67725.0 ;
      RECT  91925.0 69070.0 92630.0 70415.0 ;
      RECT  91925.0 71760.0 92630.0 70415.0 ;
      RECT  91925.0 71760.0 92630.0 73105.0 ;
      RECT  91925.0 74450.0 92630.0 73105.0 ;
      RECT  91925.0 74450.0 92630.0 75795.0 ;
      RECT  91925.0 77140.0 92630.0 75795.0 ;
      RECT  91925.0 77140.0 92630.0 78485.0 ;
      RECT  91925.0 79830.0 92630.0 78485.0 ;
      RECT  91925.0 79830.0 92630.0 81175.0 ;
      RECT  91925.0 82520.0 92630.0 81175.0 ;
      RECT  91925.0 82520.0 92630.0 83865.0 ;
      RECT  91925.0 85210.0 92630.0 83865.0 ;
      RECT  91925.0 85210.0 92630.0 86555.0 ;
      RECT  91925.0 87900.0 92630.0 86555.0 ;
      RECT  91925.0 87900.0 92630.0 89245.0 ;
      RECT  91925.0 90590.0 92630.0 89245.0 ;
      RECT  91925.0 90590.0 92630.0 91935.0 ;
      RECT  91925.0 93280.0 92630.0 91935.0 ;
      RECT  91925.0 93280.0 92630.0 94625.0 ;
      RECT  91925.0 95970.0 92630.0 94625.0 ;
      RECT  91925.0 95970.0 92630.0 97315.0 ;
      RECT  91925.0 98660.0 92630.0 97315.0 ;
      RECT  91925.0 98660.0 92630.0 100005.0 ;
      RECT  91925.0 101350.0 92630.0 100005.0 ;
      RECT  91925.0 101350.0 92630.0 102695.0 ;
      RECT  91925.0 104040.0 92630.0 102695.0 ;
      RECT  91925.0 104040.0 92630.0 105385.0 ;
      RECT  91925.0 106730.0 92630.0 105385.0 ;
      RECT  91925.0 106730.0 92630.0 108075.0 ;
      RECT  91925.0 109420.0 92630.0 108075.0 ;
      RECT  91925.0 109420.0 92630.0 110765.0 ;
      RECT  91925.0 112110.0 92630.0 110765.0 ;
      RECT  91925.0 112110.0 92630.0 113455.0 ;
      RECT  91925.0 114800.0 92630.0 113455.0 ;
      RECT  91925.0 114800.0 92630.0 116145.0 ;
      RECT  91925.0 117490.0 92630.0 116145.0 ;
      RECT  91925.0 117490.0 92630.0 118835.0 ;
      RECT  91925.0 120180.0 92630.0 118835.0 ;
      RECT  91925.0 120180.0 92630.0 121525.0 ;
      RECT  91925.0 122870.0 92630.0 121525.0 ;
      RECT  91925.0 122870.0 92630.0 124215.0 ;
      RECT  91925.0 125560.0 92630.0 124215.0 ;
      RECT  91925.0 125560.0 92630.0 126905.0 ;
      RECT  91925.0 128250.0 92630.0 126905.0 ;
      RECT  91925.0 128250.0 92630.0 129595.0 ;
      RECT  91925.0 130940.0 92630.0 129595.0 ;
      RECT  91925.0 130940.0 92630.0 132285.0 ;
      RECT  91925.0 133630.0 92630.0 132285.0 ;
      RECT  91925.0 133630.0 92630.0 134975.0 ;
      RECT  91925.0 136320.0 92630.0 134975.0 ;
      RECT  91925.0 136320.0 92630.0 137665.0 ;
      RECT  91925.0 139010.0 92630.0 137665.0 ;
      RECT  91925.0 139010.0 92630.0 140355.0 ;
      RECT  91925.0 141700.0 92630.0 140355.0 ;
      RECT  91925.0 141700.0 92630.0 143045.0 ;
      RECT  91925.0 144390.0 92630.0 143045.0 ;
      RECT  91925.0 144390.0 92630.0 145735.0 ;
      RECT  91925.0 147080.0 92630.0 145735.0 ;
      RECT  91925.0 147080.0 92630.0 148425.0 ;
      RECT  91925.0 149770.0 92630.0 148425.0 ;
      RECT  91925.0 149770.0 92630.0 151115.0 ;
      RECT  91925.0 152460.0 92630.0 151115.0 ;
      RECT  91925.0 152460.0 92630.0 153805.0 ;
      RECT  91925.0 155150.0 92630.0 153805.0 ;
      RECT  91925.0 155150.0 92630.0 156495.0 ;
      RECT  91925.0 157840.0 92630.0 156495.0 ;
      RECT  91925.0 157840.0 92630.0 159185.0 ;
      RECT  91925.0 160530.0 92630.0 159185.0 ;
      RECT  91925.0 160530.0 92630.0 161875.0 ;
      RECT  91925.0 163220.0 92630.0 161875.0 ;
      RECT  91925.0 163220.0 92630.0 164565.0 ;
      RECT  91925.0 165910.0 92630.0 164565.0 ;
      RECT  91925.0 165910.0 92630.0 167255.0 ;
      RECT  91925.0 168600.0 92630.0 167255.0 ;
      RECT  91925.0 168600.0 92630.0 169945.0 ;
      RECT  91925.0 171290.0 92630.0 169945.0 ;
      RECT  91925.0 171290.0 92630.0 172635.0 ;
      RECT  91925.0 173980.0 92630.0 172635.0 ;
      RECT  91925.0 173980.0 92630.0 175325.0 ;
      RECT  91925.0 176670.0 92630.0 175325.0 ;
      RECT  91925.0 176670.0 92630.0 178015.0 ;
      RECT  91925.0 179360.0 92630.0 178015.0 ;
      RECT  91925.0 179360.0 92630.0 180705.0 ;
      RECT  91925.0 182050.0 92630.0 180705.0 ;
      RECT  91925.0 182050.0 92630.0 183395.0 ;
      RECT  91925.0 184740.0 92630.0 183395.0 ;
      RECT  91925.0 184740.0 92630.0 186085.0 ;
      RECT  91925.0 187430.0 92630.0 186085.0 ;
      RECT  91925.0 187430.0 92630.0 188775.0 ;
      RECT  91925.0 190120.0 92630.0 188775.0 ;
      RECT  91925.0 190120.0 92630.0 191465.0 ;
      RECT  91925.0 192810.0 92630.0 191465.0 ;
      RECT  91925.0 192810.0 92630.0 194155.0 ;
      RECT  91925.0 195500.0 92630.0 194155.0 ;
      RECT  91925.0 195500.0 92630.0 196845.0 ;
      RECT  91925.0 198190.0 92630.0 196845.0 ;
      RECT  91925.0 198190.0 92630.0 199535.0 ;
      RECT  91925.0 200880.0 92630.0 199535.0 ;
      RECT  91925.0 200880.0 92630.0 202225.0 ;
      RECT  91925.0 203570.0 92630.0 202225.0 ;
      RECT  91925.0 203570.0 92630.0 204915.0 ;
      RECT  91925.0 206260.0 92630.0 204915.0 ;
      RECT  92630.0 34100.0 93335.0 35445.0 ;
      RECT  92630.0 36790.0 93335.0 35445.0 ;
      RECT  92630.0 36790.0 93335.0 38135.0 ;
      RECT  92630.0 39480.0 93335.0 38135.0 ;
      RECT  92630.0 39480.0 93335.0 40825.0 ;
      RECT  92630.0 42170.0 93335.0 40825.0 ;
      RECT  92630.0 42170.0 93335.0 43515.0 ;
      RECT  92630.0 44860.0 93335.0 43515.0 ;
      RECT  92630.0 44860.0 93335.0 46205.0 ;
      RECT  92630.0 47550.0 93335.0 46205.0 ;
      RECT  92630.0 47550.0 93335.0 48895.0 ;
      RECT  92630.0 50240.0 93335.0 48895.0 ;
      RECT  92630.0 50240.0 93335.0 51585.0 ;
      RECT  92630.0 52930.0 93335.0 51585.0 ;
      RECT  92630.0 52930.0 93335.0 54275.0 ;
      RECT  92630.0 55620.0 93335.0 54275.0 ;
      RECT  92630.0 55620.0 93335.0 56965.0 ;
      RECT  92630.0 58310.0 93335.0 56965.0 ;
      RECT  92630.0 58310.0 93335.0 59655.0 ;
      RECT  92630.0 61000.0 93335.0 59655.0 ;
      RECT  92630.0 61000.0 93335.0 62345.0 ;
      RECT  92630.0 63690.0 93335.0 62345.0 ;
      RECT  92630.0 63690.0 93335.0 65035.0 ;
      RECT  92630.0 66380.0 93335.0 65035.0 ;
      RECT  92630.0 66380.0 93335.0 67725.0 ;
      RECT  92630.0 69070.0 93335.0 67725.0 ;
      RECT  92630.0 69070.0 93335.0 70415.0 ;
      RECT  92630.0 71760.0 93335.0 70415.0 ;
      RECT  92630.0 71760.0 93335.0 73105.0 ;
      RECT  92630.0 74450.0 93335.0 73105.0 ;
      RECT  92630.0 74450.0 93335.0 75795.0 ;
      RECT  92630.0 77140.0 93335.0 75795.0 ;
      RECT  92630.0 77140.0 93335.0 78485.0 ;
      RECT  92630.0 79830.0 93335.0 78485.0 ;
      RECT  92630.0 79830.0 93335.0 81175.0 ;
      RECT  92630.0 82520.0 93335.0 81175.0 ;
      RECT  92630.0 82520.0 93335.0 83865.0 ;
      RECT  92630.0 85210.0 93335.0 83865.0 ;
      RECT  92630.0 85210.0 93335.0 86555.0 ;
      RECT  92630.0 87900.0 93335.0 86555.0 ;
      RECT  92630.0 87900.0 93335.0 89245.0 ;
      RECT  92630.0 90590.0 93335.0 89245.0 ;
      RECT  92630.0 90590.0 93335.0 91935.0 ;
      RECT  92630.0 93280.0 93335.0 91935.0 ;
      RECT  92630.0 93280.0 93335.0 94625.0 ;
      RECT  92630.0 95970.0 93335.0 94625.0 ;
      RECT  92630.0 95970.0 93335.0 97315.0 ;
      RECT  92630.0 98660.0 93335.0 97315.0 ;
      RECT  92630.0 98660.0 93335.0 100005.0 ;
      RECT  92630.0 101350.0 93335.0 100005.0 ;
      RECT  92630.0 101350.0 93335.0 102695.0 ;
      RECT  92630.0 104040.0 93335.0 102695.0 ;
      RECT  92630.0 104040.0 93335.0 105385.0 ;
      RECT  92630.0 106730.0 93335.0 105385.0 ;
      RECT  92630.0 106730.0 93335.0 108075.0 ;
      RECT  92630.0 109420.0 93335.0 108075.0 ;
      RECT  92630.0 109420.0 93335.0 110765.0 ;
      RECT  92630.0 112110.0 93335.0 110765.0 ;
      RECT  92630.0 112110.0 93335.0 113455.0 ;
      RECT  92630.0 114800.0 93335.0 113455.0 ;
      RECT  92630.0 114800.0 93335.0 116145.0 ;
      RECT  92630.0 117490.0 93335.0 116145.0 ;
      RECT  92630.0 117490.0 93335.0 118835.0 ;
      RECT  92630.0 120180.0 93335.0 118835.0 ;
      RECT  92630.0 120180.0 93335.0 121525.0 ;
      RECT  92630.0 122870.0 93335.0 121525.0 ;
      RECT  92630.0 122870.0 93335.0 124215.0 ;
      RECT  92630.0 125560.0 93335.0 124215.0 ;
      RECT  92630.0 125560.0 93335.0 126905.0 ;
      RECT  92630.0 128250.0 93335.0 126905.0 ;
      RECT  92630.0 128250.0 93335.0 129595.0 ;
      RECT  92630.0 130940.0 93335.0 129595.0 ;
      RECT  92630.0 130940.0 93335.0 132285.0 ;
      RECT  92630.0 133630.0 93335.0 132285.0 ;
      RECT  92630.0 133630.0 93335.0 134975.0 ;
      RECT  92630.0 136320.0 93335.0 134975.0 ;
      RECT  92630.0 136320.0 93335.0 137665.0 ;
      RECT  92630.0 139010.0 93335.0 137665.0 ;
      RECT  92630.0 139010.0 93335.0 140355.0 ;
      RECT  92630.0 141700.0 93335.0 140355.0 ;
      RECT  92630.0 141700.0 93335.0 143045.0 ;
      RECT  92630.0 144390.0 93335.0 143045.0 ;
      RECT  92630.0 144390.0 93335.0 145735.0 ;
      RECT  92630.0 147080.0 93335.0 145735.0 ;
      RECT  92630.0 147080.0 93335.0 148425.0 ;
      RECT  92630.0 149770.0 93335.0 148425.0 ;
      RECT  92630.0 149770.0 93335.0 151115.0 ;
      RECT  92630.0 152460.0 93335.0 151115.0 ;
      RECT  92630.0 152460.0 93335.0 153805.0 ;
      RECT  92630.0 155150.0 93335.0 153805.0 ;
      RECT  92630.0 155150.0 93335.0 156495.0 ;
      RECT  92630.0 157840.0 93335.0 156495.0 ;
      RECT  92630.0 157840.0 93335.0 159185.0 ;
      RECT  92630.0 160530.0 93335.0 159185.0 ;
      RECT  92630.0 160530.0 93335.0 161875.0 ;
      RECT  92630.0 163220.0 93335.0 161875.0 ;
      RECT  92630.0 163220.0 93335.0 164565.0 ;
      RECT  92630.0 165910.0 93335.0 164565.0 ;
      RECT  92630.0 165910.0 93335.0 167255.0 ;
      RECT  92630.0 168600.0 93335.0 167255.0 ;
      RECT  92630.0 168600.0 93335.0 169945.0 ;
      RECT  92630.0 171290.0 93335.0 169945.0 ;
      RECT  92630.0 171290.0 93335.0 172635.0 ;
      RECT  92630.0 173980.0 93335.0 172635.0 ;
      RECT  92630.0 173980.0 93335.0 175325.0 ;
      RECT  92630.0 176670.0 93335.0 175325.0 ;
      RECT  92630.0 176670.0 93335.0 178015.0 ;
      RECT  92630.0 179360.0 93335.0 178015.0 ;
      RECT  92630.0 179360.0 93335.0 180705.0 ;
      RECT  92630.0 182050.0 93335.0 180705.0 ;
      RECT  92630.0 182050.0 93335.0 183395.0 ;
      RECT  92630.0 184740.0 93335.0 183395.0 ;
      RECT  92630.0 184740.0 93335.0 186085.0 ;
      RECT  92630.0 187430.0 93335.0 186085.0 ;
      RECT  92630.0 187430.0 93335.0 188775.0 ;
      RECT  92630.0 190120.0 93335.0 188775.0 ;
      RECT  92630.0 190120.0 93335.0 191465.0 ;
      RECT  92630.0 192810.0 93335.0 191465.0 ;
      RECT  92630.0 192810.0 93335.0 194155.0 ;
      RECT  92630.0 195500.0 93335.0 194155.0 ;
      RECT  92630.0 195500.0 93335.0 196845.0 ;
      RECT  92630.0 198190.0 93335.0 196845.0 ;
      RECT  92630.0 198190.0 93335.0 199535.0 ;
      RECT  92630.0 200880.0 93335.0 199535.0 ;
      RECT  92630.0 200880.0 93335.0 202225.0 ;
      RECT  92630.0 203570.0 93335.0 202225.0 ;
      RECT  92630.0 203570.0 93335.0 204915.0 ;
      RECT  92630.0 206260.0 93335.0 204915.0 ;
      RECT  93335.0 34100.0 94040.0 35445.0 ;
      RECT  93335.0 36790.0 94040.0 35445.0 ;
      RECT  93335.0 36790.0 94040.0 38135.0 ;
      RECT  93335.0 39480.0 94040.0 38135.0 ;
      RECT  93335.0 39480.0 94040.0 40825.0 ;
      RECT  93335.0 42170.0 94040.0 40825.0 ;
      RECT  93335.0 42170.0 94040.0 43515.0 ;
      RECT  93335.0 44860.0 94040.0 43515.0 ;
      RECT  93335.0 44860.0 94040.0 46205.0 ;
      RECT  93335.0 47550.0 94040.0 46205.0 ;
      RECT  93335.0 47550.0 94040.0 48895.0 ;
      RECT  93335.0 50240.0 94040.0 48895.0 ;
      RECT  93335.0 50240.0 94040.0 51585.0 ;
      RECT  93335.0 52930.0 94040.0 51585.0 ;
      RECT  93335.0 52930.0 94040.0 54275.0 ;
      RECT  93335.0 55620.0 94040.0 54275.0 ;
      RECT  93335.0 55620.0 94040.0 56965.0 ;
      RECT  93335.0 58310.0 94040.0 56965.0 ;
      RECT  93335.0 58310.0 94040.0 59655.0 ;
      RECT  93335.0 61000.0 94040.0 59655.0 ;
      RECT  93335.0 61000.0 94040.0 62345.0 ;
      RECT  93335.0 63690.0 94040.0 62345.0 ;
      RECT  93335.0 63690.0 94040.0 65035.0 ;
      RECT  93335.0 66380.0 94040.0 65035.0 ;
      RECT  93335.0 66380.0 94040.0 67725.0 ;
      RECT  93335.0 69070.0 94040.0 67725.0 ;
      RECT  93335.0 69070.0 94040.0 70415.0 ;
      RECT  93335.0 71760.0 94040.0 70415.0 ;
      RECT  93335.0 71760.0 94040.0 73105.0 ;
      RECT  93335.0 74450.0 94040.0 73105.0 ;
      RECT  93335.0 74450.0 94040.0 75795.0 ;
      RECT  93335.0 77140.0 94040.0 75795.0 ;
      RECT  93335.0 77140.0 94040.0 78485.0 ;
      RECT  93335.0 79830.0 94040.0 78485.0 ;
      RECT  93335.0 79830.0 94040.0 81175.0 ;
      RECT  93335.0 82520.0 94040.0 81175.0 ;
      RECT  93335.0 82520.0 94040.0 83865.0 ;
      RECT  93335.0 85210.0 94040.0 83865.0 ;
      RECT  93335.0 85210.0 94040.0 86555.0 ;
      RECT  93335.0 87900.0 94040.0 86555.0 ;
      RECT  93335.0 87900.0 94040.0 89245.0 ;
      RECT  93335.0 90590.0 94040.0 89245.0 ;
      RECT  93335.0 90590.0 94040.0 91935.0 ;
      RECT  93335.0 93280.0 94040.0 91935.0 ;
      RECT  93335.0 93280.0 94040.0 94625.0 ;
      RECT  93335.0 95970.0 94040.0 94625.0 ;
      RECT  93335.0 95970.0 94040.0 97315.0 ;
      RECT  93335.0 98660.0 94040.0 97315.0 ;
      RECT  93335.0 98660.0 94040.0 100005.0 ;
      RECT  93335.0 101350.0 94040.0 100005.0 ;
      RECT  93335.0 101350.0 94040.0 102695.0 ;
      RECT  93335.0 104040.0 94040.0 102695.0 ;
      RECT  93335.0 104040.0 94040.0 105385.0 ;
      RECT  93335.0 106730.0 94040.0 105385.0 ;
      RECT  93335.0 106730.0 94040.0 108075.0 ;
      RECT  93335.0 109420.0 94040.0 108075.0 ;
      RECT  93335.0 109420.0 94040.0 110765.0 ;
      RECT  93335.0 112110.0 94040.0 110765.0 ;
      RECT  93335.0 112110.0 94040.0 113455.0 ;
      RECT  93335.0 114800.0 94040.0 113455.0 ;
      RECT  93335.0 114800.0 94040.0 116145.0 ;
      RECT  93335.0 117490.0 94040.0 116145.0 ;
      RECT  93335.0 117490.0 94040.0 118835.0 ;
      RECT  93335.0 120180.0 94040.0 118835.0 ;
      RECT  93335.0 120180.0 94040.0 121525.0 ;
      RECT  93335.0 122870.0 94040.0 121525.0 ;
      RECT  93335.0 122870.0 94040.0 124215.0 ;
      RECT  93335.0 125560.0 94040.0 124215.0 ;
      RECT  93335.0 125560.0 94040.0 126905.0 ;
      RECT  93335.0 128250.0 94040.0 126905.0 ;
      RECT  93335.0 128250.0 94040.0 129595.0 ;
      RECT  93335.0 130940.0 94040.0 129595.0 ;
      RECT  93335.0 130940.0 94040.0 132285.0 ;
      RECT  93335.0 133630.0 94040.0 132285.0 ;
      RECT  93335.0 133630.0 94040.0 134975.0 ;
      RECT  93335.0 136320.0 94040.0 134975.0 ;
      RECT  93335.0 136320.0 94040.0 137665.0 ;
      RECT  93335.0 139010.0 94040.0 137665.0 ;
      RECT  93335.0 139010.0 94040.0 140355.0 ;
      RECT  93335.0 141700.0 94040.0 140355.0 ;
      RECT  93335.0 141700.0 94040.0 143045.0 ;
      RECT  93335.0 144390.0 94040.0 143045.0 ;
      RECT  93335.0 144390.0 94040.0 145735.0 ;
      RECT  93335.0 147080.0 94040.0 145735.0 ;
      RECT  93335.0 147080.0 94040.0 148425.0 ;
      RECT  93335.0 149770.0 94040.0 148425.0 ;
      RECT  93335.0 149770.0 94040.0 151115.0 ;
      RECT  93335.0 152460.0 94040.0 151115.0 ;
      RECT  93335.0 152460.0 94040.0 153805.0 ;
      RECT  93335.0 155150.0 94040.0 153805.0 ;
      RECT  93335.0 155150.0 94040.0 156495.0 ;
      RECT  93335.0 157840.0 94040.0 156495.0 ;
      RECT  93335.0 157840.0 94040.0 159185.0 ;
      RECT  93335.0 160530.0 94040.0 159185.0 ;
      RECT  93335.0 160530.0 94040.0 161875.0 ;
      RECT  93335.0 163220.0 94040.0 161875.0 ;
      RECT  93335.0 163220.0 94040.0 164565.0 ;
      RECT  93335.0 165910.0 94040.0 164565.0 ;
      RECT  93335.0 165910.0 94040.0 167255.0 ;
      RECT  93335.0 168600.0 94040.0 167255.0 ;
      RECT  93335.0 168600.0 94040.0 169945.0 ;
      RECT  93335.0 171290.0 94040.0 169945.0 ;
      RECT  93335.0 171290.0 94040.0 172635.0 ;
      RECT  93335.0 173980.0 94040.0 172635.0 ;
      RECT  93335.0 173980.0 94040.0 175325.0 ;
      RECT  93335.0 176670.0 94040.0 175325.0 ;
      RECT  93335.0 176670.0 94040.0 178015.0 ;
      RECT  93335.0 179360.0 94040.0 178015.0 ;
      RECT  93335.0 179360.0 94040.0 180705.0 ;
      RECT  93335.0 182050.0 94040.0 180705.0 ;
      RECT  93335.0 182050.0 94040.0 183395.0 ;
      RECT  93335.0 184740.0 94040.0 183395.0 ;
      RECT  93335.0 184740.0 94040.0 186085.0 ;
      RECT  93335.0 187430.0 94040.0 186085.0 ;
      RECT  93335.0 187430.0 94040.0 188775.0 ;
      RECT  93335.0 190120.0 94040.0 188775.0 ;
      RECT  93335.0 190120.0 94040.0 191465.0 ;
      RECT  93335.0 192810.0 94040.0 191465.0 ;
      RECT  93335.0 192810.0 94040.0 194155.0 ;
      RECT  93335.0 195500.0 94040.0 194155.0 ;
      RECT  93335.0 195500.0 94040.0 196845.0 ;
      RECT  93335.0 198190.0 94040.0 196845.0 ;
      RECT  93335.0 198190.0 94040.0 199535.0 ;
      RECT  93335.0 200880.0 94040.0 199535.0 ;
      RECT  93335.0 200880.0 94040.0 202225.0 ;
      RECT  93335.0 203570.0 94040.0 202225.0 ;
      RECT  93335.0 203570.0 94040.0 204915.0 ;
      RECT  93335.0 206260.0 94040.0 204915.0 ;
      RECT  94040.0 34100.0 94745.0 35445.0 ;
      RECT  94040.0 36790.0 94745.0 35445.0 ;
      RECT  94040.0 36790.0 94745.0 38135.0 ;
      RECT  94040.0 39480.0 94745.0 38135.0 ;
      RECT  94040.0 39480.0 94745.0 40825.0 ;
      RECT  94040.0 42170.0 94745.0 40825.0 ;
      RECT  94040.0 42170.0 94745.0 43515.0 ;
      RECT  94040.0 44860.0 94745.0 43515.0 ;
      RECT  94040.0 44860.0 94745.0 46205.0 ;
      RECT  94040.0 47550.0 94745.0 46205.0 ;
      RECT  94040.0 47550.0 94745.0 48895.0 ;
      RECT  94040.0 50240.0 94745.0 48895.0 ;
      RECT  94040.0 50240.0 94745.0 51585.0 ;
      RECT  94040.0 52930.0 94745.0 51585.0 ;
      RECT  94040.0 52930.0 94745.0 54275.0 ;
      RECT  94040.0 55620.0 94745.0 54275.0 ;
      RECT  94040.0 55620.0 94745.0 56965.0 ;
      RECT  94040.0 58310.0 94745.0 56965.0 ;
      RECT  94040.0 58310.0 94745.0 59655.0 ;
      RECT  94040.0 61000.0 94745.0 59655.0 ;
      RECT  94040.0 61000.0 94745.0 62345.0 ;
      RECT  94040.0 63690.0 94745.0 62345.0 ;
      RECT  94040.0 63690.0 94745.0 65035.0 ;
      RECT  94040.0 66380.0 94745.0 65035.0 ;
      RECT  94040.0 66380.0 94745.0 67725.0 ;
      RECT  94040.0 69070.0 94745.0 67725.0 ;
      RECT  94040.0 69070.0 94745.0 70415.0 ;
      RECT  94040.0 71760.0 94745.0 70415.0 ;
      RECT  94040.0 71760.0 94745.0 73105.0 ;
      RECT  94040.0 74450.0 94745.0 73105.0 ;
      RECT  94040.0 74450.0 94745.0 75795.0 ;
      RECT  94040.0 77140.0 94745.0 75795.0 ;
      RECT  94040.0 77140.0 94745.0 78485.0 ;
      RECT  94040.0 79830.0 94745.0 78485.0 ;
      RECT  94040.0 79830.0 94745.0 81175.0 ;
      RECT  94040.0 82520.0 94745.0 81175.0 ;
      RECT  94040.0 82520.0 94745.0 83865.0 ;
      RECT  94040.0 85210.0 94745.0 83865.0 ;
      RECT  94040.0 85210.0 94745.0 86555.0 ;
      RECT  94040.0 87900.0 94745.0 86555.0 ;
      RECT  94040.0 87900.0 94745.0 89245.0 ;
      RECT  94040.0 90590.0 94745.0 89245.0 ;
      RECT  94040.0 90590.0 94745.0 91935.0 ;
      RECT  94040.0 93280.0 94745.0 91935.0 ;
      RECT  94040.0 93280.0 94745.0 94625.0 ;
      RECT  94040.0 95970.0 94745.0 94625.0 ;
      RECT  94040.0 95970.0 94745.0 97315.0 ;
      RECT  94040.0 98660.0 94745.0 97315.0 ;
      RECT  94040.0 98660.0 94745.0 100005.0 ;
      RECT  94040.0 101350.0 94745.0 100005.0 ;
      RECT  94040.0 101350.0 94745.0 102695.0 ;
      RECT  94040.0 104040.0 94745.0 102695.0 ;
      RECT  94040.0 104040.0 94745.0 105385.0 ;
      RECT  94040.0 106730.0 94745.0 105385.0 ;
      RECT  94040.0 106730.0 94745.0 108075.0 ;
      RECT  94040.0 109420.0 94745.0 108075.0 ;
      RECT  94040.0 109420.0 94745.0 110765.0 ;
      RECT  94040.0 112110.0 94745.0 110765.0 ;
      RECT  94040.0 112110.0 94745.0 113455.0 ;
      RECT  94040.0 114800.0 94745.0 113455.0 ;
      RECT  94040.0 114800.0 94745.0 116145.0 ;
      RECT  94040.0 117490.0 94745.0 116145.0 ;
      RECT  94040.0 117490.0 94745.0 118835.0 ;
      RECT  94040.0 120180.0 94745.0 118835.0 ;
      RECT  94040.0 120180.0 94745.0 121525.0 ;
      RECT  94040.0 122870.0 94745.0 121525.0 ;
      RECT  94040.0 122870.0 94745.0 124215.0 ;
      RECT  94040.0 125560.0 94745.0 124215.0 ;
      RECT  94040.0 125560.0 94745.0 126905.0 ;
      RECT  94040.0 128250.0 94745.0 126905.0 ;
      RECT  94040.0 128250.0 94745.0 129595.0 ;
      RECT  94040.0 130940.0 94745.0 129595.0 ;
      RECT  94040.0 130940.0 94745.0 132285.0 ;
      RECT  94040.0 133630.0 94745.0 132285.0 ;
      RECT  94040.0 133630.0 94745.0 134975.0 ;
      RECT  94040.0 136320.0 94745.0 134975.0 ;
      RECT  94040.0 136320.0 94745.0 137665.0 ;
      RECT  94040.0 139010.0 94745.0 137665.0 ;
      RECT  94040.0 139010.0 94745.0 140355.0 ;
      RECT  94040.0 141700.0 94745.0 140355.0 ;
      RECT  94040.0 141700.0 94745.0 143045.0 ;
      RECT  94040.0 144390.0 94745.0 143045.0 ;
      RECT  94040.0 144390.0 94745.0 145735.0 ;
      RECT  94040.0 147080.0 94745.0 145735.0 ;
      RECT  94040.0 147080.0 94745.0 148425.0 ;
      RECT  94040.0 149770.0 94745.0 148425.0 ;
      RECT  94040.0 149770.0 94745.0 151115.0 ;
      RECT  94040.0 152460.0 94745.0 151115.0 ;
      RECT  94040.0 152460.0 94745.0 153805.0 ;
      RECT  94040.0 155150.0 94745.0 153805.0 ;
      RECT  94040.0 155150.0 94745.0 156495.0 ;
      RECT  94040.0 157840.0 94745.0 156495.0 ;
      RECT  94040.0 157840.0 94745.0 159185.0 ;
      RECT  94040.0 160530.0 94745.0 159185.0 ;
      RECT  94040.0 160530.0 94745.0 161875.0 ;
      RECT  94040.0 163220.0 94745.0 161875.0 ;
      RECT  94040.0 163220.0 94745.0 164565.0 ;
      RECT  94040.0 165910.0 94745.0 164565.0 ;
      RECT  94040.0 165910.0 94745.0 167255.0 ;
      RECT  94040.0 168600.0 94745.0 167255.0 ;
      RECT  94040.0 168600.0 94745.0 169945.0 ;
      RECT  94040.0 171290.0 94745.0 169945.0 ;
      RECT  94040.0 171290.0 94745.0 172635.0 ;
      RECT  94040.0 173980.0 94745.0 172635.0 ;
      RECT  94040.0 173980.0 94745.0 175325.0 ;
      RECT  94040.0 176670.0 94745.0 175325.0 ;
      RECT  94040.0 176670.0 94745.0 178015.0 ;
      RECT  94040.0 179360.0 94745.0 178015.0 ;
      RECT  94040.0 179360.0 94745.0 180705.0 ;
      RECT  94040.0 182050.0 94745.0 180705.0 ;
      RECT  94040.0 182050.0 94745.0 183395.0 ;
      RECT  94040.0 184740.0 94745.0 183395.0 ;
      RECT  94040.0 184740.0 94745.0 186085.0 ;
      RECT  94040.0 187430.0 94745.0 186085.0 ;
      RECT  94040.0 187430.0 94745.0 188775.0 ;
      RECT  94040.0 190120.0 94745.0 188775.0 ;
      RECT  94040.0 190120.0 94745.0 191465.0 ;
      RECT  94040.0 192810.0 94745.0 191465.0 ;
      RECT  94040.0 192810.0 94745.0 194155.0 ;
      RECT  94040.0 195500.0 94745.0 194155.0 ;
      RECT  94040.0 195500.0 94745.0 196845.0 ;
      RECT  94040.0 198190.0 94745.0 196845.0 ;
      RECT  94040.0 198190.0 94745.0 199535.0 ;
      RECT  94040.0 200880.0 94745.0 199535.0 ;
      RECT  94040.0 200880.0 94745.0 202225.0 ;
      RECT  94040.0 203570.0 94745.0 202225.0 ;
      RECT  94040.0 203570.0 94745.0 204915.0 ;
      RECT  94040.0 206260.0 94745.0 204915.0 ;
      RECT  94745.0 34100.0 95450.0 35445.0 ;
      RECT  94745.0 36790.0 95450.0 35445.0 ;
      RECT  94745.0 36790.0 95450.0 38135.0 ;
      RECT  94745.0 39480.0 95450.0 38135.0 ;
      RECT  94745.0 39480.0 95450.0 40825.0 ;
      RECT  94745.0 42170.0 95450.0 40825.0 ;
      RECT  94745.0 42170.0 95450.0 43515.0 ;
      RECT  94745.0 44860.0 95450.0 43515.0 ;
      RECT  94745.0 44860.0 95450.0 46205.0 ;
      RECT  94745.0 47550.0 95450.0 46205.0 ;
      RECT  94745.0 47550.0 95450.0 48895.0 ;
      RECT  94745.0 50240.0 95450.0 48895.0 ;
      RECT  94745.0 50240.0 95450.0 51585.0 ;
      RECT  94745.0 52930.0 95450.0 51585.0 ;
      RECT  94745.0 52930.0 95450.0 54275.0 ;
      RECT  94745.0 55620.0 95450.0 54275.0 ;
      RECT  94745.0 55620.0 95450.0 56965.0 ;
      RECT  94745.0 58310.0 95450.0 56965.0 ;
      RECT  94745.0 58310.0 95450.0 59655.0 ;
      RECT  94745.0 61000.0 95450.0 59655.0 ;
      RECT  94745.0 61000.0 95450.0 62345.0 ;
      RECT  94745.0 63690.0 95450.0 62345.0 ;
      RECT  94745.0 63690.0 95450.0 65035.0 ;
      RECT  94745.0 66380.0 95450.0 65035.0 ;
      RECT  94745.0 66380.0 95450.0 67725.0 ;
      RECT  94745.0 69070.0 95450.0 67725.0 ;
      RECT  94745.0 69070.0 95450.0 70415.0 ;
      RECT  94745.0 71760.0 95450.0 70415.0 ;
      RECT  94745.0 71760.0 95450.0 73105.0 ;
      RECT  94745.0 74450.0 95450.0 73105.0 ;
      RECT  94745.0 74450.0 95450.0 75795.0 ;
      RECT  94745.0 77140.0 95450.0 75795.0 ;
      RECT  94745.0 77140.0 95450.0 78485.0 ;
      RECT  94745.0 79830.0 95450.0 78485.0 ;
      RECT  94745.0 79830.0 95450.0 81175.0 ;
      RECT  94745.0 82520.0 95450.0 81175.0 ;
      RECT  94745.0 82520.0 95450.0 83865.0 ;
      RECT  94745.0 85210.0 95450.0 83865.0 ;
      RECT  94745.0 85210.0 95450.0 86555.0 ;
      RECT  94745.0 87900.0 95450.0 86555.0 ;
      RECT  94745.0 87900.0 95450.0 89245.0 ;
      RECT  94745.0 90590.0 95450.0 89245.0 ;
      RECT  94745.0 90590.0 95450.0 91935.0 ;
      RECT  94745.0 93280.0 95450.0 91935.0 ;
      RECT  94745.0 93280.0 95450.0 94625.0 ;
      RECT  94745.0 95970.0 95450.0 94625.0 ;
      RECT  94745.0 95970.0 95450.0 97315.0 ;
      RECT  94745.0 98660.0 95450.0 97315.0 ;
      RECT  94745.0 98660.0 95450.0 100005.0 ;
      RECT  94745.0 101350.0 95450.0 100005.0 ;
      RECT  94745.0 101350.0 95450.0 102695.0 ;
      RECT  94745.0 104040.0 95450.0 102695.0 ;
      RECT  94745.0 104040.0 95450.0 105385.0 ;
      RECT  94745.0 106730.0 95450.0 105385.0 ;
      RECT  94745.0 106730.0 95450.0 108075.0 ;
      RECT  94745.0 109420.0 95450.0 108075.0 ;
      RECT  94745.0 109420.0 95450.0 110765.0 ;
      RECT  94745.0 112110.0 95450.0 110765.0 ;
      RECT  94745.0 112110.0 95450.0 113455.0 ;
      RECT  94745.0 114800.0 95450.0 113455.0 ;
      RECT  94745.0 114800.0 95450.0 116145.0 ;
      RECT  94745.0 117490.0 95450.0 116145.0 ;
      RECT  94745.0 117490.0 95450.0 118835.0 ;
      RECT  94745.0 120180.0 95450.0 118835.0 ;
      RECT  94745.0 120180.0 95450.0 121525.0 ;
      RECT  94745.0 122870.0 95450.0 121525.0 ;
      RECT  94745.0 122870.0 95450.0 124215.0 ;
      RECT  94745.0 125560.0 95450.0 124215.0 ;
      RECT  94745.0 125560.0 95450.0 126905.0 ;
      RECT  94745.0 128250.0 95450.0 126905.0 ;
      RECT  94745.0 128250.0 95450.0 129595.0 ;
      RECT  94745.0 130940.0 95450.0 129595.0 ;
      RECT  94745.0 130940.0 95450.0 132285.0 ;
      RECT  94745.0 133630.0 95450.0 132285.0 ;
      RECT  94745.0 133630.0 95450.0 134975.0 ;
      RECT  94745.0 136320.0 95450.0 134975.0 ;
      RECT  94745.0 136320.0 95450.0 137665.0 ;
      RECT  94745.0 139010.0 95450.0 137665.0 ;
      RECT  94745.0 139010.0 95450.0 140355.0 ;
      RECT  94745.0 141700.0 95450.0 140355.0 ;
      RECT  94745.0 141700.0 95450.0 143045.0 ;
      RECT  94745.0 144390.0 95450.0 143045.0 ;
      RECT  94745.0 144390.0 95450.0 145735.0 ;
      RECT  94745.0 147080.0 95450.0 145735.0 ;
      RECT  94745.0 147080.0 95450.0 148425.0 ;
      RECT  94745.0 149770.0 95450.0 148425.0 ;
      RECT  94745.0 149770.0 95450.0 151115.0 ;
      RECT  94745.0 152460.0 95450.0 151115.0 ;
      RECT  94745.0 152460.0 95450.0 153805.0 ;
      RECT  94745.0 155150.0 95450.0 153805.0 ;
      RECT  94745.0 155150.0 95450.0 156495.0 ;
      RECT  94745.0 157840.0 95450.0 156495.0 ;
      RECT  94745.0 157840.0 95450.0 159185.0 ;
      RECT  94745.0 160530.0 95450.0 159185.0 ;
      RECT  94745.0 160530.0 95450.0 161875.0 ;
      RECT  94745.0 163220.0 95450.0 161875.0 ;
      RECT  94745.0 163220.0 95450.0 164565.0 ;
      RECT  94745.0 165910.0 95450.0 164565.0 ;
      RECT  94745.0 165910.0 95450.0 167255.0 ;
      RECT  94745.0 168600.0 95450.0 167255.0 ;
      RECT  94745.0 168600.0 95450.0 169945.0 ;
      RECT  94745.0 171290.0 95450.0 169945.0 ;
      RECT  94745.0 171290.0 95450.0 172635.0 ;
      RECT  94745.0 173980.0 95450.0 172635.0 ;
      RECT  94745.0 173980.0 95450.0 175325.0 ;
      RECT  94745.0 176670.0 95450.0 175325.0 ;
      RECT  94745.0 176670.0 95450.0 178015.0 ;
      RECT  94745.0 179360.0 95450.0 178015.0 ;
      RECT  94745.0 179360.0 95450.0 180705.0 ;
      RECT  94745.0 182050.0 95450.0 180705.0 ;
      RECT  94745.0 182050.0 95450.0 183395.0 ;
      RECT  94745.0 184740.0 95450.0 183395.0 ;
      RECT  94745.0 184740.0 95450.0 186085.0 ;
      RECT  94745.0 187430.0 95450.0 186085.0 ;
      RECT  94745.0 187430.0 95450.0 188775.0 ;
      RECT  94745.0 190120.0 95450.0 188775.0 ;
      RECT  94745.0 190120.0 95450.0 191465.0 ;
      RECT  94745.0 192810.0 95450.0 191465.0 ;
      RECT  94745.0 192810.0 95450.0 194155.0 ;
      RECT  94745.0 195500.0 95450.0 194155.0 ;
      RECT  94745.0 195500.0 95450.0 196845.0 ;
      RECT  94745.0 198190.0 95450.0 196845.0 ;
      RECT  94745.0 198190.0 95450.0 199535.0 ;
      RECT  94745.0 200880.0 95450.0 199535.0 ;
      RECT  94745.0 200880.0 95450.0 202225.0 ;
      RECT  94745.0 203570.0 95450.0 202225.0 ;
      RECT  94745.0 203570.0 95450.0 204915.0 ;
      RECT  94745.0 206260.0 95450.0 204915.0 ;
      RECT  95450.0 34100.0 96155.0 35445.0 ;
      RECT  95450.0 36790.0 96155.0 35445.0 ;
      RECT  95450.0 36790.0 96155.0 38135.0 ;
      RECT  95450.0 39480.0 96155.0 38135.0 ;
      RECT  95450.0 39480.0 96155.0 40825.0 ;
      RECT  95450.0 42170.0 96155.0 40825.0 ;
      RECT  95450.0 42170.0 96155.0 43515.0 ;
      RECT  95450.0 44860.0 96155.0 43515.0 ;
      RECT  95450.0 44860.0 96155.0 46205.0 ;
      RECT  95450.0 47550.0 96155.0 46205.0 ;
      RECT  95450.0 47550.0 96155.0 48895.0 ;
      RECT  95450.0 50240.0 96155.0 48895.0 ;
      RECT  95450.0 50240.0 96155.0 51585.0 ;
      RECT  95450.0 52930.0 96155.0 51585.0 ;
      RECT  95450.0 52930.0 96155.0 54275.0 ;
      RECT  95450.0 55620.0 96155.0 54275.0 ;
      RECT  95450.0 55620.0 96155.0 56965.0 ;
      RECT  95450.0 58310.0 96155.0 56965.0 ;
      RECT  95450.0 58310.0 96155.0 59655.0 ;
      RECT  95450.0 61000.0 96155.0 59655.0 ;
      RECT  95450.0 61000.0 96155.0 62345.0 ;
      RECT  95450.0 63690.0 96155.0 62345.0 ;
      RECT  95450.0 63690.0 96155.0 65035.0 ;
      RECT  95450.0 66380.0 96155.0 65035.0 ;
      RECT  95450.0 66380.0 96155.0 67725.0 ;
      RECT  95450.0 69070.0 96155.0 67725.0 ;
      RECT  95450.0 69070.0 96155.0 70415.0 ;
      RECT  95450.0 71760.0 96155.0 70415.0 ;
      RECT  95450.0 71760.0 96155.0 73105.0 ;
      RECT  95450.0 74450.0 96155.0 73105.0 ;
      RECT  95450.0 74450.0 96155.0 75795.0 ;
      RECT  95450.0 77140.0 96155.0 75795.0 ;
      RECT  95450.0 77140.0 96155.0 78485.0 ;
      RECT  95450.0 79830.0 96155.0 78485.0 ;
      RECT  95450.0 79830.0 96155.0 81175.0 ;
      RECT  95450.0 82520.0 96155.0 81175.0 ;
      RECT  95450.0 82520.0 96155.0 83865.0 ;
      RECT  95450.0 85210.0 96155.0 83865.0 ;
      RECT  95450.0 85210.0 96155.0 86555.0 ;
      RECT  95450.0 87900.0 96155.0 86555.0 ;
      RECT  95450.0 87900.0 96155.0 89245.0 ;
      RECT  95450.0 90590.0 96155.0 89245.0 ;
      RECT  95450.0 90590.0 96155.0 91935.0 ;
      RECT  95450.0 93280.0 96155.0 91935.0 ;
      RECT  95450.0 93280.0 96155.0 94625.0 ;
      RECT  95450.0 95970.0 96155.0 94625.0 ;
      RECT  95450.0 95970.0 96155.0 97315.0 ;
      RECT  95450.0 98660.0 96155.0 97315.0 ;
      RECT  95450.0 98660.0 96155.0 100005.0 ;
      RECT  95450.0 101350.0 96155.0 100005.0 ;
      RECT  95450.0 101350.0 96155.0 102695.0 ;
      RECT  95450.0 104040.0 96155.0 102695.0 ;
      RECT  95450.0 104040.0 96155.0 105385.0 ;
      RECT  95450.0 106730.0 96155.0 105385.0 ;
      RECT  95450.0 106730.0 96155.0 108075.0 ;
      RECT  95450.0 109420.0 96155.0 108075.0 ;
      RECT  95450.0 109420.0 96155.0 110765.0 ;
      RECT  95450.0 112110.0 96155.0 110765.0 ;
      RECT  95450.0 112110.0 96155.0 113455.0 ;
      RECT  95450.0 114800.0 96155.0 113455.0 ;
      RECT  95450.0 114800.0 96155.0 116145.0 ;
      RECT  95450.0 117490.0 96155.0 116145.0 ;
      RECT  95450.0 117490.0 96155.0 118835.0 ;
      RECT  95450.0 120180.0 96155.0 118835.0 ;
      RECT  95450.0 120180.0 96155.0 121525.0 ;
      RECT  95450.0 122870.0 96155.0 121525.0 ;
      RECT  95450.0 122870.0 96155.0 124215.0 ;
      RECT  95450.0 125560.0 96155.0 124215.0 ;
      RECT  95450.0 125560.0 96155.0 126905.0 ;
      RECT  95450.0 128250.0 96155.0 126905.0 ;
      RECT  95450.0 128250.0 96155.0 129595.0 ;
      RECT  95450.0 130940.0 96155.0 129595.0 ;
      RECT  95450.0 130940.0 96155.0 132285.0 ;
      RECT  95450.0 133630.0 96155.0 132285.0 ;
      RECT  95450.0 133630.0 96155.0 134975.0 ;
      RECT  95450.0 136320.0 96155.0 134975.0 ;
      RECT  95450.0 136320.0 96155.0 137665.0 ;
      RECT  95450.0 139010.0 96155.0 137665.0 ;
      RECT  95450.0 139010.0 96155.0 140355.0 ;
      RECT  95450.0 141700.0 96155.0 140355.0 ;
      RECT  95450.0 141700.0 96155.0 143045.0 ;
      RECT  95450.0 144390.0 96155.0 143045.0 ;
      RECT  95450.0 144390.0 96155.0 145735.0 ;
      RECT  95450.0 147080.0 96155.0 145735.0 ;
      RECT  95450.0 147080.0 96155.0 148425.0 ;
      RECT  95450.0 149770.0 96155.0 148425.0 ;
      RECT  95450.0 149770.0 96155.0 151115.0 ;
      RECT  95450.0 152460.0 96155.0 151115.0 ;
      RECT  95450.0 152460.0 96155.0 153805.0 ;
      RECT  95450.0 155150.0 96155.0 153805.0 ;
      RECT  95450.0 155150.0 96155.0 156495.0 ;
      RECT  95450.0 157840.0 96155.0 156495.0 ;
      RECT  95450.0 157840.0 96155.0 159185.0 ;
      RECT  95450.0 160530.0 96155.0 159185.0 ;
      RECT  95450.0 160530.0 96155.0 161875.0 ;
      RECT  95450.0 163220.0 96155.0 161875.0 ;
      RECT  95450.0 163220.0 96155.0 164565.0 ;
      RECT  95450.0 165910.0 96155.0 164565.0 ;
      RECT  95450.0 165910.0 96155.0 167255.0 ;
      RECT  95450.0 168600.0 96155.0 167255.0 ;
      RECT  95450.0 168600.0 96155.0 169945.0 ;
      RECT  95450.0 171290.0 96155.0 169945.0 ;
      RECT  95450.0 171290.0 96155.0 172635.0 ;
      RECT  95450.0 173980.0 96155.0 172635.0 ;
      RECT  95450.0 173980.0 96155.0 175325.0 ;
      RECT  95450.0 176670.0 96155.0 175325.0 ;
      RECT  95450.0 176670.0 96155.0 178015.0 ;
      RECT  95450.0 179360.0 96155.0 178015.0 ;
      RECT  95450.0 179360.0 96155.0 180705.0 ;
      RECT  95450.0 182050.0 96155.0 180705.0 ;
      RECT  95450.0 182050.0 96155.0 183395.0 ;
      RECT  95450.0 184740.0 96155.0 183395.0 ;
      RECT  95450.0 184740.0 96155.0 186085.0 ;
      RECT  95450.0 187430.0 96155.0 186085.0 ;
      RECT  95450.0 187430.0 96155.0 188775.0 ;
      RECT  95450.0 190120.0 96155.0 188775.0 ;
      RECT  95450.0 190120.0 96155.0 191465.0 ;
      RECT  95450.0 192810.0 96155.0 191465.0 ;
      RECT  95450.0 192810.0 96155.0 194155.0 ;
      RECT  95450.0 195500.0 96155.0 194155.0 ;
      RECT  95450.0 195500.0 96155.0 196845.0 ;
      RECT  95450.0 198190.0 96155.0 196845.0 ;
      RECT  95450.0 198190.0 96155.0 199535.0 ;
      RECT  95450.0 200880.0 96155.0 199535.0 ;
      RECT  95450.0 200880.0 96155.0 202225.0 ;
      RECT  95450.0 203570.0 96155.0 202225.0 ;
      RECT  95450.0 203570.0 96155.0 204915.0 ;
      RECT  95450.0 206260.0 96155.0 204915.0 ;
      RECT  96155.0 34100.0 96860.0 35445.0 ;
      RECT  96155.0 36790.0 96860.0 35445.0 ;
      RECT  96155.0 36790.0 96860.0 38135.0 ;
      RECT  96155.0 39480.0 96860.0 38135.0 ;
      RECT  96155.0 39480.0 96860.0 40825.0 ;
      RECT  96155.0 42170.0 96860.0 40825.0 ;
      RECT  96155.0 42170.0 96860.0 43515.0 ;
      RECT  96155.0 44860.0 96860.0 43515.0 ;
      RECT  96155.0 44860.0 96860.0 46205.0 ;
      RECT  96155.0 47550.0 96860.0 46205.0 ;
      RECT  96155.0 47550.0 96860.0 48895.0 ;
      RECT  96155.0 50240.0 96860.0 48895.0 ;
      RECT  96155.0 50240.0 96860.0 51585.0 ;
      RECT  96155.0 52930.0 96860.0 51585.0 ;
      RECT  96155.0 52930.0 96860.0 54275.0 ;
      RECT  96155.0 55620.0 96860.0 54275.0 ;
      RECT  96155.0 55620.0 96860.0 56965.0 ;
      RECT  96155.0 58310.0 96860.0 56965.0 ;
      RECT  96155.0 58310.0 96860.0 59655.0 ;
      RECT  96155.0 61000.0 96860.0 59655.0 ;
      RECT  96155.0 61000.0 96860.0 62345.0 ;
      RECT  96155.0 63690.0 96860.0 62345.0 ;
      RECT  96155.0 63690.0 96860.0 65035.0 ;
      RECT  96155.0 66380.0 96860.0 65035.0 ;
      RECT  96155.0 66380.0 96860.0 67725.0 ;
      RECT  96155.0 69070.0 96860.0 67725.0 ;
      RECT  96155.0 69070.0 96860.0 70415.0 ;
      RECT  96155.0 71760.0 96860.0 70415.0 ;
      RECT  96155.0 71760.0 96860.0 73105.0 ;
      RECT  96155.0 74450.0 96860.0 73105.0 ;
      RECT  96155.0 74450.0 96860.0 75795.0 ;
      RECT  96155.0 77140.0 96860.0 75795.0 ;
      RECT  96155.0 77140.0 96860.0 78485.0 ;
      RECT  96155.0 79830.0 96860.0 78485.0 ;
      RECT  96155.0 79830.0 96860.0 81175.0 ;
      RECT  96155.0 82520.0 96860.0 81175.0 ;
      RECT  96155.0 82520.0 96860.0 83865.0 ;
      RECT  96155.0 85210.0 96860.0 83865.0 ;
      RECT  96155.0 85210.0 96860.0 86555.0 ;
      RECT  96155.0 87900.0 96860.0 86555.0 ;
      RECT  96155.0 87900.0 96860.0 89245.0 ;
      RECT  96155.0 90590.0 96860.0 89245.0 ;
      RECT  96155.0 90590.0 96860.0 91935.0 ;
      RECT  96155.0 93280.0 96860.0 91935.0 ;
      RECT  96155.0 93280.0 96860.0 94625.0 ;
      RECT  96155.0 95970.0 96860.0 94625.0 ;
      RECT  96155.0 95970.0 96860.0 97315.0 ;
      RECT  96155.0 98660.0 96860.0 97315.0 ;
      RECT  96155.0 98660.0 96860.0 100005.0 ;
      RECT  96155.0 101350.0 96860.0 100005.0 ;
      RECT  96155.0 101350.0 96860.0 102695.0 ;
      RECT  96155.0 104040.0 96860.0 102695.0 ;
      RECT  96155.0 104040.0 96860.0 105385.0 ;
      RECT  96155.0 106730.0 96860.0 105385.0 ;
      RECT  96155.0 106730.0 96860.0 108075.0 ;
      RECT  96155.0 109420.0 96860.0 108075.0 ;
      RECT  96155.0 109420.0 96860.0 110765.0 ;
      RECT  96155.0 112110.0 96860.0 110765.0 ;
      RECT  96155.0 112110.0 96860.0 113455.0 ;
      RECT  96155.0 114800.0 96860.0 113455.0 ;
      RECT  96155.0 114800.0 96860.0 116145.0 ;
      RECT  96155.0 117490.0 96860.0 116145.0 ;
      RECT  96155.0 117490.0 96860.0 118835.0 ;
      RECT  96155.0 120180.0 96860.0 118835.0 ;
      RECT  96155.0 120180.0 96860.0 121525.0 ;
      RECT  96155.0 122870.0 96860.0 121525.0 ;
      RECT  96155.0 122870.0 96860.0 124215.0 ;
      RECT  96155.0 125560.0 96860.0 124215.0 ;
      RECT  96155.0 125560.0 96860.0 126905.0 ;
      RECT  96155.0 128250.0 96860.0 126905.0 ;
      RECT  96155.0 128250.0 96860.0 129595.0 ;
      RECT  96155.0 130940.0 96860.0 129595.0 ;
      RECT  96155.0 130940.0 96860.0 132285.0 ;
      RECT  96155.0 133630.0 96860.0 132285.0 ;
      RECT  96155.0 133630.0 96860.0 134975.0 ;
      RECT  96155.0 136320.0 96860.0 134975.0 ;
      RECT  96155.0 136320.0 96860.0 137665.0 ;
      RECT  96155.0 139010.0 96860.0 137665.0 ;
      RECT  96155.0 139010.0 96860.0 140355.0 ;
      RECT  96155.0 141700.0 96860.0 140355.0 ;
      RECT  96155.0 141700.0 96860.0 143045.0 ;
      RECT  96155.0 144390.0 96860.0 143045.0 ;
      RECT  96155.0 144390.0 96860.0 145735.0 ;
      RECT  96155.0 147080.0 96860.0 145735.0 ;
      RECT  96155.0 147080.0 96860.0 148425.0 ;
      RECT  96155.0 149770.0 96860.0 148425.0 ;
      RECT  96155.0 149770.0 96860.0 151115.0 ;
      RECT  96155.0 152460.0 96860.0 151115.0 ;
      RECT  96155.0 152460.0 96860.0 153805.0 ;
      RECT  96155.0 155150.0 96860.0 153805.0 ;
      RECT  96155.0 155150.0 96860.0 156495.0 ;
      RECT  96155.0 157840.0 96860.0 156495.0 ;
      RECT  96155.0 157840.0 96860.0 159185.0 ;
      RECT  96155.0 160530.0 96860.0 159185.0 ;
      RECT  96155.0 160530.0 96860.0 161875.0 ;
      RECT  96155.0 163220.0 96860.0 161875.0 ;
      RECT  96155.0 163220.0 96860.0 164565.0 ;
      RECT  96155.0 165910.0 96860.0 164565.0 ;
      RECT  96155.0 165910.0 96860.0 167255.0 ;
      RECT  96155.0 168600.0 96860.0 167255.0 ;
      RECT  96155.0 168600.0 96860.0 169945.0 ;
      RECT  96155.0 171290.0 96860.0 169945.0 ;
      RECT  96155.0 171290.0 96860.0 172635.0 ;
      RECT  96155.0 173980.0 96860.0 172635.0 ;
      RECT  96155.0 173980.0 96860.0 175325.0 ;
      RECT  96155.0 176670.0 96860.0 175325.0 ;
      RECT  96155.0 176670.0 96860.0 178015.0 ;
      RECT  96155.0 179360.0 96860.0 178015.0 ;
      RECT  96155.0 179360.0 96860.0 180705.0 ;
      RECT  96155.0 182050.0 96860.0 180705.0 ;
      RECT  96155.0 182050.0 96860.0 183395.0 ;
      RECT  96155.0 184740.0 96860.0 183395.0 ;
      RECT  96155.0 184740.0 96860.0 186085.0 ;
      RECT  96155.0 187430.0 96860.0 186085.0 ;
      RECT  96155.0 187430.0 96860.0 188775.0 ;
      RECT  96155.0 190120.0 96860.0 188775.0 ;
      RECT  96155.0 190120.0 96860.0 191465.0 ;
      RECT  96155.0 192810.0 96860.0 191465.0 ;
      RECT  96155.0 192810.0 96860.0 194155.0 ;
      RECT  96155.0 195500.0 96860.0 194155.0 ;
      RECT  96155.0 195500.0 96860.0 196845.0 ;
      RECT  96155.0 198190.0 96860.0 196845.0 ;
      RECT  96155.0 198190.0 96860.0 199535.0 ;
      RECT  96155.0 200880.0 96860.0 199535.0 ;
      RECT  96155.0 200880.0 96860.0 202225.0 ;
      RECT  96155.0 203570.0 96860.0 202225.0 ;
      RECT  96155.0 203570.0 96860.0 204915.0 ;
      RECT  96155.0 206260.0 96860.0 204915.0 ;
      RECT  96860.0 34100.0 97565.0 35445.0 ;
      RECT  96860.0 36790.0 97565.0 35445.0 ;
      RECT  96860.0 36790.0 97565.0 38135.0 ;
      RECT  96860.0 39480.0 97565.0 38135.0 ;
      RECT  96860.0 39480.0 97565.0 40825.0 ;
      RECT  96860.0 42170.0 97565.0 40825.0 ;
      RECT  96860.0 42170.0 97565.0 43515.0 ;
      RECT  96860.0 44860.0 97565.0 43515.0 ;
      RECT  96860.0 44860.0 97565.0 46205.0 ;
      RECT  96860.0 47550.0 97565.0 46205.0 ;
      RECT  96860.0 47550.0 97565.0 48895.0 ;
      RECT  96860.0 50240.0 97565.0 48895.0 ;
      RECT  96860.0 50240.0 97565.0 51585.0 ;
      RECT  96860.0 52930.0 97565.0 51585.0 ;
      RECT  96860.0 52930.0 97565.0 54275.0 ;
      RECT  96860.0 55620.0 97565.0 54275.0 ;
      RECT  96860.0 55620.0 97565.0 56965.0 ;
      RECT  96860.0 58310.0 97565.0 56965.0 ;
      RECT  96860.0 58310.0 97565.0 59655.0 ;
      RECT  96860.0 61000.0 97565.0 59655.0 ;
      RECT  96860.0 61000.0 97565.0 62345.0 ;
      RECT  96860.0 63690.0 97565.0 62345.0 ;
      RECT  96860.0 63690.0 97565.0 65035.0 ;
      RECT  96860.0 66380.0 97565.0 65035.0 ;
      RECT  96860.0 66380.0 97565.0 67725.0 ;
      RECT  96860.0 69070.0 97565.0 67725.0 ;
      RECT  96860.0 69070.0 97565.0 70415.0 ;
      RECT  96860.0 71760.0 97565.0 70415.0 ;
      RECT  96860.0 71760.0 97565.0 73105.0 ;
      RECT  96860.0 74450.0 97565.0 73105.0 ;
      RECT  96860.0 74450.0 97565.0 75795.0 ;
      RECT  96860.0 77140.0 97565.0 75795.0 ;
      RECT  96860.0 77140.0 97565.0 78485.0 ;
      RECT  96860.0 79830.0 97565.0 78485.0 ;
      RECT  96860.0 79830.0 97565.0 81175.0 ;
      RECT  96860.0 82520.0 97565.0 81175.0 ;
      RECT  96860.0 82520.0 97565.0 83865.0 ;
      RECT  96860.0 85210.0 97565.0 83865.0 ;
      RECT  96860.0 85210.0 97565.0 86555.0 ;
      RECT  96860.0 87900.0 97565.0 86555.0 ;
      RECT  96860.0 87900.0 97565.0 89245.0 ;
      RECT  96860.0 90590.0 97565.0 89245.0 ;
      RECT  96860.0 90590.0 97565.0 91935.0 ;
      RECT  96860.0 93280.0 97565.0 91935.0 ;
      RECT  96860.0 93280.0 97565.0 94625.0 ;
      RECT  96860.0 95970.0 97565.0 94625.0 ;
      RECT  96860.0 95970.0 97565.0 97315.0 ;
      RECT  96860.0 98660.0 97565.0 97315.0 ;
      RECT  96860.0 98660.0 97565.0 100005.0 ;
      RECT  96860.0 101350.0 97565.0 100005.0 ;
      RECT  96860.0 101350.0 97565.0 102695.0 ;
      RECT  96860.0 104040.0 97565.0 102695.0 ;
      RECT  96860.0 104040.0 97565.0 105385.0 ;
      RECT  96860.0 106730.0 97565.0 105385.0 ;
      RECT  96860.0 106730.0 97565.0 108075.0 ;
      RECT  96860.0 109420.0 97565.0 108075.0 ;
      RECT  96860.0 109420.0 97565.0 110765.0 ;
      RECT  96860.0 112110.0 97565.0 110765.0 ;
      RECT  96860.0 112110.0 97565.0 113455.0 ;
      RECT  96860.0 114800.0 97565.0 113455.0 ;
      RECT  96860.0 114800.0 97565.0 116145.0 ;
      RECT  96860.0 117490.0 97565.0 116145.0 ;
      RECT  96860.0 117490.0 97565.0 118835.0 ;
      RECT  96860.0 120180.0 97565.0 118835.0 ;
      RECT  96860.0 120180.0 97565.0 121525.0 ;
      RECT  96860.0 122870.0 97565.0 121525.0 ;
      RECT  96860.0 122870.0 97565.0 124215.0 ;
      RECT  96860.0 125560.0 97565.0 124215.0 ;
      RECT  96860.0 125560.0 97565.0 126905.0 ;
      RECT  96860.0 128250.0 97565.0 126905.0 ;
      RECT  96860.0 128250.0 97565.0 129595.0 ;
      RECT  96860.0 130940.0 97565.0 129595.0 ;
      RECT  96860.0 130940.0 97565.0 132285.0 ;
      RECT  96860.0 133630.0 97565.0 132285.0 ;
      RECT  96860.0 133630.0 97565.0 134975.0 ;
      RECT  96860.0 136320.0 97565.0 134975.0 ;
      RECT  96860.0 136320.0 97565.0 137665.0 ;
      RECT  96860.0 139010.0 97565.0 137665.0 ;
      RECT  96860.0 139010.0 97565.0 140355.0 ;
      RECT  96860.0 141700.0 97565.0 140355.0 ;
      RECT  96860.0 141700.0 97565.0 143045.0 ;
      RECT  96860.0 144390.0 97565.0 143045.0 ;
      RECT  96860.0 144390.0 97565.0 145735.0 ;
      RECT  96860.0 147080.0 97565.0 145735.0 ;
      RECT  96860.0 147080.0 97565.0 148425.0 ;
      RECT  96860.0 149770.0 97565.0 148425.0 ;
      RECT  96860.0 149770.0 97565.0 151115.0 ;
      RECT  96860.0 152460.0 97565.0 151115.0 ;
      RECT  96860.0 152460.0 97565.0 153805.0 ;
      RECT  96860.0 155150.0 97565.0 153805.0 ;
      RECT  96860.0 155150.0 97565.0 156495.0 ;
      RECT  96860.0 157840.0 97565.0 156495.0 ;
      RECT  96860.0 157840.0 97565.0 159185.0 ;
      RECT  96860.0 160530.0 97565.0 159185.0 ;
      RECT  96860.0 160530.0 97565.0 161875.0 ;
      RECT  96860.0 163220.0 97565.0 161875.0 ;
      RECT  96860.0 163220.0 97565.0 164565.0 ;
      RECT  96860.0 165910.0 97565.0 164565.0 ;
      RECT  96860.0 165910.0 97565.0 167255.0 ;
      RECT  96860.0 168600.0 97565.0 167255.0 ;
      RECT  96860.0 168600.0 97565.0 169945.0 ;
      RECT  96860.0 171290.0 97565.0 169945.0 ;
      RECT  96860.0 171290.0 97565.0 172635.0 ;
      RECT  96860.0 173980.0 97565.0 172635.0 ;
      RECT  96860.0 173980.0 97565.0 175325.0 ;
      RECT  96860.0 176670.0 97565.0 175325.0 ;
      RECT  96860.0 176670.0 97565.0 178015.0 ;
      RECT  96860.0 179360.0 97565.0 178015.0 ;
      RECT  96860.0 179360.0 97565.0 180705.0 ;
      RECT  96860.0 182050.0 97565.0 180705.0 ;
      RECT  96860.0 182050.0 97565.0 183395.0 ;
      RECT  96860.0 184740.0 97565.0 183395.0 ;
      RECT  96860.0 184740.0 97565.0 186085.0 ;
      RECT  96860.0 187430.0 97565.0 186085.0 ;
      RECT  96860.0 187430.0 97565.0 188775.0 ;
      RECT  96860.0 190120.0 97565.0 188775.0 ;
      RECT  96860.0 190120.0 97565.0 191465.0 ;
      RECT  96860.0 192810.0 97565.0 191465.0 ;
      RECT  96860.0 192810.0 97565.0 194155.0 ;
      RECT  96860.0 195500.0 97565.0 194155.0 ;
      RECT  96860.0 195500.0 97565.0 196845.0 ;
      RECT  96860.0 198190.0 97565.0 196845.0 ;
      RECT  96860.0 198190.0 97565.0 199535.0 ;
      RECT  96860.0 200880.0 97565.0 199535.0 ;
      RECT  96860.0 200880.0 97565.0 202225.0 ;
      RECT  96860.0 203570.0 97565.0 202225.0 ;
      RECT  96860.0 203570.0 97565.0 204915.0 ;
      RECT  96860.0 206260.0 97565.0 204915.0 ;
      RECT  97565.0 34100.0 98270.0 35445.0 ;
      RECT  97565.0 36790.0 98270.0 35445.0 ;
      RECT  97565.0 36790.0 98270.0 38135.0 ;
      RECT  97565.0 39480.0 98270.0 38135.0 ;
      RECT  97565.0 39480.0 98270.0 40825.0 ;
      RECT  97565.0 42170.0 98270.0 40825.0 ;
      RECT  97565.0 42170.0 98270.0 43515.0 ;
      RECT  97565.0 44860.0 98270.0 43515.0 ;
      RECT  97565.0 44860.0 98270.0 46205.0 ;
      RECT  97565.0 47550.0 98270.0 46205.0 ;
      RECT  97565.0 47550.0 98270.0 48895.0 ;
      RECT  97565.0 50240.0 98270.0 48895.0 ;
      RECT  97565.0 50240.0 98270.0 51585.0 ;
      RECT  97565.0 52930.0 98270.0 51585.0 ;
      RECT  97565.0 52930.0 98270.0 54275.0 ;
      RECT  97565.0 55620.0 98270.0 54275.0 ;
      RECT  97565.0 55620.0 98270.0 56965.0 ;
      RECT  97565.0 58310.0 98270.0 56965.0 ;
      RECT  97565.0 58310.0 98270.0 59655.0 ;
      RECT  97565.0 61000.0 98270.0 59655.0 ;
      RECT  97565.0 61000.0 98270.0 62345.0 ;
      RECT  97565.0 63690.0 98270.0 62345.0 ;
      RECT  97565.0 63690.0 98270.0 65035.0 ;
      RECT  97565.0 66380.0 98270.0 65035.0 ;
      RECT  97565.0 66380.0 98270.0 67725.0 ;
      RECT  97565.0 69070.0 98270.0 67725.0 ;
      RECT  97565.0 69070.0 98270.0 70415.0 ;
      RECT  97565.0 71760.0 98270.0 70415.0 ;
      RECT  97565.0 71760.0 98270.0 73105.0 ;
      RECT  97565.0 74450.0 98270.0 73105.0 ;
      RECT  97565.0 74450.0 98270.0 75795.0 ;
      RECT  97565.0 77140.0 98270.0 75795.0 ;
      RECT  97565.0 77140.0 98270.0 78485.0 ;
      RECT  97565.0 79830.0 98270.0 78485.0 ;
      RECT  97565.0 79830.0 98270.0 81175.0 ;
      RECT  97565.0 82520.0 98270.0 81175.0 ;
      RECT  97565.0 82520.0 98270.0 83865.0 ;
      RECT  97565.0 85210.0 98270.0 83865.0 ;
      RECT  97565.0 85210.0 98270.0 86555.0 ;
      RECT  97565.0 87900.0 98270.0 86555.0 ;
      RECT  97565.0 87900.0 98270.0 89245.0 ;
      RECT  97565.0 90590.0 98270.0 89245.0 ;
      RECT  97565.0 90590.0 98270.0 91935.0 ;
      RECT  97565.0 93280.0 98270.0 91935.0 ;
      RECT  97565.0 93280.0 98270.0 94625.0 ;
      RECT  97565.0 95970.0 98270.0 94625.0 ;
      RECT  97565.0 95970.0 98270.0 97315.0 ;
      RECT  97565.0 98660.0 98270.0 97315.0 ;
      RECT  97565.0 98660.0 98270.0 100005.0 ;
      RECT  97565.0 101350.0 98270.0 100005.0 ;
      RECT  97565.0 101350.0 98270.0 102695.0 ;
      RECT  97565.0 104040.0 98270.0 102695.0 ;
      RECT  97565.0 104040.0 98270.0 105385.0 ;
      RECT  97565.0 106730.0 98270.0 105385.0 ;
      RECT  97565.0 106730.0 98270.0 108075.0 ;
      RECT  97565.0 109420.0 98270.0 108075.0 ;
      RECT  97565.0 109420.0 98270.0 110765.0 ;
      RECT  97565.0 112110.0 98270.0 110765.0 ;
      RECT  97565.0 112110.0 98270.0 113455.0 ;
      RECT  97565.0 114800.0 98270.0 113455.0 ;
      RECT  97565.0 114800.0 98270.0 116145.0 ;
      RECT  97565.0 117490.0 98270.0 116145.0 ;
      RECT  97565.0 117490.0 98270.0 118835.0 ;
      RECT  97565.0 120180.0 98270.0 118835.0 ;
      RECT  97565.0 120180.0 98270.0 121525.0 ;
      RECT  97565.0 122870.0 98270.0 121525.0 ;
      RECT  97565.0 122870.0 98270.0 124215.0 ;
      RECT  97565.0 125560.0 98270.0 124215.0 ;
      RECT  97565.0 125560.0 98270.0 126905.0 ;
      RECT  97565.0 128250.0 98270.0 126905.0 ;
      RECT  97565.0 128250.0 98270.0 129595.0 ;
      RECT  97565.0 130940.0 98270.0 129595.0 ;
      RECT  97565.0 130940.0 98270.0 132285.0 ;
      RECT  97565.0 133630.0 98270.0 132285.0 ;
      RECT  97565.0 133630.0 98270.0 134975.0 ;
      RECT  97565.0 136320.0 98270.0 134975.0 ;
      RECT  97565.0 136320.0 98270.0 137665.0 ;
      RECT  97565.0 139010.0 98270.0 137665.0 ;
      RECT  97565.0 139010.0 98270.0 140355.0 ;
      RECT  97565.0 141700.0 98270.0 140355.0 ;
      RECT  97565.0 141700.0 98270.0 143045.0 ;
      RECT  97565.0 144390.0 98270.0 143045.0 ;
      RECT  97565.0 144390.0 98270.0 145735.0 ;
      RECT  97565.0 147080.0 98270.0 145735.0 ;
      RECT  97565.0 147080.0 98270.0 148425.0 ;
      RECT  97565.0 149770.0 98270.0 148425.0 ;
      RECT  97565.0 149770.0 98270.0 151115.0 ;
      RECT  97565.0 152460.0 98270.0 151115.0 ;
      RECT  97565.0 152460.0 98270.0 153805.0 ;
      RECT  97565.0 155150.0 98270.0 153805.0 ;
      RECT  97565.0 155150.0 98270.0 156495.0 ;
      RECT  97565.0 157840.0 98270.0 156495.0 ;
      RECT  97565.0 157840.0 98270.0 159185.0 ;
      RECT  97565.0 160530.0 98270.0 159185.0 ;
      RECT  97565.0 160530.0 98270.0 161875.0 ;
      RECT  97565.0 163220.0 98270.0 161875.0 ;
      RECT  97565.0 163220.0 98270.0 164565.0 ;
      RECT  97565.0 165910.0 98270.0 164565.0 ;
      RECT  97565.0 165910.0 98270.0 167255.0 ;
      RECT  97565.0 168600.0 98270.0 167255.0 ;
      RECT  97565.0 168600.0 98270.0 169945.0 ;
      RECT  97565.0 171290.0 98270.0 169945.0 ;
      RECT  97565.0 171290.0 98270.0 172635.0 ;
      RECT  97565.0 173980.0 98270.0 172635.0 ;
      RECT  97565.0 173980.0 98270.0 175325.0 ;
      RECT  97565.0 176670.0 98270.0 175325.0 ;
      RECT  97565.0 176670.0 98270.0 178015.0 ;
      RECT  97565.0 179360.0 98270.0 178015.0 ;
      RECT  97565.0 179360.0 98270.0 180705.0 ;
      RECT  97565.0 182050.0 98270.0 180705.0 ;
      RECT  97565.0 182050.0 98270.0 183395.0 ;
      RECT  97565.0 184740.0 98270.0 183395.0 ;
      RECT  97565.0 184740.0 98270.0 186085.0 ;
      RECT  97565.0 187430.0 98270.0 186085.0 ;
      RECT  97565.0 187430.0 98270.0 188775.0 ;
      RECT  97565.0 190120.0 98270.0 188775.0 ;
      RECT  97565.0 190120.0 98270.0 191465.0 ;
      RECT  97565.0 192810.0 98270.0 191465.0 ;
      RECT  97565.0 192810.0 98270.0 194155.0 ;
      RECT  97565.0 195500.0 98270.0 194155.0 ;
      RECT  97565.0 195500.0 98270.0 196845.0 ;
      RECT  97565.0 198190.0 98270.0 196845.0 ;
      RECT  97565.0 198190.0 98270.0 199535.0 ;
      RECT  97565.0 200880.0 98270.0 199535.0 ;
      RECT  97565.0 200880.0 98270.0 202225.0 ;
      RECT  97565.0 203570.0 98270.0 202225.0 ;
      RECT  97565.0 203570.0 98270.0 204915.0 ;
      RECT  97565.0 206260.0 98270.0 204915.0 ;
      RECT  98270.0 34100.0 98975.0 35445.0 ;
      RECT  98270.0 36790.0 98975.0 35445.0 ;
      RECT  98270.0 36790.0 98975.0 38135.0 ;
      RECT  98270.0 39480.0 98975.0 38135.0 ;
      RECT  98270.0 39480.0 98975.0 40825.0 ;
      RECT  98270.0 42170.0 98975.0 40825.0 ;
      RECT  98270.0 42170.0 98975.0 43515.0 ;
      RECT  98270.0 44860.0 98975.0 43515.0 ;
      RECT  98270.0 44860.0 98975.0 46205.0 ;
      RECT  98270.0 47550.0 98975.0 46205.0 ;
      RECT  98270.0 47550.0 98975.0 48895.0 ;
      RECT  98270.0 50240.0 98975.0 48895.0 ;
      RECT  98270.0 50240.0 98975.0 51585.0 ;
      RECT  98270.0 52930.0 98975.0 51585.0 ;
      RECT  98270.0 52930.0 98975.0 54275.0 ;
      RECT  98270.0 55620.0 98975.0 54275.0 ;
      RECT  98270.0 55620.0 98975.0 56965.0 ;
      RECT  98270.0 58310.0 98975.0 56965.0 ;
      RECT  98270.0 58310.0 98975.0 59655.0 ;
      RECT  98270.0 61000.0 98975.0 59655.0 ;
      RECT  98270.0 61000.0 98975.0 62345.0 ;
      RECT  98270.0 63690.0 98975.0 62345.0 ;
      RECT  98270.0 63690.0 98975.0 65035.0 ;
      RECT  98270.0 66380.0 98975.0 65035.0 ;
      RECT  98270.0 66380.0 98975.0 67725.0 ;
      RECT  98270.0 69070.0 98975.0 67725.0 ;
      RECT  98270.0 69070.0 98975.0 70415.0 ;
      RECT  98270.0 71760.0 98975.0 70415.0 ;
      RECT  98270.0 71760.0 98975.0 73105.0 ;
      RECT  98270.0 74450.0 98975.0 73105.0 ;
      RECT  98270.0 74450.0 98975.0 75795.0 ;
      RECT  98270.0 77140.0 98975.0 75795.0 ;
      RECT  98270.0 77140.0 98975.0 78485.0 ;
      RECT  98270.0 79830.0 98975.0 78485.0 ;
      RECT  98270.0 79830.0 98975.0 81175.0 ;
      RECT  98270.0 82520.0 98975.0 81175.0 ;
      RECT  98270.0 82520.0 98975.0 83865.0 ;
      RECT  98270.0 85210.0 98975.0 83865.0 ;
      RECT  98270.0 85210.0 98975.0 86555.0 ;
      RECT  98270.0 87900.0 98975.0 86555.0 ;
      RECT  98270.0 87900.0 98975.0 89245.0 ;
      RECT  98270.0 90590.0 98975.0 89245.0 ;
      RECT  98270.0 90590.0 98975.0 91935.0 ;
      RECT  98270.0 93280.0 98975.0 91935.0 ;
      RECT  98270.0 93280.0 98975.0 94625.0 ;
      RECT  98270.0 95970.0 98975.0 94625.0 ;
      RECT  98270.0 95970.0 98975.0 97315.0 ;
      RECT  98270.0 98660.0 98975.0 97315.0 ;
      RECT  98270.0 98660.0 98975.0 100005.0 ;
      RECT  98270.0 101350.0 98975.0 100005.0 ;
      RECT  98270.0 101350.0 98975.0 102695.0 ;
      RECT  98270.0 104040.0 98975.0 102695.0 ;
      RECT  98270.0 104040.0 98975.0 105385.0 ;
      RECT  98270.0 106730.0 98975.0 105385.0 ;
      RECT  98270.0 106730.0 98975.0 108075.0 ;
      RECT  98270.0 109420.0 98975.0 108075.0 ;
      RECT  98270.0 109420.0 98975.0 110765.0 ;
      RECT  98270.0 112110.0 98975.0 110765.0 ;
      RECT  98270.0 112110.0 98975.0 113455.0 ;
      RECT  98270.0 114800.0 98975.0 113455.0 ;
      RECT  98270.0 114800.0 98975.0 116145.0 ;
      RECT  98270.0 117490.0 98975.0 116145.0 ;
      RECT  98270.0 117490.0 98975.0 118835.0 ;
      RECT  98270.0 120180.0 98975.0 118835.0 ;
      RECT  98270.0 120180.0 98975.0 121525.0 ;
      RECT  98270.0 122870.0 98975.0 121525.0 ;
      RECT  98270.0 122870.0 98975.0 124215.0 ;
      RECT  98270.0 125560.0 98975.0 124215.0 ;
      RECT  98270.0 125560.0 98975.0 126905.0 ;
      RECT  98270.0 128250.0 98975.0 126905.0 ;
      RECT  98270.0 128250.0 98975.0 129595.0 ;
      RECT  98270.0 130940.0 98975.0 129595.0 ;
      RECT  98270.0 130940.0 98975.0 132285.0 ;
      RECT  98270.0 133630.0 98975.0 132285.0 ;
      RECT  98270.0 133630.0 98975.0 134975.0 ;
      RECT  98270.0 136320.0 98975.0 134975.0 ;
      RECT  98270.0 136320.0 98975.0 137665.0 ;
      RECT  98270.0 139010.0 98975.0 137665.0 ;
      RECT  98270.0 139010.0 98975.0 140355.0 ;
      RECT  98270.0 141700.0 98975.0 140355.0 ;
      RECT  98270.0 141700.0 98975.0 143045.0 ;
      RECT  98270.0 144390.0 98975.0 143045.0 ;
      RECT  98270.0 144390.0 98975.0 145735.0 ;
      RECT  98270.0 147080.0 98975.0 145735.0 ;
      RECT  98270.0 147080.0 98975.0 148425.0 ;
      RECT  98270.0 149770.0 98975.0 148425.0 ;
      RECT  98270.0 149770.0 98975.0 151115.0 ;
      RECT  98270.0 152460.0 98975.0 151115.0 ;
      RECT  98270.0 152460.0 98975.0 153805.0 ;
      RECT  98270.0 155150.0 98975.0 153805.0 ;
      RECT  98270.0 155150.0 98975.0 156495.0 ;
      RECT  98270.0 157840.0 98975.0 156495.0 ;
      RECT  98270.0 157840.0 98975.0 159185.0 ;
      RECT  98270.0 160530.0 98975.0 159185.0 ;
      RECT  98270.0 160530.0 98975.0 161875.0 ;
      RECT  98270.0 163220.0 98975.0 161875.0 ;
      RECT  98270.0 163220.0 98975.0 164565.0 ;
      RECT  98270.0 165910.0 98975.0 164565.0 ;
      RECT  98270.0 165910.0 98975.0 167255.0 ;
      RECT  98270.0 168600.0 98975.0 167255.0 ;
      RECT  98270.0 168600.0 98975.0 169945.0 ;
      RECT  98270.0 171290.0 98975.0 169945.0 ;
      RECT  98270.0 171290.0 98975.0 172635.0 ;
      RECT  98270.0 173980.0 98975.0 172635.0 ;
      RECT  98270.0 173980.0 98975.0 175325.0 ;
      RECT  98270.0 176670.0 98975.0 175325.0 ;
      RECT  98270.0 176670.0 98975.0 178015.0 ;
      RECT  98270.0 179360.0 98975.0 178015.0 ;
      RECT  98270.0 179360.0 98975.0 180705.0 ;
      RECT  98270.0 182050.0 98975.0 180705.0 ;
      RECT  98270.0 182050.0 98975.0 183395.0 ;
      RECT  98270.0 184740.0 98975.0 183395.0 ;
      RECT  98270.0 184740.0 98975.0 186085.0 ;
      RECT  98270.0 187430.0 98975.0 186085.0 ;
      RECT  98270.0 187430.0 98975.0 188775.0 ;
      RECT  98270.0 190120.0 98975.0 188775.0 ;
      RECT  98270.0 190120.0 98975.0 191465.0 ;
      RECT  98270.0 192810.0 98975.0 191465.0 ;
      RECT  98270.0 192810.0 98975.0 194155.0 ;
      RECT  98270.0 195500.0 98975.0 194155.0 ;
      RECT  98270.0 195500.0 98975.0 196845.0 ;
      RECT  98270.0 198190.0 98975.0 196845.0 ;
      RECT  98270.0 198190.0 98975.0 199535.0 ;
      RECT  98270.0 200880.0 98975.0 199535.0 ;
      RECT  98270.0 200880.0 98975.0 202225.0 ;
      RECT  98270.0 203570.0 98975.0 202225.0 ;
      RECT  98270.0 203570.0 98975.0 204915.0 ;
      RECT  98270.0 206260.0 98975.0 204915.0 ;
      RECT  98975.0 34100.0 99680.0 35445.0 ;
      RECT  98975.0 36790.0 99680.0 35445.0 ;
      RECT  98975.0 36790.0 99680.0 38135.0 ;
      RECT  98975.0 39480.0 99680.0 38135.0 ;
      RECT  98975.0 39480.0 99680.0 40825.0 ;
      RECT  98975.0 42170.0 99680.0 40825.0 ;
      RECT  98975.0 42170.0 99680.0 43515.0 ;
      RECT  98975.0 44860.0 99680.0 43515.0 ;
      RECT  98975.0 44860.0 99680.0 46205.0 ;
      RECT  98975.0 47550.0 99680.0 46205.0 ;
      RECT  98975.0 47550.0 99680.0 48895.0 ;
      RECT  98975.0 50240.0 99680.0 48895.0 ;
      RECT  98975.0 50240.0 99680.0 51585.0 ;
      RECT  98975.0 52930.0 99680.0 51585.0 ;
      RECT  98975.0 52930.0 99680.0 54275.0 ;
      RECT  98975.0 55620.0 99680.0 54275.0 ;
      RECT  98975.0 55620.0 99680.0 56965.0 ;
      RECT  98975.0 58310.0 99680.0 56965.0 ;
      RECT  98975.0 58310.0 99680.0 59655.0 ;
      RECT  98975.0 61000.0 99680.0 59655.0 ;
      RECT  98975.0 61000.0 99680.0 62345.0 ;
      RECT  98975.0 63690.0 99680.0 62345.0 ;
      RECT  98975.0 63690.0 99680.0 65035.0 ;
      RECT  98975.0 66380.0 99680.0 65035.0 ;
      RECT  98975.0 66380.0 99680.0 67725.0 ;
      RECT  98975.0 69070.0 99680.0 67725.0 ;
      RECT  98975.0 69070.0 99680.0 70415.0 ;
      RECT  98975.0 71760.0 99680.0 70415.0 ;
      RECT  98975.0 71760.0 99680.0 73105.0 ;
      RECT  98975.0 74450.0 99680.0 73105.0 ;
      RECT  98975.0 74450.0 99680.0 75795.0 ;
      RECT  98975.0 77140.0 99680.0 75795.0 ;
      RECT  98975.0 77140.0 99680.0 78485.0 ;
      RECT  98975.0 79830.0 99680.0 78485.0 ;
      RECT  98975.0 79830.0 99680.0 81175.0 ;
      RECT  98975.0 82520.0 99680.0 81175.0 ;
      RECT  98975.0 82520.0 99680.0 83865.0 ;
      RECT  98975.0 85210.0 99680.0 83865.0 ;
      RECT  98975.0 85210.0 99680.0 86555.0 ;
      RECT  98975.0 87900.0 99680.0 86555.0 ;
      RECT  98975.0 87900.0 99680.0 89245.0 ;
      RECT  98975.0 90590.0 99680.0 89245.0 ;
      RECT  98975.0 90590.0 99680.0 91935.0 ;
      RECT  98975.0 93280.0 99680.0 91935.0 ;
      RECT  98975.0 93280.0 99680.0 94625.0 ;
      RECT  98975.0 95970.0 99680.0 94625.0 ;
      RECT  98975.0 95970.0 99680.0 97315.0 ;
      RECT  98975.0 98660.0 99680.0 97315.0 ;
      RECT  98975.0 98660.0 99680.0 100005.0 ;
      RECT  98975.0 101350.0 99680.0 100005.0 ;
      RECT  98975.0 101350.0 99680.0 102695.0 ;
      RECT  98975.0 104040.0 99680.0 102695.0 ;
      RECT  98975.0 104040.0 99680.0 105385.0 ;
      RECT  98975.0 106730.0 99680.0 105385.0 ;
      RECT  98975.0 106730.0 99680.0 108075.0 ;
      RECT  98975.0 109420.0 99680.0 108075.0 ;
      RECT  98975.0 109420.0 99680.0 110765.0 ;
      RECT  98975.0 112110.0 99680.0 110765.0 ;
      RECT  98975.0 112110.0 99680.0 113455.0 ;
      RECT  98975.0 114800.0 99680.0 113455.0 ;
      RECT  98975.0 114800.0 99680.0 116145.0 ;
      RECT  98975.0 117490.0 99680.0 116145.0 ;
      RECT  98975.0 117490.0 99680.0 118835.0 ;
      RECT  98975.0 120180.0 99680.0 118835.0 ;
      RECT  98975.0 120180.0 99680.0 121525.0 ;
      RECT  98975.0 122870.0 99680.0 121525.0 ;
      RECT  98975.0 122870.0 99680.0 124215.0 ;
      RECT  98975.0 125560.0 99680.0 124215.0 ;
      RECT  98975.0 125560.0 99680.0 126905.0 ;
      RECT  98975.0 128250.0 99680.0 126905.0 ;
      RECT  98975.0 128250.0 99680.0 129595.0 ;
      RECT  98975.0 130940.0 99680.0 129595.0 ;
      RECT  98975.0 130940.0 99680.0 132285.0 ;
      RECT  98975.0 133630.0 99680.0 132285.0 ;
      RECT  98975.0 133630.0 99680.0 134975.0 ;
      RECT  98975.0 136320.0 99680.0 134975.0 ;
      RECT  98975.0 136320.0 99680.0 137665.0 ;
      RECT  98975.0 139010.0 99680.0 137665.0 ;
      RECT  98975.0 139010.0 99680.0 140355.0 ;
      RECT  98975.0 141700.0 99680.0 140355.0 ;
      RECT  98975.0 141700.0 99680.0 143045.0 ;
      RECT  98975.0 144390.0 99680.0 143045.0 ;
      RECT  98975.0 144390.0 99680.0 145735.0 ;
      RECT  98975.0 147080.0 99680.0 145735.0 ;
      RECT  98975.0 147080.0 99680.0 148425.0 ;
      RECT  98975.0 149770.0 99680.0 148425.0 ;
      RECT  98975.0 149770.0 99680.0 151115.0 ;
      RECT  98975.0 152460.0 99680.0 151115.0 ;
      RECT  98975.0 152460.0 99680.0 153805.0 ;
      RECT  98975.0 155150.0 99680.0 153805.0 ;
      RECT  98975.0 155150.0 99680.0 156495.0 ;
      RECT  98975.0 157840.0 99680.0 156495.0 ;
      RECT  98975.0 157840.0 99680.0 159185.0 ;
      RECT  98975.0 160530.0 99680.0 159185.0 ;
      RECT  98975.0 160530.0 99680.0 161875.0 ;
      RECT  98975.0 163220.0 99680.0 161875.0 ;
      RECT  98975.0 163220.0 99680.0 164565.0 ;
      RECT  98975.0 165910.0 99680.0 164565.0 ;
      RECT  98975.0 165910.0 99680.0 167255.0 ;
      RECT  98975.0 168600.0 99680.0 167255.0 ;
      RECT  98975.0 168600.0 99680.0 169945.0 ;
      RECT  98975.0 171290.0 99680.0 169945.0 ;
      RECT  98975.0 171290.0 99680.0 172635.0 ;
      RECT  98975.0 173980.0 99680.0 172635.0 ;
      RECT  98975.0 173980.0 99680.0 175325.0 ;
      RECT  98975.0 176670.0 99680.0 175325.0 ;
      RECT  98975.0 176670.0 99680.0 178015.0 ;
      RECT  98975.0 179360.0 99680.0 178015.0 ;
      RECT  98975.0 179360.0 99680.0 180705.0 ;
      RECT  98975.0 182050.0 99680.0 180705.0 ;
      RECT  98975.0 182050.0 99680.0 183395.0 ;
      RECT  98975.0 184740.0 99680.0 183395.0 ;
      RECT  98975.0 184740.0 99680.0 186085.0 ;
      RECT  98975.0 187430.0 99680.0 186085.0 ;
      RECT  98975.0 187430.0 99680.0 188775.0 ;
      RECT  98975.0 190120.0 99680.0 188775.0 ;
      RECT  98975.0 190120.0 99680.0 191465.0 ;
      RECT  98975.0 192810.0 99680.0 191465.0 ;
      RECT  98975.0 192810.0 99680.0 194155.0 ;
      RECT  98975.0 195500.0 99680.0 194155.0 ;
      RECT  98975.0 195500.0 99680.0 196845.0 ;
      RECT  98975.0 198190.0 99680.0 196845.0 ;
      RECT  98975.0 198190.0 99680.0 199535.0 ;
      RECT  98975.0 200880.0 99680.0 199535.0 ;
      RECT  98975.0 200880.0 99680.0 202225.0 ;
      RECT  98975.0 203570.0 99680.0 202225.0 ;
      RECT  98975.0 203570.0 99680.0 204915.0 ;
      RECT  98975.0 206260.0 99680.0 204915.0 ;
      RECT  99680.0 34100.0 100385.0 35445.0 ;
      RECT  99680.0 36790.0 100385.0 35445.0 ;
      RECT  99680.0 36790.0 100385.0 38135.0 ;
      RECT  99680.0 39480.0 100385.0 38135.0 ;
      RECT  99680.0 39480.0 100385.0 40825.0 ;
      RECT  99680.0 42170.0 100385.0 40825.0 ;
      RECT  99680.0 42170.0 100385.0 43515.0 ;
      RECT  99680.0 44860.0 100385.0 43515.0 ;
      RECT  99680.0 44860.0 100385.0 46205.0 ;
      RECT  99680.0 47550.0 100385.0 46205.0 ;
      RECT  99680.0 47550.0 100385.0 48895.0 ;
      RECT  99680.0 50240.0 100385.0 48895.0 ;
      RECT  99680.0 50240.0 100385.0 51585.0 ;
      RECT  99680.0 52930.0 100385.0 51585.0 ;
      RECT  99680.0 52930.0 100385.0 54275.0 ;
      RECT  99680.0 55620.0 100385.0 54275.0 ;
      RECT  99680.0 55620.0 100385.0 56965.0 ;
      RECT  99680.0 58310.0 100385.0 56965.0 ;
      RECT  99680.0 58310.0 100385.0 59655.0 ;
      RECT  99680.0 61000.0 100385.0 59655.0 ;
      RECT  99680.0 61000.0 100385.0 62345.0 ;
      RECT  99680.0 63690.0 100385.0 62345.0 ;
      RECT  99680.0 63690.0 100385.0 65035.0 ;
      RECT  99680.0 66380.0 100385.0 65035.0 ;
      RECT  99680.0 66380.0 100385.0 67725.0 ;
      RECT  99680.0 69070.0 100385.0 67725.0 ;
      RECT  99680.0 69070.0 100385.0 70415.0 ;
      RECT  99680.0 71760.0 100385.0 70415.0 ;
      RECT  99680.0 71760.0 100385.0 73105.0 ;
      RECT  99680.0 74450.0 100385.0 73105.0 ;
      RECT  99680.0 74450.0 100385.0 75795.0 ;
      RECT  99680.0 77140.0 100385.0 75795.0 ;
      RECT  99680.0 77140.0 100385.0 78485.0 ;
      RECT  99680.0 79830.0 100385.0 78485.0 ;
      RECT  99680.0 79830.0 100385.0 81175.0 ;
      RECT  99680.0 82520.0 100385.0 81175.0 ;
      RECT  99680.0 82520.0 100385.0 83865.0 ;
      RECT  99680.0 85210.0 100385.0 83865.0 ;
      RECT  99680.0 85210.0 100385.0 86555.0 ;
      RECT  99680.0 87900.0 100385.0 86555.0 ;
      RECT  99680.0 87900.0 100385.0 89245.0 ;
      RECT  99680.0 90590.0 100385.0 89245.0 ;
      RECT  99680.0 90590.0 100385.0 91935.0 ;
      RECT  99680.0 93280.0 100385.0 91935.0 ;
      RECT  99680.0 93280.0 100385.0 94625.0 ;
      RECT  99680.0 95970.0 100385.0 94625.0 ;
      RECT  99680.0 95970.0 100385.0 97315.0 ;
      RECT  99680.0 98660.0 100385.0 97315.0 ;
      RECT  99680.0 98660.0 100385.0 100005.0 ;
      RECT  99680.0 101350.0 100385.0 100005.0 ;
      RECT  99680.0 101350.0 100385.0 102695.0 ;
      RECT  99680.0 104040.0 100385.0 102695.0 ;
      RECT  99680.0 104040.0 100385.0 105385.0 ;
      RECT  99680.0 106730.0 100385.0 105385.0 ;
      RECT  99680.0 106730.0 100385.0 108075.0 ;
      RECT  99680.0 109420.0 100385.0 108075.0 ;
      RECT  99680.0 109420.0 100385.0 110765.0 ;
      RECT  99680.0 112110.0 100385.0 110765.0 ;
      RECT  99680.0 112110.0 100385.0 113455.0 ;
      RECT  99680.0 114800.0 100385.0 113455.0 ;
      RECT  99680.0 114800.0 100385.0 116145.0 ;
      RECT  99680.0 117490.0 100385.0 116145.0 ;
      RECT  99680.0 117490.0 100385.0 118835.0 ;
      RECT  99680.0 120180.0 100385.0 118835.0 ;
      RECT  99680.0 120180.0 100385.0 121525.0 ;
      RECT  99680.0 122870.0 100385.0 121525.0 ;
      RECT  99680.0 122870.0 100385.0 124215.0 ;
      RECT  99680.0 125560.0 100385.0 124215.0 ;
      RECT  99680.0 125560.0 100385.0 126905.0 ;
      RECT  99680.0 128250.0 100385.0 126905.0 ;
      RECT  99680.0 128250.0 100385.0 129595.0 ;
      RECT  99680.0 130940.0 100385.0 129595.0 ;
      RECT  99680.0 130940.0 100385.0 132285.0 ;
      RECT  99680.0 133630.0 100385.0 132285.0 ;
      RECT  99680.0 133630.0 100385.0 134975.0 ;
      RECT  99680.0 136320.0 100385.0 134975.0 ;
      RECT  99680.0 136320.0 100385.0 137665.0 ;
      RECT  99680.0 139010.0 100385.0 137665.0 ;
      RECT  99680.0 139010.0 100385.0 140355.0 ;
      RECT  99680.0 141700.0 100385.0 140355.0 ;
      RECT  99680.0 141700.0 100385.0 143045.0 ;
      RECT  99680.0 144390.0 100385.0 143045.0 ;
      RECT  99680.0 144390.0 100385.0 145735.0 ;
      RECT  99680.0 147080.0 100385.0 145735.0 ;
      RECT  99680.0 147080.0 100385.0 148425.0 ;
      RECT  99680.0 149770.0 100385.0 148425.0 ;
      RECT  99680.0 149770.0 100385.0 151115.0 ;
      RECT  99680.0 152460.0 100385.0 151115.0 ;
      RECT  99680.0 152460.0 100385.0 153805.0 ;
      RECT  99680.0 155150.0 100385.0 153805.0 ;
      RECT  99680.0 155150.0 100385.0 156495.0 ;
      RECT  99680.0 157840.0 100385.0 156495.0 ;
      RECT  99680.0 157840.0 100385.0 159185.0 ;
      RECT  99680.0 160530.0 100385.0 159185.0 ;
      RECT  99680.0 160530.0 100385.0 161875.0 ;
      RECT  99680.0 163220.0 100385.0 161875.0 ;
      RECT  99680.0 163220.0 100385.0 164565.0 ;
      RECT  99680.0 165910.0 100385.0 164565.0 ;
      RECT  99680.0 165910.0 100385.0 167255.0 ;
      RECT  99680.0 168600.0 100385.0 167255.0 ;
      RECT  99680.0 168600.0 100385.0 169945.0 ;
      RECT  99680.0 171290.0 100385.0 169945.0 ;
      RECT  99680.0 171290.0 100385.0 172635.0 ;
      RECT  99680.0 173980.0 100385.0 172635.0 ;
      RECT  99680.0 173980.0 100385.0 175325.0 ;
      RECT  99680.0 176670.0 100385.0 175325.0 ;
      RECT  99680.0 176670.0 100385.0 178015.0 ;
      RECT  99680.0 179360.0 100385.0 178015.0 ;
      RECT  99680.0 179360.0 100385.0 180705.0 ;
      RECT  99680.0 182050.0 100385.0 180705.0 ;
      RECT  99680.0 182050.0 100385.0 183395.0 ;
      RECT  99680.0 184740.0 100385.0 183395.0 ;
      RECT  99680.0 184740.0 100385.0 186085.0 ;
      RECT  99680.0 187430.0 100385.0 186085.0 ;
      RECT  99680.0 187430.0 100385.0 188775.0 ;
      RECT  99680.0 190120.0 100385.0 188775.0 ;
      RECT  99680.0 190120.0 100385.0 191465.0 ;
      RECT  99680.0 192810.0 100385.0 191465.0 ;
      RECT  99680.0 192810.0 100385.0 194155.0 ;
      RECT  99680.0 195500.0 100385.0 194155.0 ;
      RECT  99680.0 195500.0 100385.0 196845.0 ;
      RECT  99680.0 198190.0 100385.0 196845.0 ;
      RECT  99680.0 198190.0 100385.0 199535.0 ;
      RECT  99680.0 200880.0 100385.0 199535.0 ;
      RECT  99680.0 200880.0 100385.0 202225.0 ;
      RECT  99680.0 203570.0 100385.0 202225.0 ;
      RECT  99680.0 203570.0 100385.0 204915.0 ;
      RECT  99680.0 206260.0 100385.0 204915.0 ;
      RECT  100385.0 34100.0 101090.0 35445.0 ;
      RECT  100385.0 36790.0 101090.0 35445.0 ;
      RECT  100385.0 36790.0 101090.0 38135.0 ;
      RECT  100385.0 39480.0 101090.0 38135.0 ;
      RECT  100385.0 39480.0 101090.0 40825.0 ;
      RECT  100385.0 42170.0 101090.0 40825.0 ;
      RECT  100385.0 42170.0 101090.0 43515.0 ;
      RECT  100385.0 44860.0 101090.0 43515.0 ;
      RECT  100385.0 44860.0 101090.0 46205.0 ;
      RECT  100385.0 47550.0 101090.0 46205.0 ;
      RECT  100385.0 47550.0 101090.0 48895.0 ;
      RECT  100385.0 50240.0 101090.0 48895.0 ;
      RECT  100385.0 50240.0 101090.0 51585.0 ;
      RECT  100385.0 52930.0 101090.0 51585.0 ;
      RECT  100385.0 52930.0 101090.0 54275.0 ;
      RECT  100385.0 55620.0 101090.0 54275.0 ;
      RECT  100385.0 55620.0 101090.0 56965.0 ;
      RECT  100385.0 58310.0 101090.0 56965.0 ;
      RECT  100385.0 58310.0 101090.0 59655.0 ;
      RECT  100385.0 61000.0 101090.0 59655.0 ;
      RECT  100385.0 61000.0 101090.0 62345.0 ;
      RECT  100385.0 63690.0 101090.0 62345.0 ;
      RECT  100385.0 63690.0 101090.0 65035.0 ;
      RECT  100385.0 66380.0 101090.0 65035.0 ;
      RECT  100385.0 66380.0 101090.0 67725.0 ;
      RECT  100385.0 69070.0 101090.0 67725.0 ;
      RECT  100385.0 69070.0 101090.0 70415.0 ;
      RECT  100385.0 71760.0 101090.0 70415.0 ;
      RECT  100385.0 71760.0 101090.0 73105.0 ;
      RECT  100385.0 74450.0 101090.0 73105.0 ;
      RECT  100385.0 74450.0 101090.0 75795.0 ;
      RECT  100385.0 77140.0 101090.0 75795.0 ;
      RECT  100385.0 77140.0 101090.0 78485.0 ;
      RECT  100385.0 79830.0 101090.0 78485.0 ;
      RECT  100385.0 79830.0 101090.0 81175.0 ;
      RECT  100385.0 82520.0 101090.0 81175.0 ;
      RECT  100385.0 82520.0 101090.0 83865.0 ;
      RECT  100385.0 85210.0 101090.0 83865.0 ;
      RECT  100385.0 85210.0 101090.0 86555.0 ;
      RECT  100385.0 87900.0 101090.0 86555.0 ;
      RECT  100385.0 87900.0 101090.0 89245.0 ;
      RECT  100385.0 90590.0 101090.0 89245.0 ;
      RECT  100385.0 90590.0 101090.0 91935.0 ;
      RECT  100385.0 93280.0 101090.0 91935.0 ;
      RECT  100385.0 93280.0 101090.0 94625.0 ;
      RECT  100385.0 95970.0 101090.0 94625.0 ;
      RECT  100385.0 95970.0 101090.0 97315.0 ;
      RECT  100385.0 98660.0 101090.0 97315.0 ;
      RECT  100385.0 98660.0 101090.0 100005.0 ;
      RECT  100385.0 101350.0 101090.0 100005.0 ;
      RECT  100385.0 101350.0 101090.0 102695.0 ;
      RECT  100385.0 104040.0 101090.0 102695.0 ;
      RECT  100385.0 104040.0 101090.0 105385.0 ;
      RECT  100385.0 106730.0 101090.0 105385.0 ;
      RECT  100385.0 106730.0 101090.0 108075.0 ;
      RECT  100385.0 109420.0 101090.0 108075.0 ;
      RECT  100385.0 109420.0 101090.0 110765.0 ;
      RECT  100385.0 112110.0 101090.0 110765.0 ;
      RECT  100385.0 112110.0 101090.0 113455.0 ;
      RECT  100385.0 114800.0 101090.0 113455.0 ;
      RECT  100385.0 114800.0 101090.0 116145.0 ;
      RECT  100385.0 117490.0 101090.0 116145.0 ;
      RECT  100385.0 117490.0 101090.0 118835.0 ;
      RECT  100385.0 120180.0 101090.0 118835.0 ;
      RECT  100385.0 120180.0 101090.0 121525.0 ;
      RECT  100385.0 122870.0 101090.0 121525.0 ;
      RECT  100385.0 122870.0 101090.0 124215.0 ;
      RECT  100385.0 125560.0 101090.0 124215.0 ;
      RECT  100385.0 125560.0 101090.0 126905.0 ;
      RECT  100385.0 128250.0 101090.0 126905.0 ;
      RECT  100385.0 128250.0 101090.0 129595.0 ;
      RECT  100385.0 130940.0 101090.0 129595.0 ;
      RECT  100385.0 130940.0 101090.0 132285.0 ;
      RECT  100385.0 133630.0 101090.0 132285.0 ;
      RECT  100385.0 133630.0 101090.0 134975.0 ;
      RECT  100385.0 136320.0 101090.0 134975.0 ;
      RECT  100385.0 136320.0 101090.0 137665.0 ;
      RECT  100385.0 139010.0 101090.0 137665.0 ;
      RECT  100385.0 139010.0 101090.0 140355.0 ;
      RECT  100385.0 141700.0 101090.0 140355.0 ;
      RECT  100385.0 141700.0 101090.0 143045.0 ;
      RECT  100385.0 144390.0 101090.0 143045.0 ;
      RECT  100385.0 144390.0 101090.0 145735.0 ;
      RECT  100385.0 147080.0 101090.0 145735.0 ;
      RECT  100385.0 147080.0 101090.0 148425.0 ;
      RECT  100385.0 149770.0 101090.0 148425.0 ;
      RECT  100385.0 149770.0 101090.0 151115.0 ;
      RECT  100385.0 152460.0 101090.0 151115.0 ;
      RECT  100385.0 152460.0 101090.0 153805.0 ;
      RECT  100385.0 155150.0 101090.0 153805.0 ;
      RECT  100385.0 155150.0 101090.0 156495.0 ;
      RECT  100385.0 157840.0 101090.0 156495.0 ;
      RECT  100385.0 157840.0 101090.0 159185.0 ;
      RECT  100385.0 160530.0 101090.0 159185.0 ;
      RECT  100385.0 160530.0 101090.0 161875.0 ;
      RECT  100385.0 163220.0 101090.0 161875.0 ;
      RECT  100385.0 163220.0 101090.0 164565.0 ;
      RECT  100385.0 165910.0 101090.0 164565.0 ;
      RECT  100385.0 165910.0 101090.0 167255.0 ;
      RECT  100385.0 168600.0 101090.0 167255.0 ;
      RECT  100385.0 168600.0 101090.0 169945.0 ;
      RECT  100385.0 171290.0 101090.0 169945.0 ;
      RECT  100385.0 171290.0 101090.0 172635.0 ;
      RECT  100385.0 173980.0 101090.0 172635.0 ;
      RECT  100385.0 173980.0 101090.0 175325.0 ;
      RECT  100385.0 176670.0 101090.0 175325.0 ;
      RECT  100385.0 176670.0 101090.0 178015.0 ;
      RECT  100385.0 179360.0 101090.0 178015.0 ;
      RECT  100385.0 179360.0 101090.0 180705.0 ;
      RECT  100385.0 182050.0 101090.0 180705.0 ;
      RECT  100385.0 182050.0 101090.0 183395.0 ;
      RECT  100385.0 184740.0 101090.0 183395.0 ;
      RECT  100385.0 184740.0 101090.0 186085.0 ;
      RECT  100385.0 187430.0 101090.0 186085.0 ;
      RECT  100385.0 187430.0 101090.0 188775.0 ;
      RECT  100385.0 190120.0 101090.0 188775.0 ;
      RECT  100385.0 190120.0 101090.0 191465.0 ;
      RECT  100385.0 192810.0 101090.0 191465.0 ;
      RECT  100385.0 192810.0 101090.0 194155.0 ;
      RECT  100385.0 195500.0 101090.0 194155.0 ;
      RECT  100385.0 195500.0 101090.0 196845.0 ;
      RECT  100385.0 198190.0 101090.0 196845.0 ;
      RECT  100385.0 198190.0 101090.0 199535.0 ;
      RECT  100385.0 200880.0 101090.0 199535.0 ;
      RECT  100385.0 200880.0 101090.0 202225.0 ;
      RECT  100385.0 203570.0 101090.0 202225.0 ;
      RECT  100385.0 203570.0 101090.0 204915.0 ;
      RECT  100385.0 206260.0 101090.0 204915.0 ;
      RECT  101090.0 34100.0 101795.0 35445.0 ;
      RECT  101090.0 36790.0 101795.0 35445.0 ;
      RECT  101090.0 36790.0 101795.0 38135.0 ;
      RECT  101090.0 39480.0 101795.0 38135.0 ;
      RECT  101090.0 39480.0 101795.0 40825.0 ;
      RECT  101090.0 42170.0 101795.0 40825.0 ;
      RECT  101090.0 42170.0 101795.0 43515.0 ;
      RECT  101090.0 44860.0 101795.0 43515.0 ;
      RECT  101090.0 44860.0 101795.0 46205.0 ;
      RECT  101090.0 47550.0 101795.0 46205.0 ;
      RECT  101090.0 47550.0 101795.0 48895.0 ;
      RECT  101090.0 50240.0 101795.0 48895.0 ;
      RECT  101090.0 50240.0 101795.0 51585.0 ;
      RECT  101090.0 52930.0 101795.0 51585.0 ;
      RECT  101090.0 52930.0 101795.0 54275.0 ;
      RECT  101090.0 55620.0 101795.0 54275.0 ;
      RECT  101090.0 55620.0 101795.0 56965.0 ;
      RECT  101090.0 58310.0 101795.0 56965.0 ;
      RECT  101090.0 58310.0 101795.0 59655.0 ;
      RECT  101090.0 61000.0 101795.0 59655.0 ;
      RECT  101090.0 61000.0 101795.0 62345.0 ;
      RECT  101090.0 63690.0 101795.0 62345.0 ;
      RECT  101090.0 63690.0 101795.0 65035.0 ;
      RECT  101090.0 66380.0 101795.0 65035.0 ;
      RECT  101090.0 66380.0 101795.0 67725.0 ;
      RECT  101090.0 69070.0 101795.0 67725.0 ;
      RECT  101090.0 69070.0 101795.0 70415.0 ;
      RECT  101090.0 71760.0 101795.0 70415.0 ;
      RECT  101090.0 71760.0 101795.0 73105.0 ;
      RECT  101090.0 74450.0 101795.0 73105.0 ;
      RECT  101090.0 74450.0 101795.0 75795.0 ;
      RECT  101090.0 77140.0 101795.0 75795.0 ;
      RECT  101090.0 77140.0 101795.0 78485.0 ;
      RECT  101090.0 79830.0 101795.0 78485.0 ;
      RECT  101090.0 79830.0 101795.0 81175.0 ;
      RECT  101090.0 82520.0 101795.0 81175.0 ;
      RECT  101090.0 82520.0 101795.0 83865.0 ;
      RECT  101090.0 85210.0 101795.0 83865.0 ;
      RECT  101090.0 85210.0 101795.0 86555.0 ;
      RECT  101090.0 87900.0 101795.0 86555.0 ;
      RECT  101090.0 87900.0 101795.0 89245.0 ;
      RECT  101090.0 90590.0 101795.0 89245.0 ;
      RECT  101090.0 90590.0 101795.0 91935.0 ;
      RECT  101090.0 93280.0 101795.0 91935.0 ;
      RECT  101090.0 93280.0 101795.0 94625.0 ;
      RECT  101090.0 95970.0 101795.0 94625.0 ;
      RECT  101090.0 95970.0 101795.0 97315.0 ;
      RECT  101090.0 98660.0 101795.0 97315.0 ;
      RECT  101090.0 98660.0 101795.0 100005.0 ;
      RECT  101090.0 101350.0 101795.0 100005.0 ;
      RECT  101090.0 101350.0 101795.0 102695.0 ;
      RECT  101090.0 104040.0 101795.0 102695.0 ;
      RECT  101090.0 104040.0 101795.0 105385.0 ;
      RECT  101090.0 106730.0 101795.0 105385.0 ;
      RECT  101090.0 106730.0 101795.0 108075.0 ;
      RECT  101090.0 109420.0 101795.0 108075.0 ;
      RECT  101090.0 109420.0 101795.0 110765.0 ;
      RECT  101090.0 112110.0 101795.0 110765.0 ;
      RECT  101090.0 112110.0 101795.0 113455.0 ;
      RECT  101090.0 114800.0 101795.0 113455.0 ;
      RECT  101090.0 114800.0 101795.0 116145.0 ;
      RECT  101090.0 117490.0 101795.0 116145.0 ;
      RECT  101090.0 117490.0 101795.0 118835.0 ;
      RECT  101090.0 120180.0 101795.0 118835.0 ;
      RECT  101090.0 120180.0 101795.0 121525.0 ;
      RECT  101090.0 122870.0 101795.0 121525.0 ;
      RECT  101090.0 122870.0 101795.0 124215.0 ;
      RECT  101090.0 125560.0 101795.0 124215.0 ;
      RECT  101090.0 125560.0 101795.0 126905.0 ;
      RECT  101090.0 128250.0 101795.0 126905.0 ;
      RECT  101090.0 128250.0 101795.0 129595.0 ;
      RECT  101090.0 130940.0 101795.0 129595.0 ;
      RECT  101090.0 130940.0 101795.0 132285.0 ;
      RECT  101090.0 133630.0 101795.0 132285.0 ;
      RECT  101090.0 133630.0 101795.0 134975.0 ;
      RECT  101090.0 136320.0 101795.0 134975.0 ;
      RECT  101090.0 136320.0 101795.0 137665.0 ;
      RECT  101090.0 139010.0 101795.0 137665.0 ;
      RECT  101090.0 139010.0 101795.0 140355.0 ;
      RECT  101090.0 141700.0 101795.0 140355.0 ;
      RECT  101090.0 141700.0 101795.0 143045.0 ;
      RECT  101090.0 144390.0 101795.0 143045.0 ;
      RECT  101090.0 144390.0 101795.0 145735.0 ;
      RECT  101090.0 147080.0 101795.0 145735.0 ;
      RECT  101090.0 147080.0 101795.0 148425.0 ;
      RECT  101090.0 149770.0 101795.0 148425.0 ;
      RECT  101090.0 149770.0 101795.0 151115.0 ;
      RECT  101090.0 152460.0 101795.0 151115.0 ;
      RECT  101090.0 152460.0 101795.0 153805.0 ;
      RECT  101090.0 155150.0 101795.0 153805.0 ;
      RECT  101090.0 155150.0 101795.0 156495.0 ;
      RECT  101090.0 157840.0 101795.0 156495.0 ;
      RECT  101090.0 157840.0 101795.0 159185.0 ;
      RECT  101090.0 160530.0 101795.0 159185.0 ;
      RECT  101090.0 160530.0 101795.0 161875.0 ;
      RECT  101090.0 163220.0 101795.0 161875.0 ;
      RECT  101090.0 163220.0 101795.0 164565.0 ;
      RECT  101090.0 165910.0 101795.0 164565.0 ;
      RECT  101090.0 165910.0 101795.0 167255.0 ;
      RECT  101090.0 168600.0 101795.0 167255.0 ;
      RECT  101090.0 168600.0 101795.0 169945.0 ;
      RECT  101090.0 171290.0 101795.0 169945.0 ;
      RECT  101090.0 171290.0 101795.0 172635.0 ;
      RECT  101090.0 173980.0 101795.0 172635.0 ;
      RECT  101090.0 173980.0 101795.0 175325.0 ;
      RECT  101090.0 176670.0 101795.0 175325.0 ;
      RECT  101090.0 176670.0 101795.0 178015.0 ;
      RECT  101090.0 179360.0 101795.0 178015.0 ;
      RECT  101090.0 179360.0 101795.0 180705.0 ;
      RECT  101090.0 182050.0 101795.0 180705.0 ;
      RECT  101090.0 182050.0 101795.0 183395.0 ;
      RECT  101090.0 184740.0 101795.0 183395.0 ;
      RECT  101090.0 184740.0 101795.0 186085.0 ;
      RECT  101090.0 187430.0 101795.0 186085.0 ;
      RECT  101090.0 187430.0 101795.0 188775.0 ;
      RECT  101090.0 190120.0 101795.0 188775.0 ;
      RECT  101090.0 190120.0 101795.0 191465.0 ;
      RECT  101090.0 192810.0 101795.0 191465.0 ;
      RECT  101090.0 192810.0 101795.0 194155.0 ;
      RECT  101090.0 195500.0 101795.0 194155.0 ;
      RECT  101090.0 195500.0 101795.0 196845.0 ;
      RECT  101090.0 198190.0 101795.0 196845.0 ;
      RECT  101090.0 198190.0 101795.0 199535.0 ;
      RECT  101090.0 200880.0 101795.0 199535.0 ;
      RECT  101090.0 200880.0 101795.0 202225.0 ;
      RECT  101090.0 203570.0 101795.0 202225.0 ;
      RECT  101090.0 203570.0 101795.0 204915.0 ;
      RECT  101090.0 206260.0 101795.0 204915.0 ;
      RECT  101795.0 34100.0 102500.0 35445.0 ;
      RECT  101795.0 36790.0 102500.0 35445.0 ;
      RECT  101795.0 36790.0 102500.0 38135.0 ;
      RECT  101795.0 39480.0 102500.0 38135.0 ;
      RECT  101795.0 39480.0 102500.0 40825.0 ;
      RECT  101795.0 42170.0 102500.0 40825.0 ;
      RECT  101795.0 42170.0 102500.0 43515.0 ;
      RECT  101795.0 44860.0 102500.0 43515.0 ;
      RECT  101795.0 44860.0 102500.0 46205.0 ;
      RECT  101795.0 47550.0 102500.0 46205.0 ;
      RECT  101795.0 47550.0 102500.0 48895.0 ;
      RECT  101795.0 50240.0 102500.0 48895.0 ;
      RECT  101795.0 50240.0 102500.0 51585.0 ;
      RECT  101795.0 52930.0 102500.0 51585.0 ;
      RECT  101795.0 52930.0 102500.0 54275.0 ;
      RECT  101795.0 55620.0 102500.0 54275.0 ;
      RECT  101795.0 55620.0 102500.0 56965.0 ;
      RECT  101795.0 58310.0 102500.0 56965.0 ;
      RECT  101795.0 58310.0 102500.0 59655.0 ;
      RECT  101795.0 61000.0 102500.0 59655.0 ;
      RECT  101795.0 61000.0 102500.0 62345.0 ;
      RECT  101795.0 63690.0 102500.0 62345.0 ;
      RECT  101795.0 63690.0 102500.0 65035.0 ;
      RECT  101795.0 66380.0 102500.0 65035.0 ;
      RECT  101795.0 66380.0 102500.0 67725.0 ;
      RECT  101795.0 69070.0 102500.0 67725.0 ;
      RECT  101795.0 69070.0 102500.0 70415.0 ;
      RECT  101795.0 71760.0 102500.0 70415.0 ;
      RECT  101795.0 71760.0 102500.0 73105.0 ;
      RECT  101795.0 74450.0 102500.0 73105.0 ;
      RECT  101795.0 74450.0 102500.0 75795.0 ;
      RECT  101795.0 77140.0 102500.0 75795.0 ;
      RECT  101795.0 77140.0 102500.0 78485.0 ;
      RECT  101795.0 79830.0 102500.0 78485.0 ;
      RECT  101795.0 79830.0 102500.0 81175.0 ;
      RECT  101795.0 82520.0 102500.0 81175.0 ;
      RECT  101795.0 82520.0 102500.0 83865.0 ;
      RECT  101795.0 85210.0 102500.0 83865.0 ;
      RECT  101795.0 85210.0 102500.0 86555.0 ;
      RECT  101795.0 87900.0 102500.0 86555.0 ;
      RECT  101795.0 87900.0 102500.0 89245.0 ;
      RECT  101795.0 90590.0 102500.0 89245.0 ;
      RECT  101795.0 90590.0 102500.0 91935.0 ;
      RECT  101795.0 93280.0 102500.0 91935.0 ;
      RECT  101795.0 93280.0 102500.0 94625.0 ;
      RECT  101795.0 95970.0 102500.0 94625.0 ;
      RECT  101795.0 95970.0 102500.0 97315.0 ;
      RECT  101795.0 98660.0 102500.0 97315.0 ;
      RECT  101795.0 98660.0 102500.0 100005.0 ;
      RECT  101795.0 101350.0 102500.0 100005.0 ;
      RECT  101795.0 101350.0 102500.0 102695.0 ;
      RECT  101795.0 104040.0 102500.0 102695.0 ;
      RECT  101795.0 104040.0 102500.0 105385.0 ;
      RECT  101795.0 106730.0 102500.0 105385.0 ;
      RECT  101795.0 106730.0 102500.0 108075.0 ;
      RECT  101795.0 109420.0 102500.0 108075.0 ;
      RECT  101795.0 109420.0 102500.0 110765.0 ;
      RECT  101795.0 112110.0 102500.0 110765.0 ;
      RECT  101795.0 112110.0 102500.0 113455.0 ;
      RECT  101795.0 114800.0 102500.0 113455.0 ;
      RECT  101795.0 114800.0 102500.0 116145.0 ;
      RECT  101795.0 117490.0 102500.0 116145.0 ;
      RECT  101795.0 117490.0 102500.0 118835.0 ;
      RECT  101795.0 120180.0 102500.0 118835.0 ;
      RECT  101795.0 120180.0 102500.0 121525.0 ;
      RECT  101795.0 122870.0 102500.0 121525.0 ;
      RECT  101795.0 122870.0 102500.0 124215.0 ;
      RECT  101795.0 125560.0 102500.0 124215.0 ;
      RECT  101795.0 125560.0 102500.0 126905.0 ;
      RECT  101795.0 128250.0 102500.0 126905.0 ;
      RECT  101795.0 128250.0 102500.0 129595.0 ;
      RECT  101795.0 130940.0 102500.0 129595.0 ;
      RECT  101795.0 130940.0 102500.0 132285.0 ;
      RECT  101795.0 133630.0 102500.0 132285.0 ;
      RECT  101795.0 133630.0 102500.0 134975.0 ;
      RECT  101795.0 136320.0 102500.0 134975.0 ;
      RECT  101795.0 136320.0 102500.0 137665.0 ;
      RECT  101795.0 139010.0 102500.0 137665.0 ;
      RECT  101795.0 139010.0 102500.0 140355.0 ;
      RECT  101795.0 141700.0 102500.0 140355.0 ;
      RECT  101795.0 141700.0 102500.0 143045.0 ;
      RECT  101795.0 144390.0 102500.0 143045.0 ;
      RECT  101795.0 144390.0 102500.0 145735.0 ;
      RECT  101795.0 147080.0 102500.0 145735.0 ;
      RECT  101795.0 147080.0 102500.0 148425.0 ;
      RECT  101795.0 149770.0 102500.0 148425.0 ;
      RECT  101795.0 149770.0 102500.0 151115.0 ;
      RECT  101795.0 152460.0 102500.0 151115.0 ;
      RECT  101795.0 152460.0 102500.0 153805.0 ;
      RECT  101795.0 155150.0 102500.0 153805.0 ;
      RECT  101795.0 155150.0 102500.0 156495.0 ;
      RECT  101795.0 157840.0 102500.0 156495.0 ;
      RECT  101795.0 157840.0 102500.0 159185.0 ;
      RECT  101795.0 160530.0 102500.0 159185.0 ;
      RECT  101795.0 160530.0 102500.0 161875.0 ;
      RECT  101795.0 163220.0 102500.0 161875.0 ;
      RECT  101795.0 163220.0 102500.0 164565.0 ;
      RECT  101795.0 165910.0 102500.0 164565.0 ;
      RECT  101795.0 165910.0 102500.0 167255.0 ;
      RECT  101795.0 168600.0 102500.0 167255.0 ;
      RECT  101795.0 168600.0 102500.0 169945.0 ;
      RECT  101795.0 171290.0 102500.0 169945.0 ;
      RECT  101795.0 171290.0 102500.0 172635.0 ;
      RECT  101795.0 173980.0 102500.0 172635.0 ;
      RECT  101795.0 173980.0 102500.0 175325.0 ;
      RECT  101795.0 176670.0 102500.0 175325.0 ;
      RECT  101795.0 176670.0 102500.0 178015.0 ;
      RECT  101795.0 179360.0 102500.0 178015.0 ;
      RECT  101795.0 179360.0 102500.0 180705.0 ;
      RECT  101795.0 182050.0 102500.0 180705.0 ;
      RECT  101795.0 182050.0 102500.0 183395.0 ;
      RECT  101795.0 184740.0 102500.0 183395.0 ;
      RECT  101795.0 184740.0 102500.0 186085.0 ;
      RECT  101795.0 187430.0 102500.0 186085.0 ;
      RECT  101795.0 187430.0 102500.0 188775.0 ;
      RECT  101795.0 190120.0 102500.0 188775.0 ;
      RECT  101795.0 190120.0 102500.0 191465.0 ;
      RECT  101795.0 192810.0 102500.0 191465.0 ;
      RECT  101795.0 192810.0 102500.0 194155.0 ;
      RECT  101795.0 195500.0 102500.0 194155.0 ;
      RECT  101795.0 195500.0 102500.0 196845.0 ;
      RECT  101795.0 198190.0 102500.0 196845.0 ;
      RECT  101795.0 198190.0 102500.0 199535.0 ;
      RECT  101795.0 200880.0 102500.0 199535.0 ;
      RECT  101795.0 200880.0 102500.0 202225.0 ;
      RECT  101795.0 203570.0 102500.0 202225.0 ;
      RECT  101795.0 203570.0 102500.0 204915.0 ;
      RECT  101795.0 206260.0 102500.0 204915.0 ;
      RECT  102500.0 34100.0 103205.0 35445.0 ;
      RECT  102500.0 36790.0 103205.0 35445.0 ;
      RECT  102500.0 36790.0 103205.0 38135.0 ;
      RECT  102500.0 39480.0 103205.0 38135.0 ;
      RECT  102500.0 39480.0 103205.0 40825.0 ;
      RECT  102500.0 42170.0 103205.0 40825.0 ;
      RECT  102500.0 42170.0 103205.0 43515.0 ;
      RECT  102500.0 44860.0 103205.0 43515.0 ;
      RECT  102500.0 44860.0 103205.0 46205.0 ;
      RECT  102500.0 47550.0 103205.0 46205.0 ;
      RECT  102500.0 47550.0 103205.0 48895.0 ;
      RECT  102500.0 50240.0 103205.0 48895.0 ;
      RECT  102500.0 50240.0 103205.0 51585.0 ;
      RECT  102500.0 52930.0 103205.0 51585.0 ;
      RECT  102500.0 52930.0 103205.0 54275.0 ;
      RECT  102500.0 55620.0 103205.0 54275.0 ;
      RECT  102500.0 55620.0 103205.0 56965.0 ;
      RECT  102500.0 58310.0 103205.0 56965.0 ;
      RECT  102500.0 58310.0 103205.0 59655.0 ;
      RECT  102500.0 61000.0 103205.0 59655.0 ;
      RECT  102500.0 61000.0 103205.0 62345.0 ;
      RECT  102500.0 63690.0 103205.0 62345.0 ;
      RECT  102500.0 63690.0 103205.0 65035.0 ;
      RECT  102500.0 66380.0 103205.0 65035.0 ;
      RECT  102500.0 66380.0 103205.0 67725.0 ;
      RECT  102500.0 69070.0 103205.0 67725.0 ;
      RECT  102500.0 69070.0 103205.0 70415.0 ;
      RECT  102500.0 71760.0 103205.0 70415.0 ;
      RECT  102500.0 71760.0 103205.0 73105.0 ;
      RECT  102500.0 74450.0 103205.0 73105.0 ;
      RECT  102500.0 74450.0 103205.0 75795.0 ;
      RECT  102500.0 77140.0 103205.0 75795.0 ;
      RECT  102500.0 77140.0 103205.0 78485.0 ;
      RECT  102500.0 79830.0 103205.0 78485.0 ;
      RECT  102500.0 79830.0 103205.0 81175.0 ;
      RECT  102500.0 82520.0 103205.0 81175.0 ;
      RECT  102500.0 82520.0 103205.0 83865.0 ;
      RECT  102500.0 85210.0 103205.0 83865.0 ;
      RECT  102500.0 85210.0 103205.0 86555.0 ;
      RECT  102500.0 87900.0 103205.0 86555.0 ;
      RECT  102500.0 87900.0 103205.0 89245.0 ;
      RECT  102500.0 90590.0 103205.0 89245.0 ;
      RECT  102500.0 90590.0 103205.0 91935.0 ;
      RECT  102500.0 93280.0 103205.0 91935.0 ;
      RECT  102500.0 93280.0 103205.0 94625.0 ;
      RECT  102500.0 95970.0 103205.0 94625.0 ;
      RECT  102500.0 95970.0 103205.0 97315.0 ;
      RECT  102500.0 98660.0 103205.0 97315.0 ;
      RECT  102500.0 98660.0 103205.0 100005.0 ;
      RECT  102500.0 101350.0 103205.0 100005.0 ;
      RECT  102500.0 101350.0 103205.0 102695.0 ;
      RECT  102500.0 104040.0 103205.0 102695.0 ;
      RECT  102500.0 104040.0 103205.0 105385.0 ;
      RECT  102500.0 106730.0 103205.0 105385.0 ;
      RECT  102500.0 106730.0 103205.0 108075.0 ;
      RECT  102500.0 109420.0 103205.0 108075.0 ;
      RECT  102500.0 109420.0 103205.0 110765.0 ;
      RECT  102500.0 112110.0 103205.0 110765.0 ;
      RECT  102500.0 112110.0 103205.0 113455.0 ;
      RECT  102500.0 114800.0 103205.0 113455.0 ;
      RECT  102500.0 114800.0 103205.0 116145.0 ;
      RECT  102500.0 117490.0 103205.0 116145.0 ;
      RECT  102500.0 117490.0 103205.0 118835.0 ;
      RECT  102500.0 120180.0 103205.0 118835.0 ;
      RECT  102500.0 120180.0 103205.0 121525.0 ;
      RECT  102500.0 122870.0 103205.0 121525.0 ;
      RECT  102500.0 122870.0 103205.0 124215.0 ;
      RECT  102500.0 125560.0 103205.0 124215.0 ;
      RECT  102500.0 125560.0 103205.0 126905.0 ;
      RECT  102500.0 128250.0 103205.0 126905.0 ;
      RECT  102500.0 128250.0 103205.0 129595.0 ;
      RECT  102500.0 130940.0 103205.0 129595.0 ;
      RECT  102500.0 130940.0 103205.0 132285.0 ;
      RECT  102500.0 133630.0 103205.0 132285.0 ;
      RECT  102500.0 133630.0 103205.0 134975.0 ;
      RECT  102500.0 136320.0 103205.0 134975.0 ;
      RECT  102500.0 136320.0 103205.0 137665.0 ;
      RECT  102500.0 139010.0 103205.0 137665.0 ;
      RECT  102500.0 139010.0 103205.0 140355.0 ;
      RECT  102500.0 141700.0 103205.0 140355.0 ;
      RECT  102500.0 141700.0 103205.0 143045.0 ;
      RECT  102500.0 144390.0 103205.0 143045.0 ;
      RECT  102500.0 144390.0 103205.0 145735.0 ;
      RECT  102500.0 147080.0 103205.0 145735.0 ;
      RECT  102500.0 147080.0 103205.0 148425.0 ;
      RECT  102500.0 149770.0 103205.0 148425.0 ;
      RECT  102500.0 149770.0 103205.0 151115.0 ;
      RECT  102500.0 152460.0 103205.0 151115.0 ;
      RECT  102500.0 152460.0 103205.0 153805.0 ;
      RECT  102500.0 155150.0 103205.0 153805.0 ;
      RECT  102500.0 155150.0 103205.0 156495.0 ;
      RECT  102500.0 157840.0 103205.0 156495.0 ;
      RECT  102500.0 157840.0 103205.0 159185.0 ;
      RECT  102500.0 160530.0 103205.0 159185.0 ;
      RECT  102500.0 160530.0 103205.0 161875.0 ;
      RECT  102500.0 163220.0 103205.0 161875.0 ;
      RECT  102500.0 163220.0 103205.0 164565.0 ;
      RECT  102500.0 165910.0 103205.0 164565.0 ;
      RECT  102500.0 165910.0 103205.0 167255.0 ;
      RECT  102500.0 168600.0 103205.0 167255.0 ;
      RECT  102500.0 168600.0 103205.0 169945.0 ;
      RECT  102500.0 171290.0 103205.0 169945.0 ;
      RECT  102500.0 171290.0 103205.0 172635.0 ;
      RECT  102500.0 173980.0 103205.0 172635.0 ;
      RECT  102500.0 173980.0 103205.0 175325.0 ;
      RECT  102500.0 176670.0 103205.0 175325.0 ;
      RECT  102500.0 176670.0 103205.0 178015.0 ;
      RECT  102500.0 179360.0 103205.0 178015.0 ;
      RECT  102500.0 179360.0 103205.0 180705.0 ;
      RECT  102500.0 182050.0 103205.0 180705.0 ;
      RECT  102500.0 182050.0 103205.0 183395.0 ;
      RECT  102500.0 184740.0 103205.0 183395.0 ;
      RECT  102500.0 184740.0 103205.0 186085.0 ;
      RECT  102500.0 187430.0 103205.0 186085.0 ;
      RECT  102500.0 187430.0 103205.0 188775.0 ;
      RECT  102500.0 190120.0 103205.0 188775.0 ;
      RECT  102500.0 190120.0 103205.0 191465.0 ;
      RECT  102500.0 192810.0 103205.0 191465.0 ;
      RECT  102500.0 192810.0 103205.0 194155.0 ;
      RECT  102500.0 195500.0 103205.0 194155.0 ;
      RECT  102500.0 195500.0 103205.0 196845.0 ;
      RECT  102500.0 198190.0 103205.0 196845.0 ;
      RECT  102500.0 198190.0 103205.0 199535.0 ;
      RECT  102500.0 200880.0 103205.0 199535.0 ;
      RECT  102500.0 200880.0 103205.0 202225.0 ;
      RECT  102500.0 203570.0 103205.0 202225.0 ;
      RECT  102500.0 203570.0 103205.0 204915.0 ;
      RECT  102500.0 206260.0 103205.0 204915.0 ;
      RECT  103205.0 34100.0 103910.0 35445.0 ;
      RECT  103205.0 36790.0 103910.0 35445.0 ;
      RECT  103205.0 36790.0 103910.0 38135.0 ;
      RECT  103205.0 39480.0 103910.0 38135.0 ;
      RECT  103205.0 39480.0 103910.0 40825.0 ;
      RECT  103205.0 42170.0 103910.0 40825.0 ;
      RECT  103205.0 42170.0 103910.0 43515.0 ;
      RECT  103205.0 44860.0 103910.0 43515.0 ;
      RECT  103205.0 44860.0 103910.0 46205.0 ;
      RECT  103205.0 47550.0 103910.0 46205.0 ;
      RECT  103205.0 47550.0 103910.0 48895.0 ;
      RECT  103205.0 50240.0 103910.0 48895.0 ;
      RECT  103205.0 50240.0 103910.0 51585.0 ;
      RECT  103205.0 52930.0 103910.0 51585.0 ;
      RECT  103205.0 52930.0 103910.0 54275.0 ;
      RECT  103205.0 55620.0 103910.0 54275.0 ;
      RECT  103205.0 55620.0 103910.0 56965.0 ;
      RECT  103205.0 58310.0 103910.0 56965.0 ;
      RECT  103205.0 58310.0 103910.0 59655.0 ;
      RECT  103205.0 61000.0 103910.0 59655.0 ;
      RECT  103205.0 61000.0 103910.0 62345.0 ;
      RECT  103205.0 63690.0 103910.0 62345.0 ;
      RECT  103205.0 63690.0 103910.0 65035.0 ;
      RECT  103205.0 66380.0 103910.0 65035.0 ;
      RECT  103205.0 66380.0 103910.0 67725.0 ;
      RECT  103205.0 69070.0 103910.0 67725.0 ;
      RECT  103205.0 69070.0 103910.0 70415.0 ;
      RECT  103205.0 71760.0 103910.0 70415.0 ;
      RECT  103205.0 71760.0 103910.0 73105.0 ;
      RECT  103205.0 74450.0 103910.0 73105.0 ;
      RECT  103205.0 74450.0 103910.0 75795.0 ;
      RECT  103205.0 77140.0 103910.0 75795.0 ;
      RECT  103205.0 77140.0 103910.0 78485.0 ;
      RECT  103205.0 79830.0 103910.0 78485.0 ;
      RECT  103205.0 79830.0 103910.0 81175.0 ;
      RECT  103205.0 82520.0 103910.0 81175.0 ;
      RECT  103205.0 82520.0 103910.0 83865.0 ;
      RECT  103205.0 85210.0 103910.0 83865.0 ;
      RECT  103205.0 85210.0 103910.0 86555.0 ;
      RECT  103205.0 87900.0 103910.0 86555.0 ;
      RECT  103205.0 87900.0 103910.0 89245.0 ;
      RECT  103205.0 90590.0 103910.0 89245.0 ;
      RECT  103205.0 90590.0 103910.0 91935.0 ;
      RECT  103205.0 93280.0 103910.0 91935.0 ;
      RECT  103205.0 93280.0 103910.0 94625.0 ;
      RECT  103205.0 95970.0 103910.0 94625.0 ;
      RECT  103205.0 95970.0 103910.0 97315.0 ;
      RECT  103205.0 98660.0 103910.0 97315.0 ;
      RECT  103205.0 98660.0 103910.0 100005.0 ;
      RECT  103205.0 101350.0 103910.0 100005.0 ;
      RECT  103205.0 101350.0 103910.0 102695.0 ;
      RECT  103205.0 104040.0 103910.0 102695.0 ;
      RECT  103205.0 104040.0 103910.0 105385.0 ;
      RECT  103205.0 106730.0 103910.0 105385.0 ;
      RECT  103205.0 106730.0 103910.0 108075.0 ;
      RECT  103205.0 109420.0 103910.0 108075.0 ;
      RECT  103205.0 109420.0 103910.0 110765.0 ;
      RECT  103205.0 112110.0 103910.0 110765.0 ;
      RECT  103205.0 112110.0 103910.0 113455.0 ;
      RECT  103205.0 114800.0 103910.0 113455.0 ;
      RECT  103205.0 114800.0 103910.0 116145.0 ;
      RECT  103205.0 117490.0 103910.0 116145.0 ;
      RECT  103205.0 117490.0 103910.0 118835.0 ;
      RECT  103205.0 120180.0 103910.0 118835.0 ;
      RECT  103205.0 120180.0 103910.0 121525.0 ;
      RECT  103205.0 122870.0 103910.0 121525.0 ;
      RECT  103205.0 122870.0 103910.0 124215.0 ;
      RECT  103205.0 125560.0 103910.0 124215.0 ;
      RECT  103205.0 125560.0 103910.0 126905.0 ;
      RECT  103205.0 128250.0 103910.0 126905.0 ;
      RECT  103205.0 128250.0 103910.0 129595.0 ;
      RECT  103205.0 130940.0 103910.0 129595.0 ;
      RECT  103205.0 130940.0 103910.0 132285.0 ;
      RECT  103205.0 133630.0 103910.0 132285.0 ;
      RECT  103205.0 133630.0 103910.0 134975.0 ;
      RECT  103205.0 136320.0 103910.0 134975.0 ;
      RECT  103205.0 136320.0 103910.0 137665.0 ;
      RECT  103205.0 139010.0 103910.0 137665.0 ;
      RECT  103205.0 139010.0 103910.0 140355.0 ;
      RECT  103205.0 141700.0 103910.0 140355.0 ;
      RECT  103205.0 141700.0 103910.0 143045.0 ;
      RECT  103205.0 144390.0 103910.0 143045.0 ;
      RECT  103205.0 144390.0 103910.0 145735.0 ;
      RECT  103205.0 147080.0 103910.0 145735.0 ;
      RECT  103205.0 147080.0 103910.0 148425.0 ;
      RECT  103205.0 149770.0 103910.0 148425.0 ;
      RECT  103205.0 149770.0 103910.0 151115.0 ;
      RECT  103205.0 152460.0 103910.0 151115.0 ;
      RECT  103205.0 152460.0 103910.0 153805.0 ;
      RECT  103205.0 155150.0 103910.0 153805.0 ;
      RECT  103205.0 155150.0 103910.0 156495.0 ;
      RECT  103205.0 157840.0 103910.0 156495.0 ;
      RECT  103205.0 157840.0 103910.0 159185.0 ;
      RECT  103205.0 160530.0 103910.0 159185.0 ;
      RECT  103205.0 160530.0 103910.0 161875.0 ;
      RECT  103205.0 163220.0 103910.0 161875.0 ;
      RECT  103205.0 163220.0 103910.0 164565.0 ;
      RECT  103205.0 165910.0 103910.0 164565.0 ;
      RECT  103205.0 165910.0 103910.0 167255.0 ;
      RECT  103205.0 168600.0 103910.0 167255.0 ;
      RECT  103205.0 168600.0 103910.0 169945.0 ;
      RECT  103205.0 171290.0 103910.0 169945.0 ;
      RECT  103205.0 171290.0 103910.0 172635.0 ;
      RECT  103205.0 173980.0 103910.0 172635.0 ;
      RECT  103205.0 173980.0 103910.0 175325.0 ;
      RECT  103205.0 176670.0 103910.0 175325.0 ;
      RECT  103205.0 176670.0 103910.0 178015.0 ;
      RECT  103205.0 179360.0 103910.0 178015.0 ;
      RECT  103205.0 179360.0 103910.0 180705.0 ;
      RECT  103205.0 182050.0 103910.0 180705.0 ;
      RECT  103205.0 182050.0 103910.0 183395.0 ;
      RECT  103205.0 184740.0 103910.0 183395.0 ;
      RECT  103205.0 184740.0 103910.0 186085.0 ;
      RECT  103205.0 187430.0 103910.0 186085.0 ;
      RECT  103205.0 187430.0 103910.0 188775.0 ;
      RECT  103205.0 190120.0 103910.0 188775.0 ;
      RECT  103205.0 190120.0 103910.0 191465.0 ;
      RECT  103205.0 192810.0 103910.0 191465.0 ;
      RECT  103205.0 192810.0 103910.0 194155.0 ;
      RECT  103205.0 195500.0 103910.0 194155.0 ;
      RECT  103205.0 195500.0 103910.0 196845.0 ;
      RECT  103205.0 198190.0 103910.0 196845.0 ;
      RECT  103205.0 198190.0 103910.0 199535.0 ;
      RECT  103205.0 200880.0 103910.0 199535.0 ;
      RECT  103205.0 200880.0 103910.0 202225.0 ;
      RECT  103205.0 203570.0 103910.0 202225.0 ;
      RECT  103205.0 203570.0 103910.0 204915.0 ;
      RECT  103205.0 206260.0 103910.0 204915.0 ;
      RECT  103910.0 34100.0 104615.0 35445.0 ;
      RECT  103910.0 36790.0 104615.0 35445.0 ;
      RECT  103910.0 36790.0 104615.0 38135.0 ;
      RECT  103910.0 39480.0 104615.0 38135.0 ;
      RECT  103910.0 39480.0 104615.0 40825.0 ;
      RECT  103910.0 42170.0 104615.0 40825.0 ;
      RECT  103910.0 42170.0 104615.0 43515.0 ;
      RECT  103910.0 44860.0 104615.0 43515.0 ;
      RECT  103910.0 44860.0 104615.0 46205.0 ;
      RECT  103910.0 47550.0 104615.0 46205.0 ;
      RECT  103910.0 47550.0 104615.0 48895.0 ;
      RECT  103910.0 50240.0 104615.0 48895.0 ;
      RECT  103910.0 50240.0 104615.0 51585.0 ;
      RECT  103910.0 52930.0 104615.0 51585.0 ;
      RECT  103910.0 52930.0 104615.0 54275.0 ;
      RECT  103910.0 55620.0 104615.0 54275.0 ;
      RECT  103910.0 55620.0 104615.0 56965.0 ;
      RECT  103910.0 58310.0 104615.0 56965.0 ;
      RECT  103910.0 58310.0 104615.0 59655.0 ;
      RECT  103910.0 61000.0 104615.0 59655.0 ;
      RECT  103910.0 61000.0 104615.0 62345.0 ;
      RECT  103910.0 63690.0 104615.0 62345.0 ;
      RECT  103910.0 63690.0 104615.0 65035.0 ;
      RECT  103910.0 66380.0 104615.0 65035.0 ;
      RECT  103910.0 66380.0 104615.0 67725.0 ;
      RECT  103910.0 69070.0 104615.0 67725.0 ;
      RECT  103910.0 69070.0 104615.0 70415.0 ;
      RECT  103910.0 71760.0 104615.0 70415.0 ;
      RECT  103910.0 71760.0 104615.0 73105.0 ;
      RECT  103910.0 74450.0 104615.0 73105.0 ;
      RECT  103910.0 74450.0 104615.0 75795.0 ;
      RECT  103910.0 77140.0 104615.0 75795.0 ;
      RECT  103910.0 77140.0 104615.0 78485.0 ;
      RECT  103910.0 79830.0 104615.0 78485.0 ;
      RECT  103910.0 79830.0 104615.0 81175.0 ;
      RECT  103910.0 82520.0 104615.0 81175.0 ;
      RECT  103910.0 82520.0 104615.0 83865.0 ;
      RECT  103910.0 85210.0 104615.0 83865.0 ;
      RECT  103910.0 85210.0 104615.0 86555.0 ;
      RECT  103910.0 87900.0 104615.0 86555.0 ;
      RECT  103910.0 87900.0 104615.0 89245.0 ;
      RECT  103910.0 90590.0 104615.0 89245.0 ;
      RECT  103910.0 90590.0 104615.0 91935.0 ;
      RECT  103910.0 93280.0 104615.0 91935.0 ;
      RECT  103910.0 93280.0 104615.0 94625.0 ;
      RECT  103910.0 95970.0 104615.0 94625.0 ;
      RECT  103910.0 95970.0 104615.0 97315.0 ;
      RECT  103910.0 98660.0 104615.0 97315.0 ;
      RECT  103910.0 98660.0 104615.0 100005.0 ;
      RECT  103910.0 101350.0 104615.0 100005.0 ;
      RECT  103910.0 101350.0 104615.0 102695.0 ;
      RECT  103910.0 104040.0 104615.0 102695.0 ;
      RECT  103910.0 104040.0 104615.0 105385.0 ;
      RECT  103910.0 106730.0 104615.0 105385.0 ;
      RECT  103910.0 106730.0 104615.0 108075.0 ;
      RECT  103910.0 109420.0 104615.0 108075.0 ;
      RECT  103910.0 109420.0 104615.0 110765.0 ;
      RECT  103910.0 112110.0 104615.0 110765.0 ;
      RECT  103910.0 112110.0 104615.0 113455.0 ;
      RECT  103910.0 114800.0 104615.0 113455.0 ;
      RECT  103910.0 114800.0 104615.0 116145.0 ;
      RECT  103910.0 117490.0 104615.0 116145.0 ;
      RECT  103910.0 117490.0 104615.0 118835.0 ;
      RECT  103910.0 120180.0 104615.0 118835.0 ;
      RECT  103910.0 120180.0 104615.0 121525.0 ;
      RECT  103910.0 122870.0 104615.0 121525.0 ;
      RECT  103910.0 122870.0 104615.0 124215.0 ;
      RECT  103910.0 125560.0 104615.0 124215.0 ;
      RECT  103910.0 125560.0 104615.0 126905.0 ;
      RECT  103910.0 128250.0 104615.0 126905.0 ;
      RECT  103910.0 128250.0 104615.0 129595.0 ;
      RECT  103910.0 130940.0 104615.0 129595.0 ;
      RECT  103910.0 130940.0 104615.0 132285.0 ;
      RECT  103910.0 133630.0 104615.0 132285.0 ;
      RECT  103910.0 133630.0 104615.0 134975.0 ;
      RECT  103910.0 136320.0 104615.0 134975.0 ;
      RECT  103910.0 136320.0 104615.0 137665.0 ;
      RECT  103910.0 139010.0 104615.0 137665.0 ;
      RECT  103910.0 139010.0 104615.0 140355.0 ;
      RECT  103910.0 141700.0 104615.0 140355.0 ;
      RECT  103910.0 141700.0 104615.0 143045.0 ;
      RECT  103910.0 144390.0 104615.0 143045.0 ;
      RECT  103910.0 144390.0 104615.0 145735.0 ;
      RECT  103910.0 147080.0 104615.0 145735.0 ;
      RECT  103910.0 147080.0 104615.0 148425.0 ;
      RECT  103910.0 149770.0 104615.0 148425.0 ;
      RECT  103910.0 149770.0 104615.0 151115.0 ;
      RECT  103910.0 152460.0 104615.0 151115.0 ;
      RECT  103910.0 152460.0 104615.0 153805.0 ;
      RECT  103910.0 155150.0 104615.0 153805.0 ;
      RECT  103910.0 155150.0 104615.0 156495.0 ;
      RECT  103910.0 157840.0 104615.0 156495.0 ;
      RECT  103910.0 157840.0 104615.0 159185.0 ;
      RECT  103910.0 160530.0 104615.0 159185.0 ;
      RECT  103910.0 160530.0 104615.0 161875.0 ;
      RECT  103910.0 163220.0 104615.0 161875.0 ;
      RECT  103910.0 163220.0 104615.0 164565.0 ;
      RECT  103910.0 165910.0 104615.0 164565.0 ;
      RECT  103910.0 165910.0 104615.0 167255.0 ;
      RECT  103910.0 168600.0 104615.0 167255.0 ;
      RECT  103910.0 168600.0 104615.0 169945.0 ;
      RECT  103910.0 171290.0 104615.0 169945.0 ;
      RECT  103910.0 171290.0 104615.0 172635.0 ;
      RECT  103910.0 173980.0 104615.0 172635.0 ;
      RECT  103910.0 173980.0 104615.0 175325.0 ;
      RECT  103910.0 176670.0 104615.0 175325.0 ;
      RECT  103910.0 176670.0 104615.0 178015.0 ;
      RECT  103910.0 179360.0 104615.0 178015.0 ;
      RECT  103910.0 179360.0 104615.0 180705.0 ;
      RECT  103910.0 182050.0 104615.0 180705.0 ;
      RECT  103910.0 182050.0 104615.0 183395.0 ;
      RECT  103910.0 184740.0 104615.0 183395.0 ;
      RECT  103910.0 184740.0 104615.0 186085.0 ;
      RECT  103910.0 187430.0 104615.0 186085.0 ;
      RECT  103910.0 187430.0 104615.0 188775.0 ;
      RECT  103910.0 190120.0 104615.0 188775.0 ;
      RECT  103910.0 190120.0 104615.0 191465.0 ;
      RECT  103910.0 192810.0 104615.0 191465.0 ;
      RECT  103910.0 192810.0 104615.0 194155.0 ;
      RECT  103910.0 195500.0 104615.0 194155.0 ;
      RECT  103910.0 195500.0 104615.0 196845.0 ;
      RECT  103910.0 198190.0 104615.0 196845.0 ;
      RECT  103910.0 198190.0 104615.0 199535.0 ;
      RECT  103910.0 200880.0 104615.0 199535.0 ;
      RECT  103910.0 200880.0 104615.0 202225.0 ;
      RECT  103910.0 203570.0 104615.0 202225.0 ;
      RECT  103910.0 203570.0 104615.0 204915.0 ;
      RECT  103910.0 206260.0 104615.0 204915.0 ;
      RECT  104615.0 34100.0 105320.0 35445.0 ;
      RECT  104615.0 36790.0 105320.0 35445.0 ;
      RECT  104615.0 36790.0 105320.0 38135.0 ;
      RECT  104615.0 39480.0 105320.0 38135.0 ;
      RECT  104615.0 39480.0 105320.0 40825.0 ;
      RECT  104615.0 42170.0 105320.0 40825.0 ;
      RECT  104615.0 42170.0 105320.0 43515.0 ;
      RECT  104615.0 44860.0 105320.0 43515.0 ;
      RECT  104615.0 44860.0 105320.0 46205.0 ;
      RECT  104615.0 47550.0 105320.0 46205.0 ;
      RECT  104615.0 47550.0 105320.0 48895.0 ;
      RECT  104615.0 50240.0 105320.0 48895.0 ;
      RECT  104615.0 50240.0 105320.0 51585.0 ;
      RECT  104615.0 52930.0 105320.0 51585.0 ;
      RECT  104615.0 52930.0 105320.0 54275.0 ;
      RECT  104615.0 55620.0 105320.0 54275.0 ;
      RECT  104615.0 55620.0 105320.0 56965.0 ;
      RECT  104615.0 58310.0 105320.0 56965.0 ;
      RECT  104615.0 58310.0 105320.0 59655.0 ;
      RECT  104615.0 61000.0 105320.0 59655.0 ;
      RECT  104615.0 61000.0 105320.0 62345.0 ;
      RECT  104615.0 63690.0 105320.0 62345.0 ;
      RECT  104615.0 63690.0 105320.0 65035.0 ;
      RECT  104615.0 66380.0 105320.0 65035.0 ;
      RECT  104615.0 66380.0 105320.0 67725.0 ;
      RECT  104615.0 69070.0 105320.0 67725.0 ;
      RECT  104615.0 69070.0 105320.0 70415.0 ;
      RECT  104615.0 71760.0 105320.0 70415.0 ;
      RECT  104615.0 71760.0 105320.0 73105.0 ;
      RECT  104615.0 74450.0 105320.0 73105.0 ;
      RECT  104615.0 74450.0 105320.0 75795.0 ;
      RECT  104615.0 77140.0 105320.0 75795.0 ;
      RECT  104615.0 77140.0 105320.0 78485.0 ;
      RECT  104615.0 79830.0 105320.0 78485.0 ;
      RECT  104615.0 79830.0 105320.0 81175.0 ;
      RECT  104615.0 82520.0 105320.0 81175.0 ;
      RECT  104615.0 82520.0 105320.0 83865.0 ;
      RECT  104615.0 85210.0 105320.0 83865.0 ;
      RECT  104615.0 85210.0 105320.0 86555.0 ;
      RECT  104615.0 87900.0 105320.0 86555.0 ;
      RECT  104615.0 87900.0 105320.0 89245.0 ;
      RECT  104615.0 90590.0 105320.0 89245.0 ;
      RECT  104615.0 90590.0 105320.0 91935.0 ;
      RECT  104615.0 93280.0 105320.0 91935.0 ;
      RECT  104615.0 93280.0 105320.0 94625.0 ;
      RECT  104615.0 95970.0 105320.0 94625.0 ;
      RECT  104615.0 95970.0 105320.0 97315.0 ;
      RECT  104615.0 98660.0 105320.0 97315.0 ;
      RECT  104615.0 98660.0 105320.0 100005.0 ;
      RECT  104615.0 101350.0 105320.0 100005.0 ;
      RECT  104615.0 101350.0 105320.0 102695.0 ;
      RECT  104615.0 104040.0 105320.0 102695.0 ;
      RECT  104615.0 104040.0 105320.0 105385.0 ;
      RECT  104615.0 106730.0 105320.0 105385.0 ;
      RECT  104615.0 106730.0 105320.0 108075.0 ;
      RECT  104615.0 109420.0 105320.0 108075.0 ;
      RECT  104615.0 109420.0 105320.0 110765.0 ;
      RECT  104615.0 112110.0 105320.0 110765.0 ;
      RECT  104615.0 112110.0 105320.0 113455.0 ;
      RECT  104615.0 114800.0 105320.0 113455.0 ;
      RECT  104615.0 114800.0 105320.0 116145.0 ;
      RECT  104615.0 117490.0 105320.0 116145.0 ;
      RECT  104615.0 117490.0 105320.0 118835.0 ;
      RECT  104615.0 120180.0 105320.0 118835.0 ;
      RECT  104615.0 120180.0 105320.0 121525.0 ;
      RECT  104615.0 122870.0 105320.0 121525.0 ;
      RECT  104615.0 122870.0 105320.0 124215.0 ;
      RECT  104615.0 125560.0 105320.0 124215.0 ;
      RECT  104615.0 125560.0 105320.0 126905.0 ;
      RECT  104615.0 128250.0 105320.0 126905.0 ;
      RECT  104615.0 128250.0 105320.0 129595.0 ;
      RECT  104615.0 130940.0 105320.0 129595.0 ;
      RECT  104615.0 130940.0 105320.0 132285.0 ;
      RECT  104615.0 133630.0 105320.0 132285.0 ;
      RECT  104615.0 133630.0 105320.0 134975.0 ;
      RECT  104615.0 136320.0 105320.0 134975.0 ;
      RECT  104615.0 136320.0 105320.0 137665.0 ;
      RECT  104615.0 139010.0 105320.0 137665.0 ;
      RECT  104615.0 139010.0 105320.0 140355.0 ;
      RECT  104615.0 141700.0 105320.0 140355.0 ;
      RECT  104615.0 141700.0 105320.0 143045.0 ;
      RECT  104615.0 144390.0 105320.0 143045.0 ;
      RECT  104615.0 144390.0 105320.0 145735.0 ;
      RECT  104615.0 147080.0 105320.0 145735.0 ;
      RECT  104615.0 147080.0 105320.0 148425.0 ;
      RECT  104615.0 149770.0 105320.0 148425.0 ;
      RECT  104615.0 149770.0 105320.0 151115.0 ;
      RECT  104615.0 152460.0 105320.0 151115.0 ;
      RECT  104615.0 152460.0 105320.0 153805.0 ;
      RECT  104615.0 155150.0 105320.0 153805.0 ;
      RECT  104615.0 155150.0 105320.0 156495.0 ;
      RECT  104615.0 157840.0 105320.0 156495.0 ;
      RECT  104615.0 157840.0 105320.0 159185.0 ;
      RECT  104615.0 160530.0 105320.0 159185.0 ;
      RECT  104615.0 160530.0 105320.0 161875.0 ;
      RECT  104615.0 163220.0 105320.0 161875.0 ;
      RECT  104615.0 163220.0 105320.0 164565.0 ;
      RECT  104615.0 165910.0 105320.0 164565.0 ;
      RECT  104615.0 165910.0 105320.0 167255.0 ;
      RECT  104615.0 168600.0 105320.0 167255.0 ;
      RECT  104615.0 168600.0 105320.0 169945.0 ;
      RECT  104615.0 171290.0 105320.0 169945.0 ;
      RECT  104615.0 171290.0 105320.0 172635.0 ;
      RECT  104615.0 173980.0 105320.0 172635.0 ;
      RECT  104615.0 173980.0 105320.0 175325.0 ;
      RECT  104615.0 176670.0 105320.0 175325.0 ;
      RECT  104615.0 176670.0 105320.0 178015.0 ;
      RECT  104615.0 179360.0 105320.0 178015.0 ;
      RECT  104615.0 179360.0 105320.0 180705.0 ;
      RECT  104615.0 182050.0 105320.0 180705.0 ;
      RECT  104615.0 182050.0 105320.0 183395.0 ;
      RECT  104615.0 184740.0 105320.0 183395.0 ;
      RECT  104615.0 184740.0 105320.0 186085.0 ;
      RECT  104615.0 187430.0 105320.0 186085.0 ;
      RECT  104615.0 187430.0 105320.0 188775.0 ;
      RECT  104615.0 190120.0 105320.0 188775.0 ;
      RECT  104615.0 190120.0 105320.0 191465.0 ;
      RECT  104615.0 192810.0 105320.0 191465.0 ;
      RECT  104615.0 192810.0 105320.0 194155.0 ;
      RECT  104615.0 195500.0 105320.0 194155.0 ;
      RECT  104615.0 195500.0 105320.0 196845.0 ;
      RECT  104615.0 198190.0 105320.0 196845.0 ;
      RECT  104615.0 198190.0 105320.0 199535.0 ;
      RECT  104615.0 200880.0 105320.0 199535.0 ;
      RECT  104615.0 200880.0 105320.0 202225.0 ;
      RECT  104615.0 203570.0 105320.0 202225.0 ;
      RECT  104615.0 203570.0 105320.0 204915.0 ;
      RECT  104615.0 206260.0 105320.0 204915.0 ;
      RECT  105320.0 34100.0 106025.0 35445.0 ;
      RECT  105320.0 36790.0 106025.0 35445.0 ;
      RECT  105320.0 36790.0 106025.0 38135.0 ;
      RECT  105320.0 39480.0 106025.0 38135.0 ;
      RECT  105320.0 39480.0 106025.0 40825.0 ;
      RECT  105320.0 42170.0 106025.0 40825.0 ;
      RECT  105320.0 42170.0 106025.0 43515.0 ;
      RECT  105320.0 44860.0 106025.0 43515.0 ;
      RECT  105320.0 44860.0 106025.0 46205.0 ;
      RECT  105320.0 47550.0 106025.0 46205.0 ;
      RECT  105320.0 47550.0 106025.0 48895.0 ;
      RECT  105320.0 50240.0 106025.0 48895.0 ;
      RECT  105320.0 50240.0 106025.0 51585.0 ;
      RECT  105320.0 52930.0 106025.0 51585.0 ;
      RECT  105320.0 52930.0 106025.0 54275.0 ;
      RECT  105320.0 55620.0 106025.0 54275.0 ;
      RECT  105320.0 55620.0 106025.0 56965.0 ;
      RECT  105320.0 58310.0 106025.0 56965.0 ;
      RECT  105320.0 58310.0 106025.0 59655.0 ;
      RECT  105320.0 61000.0 106025.0 59655.0 ;
      RECT  105320.0 61000.0 106025.0 62345.0 ;
      RECT  105320.0 63690.0 106025.0 62345.0 ;
      RECT  105320.0 63690.0 106025.0 65035.0 ;
      RECT  105320.0 66380.0 106025.0 65035.0 ;
      RECT  105320.0 66380.0 106025.0 67725.0 ;
      RECT  105320.0 69070.0 106025.0 67725.0 ;
      RECT  105320.0 69070.0 106025.0 70415.0 ;
      RECT  105320.0 71760.0 106025.0 70415.0 ;
      RECT  105320.0 71760.0 106025.0 73105.0 ;
      RECT  105320.0 74450.0 106025.0 73105.0 ;
      RECT  105320.0 74450.0 106025.0 75795.0 ;
      RECT  105320.0 77140.0 106025.0 75795.0 ;
      RECT  105320.0 77140.0 106025.0 78485.0 ;
      RECT  105320.0 79830.0 106025.0 78485.0 ;
      RECT  105320.0 79830.0 106025.0 81175.0 ;
      RECT  105320.0 82520.0 106025.0 81175.0 ;
      RECT  105320.0 82520.0 106025.0 83865.0 ;
      RECT  105320.0 85210.0 106025.0 83865.0 ;
      RECT  105320.0 85210.0 106025.0 86555.0 ;
      RECT  105320.0 87900.0 106025.0 86555.0 ;
      RECT  105320.0 87900.0 106025.0 89245.0 ;
      RECT  105320.0 90590.0 106025.0 89245.0 ;
      RECT  105320.0 90590.0 106025.0 91935.0 ;
      RECT  105320.0 93280.0 106025.0 91935.0 ;
      RECT  105320.0 93280.0 106025.0 94625.0 ;
      RECT  105320.0 95970.0 106025.0 94625.0 ;
      RECT  105320.0 95970.0 106025.0 97315.0 ;
      RECT  105320.0 98660.0 106025.0 97315.0 ;
      RECT  105320.0 98660.0 106025.0 100005.0 ;
      RECT  105320.0 101350.0 106025.0 100005.0 ;
      RECT  105320.0 101350.0 106025.0 102695.0 ;
      RECT  105320.0 104040.0 106025.0 102695.0 ;
      RECT  105320.0 104040.0 106025.0 105385.0 ;
      RECT  105320.0 106730.0 106025.0 105385.0 ;
      RECT  105320.0 106730.0 106025.0 108075.0 ;
      RECT  105320.0 109420.0 106025.0 108075.0 ;
      RECT  105320.0 109420.0 106025.0 110765.0 ;
      RECT  105320.0 112110.0 106025.0 110765.0 ;
      RECT  105320.0 112110.0 106025.0 113455.0 ;
      RECT  105320.0 114800.0 106025.0 113455.0 ;
      RECT  105320.0 114800.0 106025.0 116145.0 ;
      RECT  105320.0 117490.0 106025.0 116145.0 ;
      RECT  105320.0 117490.0 106025.0 118835.0 ;
      RECT  105320.0 120180.0 106025.0 118835.0 ;
      RECT  105320.0 120180.0 106025.0 121525.0 ;
      RECT  105320.0 122870.0 106025.0 121525.0 ;
      RECT  105320.0 122870.0 106025.0 124215.0 ;
      RECT  105320.0 125560.0 106025.0 124215.0 ;
      RECT  105320.0 125560.0 106025.0 126905.0 ;
      RECT  105320.0 128250.0 106025.0 126905.0 ;
      RECT  105320.0 128250.0 106025.0 129595.0 ;
      RECT  105320.0 130940.0 106025.0 129595.0 ;
      RECT  105320.0 130940.0 106025.0 132285.0 ;
      RECT  105320.0 133630.0 106025.0 132285.0 ;
      RECT  105320.0 133630.0 106025.0 134975.0 ;
      RECT  105320.0 136320.0 106025.0 134975.0 ;
      RECT  105320.0 136320.0 106025.0 137665.0 ;
      RECT  105320.0 139010.0 106025.0 137665.0 ;
      RECT  105320.0 139010.0 106025.0 140355.0 ;
      RECT  105320.0 141700.0 106025.0 140355.0 ;
      RECT  105320.0 141700.0 106025.0 143045.0 ;
      RECT  105320.0 144390.0 106025.0 143045.0 ;
      RECT  105320.0 144390.0 106025.0 145735.0 ;
      RECT  105320.0 147080.0 106025.0 145735.0 ;
      RECT  105320.0 147080.0 106025.0 148425.0 ;
      RECT  105320.0 149770.0 106025.0 148425.0 ;
      RECT  105320.0 149770.0 106025.0 151115.0 ;
      RECT  105320.0 152460.0 106025.0 151115.0 ;
      RECT  105320.0 152460.0 106025.0 153805.0 ;
      RECT  105320.0 155150.0 106025.0 153805.0 ;
      RECT  105320.0 155150.0 106025.0 156495.0 ;
      RECT  105320.0 157840.0 106025.0 156495.0 ;
      RECT  105320.0 157840.0 106025.0 159185.0 ;
      RECT  105320.0 160530.0 106025.0 159185.0 ;
      RECT  105320.0 160530.0 106025.0 161875.0 ;
      RECT  105320.0 163220.0 106025.0 161875.0 ;
      RECT  105320.0 163220.0 106025.0 164565.0 ;
      RECT  105320.0 165910.0 106025.0 164565.0 ;
      RECT  105320.0 165910.0 106025.0 167255.0 ;
      RECT  105320.0 168600.0 106025.0 167255.0 ;
      RECT  105320.0 168600.0 106025.0 169945.0 ;
      RECT  105320.0 171290.0 106025.0 169945.0 ;
      RECT  105320.0 171290.0 106025.0 172635.0 ;
      RECT  105320.0 173980.0 106025.0 172635.0 ;
      RECT  105320.0 173980.0 106025.0 175325.0 ;
      RECT  105320.0 176670.0 106025.0 175325.0 ;
      RECT  105320.0 176670.0 106025.0 178015.0 ;
      RECT  105320.0 179360.0 106025.0 178015.0 ;
      RECT  105320.0 179360.0 106025.0 180705.0 ;
      RECT  105320.0 182050.0 106025.0 180705.0 ;
      RECT  105320.0 182050.0 106025.0 183395.0 ;
      RECT  105320.0 184740.0 106025.0 183395.0 ;
      RECT  105320.0 184740.0 106025.0 186085.0 ;
      RECT  105320.0 187430.0 106025.0 186085.0 ;
      RECT  105320.0 187430.0 106025.0 188775.0 ;
      RECT  105320.0 190120.0 106025.0 188775.0 ;
      RECT  105320.0 190120.0 106025.0 191465.0 ;
      RECT  105320.0 192810.0 106025.0 191465.0 ;
      RECT  105320.0 192810.0 106025.0 194155.0 ;
      RECT  105320.0 195500.0 106025.0 194155.0 ;
      RECT  105320.0 195500.0 106025.0 196845.0 ;
      RECT  105320.0 198190.0 106025.0 196845.0 ;
      RECT  105320.0 198190.0 106025.0 199535.0 ;
      RECT  105320.0 200880.0 106025.0 199535.0 ;
      RECT  105320.0 200880.0 106025.0 202225.0 ;
      RECT  105320.0 203570.0 106025.0 202225.0 ;
      RECT  105320.0 203570.0 106025.0 204915.0 ;
      RECT  105320.0 206260.0 106025.0 204915.0 ;
      RECT  106025.0 34100.0 106730.0 35445.0 ;
      RECT  106025.0 36790.0 106730.0 35445.0 ;
      RECT  106025.0 36790.0 106730.0 38135.0 ;
      RECT  106025.0 39480.0 106730.0 38135.0 ;
      RECT  106025.0 39480.0 106730.0 40825.0 ;
      RECT  106025.0 42170.0 106730.0 40825.0 ;
      RECT  106025.0 42170.0 106730.0 43515.0 ;
      RECT  106025.0 44860.0 106730.0 43515.0 ;
      RECT  106025.0 44860.0 106730.0 46205.0 ;
      RECT  106025.0 47550.0 106730.0 46205.0 ;
      RECT  106025.0 47550.0 106730.0 48895.0 ;
      RECT  106025.0 50240.0 106730.0 48895.0 ;
      RECT  106025.0 50240.0 106730.0 51585.0 ;
      RECT  106025.0 52930.0 106730.0 51585.0 ;
      RECT  106025.0 52930.0 106730.0 54275.0 ;
      RECT  106025.0 55620.0 106730.0 54275.0 ;
      RECT  106025.0 55620.0 106730.0 56965.0 ;
      RECT  106025.0 58310.0 106730.0 56965.0 ;
      RECT  106025.0 58310.0 106730.0 59655.0 ;
      RECT  106025.0 61000.0 106730.0 59655.0 ;
      RECT  106025.0 61000.0 106730.0 62345.0 ;
      RECT  106025.0 63690.0 106730.0 62345.0 ;
      RECT  106025.0 63690.0 106730.0 65035.0 ;
      RECT  106025.0 66380.0 106730.0 65035.0 ;
      RECT  106025.0 66380.0 106730.0 67725.0 ;
      RECT  106025.0 69070.0 106730.0 67725.0 ;
      RECT  106025.0 69070.0 106730.0 70415.0 ;
      RECT  106025.0 71760.0 106730.0 70415.0 ;
      RECT  106025.0 71760.0 106730.0 73105.0 ;
      RECT  106025.0 74450.0 106730.0 73105.0 ;
      RECT  106025.0 74450.0 106730.0 75795.0 ;
      RECT  106025.0 77140.0 106730.0 75795.0 ;
      RECT  106025.0 77140.0 106730.0 78485.0 ;
      RECT  106025.0 79830.0 106730.0 78485.0 ;
      RECT  106025.0 79830.0 106730.0 81175.0 ;
      RECT  106025.0 82520.0 106730.0 81175.0 ;
      RECT  106025.0 82520.0 106730.0 83865.0 ;
      RECT  106025.0 85210.0 106730.0 83865.0 ;
      RECT  106025.0 85210.0 106730.0 86555.0 ;
      RECT  106025.0 87900.0 106730.0 86555.0 ;
      RECT  106025.0 87900.0 106730.0 89245.0 ;
      RECT  106025.0 90590.0 106730.0 89245.0 ;
      RECT  106025.0 90590.0 106730.0 91935.0 ;
      RECT  106025.0 93280.0 106730.0 91935.0 ;
      RECT  106025.0 93280.0 106730.0 94625.0 ;
      RECT  106025.0 95970.0 106730.0 94625.0 ;
      RECT  106025.0 95970.0 106730.0 97315.0 ;
      RECT  106025.0 98660.0 106730.0 97315.0 ;
      RECT  106025.0 98660.0 106730.0 100005.0 ;
      RECT  106025.0 101350.0 106730.0 100005.0 ;
      RECT  106025.0 101350.0 106730.0 102695.0 ;
      RECT  106025.0 104040.0 106730.0 102695.0 ;
      RECT  106025.0 104040.0 106730.0 105385.0 ;
      RECT  106025.0 106730.0 106730.0 105385.0 ;
      RECT  106025.0 106730.0 106730.0 108075.0 ;
      RECT  106025.0 109420.0 106730.0 108075.0 ;
      RECT  106025.0 109420.0 106730.0 110765.0 ;
      RECT  106025.0 112110.0 106730.0 110765.0 ;
      RECT  106025.0 112110.0 106730.0 113455.0 ;
      RECT  106025.0 114800.0 106730.0 113455.0 ;
      RECT  106025.0 114800.0 106730.0 116145.0 ;
      RECT  106025.0 117490.0 106730.0 116145.0 ;
      RECT  106025.0 117490.0 106730.0 118835.0 ;
      RECT  106025.0 120180.0 106730.0 118835.0 ;
      RECT  106025.0 120180.0 106730.0 121525.0 ;
      RECT  106025.0 122870.0 106730.0 121525.0 ;
      RECT  106025.0 122870.0 106730.0 124215.0 ;
      RECT  106025.0 125560.0 106730.0 124215.0 ;
      RECT  106025.0 125560.0 106730.0 126905.0 ;
      RECT  106025.0 128250.0 106730.0 126905.0 ;
      RECT  106025.0 128250.0 106730.0 129595.0 ;
      RECT  106025.0 130940.0 106730.0 129595.0 ;
      RECT  106025.0 130940.0 106730.0 132285.0 ;
      RECT  106025.0 133630.0 106730.0 132285.0 ;
      RECT  106025.0 133630.0 106730.0 134975.0 ;
      RECT  106025.0 136320.0 106730.0 134975.0 ;
      RECT  106025.0 136320.0 106730.0 137665.0 ;
      RECT  106025.0 139010.0 106730.0 137665.0 ;
      RECT  106025.0 139010.0 106730.0 140355.0 ;
      RECT  106025.0 141700.0 106730.0 140355.0 ;
      RECT  106025.0 141700.0 106730.0 143045.0 ;
      RECT  106025.0 144390.0 106730.0 143045.0 ;
      RECT  106025.0 144390.0 106730.0 145735.0 ;
      RECT  106025.0 147080.0 106730.0 145735.0 ;
      RECT  106025.0 147080.0 106730.0 148425.0 ;
      RECT  106025.0 149770.0 106730.0 148425.0 ;
      RECT  106025.0 149770.0 106730.0 151115.0 ;
      RECT  106025.0 152460.0 106730.0 151115.0 ;
      RECT  106025.0 152460.0 106730.0 153805.0 ;
      RECT  106025.0 155150.0 106730.0 153805.0 ;
      RECT  106025.0 155150.0 106730.0 156495.0 ;
      RECT  106025.0 157840.0 106730.0 156495.0 ;
      RECT  106025.0 157840.0 106730.0 159185.0 ;
      RECT  106025.0 160530.0 106730.0 159185.0 ;
      RECT  106025.0 160530.0 106730.0 161875.0 ;
      RECT  106025.0 163220.0 106730.0 161875.0 ;
      RECT  106025.0 163220.0 106730.0 164565.0 ;
      RECT  106025.0 165910.0 106730.0 164565.0 ;
      RECT  106025.0 165910.0 106730.0 167255.0 ;
      RECT  106025.0 168600.0 106730.0 167255.0 ;
      RECT  106025.0 168600.0 106730.0 169945.0 ;
      RECT  106025.0 171290.0 106730.0 169945.0 ;
      RECT  106025.0 171290.0 106730.0 172635.0 ;
      RECT  106025.0 173980.0 106730.0 172635.0 ;
      RECT  106025.0 173980.0 106730.0 175325.0 ;
      RECT  106025.0 176670.0 106730.0 175325.0 ;
      RECT  106025.0 176670.0 106730.0 178015.0 ;
      RECT  106025.0 179360.0 106730.0 178015.0 ;
      RECT  106025.0 179360.0 106730.0 180705.0 ;
      RECT  106025.0 182050.0 106730.0 180705.0 ;
      RECT  106025.0 182050.0 106730.0 183395.0 ;
      RECT  106025.0 184740.0 106730.0 183395.0 ;
      RECT  106025.0 184740.0 106730.0 186085.0 ;
      RECT  106025.0 187430.0 106730.0 186085.0 ;
      RECT  106025.0 187430.0 106730.0 188775.0 ;
      RECT  106025.0 190120.0 106730.0 188775.0 ;
      RECT  106025.0 190120.0 106730.0 191465.0 ;
      RECT  106025.0 192810.0 106730.0 191465.0 ;
      RECT  106025.0 192810.0 106730.0 194155.0 ;
      RECT  106025.0 195500.0 106730.0 194155.0 ;
      RECT  106025.0 195500.0 106730.0 196845.0 ;
      RECT  106025.0 198190.0 106730.0 196845.0 ;
      RECT  106025.0 198190.0 106730.0 199535.0 ;
      RECT  106025.0 200880.0 106730.0 199535.0 ;
      RECT  106025.0 200880.0 106730.0 202225.0 ;
      RECT  106025.0 203570.0 106730.0 202225.0 ;
      RECT  106025.0 203570.0 106730.0 204915.0 ;
      RECT  106025.0 206260.0 106730.0 204915.0 ;
      RECT  106730.0 34100.0 107435.0 35445.0 ;
      RECT  106730.0 36790.0 107435.0 35445.0 ;
      RECT  106730.0 36790.0 107435.0 38135.0 ;
      RECT  106730.0 39480.0 107435.0 38135.0 ;
      RECT  106730.0 39480.0 107435.0 40825.0 ;
      RECT  106730.0 42170.0 107435.0 40825.0 ;
      RECT  106730.0 42170.0 107435.0 43515.0 ;
      RECT  106730.0 44860.0 107435.0 43515.0 ;
      RECT  106730.0 44860.0 107435.0 46205.0 ;
      RECT  106730.0 47550.0 107435.0 46205.0 ;
      RECT  106730.0 47550.0 107435.0 48895.0 ;
      RECT  106730.0 50240.0 107435.0 48895.0 ;
      RECT  106730.0 50240.0 107435.0 51585.0 ;
      RECT  106730.0 52930.0 107435.0 51585.0 ;
      RECT  106730.0 52930.0 107435.0 54275.0 ;
      RECT  106730.0 55620.0 107435.0 54275.0 ;
      RECT  106730.0 55620.0 107435.0 56965.0 ;
      RECT  106730.0 58310.0 107435.0 56965.0 ;
      RECT  106730.0 58310.0 107435.0 59655.0 ;
      RECT  106730.0 61000.0 107435.0 59655.0 ;
      RECT  106730.0 61000.0 107435.0 62345.0 ;
      RECT  106730.0 63690.0 107435.0 62345.0 ;
      RECT  106730.0 63690.0 107435.0 65035.0 ;
      RECT  106730.0 66380.0 107435.0 65035.0 ;
      RECT  106730.0 66380.0 107435.0 67725.0 ;
      RECT  106730.0 69070.0 107435.0 67725.0 ;
      RECT  106730.0 69070.0 107435.0 70415.0 ;
      RECT  106730.0 71760.0 107435.0 70415.0 ;
      RECT  106730.0 71760.0 107435.0 73105.0 ;
      RECT  106730.0 74450.0 107435.0 73105.0 ;
      RECT  106730.0 74450.0 107435.0 75795.0 ;
      RECT  106730.0 77140.0 107435.0 75795.0 ;
      RECT  106730.0 77140.0 107435.0 78485.0 ;
      RECT  106730.0 79830.0 107435.0 78485.0 ;
      RECT  106730.0 79830.0 107435.0 81175.0 ;
      RECT  106730.0 82520.0 107435.0 81175.0 ;
      RECT  106730.0 82520.0 107435.0 83865.0 ;
      RECT  106730.0 85210.0 107435.0 83865.0 ;
      RECT  106730.0 85210.0 107435.0 86555.0 ;
      RECT  106730.0 87900.0 107435.0 86555.0 ;
      RECT  106730.0 87900.0 107435.0 89245.0 ;
      RECT  106730.0 90590.0 107435.0 89245.0 ;
      RECT  106730.0 90590.0 107435.0 91935.0 ;
      RECT  106730.0 93280.0 107435.0 91935.0 ;
      RECT  106730.0 93280.0 107435.0 94625.0 ;
      RECT  106730.0 95970.0 107435.0 94625.0 ;
      RECT  106730.0 95970.0 107435.0 97315.0 ;
      RECT  106730.0 98660.0 107435.0 97315.0 ;
      RECT  106730.0 98660.0 107435.0 100005.0 ;
      RECT  106730.0 101350.0 107435.0 100005.0 ;
      RECT  106730.0 101350.0 107435.0 102695.0 ;
      RECT  106730.0 104040.0 107435.0 102695.0 ;
      RECT  106730.0 104040.0 107435.0 105385.0 ;
      RECT  106730.0 106730.0 107435.0 105385.0 ;
      RECT  106730.0 106730.0 107435.0 108075.0 ;
      RECT  106730.0 109420.0 107435.0 108075.0 ;
      RECT  106730.0 109420.0 107435.0 110765.0 ;
      RECT  106730.0 112110.0 107435.0 110765.0 ;
      RECT  106730.0 112110.0 107435.0 113455.0 ;
      RECT  106730.0 114800.0 107435.0 113455.0 ;
      RECT  106730.0 114800.0 107435.0 116145.0 ;
      RECT  106730.0 117490.0 107435.0 116145.0 ;
      RECT  106730.0 117490.0 107435.0 118835.0 ;
      RECT  106730.0 120180.0 107435.0 118835.0 ;
      RECT  106730.0 120180.0 107435.0 121525.0 ;
      RECT  106730.0 122870.0 107435.0 121525.0 ;
      RECT  106730.0 122870.0 107435.0 124215.0 ;
      RECT  106730.0 125560.0 107435.0 124215.0 ;
      RECT  106730.0 125560.0 107435.0 126905.0 ;
      RECT  106730.0 128250.0 107435.0 126905.0 ;
      RECT  106730.0 128250.0 107435.0 129595.0 ;
      RECT  106730.0 130940.0 107435.0 129595.0 ;
      RECT  106730.0 130940.0 107435.0 132285.0 ;
      RECT  106730.0 133630.0 107435.0 132285.0 ;
      RECT  106730.0 133630.0 107435.0 134975.0 ;
      RECT  106730.0 136320.0 107435.0 134975.0 ;
      RECT  106730.0 136320.0 107435.0 137665.0 ;
      RECT  106730.0 139010.0 107435.0 137665.0 ;
      RECT  106730.0 139010.0 107435.0 140355.0 ;
      RECT  106730.0 141700.0 107435.0 140355.0 ;
      RECT  106730.0 141700.0 107435.0 143045.0 ;
      RECT  106730.0 144390.0 107435.0 143045.0 ;
      RECT  106730.0 144390.0 107435.0 145735.0 ;
      RECT  106730.0 147080.0 107435.0 145735.0 ;
      RECT  106730.0 147080.0 107435.0 148425.0 ;
      RECT  106730.0 149770.0 107435.0 148425.0 ;
      RECT  106730.0 149770.0 107435.0 151115.0 ;
      RECT  106730.0 152460.0 107435.0 151115.0 ;
      RECT  106730.0 152460.0 107435.0 153805.0 ;
      RECT  106730.0 155150.0 107435.0 153805.0 ;
      RECT  106730.0 155150.0 107435.0 156495.0 ;
      RECT  106730.0 157840.0 107435.0 156495.0 ;
      RECT  106730.0 157840.0 107435.0 159185.0 ;
      RECT  106730.0 160530.0 107435.0 159185.0 ;
      RECT  106730.0 160530.0 107435.0 161875.0 ;
      RECT  106730.0 163220.0 107435.0 161875.0 ;
      RECT  106730.0 163220.0 107435.0 164565.0 ;
      RECT  106730.0 165910.0 107435.0 164565.0 ;
      RECT  106730.0 165910.0 107435.0 167255.0 ;
      RECT  106730.0 168600.0 107435.0 167255.0 ;
      RECT  106730.0 168600.0 107435.0 169945.0 ;
      RECT  106730.0 171290.0 107435.0 169945.0 ;
      RECT  106730.0 171290.0 107435.0 172635.0 ;
      RECT  106730.0 173980.0 107435.0 172635.0 ;
      RECT  106730.0 173980.0 107435.0 175325.0 ;
      RECT  106730.0 176670.0 107435.0 175325.0 ;
      RECT  106730.0 176670.0 107435.0 178015.0 ;
      RECT  106730.0 179360.0 107435.0 178015.0 ;
      RECT  106730.0 179360.0 107435.0 180705.0 ;
      RECT  106730.0 182050.0 107435.0 180705.0 ;
      RECT  106730.0 182050.0 107435.0 183395.0 ;
      RECT  106730.0 184740.0 107435.0 183395.0 ;
      RECT  106730.0 184740.0 107435.0 186085.0 ;
      RECT  106730.0 187430.0 107435.0 186085.0 ;
      RECT  106730.0 187430.0 107435.0 188775.0 ;
      RECT  106730.0 190120.0 107435.0 188775.0 ;
      RECT  106730.0 190120.0 107435.0 191465.0 ;
      RECT  106730.0 192810.0 107435.0 191465.0 ;
      RECT  106730.0 192810.0 107435.0 194155.0 ;
      RECT  106730.0 195500.0 107435.0 194155.0 ;
      RECT  106730.0 195500.0 107435.0 196845.0 ;
      RECT  106730.0 198190.0 107435.0 196845.0 ;
      RECT  106730.0 198190.0 107435.0 199535.0 ;
      RECT  106730.0 200880.0 107435.0 199535.0 ;
      RECT  106730.0 200880.0 107435.0 202225.0 ;
      RECT  106730.0 203570.0 107435.0 202225.0 ;
      RECT  106730.0 203570.0 107435.0 204915.0 ;
      RECT  106730.0 206260.0 107435.0 204915.0 ;
      RECT  17345.0 34000.0 17415.0 206415.0 ;
      RECT  17680.0 34000.0 17750.0 206415.0 ;
      RECT  18050.0 34000.0 18120.0 206415.0 ;
      RECT  18385.0 34000.0 18455.0 206415.0 ;
      RECT  18755.0 34000.0 18825.0 206415.0 ;
      RECT  19090.0 34000.0 19160.0 206415.0 ;
      RECT  19460.0 34000.0 19530.0 206415.0 ;
      RECT  19795.0 34000.0 19865.0 206415.0 ;
      RECT  20165.0 34000.0 20235.0 206415.0 ;
      RECT  20500.0 34000.0 20570.0 206415.0 ;
      RECT  20870.0 34000.0 20940.0 206415.0 ;
      RECT  21205.0 34000.0 21275.0 206415.0 ;
      RECT  21575.0 34000.0 21645.0 206415.0 ;
      RECT  21910.0 34000.0 21980.0 206415.0 ;
      RECT  22280.0 34000.0 22350.0 206415.0 ;
      RECT  22615.0 34000.0 22685.0 206415.0 ;
      RECT  22985.0 34000.0 23055.0 206415.0 ;
      RECT  23320.0 34000.0 23390.0 206415.0 ;
      RECT  23690.0 34000.0 23760.0 206415.0 ;
      RECT  24025.0 34000.0 24095.0 206415.0 ;
      RECT  24395.0 34000.0 24465.0 206415.0 ;
      RECT  24730.0 34000.0 24800.0 206415.0 ;
      RECT  25100.0 34000.0 25170.0 206415.0 ;
      RECT  25435.0 34000.0 25505.0 206415.0 ;
      RECT  25805.0 34000.0 25875.0 206415.0 ;
      RECT  26140.0 34000.0 26210.0 206415.0 ;
      RECT  26510.0 34000.0 26580.0 206415.0 ;
      RECT  26845.0 34000.0 26915.0 206415.0 ;
      RECT  27215.0 34000.0 27285.0 206415.0 ;
      RECT  27550.0 34000.0 27620.0 206415.0 ;
      RECT  27920.0 34000.0 27990.0 206415.0 ;
      RECT  28255.0 34000.0 28325.0 206415.0 ;
      RECT  28625.0 34000.0 28695.0 206415.0 ;
      RECT  28960.0 34000.0 29030.0 206415.0 ;
      RECT  29330.0 34000.0 29400.0 206415.0 ;
      RECT  29665.0 34000.0 29735.0 206415.0 ;
      RECT  30035.0 34000.0 30105.0 206415.0 ;
      RECT  30370.0 34000.0 30440.0 206415.0 ;
      RECT  30740.0 34000.0 30810.0 206415.0 ;
      RECT  31075.0 34000.0 31145.0 206415.0 ;
      RECT  31445.0 34000.0 31515.0 206415.0 ;
      RECT  31780.0 34000.0 31850.0 206415.0 ;
      RECT  32150.0 34000.0 32220.0 206415.0 ;
      RECT  32485.0 34000.0 32555.0 206415.0 ;
      RECT  32855.0 34000.0 32925.0 206415.0 ;
      RECT  33190.0 34000.0 33260.0 206415.0 ;
      RECT  33560.0 34000.0 33630.0 206415.0 ;
      RECT  33895.0 34000.0 33965.0 206415.0 ;
      RECT  34265.0 34000.0 34335.0 206415.0 ;
      RECT  34600.0 34000.0 34670.0 206415.0 ;
      RECT  34970.0 34000.0 35040.0 206415.0 ;
      RECT  35305.0 34000.0 35375.0 206415.0 ;
      RECT  35675.0 34000.0 35745.0 206415.0 ;
      RECT  36010.0 34000.0 36080.0 206415.0 ;
      RECT  36380.0 34000.0 36450.0 206415.0 ;
      RECT  36715.0 34000.0 36785.0 206415.0 ;
      RECT  37085.0 34000.0 37155.0 206415.0 ;
      RECT  37420.0 34000.0 37490.0 206415.0 ;
      RECT  37790.0 34000.0 37860.0 206415.0 ;
      RECT  38125.0 34000.0 38195.0 206415.0 ;
      RECT  38495.0 34000.0 38565.0 206415.0 ;
      RECT  38830.0 34000.0 38900.0 206415.0 ;
      RECT  39200.0 34000.0 39270.0 206415.0 ;
      RECT  39535.0 34000.0 39605.0 206415.0 ;
      RECT  39905.0 34000.0 39975.0 206415.0 ;
      RECT  40240.0 34000.0 40310.0 206415.0 ;
      RECT  40610.0 34000.0 40680.0 206415.0 ;
      RECT  40945.0 34000.0 41015.0 206415.0 ;
      RECT  41315.0 34000.0 41385.0 206415.0 ;
      RECT  41650.0 34000.0 41720.0 206415.0 ;
      RECT  42020.0 34000.0 42090.0 206415.0 ;
      RECT  42355.0 34000.0 42425.0 206415.0 ;
      RECT  42725.0 34000.0 42795.0 206415.0 ;
      RECT  43060.0 34000.0 43130.0 206415.0 ;
      RECT  43430.0 34000.0 43500.0 206415.0 ;
      RECT  43765.0 34000.0 43835.0 206415.0 ;
      RECT  44135.0 34000.0 44205.0 206415.0 ;
      RECT  44470.0 34000.0 44540.0 206415.0 ;
      RECT  44840.0 34000.0 44910.0 206415.0 ;
      RECT  45175.0 34000.0 45245.0 206415.0 ;
      RECT  45545.0 34000.0 45615.0 206415.0 ;
      RECT  45880.0 34000.0 45950.0 206415.0 ;
      RECT  46250.0 34000.0 46320.0 206415.0 ;
      RECT  46585.0 34000.0 46655.0 206415.0 ;
      RECT  46955.0 34000.0 47025.0 206415.0 ;
      RECT  47290.0 34000.0 47360.0 206415.0 ;
      RECT  47660.0 34000.0 47730.0 206415.0 ;
      RECT  47995.0 34000.0 48065.0 206415.0 ;
      RECT  48365.0 34000.0 48435.0 206415.0 ;
      RECT  48700.0 34000.0 48770.0 206415.0 ;
      RECT  49070.0 34000.0 49140.0 206415.0 ;
      RECT  49405.0 34000.0 49475.0 206415.0 ;
      RECT  49775.0 34000.0 49845.0 206415.0 ;
      RECT  50110.0 34000.0 50180.0 206415.0 ;
      RECT  50480.0 34000.0 50550.0 206415.0 ;
      RECT  50815.0 34000.0 50885.0 206415.0 ;
      RECT  51185.0 34000.0 51255.0 206415.0 ;
      RECT  51520.0 34000.0 51590.0 206415.0 ;
      RECT  51890.0 34000.0 51960.0 206415.0 ;
      RECT  52225.0 34000.0 52295.0 206415.0 ;
      RECT  52595.0 34000.0 52665.0 206415.0 ;
      RECT  52930.0 34000.0 53000.0 206415.0 ;
      RECT  53300.0 34000.0 53370.0 206415.0 ;
      RECT  53635.0 34000.0 53705.0 206415.0 ;
      RECT  54005.0 34000.0 54075.0 206415.0 ;
      RECT  54340.0 34000.0 54410.0 206415.0 ;
      RECT  54710.0 34000.0 54780.0 206415.0 ;
      RECT  55045.0 34000.0 55115.0 206415.0 ;
      RECT  55415.0 34000.0 55485.0 206415.0 ;
      RECT  55750.0 34000.0 55820.0 206415.0 ;
      RECT  56120.0 34000.0 56190.0 206415.0 ;
      RECT  56455.0 34000.0 56525.0 206415.0 ;
      RECT  56825.0 34000.0 56895.0 206415.0 ;
      RECT  57160.0 34000.0 57230.0 206415.0 ;
      RECT  57530.0 34000.0 57600.0 206415.0 ;
      RECT  57865.0 34000.0 57935.0 206415.0 ;
      RECT  58235.0 34000.0 58305.0 206415.0 ;
      RECT  58570.0 34000.0 58640.0 206415.0 ;
      RECT  58940.0 34000.0 59010.0 206415.0 ;
      RECT  59275.0 34000.0 59345.0 206415.0 ;
      RECT  59645.0 34000.0 59715.0 206415.0 ;
      RECT  59980.0 34000.0 60050.0 206415.0 ;
      RECT  60350.0 34000.0 60420.0 206415.0 ;
      RECT  60685.0 34000.0 60755.0 206415.0 ;
      RECT  61055.0 34000.0 61125.0 206415.0 ;
      RECT  61390.0 34000.0 61460.0 206415.0 ;
      RECT  61760.0 34000.0 61830.0 206415.0 ;
      RECT  62095.0 34000.0 62165.0 206415.0 ;
      RECT  62465.0 34000.0 62535.0 206415.0 ;
      RECT  62800.0 34000.0 62870.0 206415.0 ;
      RECT  63170.0 34000.0 63240.0 206415.0 ;
      RECT  63505.0 34000.0 63575.0 206415.0 ;
      RECT  63875.0 34000.0 63945.0 206415.0 ;
      RECT  64210.0 34000.0 64280.0 206415.0 ;
      RECT  64580.0 34000.0 64650.0 206415.0 ;
      RECT  64915.0 34000.0 64985.0 206415.0 ;
      RECT  65285.0 34000.0 65355.0 206415.0 ;
      RECT  65620.0 34000.0 65690.0 206415.0 ;
      RECT  65990.0 34000.0 66060.0 206415.0 ;
      RECT  66325.0 34000.0 66395.0 206415.0 ;
      RECT  66695.0 34000.0 66765.0 206415.0 ;
      RECT  67030.0 34000.0 67100.0 206415.0 ;
      RECT  67400.0 34000.0 67470.0 206415.0 ;
      RECT  67735.0 34000.0 67805.0 206415.0 ;
      RECT  68105.0 34000.0 68175.0 206415.0 ;
      RECT  68440.0 34000.0 68510.0 206415.0 ;
      RECT  68810.0 34000.0 68880.0 206415.0 ;
      RECT  69145.0 34000.0 69215.0 206415.0 ;
      RECT  69515.0 34000.0 69585.0 206415.0 ;
      RECT  69850.0 34000.0 69920.0 206415.0 ;
      RECT  70220.0 34000.0 70290.0 206415.0 ;
      RECT  70555.0 34000.0 70625.0 206415.0 ;
      RECT  70925.0 34000.0 70995.0 206415.0 ;
      RECT  71260.0 34000.0 71330.0 206415.0 ;
      RECT  71630.0 34000.0 71700.0 206415.0 ;
      RECT  71965.0 34000.0 72035.0 206415.0 ;
      RECT  72335.0 34000.0 72405.0 206415.0 ;
      RECT  72670.0 34000.0 72740.0 206415.0 ;
      RECT  73040.0 34000.0 73110.0 206415.0 ;
      RECT  73375.0 34000.0 73445.0 206415.0 ;
      RECT  73745.0 34000.0 73815.0 206415.0 ;
      RECT  74080.0 34000.0 74150.0 206415.0 ;
      RECT  74450.0 34000.0 74520.0 206415.0 ;
      RECT  74785.0 34000.0 74855.0 206415.0 ;
      RECT  75155.0 34000.0 75225.0 206415.0 ;
      RECT  75490.0 34000.0 75560.0 206415.0 ;
      RECT  75860.0 34000.0 75930.0 206415.0 ;
      RECT  76195.0 34000.0 76265.0 206415.0 ;
      RECT  76565.0 34000.0 76635.0 206415.0 ;
      RECT  76900.0 34000.0 76970.0 206415.0 ;
      RECT  77270.0 34000.0 77340.0 206415.0 ;
      RECT  77605.0 34000.0 77675.0 206415.0 ;
      RECT  77975.0 34000.0 78045.0 206415.0 ;
      RECT  78310.0 34000.0 78380.0 206415.0 ;
      RECT  78680.0 34000.0 78750.0 206415.0 ;
      RECT  79015.0 34000.0 79085.0 206415.0 ;
      RECT  79385.0 34000.0 79455.0 206415.0 ;
      RECT  79720.0 34000.0 79790.0 206415.0 ;
      RECT  80090.0 34000.0 80160.0 206415.0 ;
      RECT  80425.0 34000.0 80495.0 206415.0 ;
      RECT  80795.0 34000.0 80865.0 206415.0 ;
      RECT  81130.0 34000.0 81200.0 206415.0 ;
      RECT  81500.0 34000.0 81570.0 206415.0 ;
      RECT  81835.0 34000.0 81905.0 206415.0 ;
      RECT  82205.0 34000.0 82275.0 206415.0 ;
      RECT  82540.0 34000.0 82610.0 206415.0 ;
      RECT  82910.0 34000.0 82980.0 206415.0 ;
      RECT  83245.0 34000.0 83315.0 206415.0 ;
      RECT  83615.0 34000.0 83685.0 206415.0 ;
      RECT  83950.0 34000.0 84020.0 206415.0 ;
      RECT  84320.0 34000.0 84390.0 206415.0 ;
      RECT  84655.0 34000.0 84725.0 206415.0 ;
      RECT  85025.0 34000.0 85095.0 206415.0 ;
      RECT  85360.0 34000.0 85430.0 206415.0 ;
      RECT  85730.0 34000.0 85800.0 206415.0 ;
      RECT  86065.0 34000.0 86135.0 206415.0 ;
      RECT  86435.0 34000.0 86505.0 206415.0 ;
      RECT  86770.0 34000.0 86840.0 206415.0 ;
      RECT  87140.0 34000.0 87210.0 206415.0 ;
      RECT  87475.0 34000.0 87545.0 206415.0 ;
      RECT  87845.0 34000.0 87915.0 206415.0 ;
      RECT  88180.0 34000.0 88250.0 206415.0 ;
      RECT  88550.0 34000.0 88620.0 206415.0 ;
      RECT  88885.0 34000.0 88955.0 206415.0 ;
      RECT  89255.0 34000.0 89325.0 206415.0 ;
      RECT  89590.0 34000.0 89660.0 206415.0 ;
      RECT  89960.0 34000.0 90030.0 206415.0 ;
      RECT  90295.0 34000.0 90365.0 206415.0 ;
      RECT  90665.0 34000.0 90735.0 206415.0 ;
      RECT  91000.0 34000.0 91070.0 206415.0 ;
      RECT  91370.0 34000.0 91440.0 206415.0 ;
      RECT  91705.0 34000.0 91775.0 206415.0 ;
      RECT  92075.0 34000.0 92145.0 206415.0 ;
      RECT  92410.0 34000.0 92480.0 206415.0 ;
      RECT  92780.0 34000.0 92850.0 206415.0 ;
      RECT  93115.0 34000.0 93185.0 206415.0 ;
      RECT  93485.0 34000.0 93555.0 206415.0 ;
      RECT  93820.0 34000.0 93890.0 206415.0 ;
      RECT  94190.0 34000.0 94260.0 206415.0 ;
      RECT  94525.0 34000.0 94595.0 206415.0 ;
      RECT  94895.0 34000.0 94965.0 206415.0 ;
      RECT  95230.0 34000.0 95300.0 206415.0 ;
      RECT  95600.0 34000.0 95670.0 206415.0 ;
      RECT  95935.0 34000.0 96005.0 206415.0 ;
      RECT  96305.0 34000.0 96375.0 206415.0 ;
      RECT  96640.0 34000.0 96710.0 206415.0 ;
      RECT  97010.0 34000.0 97080.0 206415.0 ;
      RECT  97345.0 34000.0 97415.0 206415.0 ;
      RECT  97715.0 34000.0 97785.0 206415.0 ;
      RECT  98050.0 34000.0 98120.0 206415.0 ;
      RECT  98420.0 34000.0 98490.0 206415.0 ;
      RECT  98755.0 34000.0 98825.0 206415.0 ;
      RECT  99125.0 34000.0 99195.0 206415.0 ;
      RECT  99460.0 34000.0 99530.0 206415.0 ;
      RECT  99830.0 34000.0 99900.0 206415.0 ;
      RECT  100165.0 34000.0 100235.0 206415.0 ;
      RECT  100535.0 34000.0 100605.0 206415.0 ;
      RECT  100870.0 34000.0 100940.0 206415.0 ;
      RECT  101240.0 34000.0 101310.0 206415.0 ;
      RECT  101575.0 34000.0 101645.0 206415.0 ;
      RECT  101945.0 34000.0 102015.0 206415.0 ;
      RECT  102280.0 34000.0 102350.0 206415.0 ;
      RECT  102650.0 34000.0 102720.0 206415.0 ;
      RECT  102985.0 34000.0 103055.0 206415.0 ;
      RECT  103355.0 34000.0 103425.0 206415.0 ;
      RECT  103690.0 34000.0 103760.0 206415.0 ;
      RECT  104060.0 34000.0 104130.0 206415.0 ;
      RECT  104395.0 34000.0 104465.0 206415.0 ;
      RECT  104765.0 34000.0 104835.0 206415.0 ;
      RECT  105100.0 34000.0 105170.0 206415.0 ;
      RECT  105470.0 34000.0 105540.0 206415.0 ;
      RECT  105805.0 34000.0 105875.0 206415.0 ;
      RECT  106175.0 34000.0 106245.0 206415.0 ;
      RECT  106510.0 34000.0 106580.0 206415.0 ;
      RECT  106880.0 34000.0 106950.0 206415.0 ;
      RECT  107215.0 34000.0 107285.0 206415.0 ;
      RECT  17160.0 34000.0 17230.0 206415.0 ;
      RECT  17865.0 34000.0 17935.0 206415.0 ;
      RECT  18570.0 34000.0 18640.0 206415.0 ;
      RECT  19275.0 34000.0 19345.0 206415.0 ;
      RECT  19980.0 34000.0 20050.0 206415.0 ;
      RECT  20685.0 34000.0 20755.0 206415.0 ;
      RECT  21390.0 34000.0 21460.0 206415.0 ;
      RECT  22095.0 34000.0 22165.0 206415.0 ;
      RECT  22800.0 34000.0 22870.0 206415.0 ;
      RECT  23505.0 34000.0 23575.0 206415.0 ;
      RECT  24210.0 34000.0 24280.0 206415.0 ;
      RECT  24915.0 34000.0 24985.0 206415.0 ;
      RECT  25620.0 34000.0 25690.0 206415.0 ;
      RECT  26325.0 34000.0 26395.0 206415.0 ;
      RECT  27030.0 34000.0 27100.0 206415.0 ;
      RECT  27735.0 34000.0 27805.0 206415.0 ;
      RECT  28440.0 34000.0 28510.0 206415.0 ;
      RECT  29145.0 34000.0 29215.0 206415.0 ;
      RECT  29850.0 34000.0 29920.0 206415.0 ;
      RECT  30555.0 34000.0 30625.0 206415.0 ;
      RECT  31260.0 34000.0 31330.0 206415.0 ;
      RECT  31965.0 34000.0 32035.0 206415.0 ;
      RECT  32670.0 34000.0 32740.0 206415.0 ;
      RECT  33375.0 34000.0 33445.0 206415.0 ;
      RECT  34080.0 34000.0 34150.0 206415.0 ;
      RECT  34785.0 34000.0 34855.0 206415.0 ;
      RECT  35490.0 34000.0 35560.0 206415.0 ;
      RECT  36195.0 34000.0 36265.0 206415.0 ;
      RECT  36900.0 34000.0 36970.0 206415.0 ;
      RECT  37605.0 34000.0 37675.0 206415.0 ;
      RECT  38310.0 34000.0 38380.0 206415.0 ;
      RECT  39015.0 34000.0 39085.0 206415.0 ;
      RECT  39720.0 34000.0 39790.0 206415.0 ;
      RECT  40425.0 34000.0 40495.0 206415.0 ;
      RECT  41130.0 34000.0 41200.0 206415.0 ;
      RECT  41835.0 34000.0 41905.0 206415.0 ;
      RECT  42540.0 34000.0 42610.0 206415.0 ;
      RECT  43245.0 34000.0 43315.0 206415.0 ;
      RECT  43950.0 34000.0 44020.0 206415.0 ;
      RECT  44655.0 34000.0 44725.0 206415.0 ;
      RECT  45360.0 34000.0 45430.0 206415.0 ;
      RECT  46065.0 34000.0 46135.0 206415.0 ;
      RECT  46770.0 34000.0 46840.0 206415.0 ;
      RECT  47475.0 34000.0 47545.0 206415.0 ;
      RECT  48180.0 34000.0 48250.0 206415.0 ;
      RECT  48885.0 34000.0 48955.0 206415.0 ;
      RECT  49590.0 34000.0 49660.0 206415.0 ;
      RECT  50295.0 34000.0 50365.0 206415.0 ;
      RECT  51000.0 34000.0 51070.0 206415.0 ;
      RECT  51705.0 34000.0 51775.0 206415.0 ;
      RECT  52410.0 34000.0 52480.0 206415.0 ;
      RECT  53115.0 34000.0 53185.0 206415.0 ;
      RECT  53820.0 34000.0 53890.0 206415.0 ;
      RECT  54525.0 34000.0 54595.0 206415.0 ;
      RECT  55230.0 34000.0 55300.0 206415.0 ;
      RECT  55935.0 34000.0 56005.0 206415.0 ;
      RECT  56640.0 34000.0 56710.0 206415.0 ;
      RECT  57345.0 34000.0 57415.0 206415.0 ;
      RECT  58050.0 34000.0 58120.0 206415.0 ;
      RECT  58755.0 34000.0 58825.0 206415.0 ;
      RECT  59460.0 34000.0 59530.0 206415.0 ;
      RECT  60165.0 34000.0 60235.0 206415.0 ;
      RECT  60870.0 34000.0 60940.0 206415.0 ;
      RECT  61575.0 34000.0 61645.0 206415.0 ;
      RECT  62280.0 34000.0 62350.0 206415.0 ;
      RECT  62985.0 34000.0 63055.0 206415.0 ;
      RECT  63690.0 34000.0 63760.0 206415.0 ;
      RECT  64395.0 34000.0 64465.0 206415.0 ;
      RECT  65100.0 34000.0 65170.0 206415.0 ;
      RECT  65805.0 34000.0 65875.0 206415.0 ;
      RECT  66510.0 34000.0 66580.0 206415.0 ;
      RECT  67215.0 34000.0 67285.0 206415.0 ;
      RECT  67920.0 34000.0 67990.0 206415.0 ;
      RECT  68625.0 34000.0 68695.0 206415.0 ;
      RECT  69330.0 34000.0 69400.0 206415.0 ;
      RECT  70035.0 34000.0 70105.0 206415.0 ;
      RECT  70740.0 34000.0 70810.0 206415.0 ;
      RECT  71445.0 34000.0 71515.0 206415.0 ;
      RECT  72150.0 34000.0 72220.0 206415.0 ;
      RECT  72855.0 34000.0 72925.0 206415.0 ;
      RECT  73560.0 34000.0 73630.0 206415.0 ;
      RECT  74265.0 34000.0 74335.0 206415.0 ;
      RECT  74970.0 34000.0 75040.0 206415.0 ;
      RECT  75675.0 34000.0 75745.0 206415.0 ;
      RECT  76380.0 34000.0 76450.0 206415.0 ;
      RECT  77085.0 34000.0 77155.0 206415.0 ;
      RECT  77790.0 34000.0 77860.0 206415.0 ;
      RECT  78495.0 34000.0 78565.0 206415.0 ;
      RECT  79200.0 34000.0 79270.0 206415.0 ;
      RECT  79905.0 34000.0 79975.0 206415.0 ;
      RECT  80610.0 34000.0 80680.0 206415.0 ;
      RECT  81315.0 34000.0 81385.0 206415.0 ;
      RECT  82020.0 34000.0 82090.0 206415.0 ;
      RECT  82725.0 34000.0 82795.0 206415.0 ;
      RECT  83430.0 34000.0 83500.0 206415.0 ;
      RECT  84135.0 34000.0 84205.0 206415.0 ;
      RECT  84840.0 34000.0 84910.0 206415.0 ;
      RECT  85545.0 34000.0 85615.0 206415.0 ;
      RECT  86250.0 34000.0 86320.0 206415.0 ;
      RECT  86955.0 34000.0 87025.0 206415.0 ;
      RECT  87660.0 34000.0 87730.0 206415.0 ;
      RECT  88365.0 34000.0 88435.0 206415.0 ;
      RECT  89070.0 34000.0 89140.0 206415.0 ;
      RECT  89775.0 34000.0 89845.0 206415.0 ;
      RECT  90480.0 34000.0 90550.0 206415.0 ;
      RECT  91185.0 34000.0 91255.0 206415.0 ;
      RECT  91890.0 34000.0 91960.0 206415.0 ;
      RECT  92595.0 34000.0 92665.0 206415.0 ;
      RECT  93300.0 34000.0 93370.0 206415.0 ;
      RECT  94005.0 34000.0 94075.0 206415.0 ;
      RECT  94710.0 34000.0 94780.0 206415.0 ;
      RECT  95415.0 34000.0 95485.0 206415.0 ;
      RECT  96120.0 34000.0 96190.0 206415.0 ;
      RECT  96825.0 34000.0 96895.0 206415.0 ;
      RECT  97530.0 34000.0 97600.0 206415.0 ;
      RECT  98235.0 34000.0 98305.0 206415.0 ;
      RECT  98940.0 34000.0 99010.0 206415.0 ;
      RECT  99645.0 34000.0 99715.0 206415.0 ;
      RECT  100350.0 34000.0 100420.0 206415.0 ;
      RECT  101055.0 34000.0 101125.0 206415.0 ;
      RECT  101760.0 34000.0 101830.0 206415.0 ;
      RECT  102465.0 34000.0 102535.0 206415.0 ;
      RECT  103170.0 34000.0 103240.0 206415.0 ;
      RECT  103875.0 34000.0 103945.0 206415.0 ;
      RECT  104580.0 34000.0 104650.0 206415.0 ;
      RECT  105285.0 34000.0 105355.0 206415.0 ;
      RECT  105990.0 34000.0 106060.0 206415.0 ;
      RECT  106695.0 34000.0 106765.0 206415.0 ;
      RECT  107400.0 34000.0 107470.0 206415.0 ;
      RECT  17345.0 206942.5 17422.5 207077.5 ;
      RECT  17547.5 206942.5 17750.0 207077.5 ;
      RECT  17345.0 207472.5 17422.5 207607.5 ;
      RECT  17680.0 207472.5 17802.5 207607.5 ;
      RECT  17355.0 206942.5 17425.0 207077.5 ;
      RECT  17545.0 206942.5 17615.0 207077.5 ;
      RECT  17355.0 207472.5 17425.0 207607.5 ;
      RECT  17735.0 207472.5 17805.0 207607.5 ;
      RECT  17345.0 206820.0 17415.0 207987.5 ;
      RECT  17680.0 206820.0 17750.0 207987.5 ;
      RECT  18050.0 206942.5 18127.5 207077.5 ;
      RECT  18252.5 206942.5 18455.0 207077.5 ;
      RECT  18050.0 207472.5 18127.5 207607.5 ;
      RECT  18385.0 207472.5 18507.5 207607.5 ;
      RECT  18060.0 206942.5 18130.0 207077.5 ;
      RECT  18250.0 206942.5 18320.0 207077.5 ;
      RECT  18060.0 207472.5 18130.0 207607.5 ;
      RECT  18440.0 207472.5 18510.0 207607.5 ;
      RECT  18050.0 206820.0 18120.0 207987.5 ;
      RECT  18385.0 206820.0 18455.0 207987.5 ;
      RECT  18755.0 206942.5 18832.5 207077.5 ;
      RECT  18957.5 206942.5 19160.0 207077.5 ;
      RECT  18755.0 207472.5 18832.5 207607.5 ;
      RECT  19090.0 207472.5 19212.5 207607.5 ;
      RECT  18765.0 206942.5 18835.0 207077.5 ;
      RECT  18955.0 206942.5 19025.0 207077.5 ;
      RECT  18765.0 207472.5 18835.0 207607.5 ;
      RECT  19145.0 207472.5 19215.0 207607.5 ;
      RECT  18755.0 206820.0 18825.0 207987.5 ;
      RECT  19090.0 206820.0 19160.0 207987.5 ;
      RECT  19460.0 206942.5 19537.5 207077.5 ;
      RECT  19662.5 206942.5 19865.0 207077.5 ;
      RECT  19460.0 207472.5 19537.5 207607.5 ;
      RECT  19795.0 207472.5 19917.5 207607.5 ;
      RECT  19470.0 206942.5 19540.0 207077.5 ;
      RECT  19660.0 206942.5 19730.0 207077.5 ;
      RECT  19470.0 207472.5 19540.0 207607.5 ;
      RECT  19850.0 207472.5 19920.0 207607.5 ;
      RECT  19460.0 206820.0 19530.0 207987.5 ;
      RECT  19795.0 206820.0 19865.0 207987.5 ;
      RECT  20165.0 206942.5 20242.5 207077.5 ;
      RECT  20367.5 206942.5 20570.0 207077.5 ;
      RECT  20165.0 207472.5 20242.5 207607.5 ;
      RECT  20500.0 207472.5 20622.5 207607.5 ;
      RECT  20175.0 206942.5 20245.0 207077.5 ;
      RECT  20365.0 206942.5 20435.0 207077.5 ;
      RECT  20175.0 207472.5 20245.0 207607.5 ;
      RECT  20555.0 207472.5 20625.0 207607.5 ;
      RECT  20165.0 206820.0 20235.0 207987.5 ;
      RECT  20500.0 206820.0 20570.0 207987.5 ;
      RECT  20870.0 206942.5 20947.5 207077.5 ;
      RECT  21072.5 206942.5 21275.0 207077.5 ;
      RECT  20870.0 207472.5 20947.5 207607.5 ;
      RECT  21205.0 207472.5 21327.5 207607.5 ;
      RECT  20880.0 206942.5 20950.0 207077.5 ;
      RECT  21070.0 206942.5 21140.0 207077.5 ;
      RECT  20880.0 207472.5 20950.0 207607.5 ;
      RECT  21260.0 207472.5 21330.0 207607.5 ;
      RECT  20870.0 206820.0 20940.0 207987.5 ;
      RECT  21205.0 206820.0 21275.0 207987.5 ;
      RECT  21575.0 206942.5 21652.5 207077.5 ;
      RECT  21777.5 206942.5 21980.0 207077.5 ;
      RECT  21575.0 207472.5 21652.5 207607.5 ;
      RECT  21910.0 207472.5 22032.5 207607.5 ;
      RECT  21585.0 206942.5 21655.0 207077.5 ;
      RECT  21775.0 206942.5 21845.0 207077.5 ;
      RECT  21585.0 207472.5 21655.0 207607.5 ;
      RECT  21965.0 207472.5 22035.0 207607.5 ;
      RECT  21575.0 206820.0 21645.0 207987.5 ;
      RECT  21910.0 206820.0 21980.0 207987.5 ;
      RECT  22280.0 206942.5 22357.5 207077.5 ;
      RECT  22482.5 206942.5 22685.0 207077.5 ;
      RECT  22280.0 207472.5 22357.5 207607.5 ;
      RECT  22615.0 207472.5 22737.5 207607.5 ;
      RECT  22290.0 206942.5 22360.0 207077.5 ;
      RECT  22480.0 206942.5 22550.0 207077.5 ;
      RECT  22290.0 207472.5 22360.0 207607.5 ;
      RECT  22670.0 207472.5 22740.0 207607.5 ;
      RECT  22280.0 206820.0 22350.0 207987.5 ;
      RECT  22615.0 206820.0 22685.0 207987.5 ;
      RECT  22985.0 206942.5 23062.5 207077.5 ;
      RECT  23187.5 206942.5 23390.0 207077.5 ;
      RECT  22985.0 207472.5 23062.5 207607.5 ;
      RECT  23320.0 207472.5 23442.5 207607.5 ;
      RECT  22995.0 206942.5 23065.0 207077.5 ;
      RECT  23185.0 206942.5 23255.0 207077.5 ;
      RECT  22995.0 207472.5 23065.0 207607.5 ;
      RECT  23375.0 207472.5 23445.0 207607.5 ;
      RECT  22985.0 206820.0 23055.0 207987.5 ;
      RECT  23320.0 206820.0 23390.0 207987.5 ;
      RECT  23690.0 206942.5 23767.5 207077.5 ;
      RECT  23892.5 206942.5 24095.0 207077.5 ;
      RECT  23690.0 207472.5 23767.5 207607.5 ;
      RECT  24025.0 207472.5 24147.5 207607.5 ;
      RECT  23700.0 206942.5 23770.0 207077.5 ;
      RECT  23890.0 206942.5 23960.0 207077.5 ;
      RECT  23700.0 207472.5 23770.0 207607.5 ;
      RECT  24080.0 207472.5 24150.0 207607.5 ;
      RECT  23690.0 206820.0 23760.0 207987.5 ;
      RECT  24025.0 206820.0 24095.0 207987.5 ;
      RECT  24395.0 206942.5 24472.5 207077.5 ;
      RECT  24597.5 206942.5 24800.0 207077.5 ;
      RECT  24395.0 207472.5 24472.5 207607.5 ;
      RECT  24730.0 207472.5 24852.5 207607.5 ;
      RECT  24405.0 206942.5 24475.0 207077.5 ;
      RECT  24595.0 206942.5 24665.0 207077.5 ;
      RECT  24405.0 207472.5 24475.0 207607.5 ;
      RECT  24785.0 207472.5 24855.0 207607.5 ;
      RECT  24395.0 206820.0 24465.0 207987.5 ;
      RECT  24730.0 206820.0 24800.0 207987.5 ;
      RECT  25100.0 206942.5 25177.5 207077.5 ;
      RECT  25302.5 206942.5 25505.0 207077.5 ;
      RECT  25100.0 207472.5 25177.5 207607.5 ;
      RECT  25435.0 207472.5 25557.5 207607.5 ;
      RECT  25110.0 206942.5 25180.0 207077.5 ;
      RECT  25300.0 206942.5 25370.0 207077.5 ;
      RECT  25110.0 207472.5 25180.0 207607.5 ;
      RECT  25490.0 207472.5 25560.0 207607.5 ;
      RECT  25100.0 206820.0 25170.0 207987.5 ;
      RECT  25435.0 206820.0 25505.0 207987.5 ;
      RECT  25805.0 206942.5 25882.5 207077.5 ;
      RECT  26007.5 206942.5 26210.0 207077.5 ;
      RECT  25805.0 207472.5 25882.5 207607.5 ;
      RECT  26140.0 207472.5 26262.5 207607.5 ;
      RECT  25815.0 206942.5 25885.0 207077.5 ;
      RECT  26005.0 206942.5 26075.0 207077.5 ;
      RECT  25815.0 207472.5 25885.0 207607.5 ;
      RECT  26195.0 207472.5 26265.0 207607.5 ;
      RECT  25805.0 206820.0 25875.0 207987.5 ;
      RECT  26140.0 206820.0 26210.0 207987.5 ;
      RECT  26510.0 206942.5 26587.5 207077.5 ;
      RECT  26712.5 206942.5 26915.0 207077.5 ;
      RECT  26510.0 207472.5 26587.5 207607.5 ;
      RECT  26845.0 207472.5 26967.5 207607.5 ;
      RECT  26520.0 206942.5 26590.0 207077.5 ;
      RECT  26710.0 206942.5 26780.0 207077.5 ;
      RECT  26520.0 207472.5 26590.0 207607.5 ;
      RECT  26900.0 207472.5 26970.0 207607.5 ;
      RECT  26510.0 206820.0 26580.0 207987.5 ;
      RECT  26845.0 206820.0 26915.0 207987.5 ;
      RECT  27215.0 206942.5 27292.5 207077.5 ;
      RECT  27417.5 206942.5 27620.0 207077.5 ;
      RECT  27215.0 207472.5 27292.5 207607.5 ;
      RECT  27550.0 207472.5 27672.5 207607.5 ;
      RECT  27225.0 206942.5 27295.0 207077.5 ;
      RECT  27415.0 206942.5 27485.0 207077.5 ;
      RECT  27225.0 207472.5 27295.0 207607.5 ;
      RECT  27605.0 207472.5 27675.0 207607.5 ;
      RECT  27215.0 206820.0 27285.0 207987.5 ;
      RECT  27550.0 206820.0 27620.0 207987.5 ;
      RECT  27920.0 206942.5 27997.5 207077.5 ;
      RECT  28122.5 206942.5 28325.0 207077.5 ;
      RECT  27920.0 207472.5 27997.5 207607.5 ;
      RECT  28255.0 207472.5 28377.5 207607.5 ;
      RECT  27930.0 206942.5 28000.0 207077.5 ;
      RECT  28120.0 206942.5 28190.0 207077.5 ;
      RECT  27930.0 207472.5 28000.0 207607.5 ;
      RECT  28310.0 207472.5 28380.0 207607.5 ;
      RECT  27920.0 206820.0 27990.0 207987.5 ;
      RECT  28255.0 206820.0 28325.0 207987.5 ;
      RECT  28625.0 206942.5 28702.5 207077.5 ;
      RECT  28827.5 206942.5 29030.0 207077.5 ;
      RECT  28625.0 207472.5 28702.5 207607.5 ;
      RECT  28960.0 207472.5 29082.5 207607.5 ;
      RECT  28635.0 206942.5 28705.0 207077.5 ;
      RECT  28825.0 206942.5 28895.0 207077.5 ;
      RECT  28635.0 207472.5 28705.0 207607.5 ;
      RECT  29015.0 207472.5 29085.0 207607.5 ;
      RECT  28625.0 206820.0 28695.0 207987.5 ;
      RECT  28960.0 206820.0 29030.0 207987.5 ;
      RECT  29330.0 206942.5 29407.5 207077.5 ;
      RECT  29532.5 206942.5 29735.0 207077.5 ;
      RECT  29330.0 207472.5 29407.5 207607.5 ;
      RECT  29665.0 207472.5 29787.5 207607.5 ;
      RECT  29340.0 206942.5 29410.0 207077.5 ;
      RECT  29530.0 206942.5 29600.0 207077.5 ;
      RECT  29340.0 207472.5 29410.0 207607.5 ;
      RECT  29720.0 207472.5 29790.0 207607.5 ;
      RECT  29330.0 206820.0 29400.0 207987.5 ;
      RECT  29665.0 206820.0 29735.0 207987.5 ;
      RECT  30035.0 206942.5 30112.5 207077.5 ;
      RECT  30237.5 206942.5 30440.0 207077.5 ;
      RECT  30035.0 207472.5 30112.5 207607.5 ;
      RECT  30370.0 207472.5 30492.5 207607.5 ;
      RECT  30045.0 206942.5 30115.0 207077.5 ;
      RECT  30235.0 206942.5 30305.0 207077.5 ;
      RECT  30045.0 207472.5 30115.0 207607.5 ;
      RECT  30425.0 207472.5 30495.0 207607.5 ;
      RECT  30035.0 206820.0 30105.0 207987.5 ;
      RECT  30370.0 206820.0 30440.0 207987.5 ;
      RECT  30740.0 206942.5 30817.5 207077.5 ;
      RECT  30942.5 206942.5 31145.0 207077.5 ;
      RECT  30740.0 207472.5 30817.5 207607.5 ;
      RECT  31075.0 207472.5 31197.5 207607.5 ;
      RECT  30750.0 206942.5 30820.0 207077.5 ;
      RECT  30940.0 206942.5 31010.0 207077.5 ;
      RECT  30750.0 207472.5 30820.0 207607.5 ;
      RECT  31130.0 207472.5 31200.0 207607.5 ;
      RECT  30740.0 206820.0 30810.0 207987.5 ;
      RECT  31075.0 206820.0 31145.0 207987.5 ;
      RECT  31445.0 206942.5 31522.5 207077.5 ;
      RECT  31647.5 206942.5 31850.0 207077.5 ;
      RECT  31445.0 207472.5 31522.5 207607.5 ;
      RECT  31780.0 207472.5 31902.5 207607.5 ;
      RECT  31455.0 206942.5 31525.0 207077.5 ;
      RECT  31645.0 206942.5 31715.0 207077.5 ;
      RECT  31455.0 207472.5 31525.0 207607.5 ;
      RECT  31835.0 207472.5 31905.0 207607.5 ;
      RECT  31445.0 206820.0 31515.0 207987.5 ;
      RECT  31780.0 206820.0 31850.0 207987.5 ;
      RECT  32150.0 206942.5 32227.5 207077.5 ;
      RECT  32352.5 206942.5 32555.0 207077.5 ;
      RECT  32150.0 207472.5 32227.5 207607.5 ;
      RECT  32485.0 207472.5 32607.5 207607.5 ;
      RECT  32160.0 206942.5 32230.0 207077.5 ;
      RECT  32350.0 206942.5 32420.0 207077.5 ;
      RECT  32160.0 207472.5 32230.0 207607.5 ;
      RECT  32540.0 207472.5 32610.0 207607.5 ;
      RECT  32150.0 206820.0 32220.0 207987.5 ;
      RECT  32485.0 206820.0 32555.0 207987.5 ;
      RECT  32855.0 206942.5 32932.5 207077.5 ;
      RECT  33057.5 206942.5 33260.0 207077.5 ;
      RECT  32855.0 207472.5 32932.5 207607.5 ;
      RECT  33190.0 207472.5 33312.5 207607.5 ;
      RECT  32865.0 206942.5 32935.0 207077.5 ;
      RECT  33055.0 206942.5 33125.0 207077.5 ;
      RECT  32865.0 207472.5 32935.0 207607.5 ;
      RECT  33245.0 207472.5 33315.0 207607.5 ;
      RECT  32855.0 206820.0 32925.0 207987.5 ;
      RECT  33190.0 206820.0 33260.0 207987.5 ;
      RECT  33560.0 206942.5 33637.5 207077.5 ;
      RECT  33762.5 206942.5 33965.0 207077.5 ;
      RECT  33560.0 207472.5 33637.5 207607.5 ;
      RECT  33895.0 207472.5 34017.5 207607.5 ;
      RECT  33570.0 206942.5 33640.0 207077.5 ;
      RECT  33760.0 206942.5 33830.0 207077.5 ;
      RECT  33570.0 207472.5 33640.0 207607.5 ;
      RECT  33950.0 207472.5 34020.0 207607.5 ;
      RECT  33560.0 206820.0 33630.0 207987.5 ;
      RECT  33895.0 206820.0 33965.0 207987.5 ;
      RECT  34265.0 206942.5 34342.5 207077.5 ;
      RECT  34467.5 206942.5 34670.0 207077.5 ;
      RECT  34265.0 207472.5 34342.5 207607.5 ;
      RECT  34600.0 207472.5 34722.5 207607.5 ;
      RECT  34275.0 206942.5 34345.0 207077.5 ;
      RECT  34465.0 206942.5 34535.0 207077.5 ;
      RECT  34275.0 207472.5 34345.0 207607.5 ;
      RECT  34655.0 207472.5 34725.0 207607.5 ;
      RECT  34265.0 206820.0 34335.0 207987.5 ;
      RECT  34600.0 206820.0 34670.0 207987.5 ;
      RECT  34970.0 206942.5 35047.5 207077.5 ;
      RECT  35172.5 206942.5 35375.0 207077.5 ;
      RECT  34970.0 207472.5 35047.5 207607.5 ;
      RECT  35305.0 207472.5 35427.5 207607.5 ;
      RECT  34980.0 206942.5 35050.0 207077.5 ;
      RECT  35170.0 206942.5 35240.0 207077.5 ;
      RECT  34980.0 207472.5 35050.0 207607.5 ;
      RECT  35360.0 207472.5 35430.0 207607.5 ;
      RECT  34970.0 206820.0 35040.0 207987.5 ;
      RECT  35305.0 206820.0 35375.0 207987.5 ;
      RECT  35675.0 206942.5 35752.5 207077.5 ;
      RECT  35877.5 206942.5 36080.0 207077.5 ;
      RECT  35675.0 207472.5 35752.5 207607.5 ;
      RECT  36010.0 207472.5 36132.5 207607.5 ;
      RECT  35685.0 206942.5 35755.0 207077.5 ;
      RECT  35875.0 206942.5 35945.0 207077.5 ;
      RECT  35685.0 207472.5 35755.0 207607.5 ;
      RECT  36065.0 207472.5 36135.0 207607.5 ;
      RECT  35675.0 206820.0 35745.0 207987.5 ;
      RECT  36010.0 206820.0 36080.0 207987.5 ;
      RECT  36380.0 206942.5 36457.5 207077.5 ;
      RECT  36582.5 206942.5 36785.0 207077.5 ;
      RECT  36380.0 207472.5 36457.5 207607.5 ;
      RECT  36715.0 207472.5 36837.5 207607.5 ;
      RECT  36390.0 206942.5 36460.0 207077.5 ;
      RECT  36580.0 206942.5 36650.0 207077.5 ;
      RECT  36390.0 207472.5 36460.0 207607.5 ;
      RECT  36770.0 207472.5 36840.0 207607.5 ;
      RECT  36380.0 206820.0 36450.0 207987.5 ;
      RECT  36715.0 206820.0 36785.0 207987.5 ;
      RECT  37085.0 206942.5 37162.5 207077.5 ;
      RECT  37287.5 206942.5 37490.0 207077.5 ;
      RECT  37085.0 207472.5 37162.5 207607.5 ;
      RECT  37420.0 207472.5 37542.5 207607.5 ;
      RECT  37095.0 206942.5 37165.0 207077.5 ;
      RECT  37285.0 206942.5 37355.0 207077.5 ;
      RECT  37095.0 207472.5 37165.0 207607.5 ;
      RECT  37475.0 207472.5 37545.0 207607.5 ;
      RECT  37085.0 206820.0 37155.0 207987.5 ;
      RECT  37420.0 206820.0 37490.0 207987.5 ;
      RECT  37790.0 206942.5 37867.5 207077.5 ;
      RECT  37992.5 206942.5 38195.0 207077.5 ;
      RECT  37790.0 207472.5 37867.5 207607.5 ;
      RECT  38125.0 207472.5 38247.5 207607.5 ;
      RECT  37800.0 206942.5 37870.0 207077.5 ;
      RECT  37990.0 206942.5 38060.0 207077.5 ;
      RECT  37800.0 207472.5 37870.0 207607.5 ;
      RECT  38180.0 207472.5 38250.0 207607.5 ;
      RECT  37790.0 206820.0 37860.0 207987.5 ;
      RECT  38125.0 206820.0 38195.0 207987.5 ;
      RECT  38495.0 206942.5 38572.5 207077.5 ;
      RECT  38697.5 206942.5 38900.0 207077.5 ;
      RECT  38495.0 207472.5 38572.5 207607.5 ;
      RECT  38830.0 207472.5 38952.5 207607.5 ;
      RECT  38505.0 206942.5 38575.0 207077.5 ;
      RECT  38695.0 206942.5 38765.0 207077.5 ;
      RECT  38505.0 207472.5 38575.0 207607.5 ;
      RECT  38885.0 207472.5 38955.0 207607.5 ;
      RECT  38495.0 206820.0 38565.0 207987.5 ;
      RECT  38830.0 206820.0 38900.0 207987.5 ;
      RECT  39200.0 206942.5 39277.5 207077.5 ;
      RECT  39402.5 206942.5 39605.0 207077.5 ;
      RECT  39200.0 207472.5 39277.5 207607.5 ;
      RECT  39535.0 207472.5 39657.5 207607.5 ;
      RECT  39210.0 206942.5 39280.0 207077.5 ;
      RECT  39400.0 206942.5 39470.0 207077.5 ;
      RECT  39210.0 207472.5 39280.0 207607.5 ;
      RECT  39590.0 207472.5 39660.0 207607.5 ;
      RECT  39200.0 206820.0 39270.0 207987.5 ;
      RECT  39535.0 206820.0 39605.0 207987.5 ;
      RECT  39905.0 206942.5 39982.5 207077.5 ;
      RECT  40107.5 206942.5 40310.0 207077.5 ;
      RECT  39905.0 207472.5 39982.5 207607.5 ;
      RECT  40240.0 207472.5 40362.5 207607.5 ;
      RECT  39915.0 206942.5 39985.0 207077.5 ;
      RECT  40105.0 206942.5 40175.0 207077.5 ;
      RECT  39915.0 207472.5 39985.0 207607.5 ;
      RECT  40295.0 207472.5 40365.0 207607.5 ;
      RECT  39905.0 206820.0 39975.0 207987.5 ;
      RECT  40240.0 206820.0 40310.0 207987.5 ;
      RECT  40610.0 206942.5 40687.5 207077.5 ;
      RECT  40812.5 206942.5 41015.0 207077.5 ;
      RECT  40610.0 207472.5 40687.5 207607.5 ;
      RECT  40945.0 207472.5 41067.5 207607.5 ;
      RECT  40620.0 206942.5 40690.0 207077.5 ;
      RECT  40810.0 206942.5 40880.0 207077.5 ;
      RECT  40620.0 207472.5 40690.0 207607.5 ;
      RECT  41000.0 207472.5 41070.0 207607.5 ;
      RECT  40610.0 206820.0 40680.0 207987.5 ;
      RECT  40945.0 206820.0 41015.0 207987.5 ;
      RECT  41315.0 206942.5 41392.5 207077.5 ;
      RECT  41517.5 206942.5 41720.0 207077.5 ;
      RECT  41315.0 207472.5 41392.5 207607.5 ;
      RECT  41650.0 207472.5 41772.5 207607.5 ;
      RECT  41325.0 206942.5 41395.0 207077.5 ;
      RECT  41515.0 206942.5 41585.0 207077.5 ;
      RECT  41325.0 207472.5 41395.0 207607.5 ;
      RECT  41705.0 207472.5 41775.0 207607.5 ;
      RECT  41315.0 206820.0 41385.0 207987.5 ;
      RECT  41650.0 206820.0 41720.0 207987.5 ;
      RECT  42020.0 206942.5 42097.5 207077.5 ;
      RECT  42222.5 206942.5 42425.0 207077.5 ;
      RECT  42020.0 207472.5 42097.5 207607.5 ;
      RECT  42355.0 207472.5 42477.5 207607.5 ;
      RECT  42030.0 206942.5 42100.0 207077.5 ;
      RECT  42220.0 206942.5 42290.0 207077.5 ;
      RECT  42030.0 207472.5 42100.0 207607.5 ;
      RECT  42410.0 207472.5 42480.0 207607.5 ;
      RECT  42020.0 206820.0 42090.0 207987.5 ;
      RECT  42355.0 206820.0 42425.0 207987.5 ;
      RECT  42725.0 206942.5 42802.5 207077.5 ;
      RECT  42927.5 206942.5 43130.0 207077.5 ;
      RECT  42725.0 207472.5 42802.5 207607.5 ;
      RECT  43060.0 207472.5 43182.5 207607.5 ;
      RECT  42735.0 206942.5 42805.0 207077.5 ;
      RECT  42925.0 206942.5 42995.0 207077.5 ;
      RECT  42735.0 207472.5 42805.0 207607.5 ;
      RECT  43115.0 207472.5 43185.0 207607.5 ;
      RECT  42725.0 206820.0 42795.0 207987.5 ;
      RECT  43060.0 206820.0 43130.0 207987.5 ;
      RECT  43430.0 206942.5 43507.5 207077.5 ;
      RECT  43632.5 206942.5 43835.0 207077.5 ;
      RECT  43430.0 207472.5 43507.5 207607.5 ;
      RECT  43765.0 207472.5 43887.5 207607.5 ;
      RECT  43440.0 206942.5 43510.0 207077.5 ;
      RECT  43630.0 206942.5 43700.0 207077.5 ;
      RECT  43440.0 207472.5 43510.0 207607.5 ;
      RECT  43820.0 207472.5 43890.0 207607.5 ;
      RECT  43430.0 206820.0 43500.0 207987.5 ;
      RECT  43765.0 206820.0 43835.0 207987.5 ;
      RECT  44135.0 206942.5 44212.5 207077.5 ;
      RECT  44337.5 206942.5 44540.0 207077.5 ;
      RECT  44135.0 207472.5 44212.5 207607.5 ;
      RECT  44470.0 207472.5 44592.5 207607.5 ;
      RECT  44145.0 206942.5 44215.0 207077.5 ;
      RECT  44335.0 206942.5 44405.0 207077.5 ;
      RECT  44145.0 207472.5 44215.0 207607.5 ;
      RECT  44525.0 207472.5 44595.0 207607.5 ;
      RECT  44135.0 206820.0 44205.0 207987.5 ;
      RECT  44470.0 206820.0 44540.0 207987.5 ;
      RECT  44840.0 206942.5 44917.5 207077.5 ;
      RECT  45042.5 206942.5 45245.0 207077.5 ;
      RECT  44840.0 207472.5 44917.5 207607.5 ;
      RECT  45175.0 207472.5 45297.5 207607.5 ;
      RECT  44850.0 206942.5 44920.0 207077.5 ;
      RECT  45040.0 206942.5 45110.0 207077.5 ;
      RECT  44850.0 207472.5 44920.0 207607.5 ;
      RECT  45230.0 207472.5 45300.0 207607.5 ;
      RECT  44840.0 206820.0 44910.0 207987.5 ;
      RECT  45175.0 206820.0 45245.0 207987.5 ;
      RECT  45545.0 206942.5 45622.5 207077.5 ;
      RECT  45747.5 206942.5 45950.0 207077.5 ;
      RECT  45545.0 207472.5 45622.5 207607.5 ;
      RECT  45880.0 207472.5 46002.5 207607.5 ;
      RECT  45555.0 206942.5 45625.0 207077.5 ;
      RECT  45745.0 206942.5 45815.0 207077.5 ;
      RECT  45555.0 207472.5 45625.0 207607.5 ;
      RECT  45935.0 207472.5 46005.0 207607.5 ;
      RECT  45545.0 206820.0 45615.0 207987.5 ;
      RECT  45880.0 206820.0 45950.0 207987.5 ;
      RECT  46250.0 206942.5 46327.5 207077.5 ;
      RECT  46452.5 206942.5 46655.0 207077.5 ;
      RECT  46250.0 207472.5 46327.5 207607.5 ;
      RECT  46585.0 207472.5 46707.5 207607.5 ;
      RECT  46260.0 206942.5 46330.0 207077.5 ;
      RECT  46450.0 206942.5 46520.0 207077.5 ;
      RECT  46260.0 207472.5 46330.0 207607.5 ;
      RECT  46640.0 207472.5 46710.0 207607.5 ;
      RECT  46250.0 206820.0 46320.0 207987.5 ;
      RECT  46585.0 206820.0 46655.0 207987.5 ;
      RECT  46955.0 206942.5 47032.5 207077.5 ;
      RECT  47157.5 206942.5 47360.0 207077.5 ;
      RECT  46955.0 207472.5 47032.5 207607.5 ;
      RECT  47290.0 207472.5 47412.5 207607.5 ;
      RECT  46965.0 206942.5 47035.0 207077.5 ;
      RECT  47155.0 206942.5 47225.0 207077.5 ;
      RECT  46965.0 207472.5 47035.0 207607.5 ;
      RECT  47345.0 207472.5 47415.0 207607.5 ;
      RECT  46955.0 206820.0 47025.0 207987.5 ;
      RECT  47290.0 206820.0 47360.0 207987.5 ;
      RECT  47660.0 206942.5 47737.5 207077.5 ;
      RECT  47862.5 206942.5 48065.0 207077.5 ;
      RECT  47660.0 207472.5 47737.5 207607.5 ;
      RECT  47995.0 207472.5 48117.5 207607.5 ;
      RECT  47670.0 206942.5 47740.0 207077.5 ;
      RECT  47860.0 206942.5 47930.0 207077.5 ;
      RECT  47670.0 207472.5 47740.0 207607.5 ;
      RECT  48050.0 207472.5 48120.0 207607.5 ;
      RECT  47660.0 206820.0 47730.0 207987.5 ;
      RECT  47995.0 206820.0 48065.0 207987.5 ;
      RECT  48365.0 206942.5 48442.5 207077.5 ;
      RECT  48567.5 206942.5 48770.0 207077.5 ;
      RECT  48365.0 207472.5 48442.5 207607.5 ;
      RECT  48700.0 207472.5 48822.5 207607.5 ;
      RECT  48375.0 206942.5 48445.0 207077.5 ;
      RECT  48565.0 206942.5 48635.0 207077.5 ;
      RECT  48375.0 207472.5 48445.0 207607.5 ;
      RECT  48755.0 207472.5 48825.0 207607.5 ;
      RECT  48365.0 206820.0 48435.0 207987.5 ;
      RECT  48700.0 206820.0 48770.0 207987.5 ;
      RECT  49070.0 206942.5 49147.5 207077.5 ;
      RECT  49272.5 206942.5 49475.0 207077.5 ;
      RECT  49070.0 207472.5 49147.5 207607.5 ;
      RECT  49405.0 207472.5 49527.5 207607.5 ;
      RECT  49080.0 206942.5 49150.0 207077.5 ;
      RECT  49270.0 206942.5 49340.0 207077.5 ;
      RECT  49080.0 207472.5 49150.0 207607.5 ;
      RECT  49460.0 207472.5 49530.0 207607.5 ;
      RECT  49070.0 206820.0 49140.0 207987.5 ;
      RECT  49405.0 206820.0 49475.0 207987.5 ;
      RECT  49775.0 206942.5 49852.5 207077.5 ;
      RECT  49977.5 206942.5 50180.0 207077.5 ;
      RECT  49775.0 207472.5 49852.5 207607.5 ;
      RECT  50110.0 207472.5 50232.5 207607.5 ;
      RECT  49785.0 206942.5 49855.0 207077.5 ;
      RECT  49975.0 206942.5 50045.0 207077.5 ;
      RECT  49785.0 207472.5 49855.0 207607.5 ;
      RECT  50165.0 207472.5 50235.0 207607.5 ;
      RECT  49775.0 206820.0 49845.0 207987.5 ;
      RECT  50110.0 206820.0 50180.0 207987.5 ;
      RECT  50480.0 206942.5 50557.5 207077.5 ;
      RECT  50682.5 206942.5 50885.0 207077.5 ;
      RECT  50480.0 207472.5 50557.5 207607.5 ;
      RECT  50815.0 207472.5 50937.5 207607.5 ;
      RECT  50490.0 206942.5 50560.0 207077.5 ;
      RECT  50680.0 206942.5 50750.0 207077.5 ;
      RECT  50490.0 207472.5 50560.0 207607.5 ;
      RECT  50870.0 207472.5 50940.0 207607.5 ;
      RECT  50480.0 206820.0 50550.0 207987.5 ;
      RECT  50815.0 206820.0 50885.0 207987.5 ;
      RECT  51185.0 206942.5 51262.5 207077.5 ;
      RECT  51387.5 206942.5 51590.0 207077.5 ;
      RECT  51185.0 207472.5 51262.5 207607.5 ;
      RECT  51520.0 207472.5 51642.5 207607.5 ;
      RECT  51195.0 206942.5 51265.0 207077.5 ;
      RECT  51385.0 206942.5 51455.0 207077.5 ;
      RECT  51195.0 207472.5 51265.0 207607.5 ;
      RECT  51575.0 207472.5 51645.0 207607.5 ;
      RECT  51185.0 206820.0 51255.0 207987.5 ;
      RECT  51520.0 206820.0 51590.0 207987.5 ;
      RECT  51890.0 206942.5 51967.5 207077.5 ;
      RECT  52092.5 206942.5 52295.0 207077.5 ;
      RECT  51890.0 207472.5 51967.5 207607.5 ;
      RECT  52225.0 207472.5 52347.5 207607.5 ;
      RECT  51900.0 206942.5 51970.0 207077.5 ;
      RECT  52090.0 206942.5 52160.0 207077.5 ;
      RECT  51900.0 207472.5 51970.0 207607.5 ;
      RECT  52280.0 207472.5 52350.0 207607.5 ;
      RECT  51890.0 206820.0 51960.0 207987.5 ;
      RECT  52225.0 206820.0 52295.0 207987.5 ;
      RECT  52595.0 206942.5 52672.5 207077.5 ;
      RECT  52797.5 206942.5 53000.0 207077.5 ;
      RECT  52595.0 207472.5 52672.5 207607.5 ;
      RECT  52930.0 207472.5 53052.5 207607.5 ;
      RECT  52605.0 206942.5 52675.0 207077.5 ;
      RECT  52795.0 206942.5 52865.0 207077.5 ;
      RECT  52605.0 207472.5 52675.0 207607.5 ;
      RECT  52985.0 207472.5 53055.0 207607.5 ;
      RECT  52595.0 206820.0 52665.0 207987.5 ;
      RECT  52930.0 206820.0 53000.0 207987.5 ;
      RECT  53300.0 206942.5 53377.5 207077.5 ;
      RECT  53502.5 206942.5 53705.0 207077.5 ;
      RECT  53300.0 207472.5 53377.5 207607.5 ;
      RECT  53635.0 207472.5 53757.5 207607.5 ;
      RECT  53310.0 206942.5 53380.0 207077.5 ;
      RECT  53500.0 206942.5 53570.0 207077.5 ;
      RECT  53310.0 207472.5 53380.0 207607.5 ;
      RECT  53690.0 207472.5 53760.0 207607.5 ;
      RECT  53300.0 206820.0 53370.0 207987.5 ;
      RECT  53635.0 206820.0 53705.0 207987.5 ;
      RECT  54005.0 206942.5 54082.5 207077.5 ;
      RECT  54207.5 206942.5 54410.0 207077.5 ;
      RECT  54005.0 207472.5 54082.5 207607.5 ;
      RECT  54340.0 207472.5 54462.5 207607.5 ;
      RECT  54015.0 206942.5 54085.0 207077.5 ;
      RECT  54205.0 206942.5 54275.0 207077.5 ;
      RECT  54015.0 207472.5 54085.0 207607.5 ;
      RECT  54395.0 207472.5 54465.0 207607.5 ;
      RECT  54005.0 206820.0 54075.0 207987.5 ;
      RECT  54340.0 206820.0 54410.0 207987.5 ;
      RECT  54710.0 206942.5 54787.5 207077.5 ;
      RECT  54912.5 206942.5 55115.0 207077.5 ;
      RECT  54710.0 207472.5 54787.5 207607.5 ;
      RECT  55045.0 207472.5 55167.5 207607.5 ;
      RECT  54720.0 206942.5 54790.0 207077.5 ;
      RECT  54910.0 206942.5 54980.0 207077.5 ;
      RECT  54720.0 207472.5 54790.0 207607.5 ;
      RECT  55100.0 207472.5 55170.0 207607.5 ;
      RECT  54710.0 206820.0 54780.0 207987.5 ;
      RECT  55045.0 206820.0 55115.0 207987.5 ;
      RECT  55415.0 206942.5 55492.5 207077.5 ;
      RECT  55617.5 206942.5 55820.0 207077.5 ;
      RECT  55415.0 207472.5 55492.5 207607.5 ;
      RECT  55750.0 207472.5 55872.5 207607.5 ;
      RECT  55425.0 206942.5 55495.0 207077.5 ;
      RECT  55615.0 206942.5 55685.0 207077.5 ;
      RECT  55425.0 207472.5 55495.0 207607.5 ;
      RECT  55805.0 207472.5 55875.0 207607.5 ;
      RECT  55415.0 206820.0 55485.0 207987.5 ;
      RECT  55750.0 206820.0 55820.0 207987.5 ;
      RECT  56120.0 206942.5 56197.5 207077.5 ;
      RECT  56322.5 206942.5 56525.0 207077.5 ;
      RECT  56120.0 207472.5 56197.5 207607.5 ;
      RECT  56455.0 207472.5 56577.5 207607.5 ;
      RECT  56130.0 206942.5 56200.0 207077.5 ;
      RECT  56320.0 206942.5 56390.0 207077.5 ;
      RECT  56130.0 207472.5 56200.0 207607.5 ;
      RECT  56510.0 207472.5 56580.0 207607.5 ;
      RECT  56120.0 206820.0 56190.0 207987.5 ;
      RECT  56455.0 206820.0 56525.0 207987.5 ;
      RECT  56825.0 206942.5 56902.5 207077.5 ;
      RECT  57027.5 206942.5 57230.0 207077.5 ;
      RECT  56825.0 207472.5 56902.5 207607.5 ;
      RECT  57160.0 207472.5 57282.5 207607.5 ;
      RECT  56835.0 206942.5 56905.0 207077.5 ;
      RECT  57025.0 206942.5 57095.0 207077.5 ;
      RECT  56835.0 207472.5 56905.0 207607.5 ;
      RECT  57215.0 207472.5 57285.0 207607.5 ;
      RECT  56825.0 206820.0 56895.0 207987.5 ;
      RECT  57160.0 206820.0 57230.0 207987.5 ;
      RECT  57530.0 206942.5 57607.5 207077.5 ;
      RECT  57732.5 206942.5 57935.0 207077.5 ;
      RECT  57530.0 207472.5 57607.5 207607.5 ;
      RECT  57865.0 207472.5 57987.5 207607.5 ;
      RECT  57540.0 206942.5 57610.0 207077.5 ;
      RECT  57730.0 206942.5 57800.0 207077.5 ;
      RECT  57540.0 207472.5 57610.0 207607.5 ;
      RECT  57920.0 207472.5 57990.0 207607.5 ;
      RECT  57530.0 206820.0 57600.0 207987.5 ;
      RECT  57865.0 206820.0 57935.0 207987.5 ;
      RECT  58235.0 206942.5 58312.5 207077.5 ;
      RECT  58437.5 206942.5 58640.0 207077.5 ;
      RECT  58235.0 207472.5 58312.5 207607.5 ;
      RECT  58570.0 207472.5 58692.5 207607.5 ;
      RECT  58245.0 206942.5 58315.0 207077.5 ;
      RECT  58435.0 206942.5 58505.0 207077.5 ;
      RECT  58245.0 207472.5 58315.0 207607.5 ;
      RECT  58625.0 207472.5 58695.0 207607.5 ;
      RECT  58235.0 206820.0 58305.0 207987.5 ;
      RECT  58570.0 206820.0 58640.0 207987.5 ;
      RECT  58940.0 206942.5 59017.5 207077.5 ;
      RECT  59142.5 206942.5 59345.0 207077.5 ;
      RECT  58940.0 207472.5 59017.5 207607.5 ;
      RECT  59275.0 207472.5 59397.5 207607.5 ;
      RECT  58950.0 206942.5 59020.0 207077.5 ;
      RECT  59140.0 206942.5 59210.0 207077.5 ;
      RECT  58950.0 207472.5 59020.0 207607.5 ;
      RECT  59330.0 207472.5 59400.0 207607.5 ;
      RECT  58940.0 206820.0 59010.0 207987.5 ;
      RECT  59275.0 206820.0 59345.0 207987.5 ;
      RECT  59645.0 206942.5 59722.5 207077.5 ;
      RECT  59847.5 206942.5 60050.0 207077.5 ;
      RECT  59645.0 207472.5 59722.5 207607.5 ;
      RECT  59980.0 207472.5 60102.5 207607.5 ;
      RECT  59655.0 206942.5 59725.0 207077.5 ;
      RECT  59845.0 206942.5 59915.0 207077.5 ;
      RECT  59655.0 207472.5 59725.0 207607.5 ;
      RECT  60035.0 207472.5 60105.0 207607.5 ;
      RECT  59645.0 206820.0 59715.0 207987.5 ;
      RECT  59980.0 206820.0 60050.0 207987.5 ;
      RECT  60350.0 206942.5 60427.5 207077.5 ;
      RECT  60552.5 206942.5 60755.0 207077.5 ;
      RECT  60350.0 207472.5 60427.5 207607.5 ;
      RECT  60685.0 207472.5 60807.5 207607.5 ;
      RECT  60360.0 206942.5 60430.0 207077.5 ;
      RECT  60550.0 206942.5 60620.0 207077.5 ;
      RECT  60360.0 207472.5 60430.0 207607.5 ;
      RECT  60740.0 207472.5 60810.0 207607.5 ;
      RECT  60350.0 206820.0 60420.0 207987.5 ;
      RECT  60685.0 206820.0 60755.0 207987.5 ;
      RECT  61055.0 206942.5 61132.5 207077.5 ;
      RECT  61257.5 206942.5 61460.0 207077.5 ;
      RECT  61055.0 207472.5 61132.5 207607.5 ;
      RECT  61390.0 207472.5 61512.5 207607.5 ;
      RECT  61065.0 206942.5 61135.0 207077.5 ;
      RECT  61255.0 206942.5 61325.0 207077.5 ;
      RECT  61065.0 207472.5 61135.0 207607.5 ;
      RECT  61445.0 207472.5 61515.0 207607.5 ;
      RECT  61055.0 206820.0 61125.0 207987.5 ;
      RECT  61390.0 206820.0 61460.0 207987.5 ;
      RECT  61760.0 206942.5 61837.5 207077.5 ;
      RECT  61962.5 206942.5 62165.0 207077.5 ;
      RECT  61760.0 207472.5 61837.5 207607.5 ;
      RECT  62095.0 207472.5 62217.5 207607.5 ;
      RECT  61770.0 206942.5 61840.0 207077.5 ;
      RECT  61960.0 206942.5 62030.0 207077.5 ;
      RECT  61770.0 207472.5 61840.0 207607.5 ;
      RECT  62150.0 207472.5 62220.0 207607.5 ;
      RECT  61760.0 206820.0 61830.0 207987.5 ;
      RECT  62095.0 206820.0 62165.0 207987.5 ;
      RECT  62465.0 206942.5 62542.5 207077.5 ;
      RECT  62667.5 206942.5 62870.0 207077.5 ;
      RECT  62465.0 207472.5 62542.5 207607.5 ;
      RECT  62800.0 207472.5 62922.5 207607.5 ;
      RECT  62475.0 206942.5 62545.0 207077.5 ;
      RECT  62665.0 206942.5 62735.0 207077.5 ;
      RECT  62475.0 207472.5 62545.0 207607.5 ;
      RECT  62855.0 207472.5 62925.0 207607.5 ;
      RECT  62465.0 206820.0 62535.0 207987.5 ;
      RECT  62800.0 206820.0 62870.0 207987.5 ;
      RECT  63170.0 206942.5 63247.5 207077.5 ;
      RECT  63372.5 206942.5 63575.0 207077.5 ;
      RECT  63170.0 207472.5 63247.5 207607.5 ;
      RECT  63505.0 207472.5 63627.5 207607.5 ;
      RECT  63180.0 206942.5 63250.0 207077.5 ;
      RECT  63370.0 206942.5 63440.0 207077.5 ;
      RECT  63180.0 207472.5 63250.0 207607.5 ;
      RECT  63560.0 207472.5 63630.0 207607.5 ;
      RECT  63170.0 206820.0 63240.0 207987.5 ;
      RECT  63505.0 206820.0 63575.0 207987.5 ;
      RECT  63875.0 206942.5 63952.5 207077.5 ;
      RECT  64077.5 206942.5 64280.0 207077.5 ;
      RECT  63875.0 207472.5 63952.5 207607.5 ;
      RECT  64210.0 207472.5 64332.5 207607.5 ;
      RECT  63885.0 206942.5 63955.0 207077.5 ;
      RECT  64075.0 206942.5 64145.0 207077.5 ;
      RECT  63885.0 207472.5 63955.0 207607.5 ;
      RECT  64265.0 207472.5 64335.0 207607.5 ;
      RECT  63875.0 206820.0 63945.0 207987.5 ;
      RECT  64210.0 206820.0 64280.0 207987.5 ;
      RECT  64580.0 206942.5 64657.5 207077.5 ;
      RECT  64782.5 206942.5 64985.0 207077.5 ;
      RECT  64580.0 207472.5 64657.5 207607.5 ;
      RECT  64915.0 207472.5 65037.5 207607.5 ;
      RECT  64590.0 206942.5 64660.0 207077.5 ;
      RECT  64780.0 206942.5 64850.0 207077.5 ;
      RECT  64590.0 207472.5 64660.0 207607.5 ;
      RECT  64970.0 207472.5 65040.0 207607.5 ;
      RECT  64580.0 206820.0 64650.0 207987.5 ;
      RECT  64915.0 206820.0 64985.0 207987.5 ;
      RECT  65285.0 206942.5 65362.5 207077.5 ;
      RECT  65487.5 206942.5 65690.0 207077.5 ;
      RECT  65285.0 207472.5 65362.5 207607.5 ;
      RECT  65620.0 207472.5 65742.5 207607.5 ;
      RECT  65295.0 206942.5 65365.0 207077.5 ;
      RECT  65485.0 206942.5 65555.0 207077.5 ;
      RECT  65295.0 207472.5 65365.0 207607.5 ;
      RECT  65675.0 207472.5 65745.0 207607.5 ;
      RECT  65285.0 206820.0 65355.0 207987.5 ;
      RECT  65620.0 206820.0 65690.0 207987.5 ;
      RECT  65990.0 206942.5 66067.5 207077.5 ;
      RECT  66192.5 206942.5 66395.0 207077.5 ;
      RECT  65990.0 207472.5 66067.5 207607.5 ;
      RECT  66325.0 207472.5 66447.5 207607.5 ;
      RECT  66000.0 206942.5 66070.0 207077.5 ;
      RECT  66190.0 206942.5 66260.0 207077.5 ;
      RECT  66000.0 207472.5 66070.0 207607.5 ;
      RECT  66380.0 207472.5 66450.0 207607.5 ;
      RECT  65990.0 206820.0 66060.0 207987.5 ;
      RECT  66325.0 206820.0 66395.0 207987.5 ;
      RECT  66695.0 206942.5 66772.5 207077.5 ;
      RECT  66897.5 206942.5 67100.0 207077.5 ;
      RECT  66695.0 207472.5 66772.5 207607.5 ;
      RECT  67030.0 207472.5 67152.5 207607.5 ;
      RECT  66705.0 206942.5 66775.0 207077.5 ;
      RECT  66895.0 206942.5 66965.0 207077.5 ;
      RECT  66705.0 207472.5 66775.0 207607.5 ;
      RECT  67085.0 207472.5 67155.0 207607.5 ;
      RECT  66695.0 206820.0 66765.0 207987.5 ;
      RECT  67030.0 206820.0 67100.0 207987.5 ;
      RECT  67400.0 206942.5 67477.5 207077.5 ;
      RECT  67602.5 206942.5 67805.0 207077.5 ;
      RECT  67400.0 207472.5 67477.5 207607.5 ;
      RECT  67735.0 207472.5 67857.5 207607.5 ;
      RECT  67410.0 206942.5 67480.0 207077.5 ;
      RECT  67600.0 206942.5 67670.0 207077.5 ;
      RECT  67410.0 207472.5 67480.0 207607.5 ;
      RECT  67790.0 207472.5 67860.0 207607.5 ;
      RECT  67400.0 206820.0 67470.0 207987.5 ;
      RECT  67735.0 206820.0 67805.0 207987.5 ;
      RECT  68105.0 206942.5 68182.5 207077.5 ;
      RECT  68307.5 206942.5 68510.0 207077.5 ;
      RECT  68105.0 207472.5 68182.5 207607.5 ;
      RECT  68440.0 207472.5 68562.5 207607.5 ;
      RECT  68115.0 206942.5 68185.0 207077.5 ;
      RECT  68305.0 206942.5 68375.0 207077.5 ;
      RECT  68115.0 207472.5 68185.0 207607.5 ;
      RECT  68495.0 207472.5 68565.0 207607.5 ;
      RECT  68105.0 206820.0 68175.0 207987.5 ;
      RECT  68440.0 206820.0 68510.0 207987.5 ;
      RECT  68810.0 206942.5 68887.5 207077.5 ;
      RECT  69012.5 206942.5 69215.0 207077.5 ;
      RECT  68810.0 207472.5 68887.5 207607.5 ;
      RECT  69145.0 207472.5 69267.5 207607.5 ;
      RECT  68820.0 206942.5 68890.0 207077.5 ;
      RECT  69010.0 206942.5 69080.0 207077.5 ;
      RECT  68820.0 207472.5 68890.0 207607.5 ;
      RECT  69200.0 207472.5 69270.0 207607.5 ;
      RECT  68810.0 206820.0 68880.0 207987.5 ;
      RECT  69145.0 206820.0 69215.0 207987.5 ;
      RECT  69515.0 206942.5 69592.5 207077.5 ;
      RECT  69717.5 206942.5 69920.0 207077.5 ;
      RECT  69515.0 207472.5 69592.5 207607.5 ;
      RECT  69850.0 207472.5 69972.5 207607.5 ;
      RECT  69525.0 206942.5 69595.0 207077.5 ;
      RECT  69715.0 206942.5 69785.0 207077.5 ;
      RECT  69525.0 207472.5 69595.0 207607.5 ;
      RECT  69905.0 207472.5 69975.0 207607.5 ;
      RECT  69515.0 206820.0 69585.0 207987.5 ;
      RECT  69850.0 206820.0 69920.0 207987.5 ;
      RECT  70220.0 206942.5 70297.5 207077.5 ;
      RECT  70422.5 206942.5 70625.0 207077.5 ;
      RECT  70220.0 207472.5 70297.5 207607.5 ;
      RECT  70555.0 207472.5 70677.5 207607.5 ;
      RECT  70230.0 206942.5 70300.0 207077.5 ;
      RECT  70420.0 206942.5 70490.0 207077.5 ;
      RECT  70230.0 207472.5 70300.0 207607.5 ;
      RECT  70610.0 207472.5 70680.0 207607.5 ;
      RECT  70220.0 206820.0 70290.0 207987.5 ;
      RECT  70555.0 206820.0 70625.0 207987.5 ;
      RECT  70925.0 206942.5 71002.5 207077.5 ;
      RECT  71127.5 206942.5 71330.0 207077.5 ;
      RECT  70925.0 207472.5 71002.5 207607.5 ;
      RECT  71260.0 207472.5 71382.5 207607.5 ;
      RECT  70935.0 206942.5 71005.0 207077.5 ;
      RECT  71125.0 206942.5 71195.0 207077.5 ;
      RECT  70935.0 207472.5 71005.0 207607.5 ;
      RECT  71315.0 207472.5 71385.0 207607.5 ;
      RECT  70925.0 206820.0 70995.0 207987.5 ;
      RECT  71260.0 206820.0 71330.0 207987.5 ;
      RECT  71630.0 206942.5 71707.5 207077.5 ;
      RECT  71832.5 206942.5 72035.0 207077.5 ;
      RECT  71630.0 207472.5 71707.5 207607.5 ;
      RECT  71965.0 207472.5 72087.5 207607.5 ;
      RECT  71640.0 206942.5 71710.0 207077.5 ;
      RECT  71830.0 206942.5 71900.0 207077.5 ;
      RECT  71640.0 207472.5 71710.0 207607.5 ;
      RECT  72020.0 207472.5 72090.0 207607.5 ;
      RECT  71630.0 206820.0 71700.0 207987.5 ;
      RECT  71965.0 206820.0 72035.0 207987.5 ;
      RECT  72335.0 206942.5 72412.5 207077.5 ;
      RECT  72537.5 206942.5 72740.0 207077.5 ;
      RECT  72335.0 207472.5 72412.5 207607.5 ;
      RECT  72670.0 207472.5 72792.5 207607.5 ;
      RECT  72345.0 206942.5 72415.0 207077.5 ;
      RECT  72535.0 206942.5 72605.0 207077.5 ;
      RECT  72345.0 207472.5 72415.0 207607.5 ;
      RECT  72725.0 207472.5 72795.0 207607.5 ;
      RECT  72335.0 206820.0 72405.0 207987.5 ;
      RECT  72670.0 206820.0 72740.0 207987.5 ;
      RECT  73040.0 206942.5 73117.5 207077.5 ;
      RECT  73242.5 206942.5 73445.0 207077.5 ;
      RECT  73040.0 207472.5 73117.5 207607.5 ;
      RECT  73375.0 207472.5 73497.5 207607.5 ;
      RECT  73050.0 206942.5 73120.0 207077.5 ;
      RECT  73240.0 206942.5 73310.0 207077.5 ;
      RECT  73050.0 207472.5 73120.0 207607.5 ;
      RECT  73430.0 207472.5 73500.0 207607.5 ;
      RECT  73040.0 206820.0 73110.0 207987.5 ;
      RECT  73375.0 206820.0 73445.0 207987.5 ;
      RECT  73745.0 206942.5 73822.5 207077.5 ;
      RECT  73947.5 206942.5 74150.0 207077.5 ;
      RECT  73745.0 207472.5 73822.5 207607.5 ;
      RECT  74080.0 207472.5 74202.5 207607.5 ;
      RECT  73755.0 206942.5 73825.0 207077.5 ;
      RECT  73945.0 206942.5 74015.0 207077.5 ;
      RECT  73755.0 207472.5 73825.0 207607.5 ;
      RECT  74135.0 207472.5 74205.0 207607.5 ;
      RECT  73745.0 206820.0 73815.0 207987.5 ;
      RECT  74080.0 206820.0 74150.0 207987.5 ;
      RECT  74450.0 206942.5 74527.5 207077.5 ;
      RECT  74652.5 206942.5 74855.0 207077.5 ;
      RECT  74450.0 207472.5 74527.5 207607.5 ;
      RECT  74785.0 207472.5 74907.5 207607.5 ;
      RECT  74460.0 206942.5 74530.0 207077.5 ;
      RECT  74650.0 206942.5 74720.0 207077.5 ;
      RECT  74460.0 207472.5 74530.0 207607.5 ;
      RECT  74840.0 207472.5 74910.0 207607.5 ;
      RECT  74450.0 206820.0 74520.0 207987.5 ;
      RECT  74785.0 206820.0 74855.0 207987.5 ;
      RECT  75155.0 206942.5 75232.5 207077.5 ;
      RECT  75357.5 206942.5 75560.0 207077.5 ;
      RECT  75155.0 207472.5 75232.5 207607.5 ;
      RECT  75490.0 207472.5 75612.5 207607.5 ;
      RECT  75165.0 206942.5 75235.0 207077.5 ;
      RECT  75355.0 206942.5 75425.0 207077.5 ;
      RECT  75165.0 207472.5 75235.0 207607.5 ;
      RECT  75545.0 207472.5 75615.0 207607.5 ;
      RECT  75155.0 206820.0 75225.0 207987.5 ;
      RECT  75490.0 206820.0 75560.0 207987.5 ;
      RECT  75860.0 206942.5 75937.5 207077.5 ;
      RECT  76062.5 206942.5 76265.0 207077.5 ;
      RECT  75860.0 207472.5 75937.5 207607.5 ;
      RECT  76195.0 207472.5 76317.5 207607.5 ;
      RECT  75870.0 206942.5 75940.0 207077.5 ;
      RECT  76060.0 206942.5 76130.0 207077.5 ;
      RECT  75870.0 207472.5 75940.0 207607.5 ;
      RECT  76250.0 207472.5 76320.0 207607.5 ;
      RECT  75860.0 206820.0 75930.0 207987.5 ;
      RECT  76195.0 206820.0 76265.0 207987.5 ;
      RECT  76565.0 206942.5 76642.5 207077.5 ;
      RECT  76767.5 206942.5 76970.0 207077.5 ;
      RECT  76565.0 207472.5 76642.5 207607.5 ;
      RECT  76900.0 207472.5 77022.5 207607.5 ;
      RECT  76575.0 206942.5 76645.0 207077.5 ;
      RECT  76765.0 206942.5 76835.0 207077.5 ;
      RECT  76575.0 207472.5 76645.0 207607.5 ;
      RECT  76955.0 207472.5 77025.0 207607.5 ;
      RECT  76565.0 206820.0 76635.0 207987.5 ;
      RECT  76900.0 206820.0 76970.0 207987.5 ;
      RECT  77270.0 206942.5 77347.5 207077.5 ;
      RECT  77472.5 206942.5 77675.0 207077.5 ;
      RECT  77270.0 207472.5 77347.5 207607.5 ;
      RECT  77605.0 207472.5 77727.5 207607.5 ;
      RECT  77280.0 206942.5 77350.0 207077.5 ;
      RECT  77470.0 206942.5 77540.0 207077.5 ;
      RECT  77280.0 207472.5 77350.0 207607.5 ;
      RECT  77660.0 207472.5 77730.0 207607.5 ;
      RECT  77270.0 206820.0 77340.0 207987.5 ;
      RECT  77605.0 206820.0 77675.0 207987.5 ;
      RECT  77975.0 206942.5 78052.5 207077.5 ;
      RECT  78177.5 206942.5 78380.0 207077.5 ;
      RECT  77975.0 207472.5 78052.5 207607.5 ;
      RECT  78310.0 207472.5 78432.5 207607.5 ;
      RECT  77985.0 206942.5 78055.0 207077.5 ;
      RECT  78175.0 206942.5 78245.0 207077.5 ;
      RECT  77985.0 207472.5 78055.0 207607.5 ;
      RECT  78365.0 207472.5 78435.0 207607.5 ;
      RECT  77975.0 206820.0 78045.0 207987.5 ;
      RECT  78310.0 206820.0 78380.0 207987.5 ;
      RECT  78680.0 206942.5 78757.5 207077.5 ;
      RECT  78882.5 206942.5 79085.0 207077.5 ;
      RECT  78680.0 207472.5 78757.5 207607.5 ;
      RECT  79015.0 207472.5 79137.5 207607.5 ;
      RECT  78690.0 206942.5 78760.0 207077.5 ;
      RECT  78880.0 206942.5 78950.0 207077.5 ;
      RECT  78690.0 207472.5 78760.0 207607.5 ;
      RECT  79070.0 207472.5 79140.0 207607.5 ;
      RECT  78680.0 206820.0 78750.0 207987.5 ;
      RECT  79015.0 206820.0 79085.0 207987.5 ;
      RECT  79385.0 206942.5 79462.5 207077.5 ;
      RECT  79587.5 206942.5 79790.0 207077.5 ;
      RECT  79385.0 207472.5 79462.5 207607.5 ;
      RECT  79720.0 207472.5 79842.5 207607.5 ;
      RECT  79395.0 206942.5 79465.0 207077.5 ;
      RECT  79585.0 206942.5 79655.0 207077.5 ;
      RECT  79395.0 207472.5 79465.0 207607.5 ;
      RECT  79775.0 207472.5 79845.0 207607.5 ;
      RECT  79385.0 206820.0 79455.0 207987.5 ;
      RECT  79720.0 206820.0 79790.0 207987.5 ;
      RECT  80090.0 206942.5 80167.5 207077.5 ;
      RECT  80292.5 206942.5 80495.0 207077.5 ;
      RECT  80090.0 207472.5 80167.5 207607.5 ;
      RECT  80425.0 207472.5 80547.5 207607.5 ;
      RECT  80100.0 206942.5 80170.0 207077.5 ;
      RECT  80290.0 206942.5 80360.0 207077.5 ;
      RECT  80100.0 207472.5 80170.0 207607.5 ;
      RECT  80480.0 207472.5 80550.0 207607.5 ;
      RECT  80090.0 206820.0 80160.0 207987.5 ;
      RECT  80425.0 206820.0 80495.0 207987.5 ;
      RECT  80795.0 206942.5 80872.5 207077.5 ;
      RECT  80997.5 206942.5 81200.0 207077.5 ;
      RECT  80795.0 207472.5 80872.5 207607.5 ;
      RECT  81130.0 207472.5 81252.5 207607.5 ;
      RECT  80805.0 206942.5 80875.0 207077.5 ;
      RECT  80995.0 206942.5 81065.0 207077.5 ;
      RECT  80805.0 207472.5 80875.0 207607.5 ;
      RECT  81185.0 207472.5 81255.0 207607.5 ;
      RECT  80795.0 206820.0 80865.0 207987.5 ;
      RECT  81130.0 206820.0 81200.0 207987.5 ;
      RECT  81500.0 206942.5 81577.5 207077.5 ;
      RECT  81702.5 206942.5 81905.0 207077.5 ;
      RECT  81500.0 207472.5 81577.5 207607.5 ;
      RECT  81835.0 207472.5 81957.5 207607.5 ;
      RECT  81510.0 206942.5 81580.0 207077.5 ;
      RECT  81700.0 206942.5 81770.0 207077.5 ;
      RECT  81510.0 207472.5 81580.0 207607.5 ;
      RECT  81890.0 207472.5 81960.0 207607.5 ;
      RECT  81500.0 206820.0 81570.0 207987.5 ;
      RECT  81835.0 206820.0 81905.0 207987.5 ;
      RECT  82205.0 206942.5 82282.5 207077.5 ;
      RECT  82407.5 206942.5 82610.0 207077.5 ;
      RECT  82205.0 207472.5 82282.5 207607.5 ;
      RECT  82540.0 207472.5 82662.5 207607.5 ;
      RECT  82215.0 206942.5 82285.0 207077.5 ;
      RECT  82405.0 206942.5 82475.0 207077.5 ;
      RECT  82215.0 207472.5 82285.0 207607.5 ;
      RECT  82595.0 207472.5 82665.0 207607.5 ;
      RECT  82205.0 206820.0 82275.0 207987.5 ;
      RECT  82540.0 206820.0 82610.0 207987.5 ;
      RECT  82910.0 206942.5 82987.5 207077.5 ;
      RECT  83112.5 206942.5 83315.0 207077.5 ;
      RECT  82910.0 207472.5 82987.5 207607.5 ;
      RECT  83245.0 207472.5 83367.5 207607.5 ;
      RECT  82920.0 206942.5 82990.0 207077.5 ;
      RECT  83110.0 206942.5 83180.0 207077.5 ;
      RECT  82920.0 207472.5 82990.0 207607.5 ;
      RECT  83300.0 207472.5 83370.0 207607.5 ;
      RECT  82910.0 206820.0 82980.0 207987.5 ;
      RECT  83245.0 206820.0 83315.0 207987.5 ;
      RECT  83615.0 206942.5 83692.5 207077.5 ;
      RECT  83817.5 206942.5 84020.0 207077.5 ;
      RECT  83615.0 207472.5 83692.5 207607.5 ;
      RECT  83950.0 207472.5 84072.5 207607.5 ;
      RECT  83625.0 206942.5 83695.0 207077.5 ;
      RECT  83815.0 206942.5 83885.0 207077.5 ;
      RECT  83625.0 207472.5 83695.0 207607.5 ;
      RECT  84005.0 207472.5 84075.0 207607.5 ;
      RECT  83615.0 206820.0 83685.0 207987.5 ;
      RECT  83950.0 206820.0 84020.0 207987.5 ;
      RECT  84320.0 206942.5 84397.5 207077.5 ;
      RECT  84522.5 206942.5 84725.0 207077.5 ;
      RECT  84320.0 207472.5 84397.5 207607.5 ;
      RECT  84655.0 207472.5 84777.5 207607.5 ;
      RECT  84330.0 206942.5 84400.0 207077.5 ;
      RECT  84520.0 206942.5 84590.0 207077.5 ;
      RECT  84330.0 207472.5 84400.0 207607.5 ;
      RECT  84710.0 207472.5 84780.0 207607.5 ;
      RECT  84320.0 206820.0 84390.0 207987.5 ;
      RECT  84655.0 206820.0 84725.0 207987.5 ;
      RECT  85025.0 206942.5 85102.5 207077.5 ;
      RECT  85227.5 206942.5 85430.0 207077.5 ;
      RECT  85025.0 207472.5 85102.5 207607.5 ;
      RECT  85360.0 207472.5 85482.5 207607.5 ;
      RECT  85035.0 206942.5 85105.0 207077.5 ;
      RECT  85225.0 206942.5 85295.0 207077.5 ;
      RECT  85035.0 207472.5 85105.0 207607.5 ;
      RECT  85415.0 207472.5 85485.0 207607.5 ;
      RECT  85025.0 206820.0 85095.0 207987.5 ;
      RECT  85360.0 206820.0 85430.0 207987.5 ;
      RECT  85730.0 206942.5 85807.5 207077.5 ;
      RECT  85932.5 206942.5 86135.0 207077.5 ;
      RECT  85730.0 207472.5 85807.5 207607.5 ;
      RECT  86065.0 207472.5 86187.5 207607.5 ;
      RECT  85740.0 206942.5 85810.0 207077.5 ;
      RECT  85930.0 206942.5 86000.0 207077.5 ;
      RECT  85740.0 207472.5 85810.0 207607.5 ;
      RECT  86120.0 207472.5 86190.0 207607.5 ;
      RECT  85730.0 206820.0 85800.0 207987.5 ;
      RECT  86065.0 206820.0 86135.0 207987.5 ;
      RECT  86435.0 206942.5 86512.5 207077.5 ;
      RECT  86637.5 206942.5 86840.0 207077.5 ;
      RECT  86435.0 207472.5 86512.5 207607.5 ;
      RECT  86770.0 207472.5 86892.5 207607.5 ;
      RECT  86445.0 206942.5 86515.0 207077.5 ;
      RECT  86635.0 206942.5 86705.0 207077.5 ;
      RECT  86445.0 207472.5 86515.0 207607.5 ;
      RECT  86825.0 207472.5 86895.0 207607.5 ;
      RECT  86435.0 206820.0 86505.0 207987.5 ;
      RECT  86770.0 206820.0 86840.0 207987.5 ;
      RECT  87140.0 206942.5 87217.5 207077.5 ;
      RECT  87342.5 206942.5 87545.0 207077.5 ;
      RECT  87140.0 207472.5 87217.5 207607.5 ;
      RECT  87475.0 207472.5 87597.5 207607.5 ;
      RECT  87150.0 206942.5 87220.0 207077.5 ;
      RECT  87340.0 206942.5 87410.0 207077.5 ;
      RECT  87150.0 207472.5 87220.0 207607.5 ;
      RECT  87530.0 207472.5 87600.0 207607.5 ;
      RECT  87140.0 206820.0 87210.0 207987.5 ;
      RECT  87475.0 206820.0 87545.0 207987.5 ;
      RECT  87845.0 206942.5 87922.5 207077.5 ;
      RECT  88047.5 206942.5 88250.0 207077.5 ;
      RECT  87845.0 207472.5 87922.5 207607.5 ;
      RECT  88180.0 207472.5 88302.5 207607.5 ;
      RECT  87855.0 206942.5 87925.0 207077.5 ;
      RECT  88045.0 206942.5 88115.0 207077.5 ;
      RECT  87855.0 207472.5 87925.0 207607.5 ;
      RECT  88235.0 207472.5 88305.0 207607.5 ;
      RECT  87845.0 206820.0 87915.0 207987.5 ;
      RECT  88180.0 206820.0 88250.0 207987.5 ;
      RECT  88550.0 206942.5 88627.5 207077.5 ;
      RECT  88752.5 206942.5 88955.0 207077.5 ;
      RECT  88550.0 207472.5 88627.5 207607.5 ;
      RECT  88885.0 207472.5 89007.5 207607.5 ;
      RECT  88560.0 206942.5 88630.0 207077.5 ;
      RECT  88750.0 206942.5 88820.0 207077.5 ;
      RECT  88560.0 207472.5 88630.0 207607.5 ;
      RECT  88940.0 207472.5 89010.0 207607.5 ;
      RECT  88550.0 206820.0 88620.0 207987.5 ;
      RECT  88885.0 206820.0 88955.0 207987.5 ;
      RECT  89255.0 206942.5 89332.5 207077.5 ;
      RECT  89457.5 206942.5 89660.0 207077.5 ;
      RECT  89255.0 207472.5 89332.5 207607.5 ;
      RECT  89590.0 207472.5 89712.5 207607.5 ;
      RECT  89265.0 206942.5 89335.0 207077.5 ;
      RECT  89455.0 206942.5 89525.0 207077.5 ;
      RECT  89265.0 207472.5 89335.0 207607.5 ;
      RECT  89645.0 207472.5 89715.0 207607.5 ;
      RECT  89255.0 206820.0 89325.0 207987.5 ;
      RECT  89590.0 206820.0 89660.0 207987.5 ;
      RECT  89960.0 206942.5 90037.5 207077.5 ;
      RECT  90162.5 206942.5 90365.0 207077.5 ;
      RECT  89960.0 207472.5 90037.5 207607.5 ;
      RECT  90295.0 207472.5 90417.5 207607.5 ;
      RECT  89970.0 206942.5 90040.0 207077.5 ;
      RECT  90160.0 206942.5 90230.0 207077.5 ;
      RECT  89970.0 207472.5 90040.0 207607.5 ;
      RECT  90350.0 207472.5 90420.0 207607.5 ;
      RECT  89960.0 206820.0 90030.0 207987.5 ;
      RECT  90295.0 206820.0 90365.0 207987.5 ;
      RECT  90665.0 206942.5 90742.5 207077.5 ;
      RECT  90867.5 206942.5 91070.0 207077.5 ;
      RECT  90665.0 207472.5 90742.5 207607.5 ;
      RECT  91000.0 207472.5 91122.5 207607.5 ;
      RECT  90675.0 206942.5 90745.0 207077.5 ;
      RECT  90865.0 206942.5 90935.0 207077.5 ;
      RECT  90675.0 207472.5 90745.0 207607.5 ;
      RECT  91055.0 207472.5 91125.0 207607.5 ;
      RECT  90665.0 206820.0 90735.0 207987.5 ;
      RECT  91000.0 206820.0 91070.0 207987.5 ;
      RECT  91370.0 206942.5 91447.5 207077.5 ;
      RECT  91572.5 206942.5 91775.0 207077.5 ;
      RECT  91370.0 207472.5 91447.5 207607.5 ;
      RECT  91705.0 207472.5 91827.5 207607.5 ;
      RECT  91380.0 206942.5 91450.0 207077.5 ;
      RECT  91570.0 206942.5 91640.0 207077.5 ;
      RECT  91380.0 207472.5 91450.0 207607.5 ;
      RECT  91760.0 207472.5 91830.0 207607.5 ;
      RECT  91370.0 206820.0 91440.0 207987.5 ;
      RECT  91705.0 206820.0 91775.0 207987.5 ;
      RECT  92075.0 206942.5 92152.5 207077.5 ;
      RECT  92277.5 206942.5 92480.0 207077.5 ;
      RECT  92075.0 207472.5 92152.5 207607.5 ;
      RECT  92410.0 207472.5 92532.5 207607.5 ;
      RECT  92085.0 206942.5 92155.0 207077.5 ;
      RECT  92275.0 206942.5 92345.0 207077.5 ;
      RECT  92085.0 207472.5 92155.0 207607.5 ;
      RECT  92465.0 207472.5 92535.0 207607.5 ;
      RECT  92075.0 206820.0 92145.0 207987.5 ;
      RECT  92410.0 206820.0 92480.0 207987.5 ;
      RECT  92780.0 206942.5 92857.5 207077.5 ;
      RECT  92982.5 206942.5 93185.0 207077.5 ;
      RECT  92780.0 207472.5 92857.5 207607.5 ;
      RECT  93115.0 207472.5 93237.5 207607.5 ;
      RECT  92790.0 206942.5 92860.0 207077.5 ;
      RECT  92980.0 206942.5 93050.0 207077.5 ;
      RECT  92790.0 207472.5 92860.0 207607.5 ;
      RECT  93170.0 207472.5 93240.0 207607.5 ;
      RECT  92780.0 206820.0 92850.0 207987.5 ;
      RECT  93115.0 206820.0 93185.0 207987.5 ;
      RECT  93485.0 206942.5 93562.5 207077.5 ;
      RECT  93687.5 206942.5 93890.0 207077.5 ;
      RECT  93485.0 207472.5 93562.5 207607.5 ;
      RECT  93820.0 207472.5 93942.5 207607.5 ;
      RECT  93495.0 206942.5 93565.0 207077.5 ;
      RECT  93685.0 206942.5 93755.0 207077.5 ;
      RECT  93495.0 207472.5 93565.0 207607.5 ;
      RECT  93875.0 207472.5 93945.0 207607.5 ;
      RECT  93485.0 206820.0 93555.0 207987.5 ;
      RECT  93820.0 206820.0 93890.0 207987.5 ;
      RECT  94190.0 206942.5 94267.5 207077.5 ;
      RECT  94392.5 206942.5 94595.0 207077.5 ;
      RECT  94190.0 207472.5 94267.5 207607.5 ;
      RECT  94525.0 207472.5 94647.5 207607.5 ;
      RECT  94200.0 206942.5 94270.0 207077.5 ;
      RECT  94390.0 206942.5 94460.0 207077.5 ;
      RECT  94200.0 207472.5 94270.0 207607.5 ;
      RECT  94580.0 207472.5 94650.0 207607.5 ;
      RECT  94190.0 206820.0 94260.0 207987.5 ;
      RECT  94525.0 206820.0 94595.0 207987.5 ;
      RECT  94895.0 206942.5 94972.5 207077.5 ;
      RECT  95097.5 206942.5 95300.0 207077.5 ;
      RECT  94895.0 207472.5 94972.5 207607.5 ;
      RECT  95230.0 207472.5 95352.5 207607.5 ;
      RECT  94905.0 206942.5 94975.0 207077.5 ;
      RECT  95095.0 206942.5 95165.0 207077.5 ;
      RECT  94905.0 207472.5 94975.0 207607.5 ;
      RECT  95285.0 207472.5 95355.0 207607.5 ;
      RECT  94895.0 206820.0 94965.0 207987.5 ;
      RECT  95230.0 206820.0 95300.0 207987.5 ;
      RECT  95600.0 206942.5 95677.5 207077.5 ;
      RECT  95802.5 206942.5 96005.0 207077.5 ;
      RECT  95600.0 207472.5 95677.5 207607.5 ;
      RECT  95935.0 207472.5 96057.5 207607.5 ;
      RECT  95610.0 206942.5 95680.0 207077.5 ;
      RECT  95800.0 206942.5 95870.0 207077.5 ;
      RECT  95610.0 207472.5 95680.0 207607.5 ;
      RECT  95990.0 207472.5 96060.0 207607.5 ;
      RECT  95600.0 206820.0 95670.0 207987.5 ;
      RECT  95935.0 206820.0 96005.0 207987.5 ;
      RECT  96305.0 206942.5 96382.5 207077.5 ;
      RECT  96507.5 206942.5 96710.0 207077.5 ;
      RECT  96305.0 207472.5 96382.5 207607.5 ;
      RECT  96640.0 207472.5 96762.5 207607.5 ;
      RECT  96315.0 206942.5 96385.0 207077.5 ;
      RECT  96505.0 206942.5 96575.0 207077.5 ;
      RECT  96315.0 207472.5 96385.0 207607.5 ;
      RECT  96695.0 207472.5 96765.0 207607.5 ;
      RECT  96305.0 206820.0 96375.0 207987.5 ;
      RECT  96640.0 206820.0 96710.0 207987.5 ;
      RECT  97010.0 206942.5 97087.5 207077.5 ;
      RECT  97212.5 206942.5 97415.0 207077.5 ;
      RECT  97010.0 207472.5 97087.5 207607.5 ;
      RECT  97345.0 207472.5 97467.5 207607.5 ;
      RECT  97020.0 206942.5 97090.0 207077.5 ;
      RECT  97210.0 206942.5 97280.0 207077.5 ;
      RECT  97020.0 207472.5 97090.0 207607.5 ;
      RECT  97400.0 207472.5 97470.0 207607.5 ;
      RECT  97010.0 206820.0 97080.0 207987.5 ;
      RECT  97345.0 206820.0 97415.0 207987.5 ;
      RECT  97715.0 206942.5 97792.5 207077.5 ;
      RECT  97917.5 206942.5 98120.0 207077.5 ;
      RECT  97715.0 207472.5 97792.5 207607.5 ;
      RECT  98050.0 207472.5 98172.5 207607.5 ;
      RECT  97725.0 206942.5 97795.0 207077.5 ;
      RECT  97915.0 206942.5 97985.0 207077.5 ;
      RECT  97725.0 207472.5 97795.0 207607.5 ;
      RECT  98105.0 207472.5 98175.0 207607.5 ;
      RECT  97715.0 206820.0 97785.0 207987.5 ;
      RECT  98050.0 206820.0 98120.0 207987.5 ;
      RECT  98420.0 206942.5 98497.5 207077.5 ;
      RECT  98622.5 206942.5 98825.0 207077.5 ;
      RECT  98420.0 207472.5 98497.5 207607.5 ;
      RECT  98755.0 207472.5 98877.5 207607.5 ;
      RECT  98430.0 206942.5 98500.0 207077.5 ;
      RECT  98620.0 206942.5 98690.0 207077.5 ;
      RECT  98430.0 207472.5 98500.0 207607.5 ;
      RECT  98810.0 207472.5 98880.0 207607.5 ;
      RECT  98420.0 206820.0 98490.0 207987.5 ;
      RECT  98755.0 206820.0 98825.0 207987.5 ;
      RECT  99125.0 206942.5 99202.5 207077.5 ;
      RECT  99327.5 206942.5 99530.0 207077.5 ;
      RECT  99125.0 207472.5 99202.5 207607.5 ;
      RECT  99460.0 207472.5 99582.5 207607.5 ;
      RECT  99135.0 206942.5 99205.0 207077.5 ;
      RECT  99325.0 206942.5 99395.0 207077.5 ;
      RECT  99135.0 207472.5 99205.0 207607.5 ;
      RECT  99515.0 207472.5 99585.0 207607.5 ;
      RECT  99125.0 206820.0 99195.0 207987.5 ;
      RECT  99460.0 206820.0 99530.0 207987.5 ;
      RECT  99830.0 206942.5 99907.5 207077.5 ;
      RECT  100032.5 206942.5 100235.0 207077.5 ;
      RECT  99830.0 207472.5 99907.5 207607.5 ;
      RECT  100165.0 207472.5 100287.5 207607.5 ;
      RECT  99840.0 206942.5 99910.0 207077.5 ;
      RECT  100030.0 206942.5 100100.0 207077.5 ;
      RECT  99840.0 207472.5 99910.0 207607.5 ;
      RECT  100220.0 207472.5 100290.0 207607.5 ;
      RECT  99830.0 206820.0 99900.0 207987.5 ;
      RECT  100165.0 206820.0 100235.0 207987.5 ;
      RECT  100535.0 206942.5 100612.5 207077.5 ;
      RECT  100737.5 206942.5 100940.0 207077.5 ;
      RECT  100535.0 207472.5 100612.5 207607.5 ;
      RECT  100870.0 207472.5 100992.5 207607.5 ;
      RECT  100545.0 206942.5 100615.0 207077.5 ;
      RECT  100735.0 206942.5 100805.0 207077.5 ;
      RECT  100545.0 207472.5 100615.0 207607.5 ;
      RECT  100925.0 207472.5 100995.0 207607.5 ;
      RECT  100535.0 206820.0 100605.0 207987.5 ;
      RECT  100870.0 206820.0 100940.0 207987.5 ;
      RECT  101240.0 206942.5 101317.5 207077.5 ;
      RECT  101442.5 206942.5 101645.0 207077.5 ;
      RECT  101240.0 207472.5 101317.5 207607.5 ;
      RECT  101575.0 207472.5 101697.5 207607.5 ;
      RECT  101250.0 206942.5 101320.0 207077.5 ;
      RECT  101440.0 206942.5 101510.0 207077.5 ;
      RECT  101250.0 207472.5 101320.0 207607.5 ;
      RECT  101630.0 207472.5 101700.0 207607.5 ;
      RECT  101240.0 206820.0 101310.0 207987.5 ;
      RECT  101575.0 206820.0 101645.0 207987.5 ;
      RECT  101945.0 206942.5 102022.5 207077.5 ;
      RECT  102147.5 206942.5 102350.0 207077.5 ;
      RECT  101945.0 207472.5 102022.5 207607.5 ;
      RECT  102280.0 207472.5 102402.5 207607.5 ;
      RECT  101955.0 206942.5 102025.0 207077.5 ;
      RECT  102145.0 206942.5 102215.0 207077.5 ;
      RECT  101955.0 207472.5 102025.0 207607.5 ;
      RECT  102335.0 207472.5 102405.0 207607.5 ;
      RECT  101945.0 206820.0 102015.0 207987.5 ;
      RECT  102280.0 206820.0 102350.0 207987.5 ;
      RECT  102650.0 206942.5 102727.5 207077.5 ;
      RECT  102852.5 206942.5 103055.0 207077.5 ;
      RECT  102650.0 207472.5 102727.5 207607.5 ;
      RECT  102985.0 207472.5 103107.5 207607.5 ;
      RECT  102660.0 206942.5 102730.0 207077.5 ;
      RECT  102850.0 206942.5 102920.0 207077.5 ;
      RECT  102660.0 207472.5 102730.0 207607.5 ;
      RECT  103040.0 207472.5 103110.0 207607.5 ;
      RECT  102650.0 206820.0 102720.0 207987.5 ;
      RECT  102985.0 206820.0 103055.0 207987.5 ;
      RECT  103355.0 206942.5 103432.5 207077.5 ;
      RECT  103557.5 206942.5 103760.0 207077.5 ;
      RECT  103355.0 207472.5 103432.5 207607.5 ;
      RECT  103690.0 207472.5 103812.5 207607.5 ;
      RECT  103365.0 206942.5 103435.0 207077.5 ;
      RECT  103555.0 206942.5 103625.0 207077.5 ;
      RECT  103365.0 207472.5 103435.0 207607.5 ;
      RECT  103745.0 207472.5 103815.0 207607.5 ;
      RECT  103355.0 206820.0 103425.0 207987.5 ;
      RECT  103690.0 206820.0 103760.0 207987.5 ;
      RECT  104060.0 206942.5 104137.5 207077.5 ;
      RECT  104262.5 206942.5 104465.0 207077.5 ;
      RECT  104060.0 207472.5 104137.5 207607.5 ;
      RECT  104395.0 207472.5 104517.5 207607.5 ;
      RECT  104070.0 206942.5 104140.0 207077.5 ;
      RECT  104260.0 206942.5 104330.0 207077.5 ;
      RECT  104070.0 207472.5 104140.0 207607.5 ;
      RECT  104450.0 207472.5 104520.0 207607.5 ;
      RECT  104060.0 206820.0 104130.0 207987.5 ;
      RECT  104395.0 206820.0 104465.0 207987.5 ;
      RECT  104765.0 206942.5 104842.5 207077.5 ;
      RECT  104967.5 206942.5 105170.0 207077.5 ;
      RECT  104765.0 207472.5 104842.5 207607.5 ;
      RECT  105100.0 207472.5 105222.5 207607.5 ;
      RECT  104775.0 206942.5 104845.0 207077.5 ;
      RECT  104965.0 206942.5 105035.0 207077.5 ;
      RECT  104775.0 207472.5 104845.0 207607.5 ;
      RECT  105155.0 207472.5 105225.0 207607.5 ;
      RECT  104765.0 206820.0 104835.0 207987.5 ;
      RECT  105100.0 206820.0 105170.0 207987.5 ;
      RECT  105470.0 206942.5 105547.5 207077.5 ;
      RECT  105672.5 206942.5 105875.0 207077.5 ;
      RECT  105470.0 207472.5 105547.5 207607.5 ;
      RECT  105805.0 207472.5 105927.5 207607.5 ;
      RECT  105480.0 206942.5 105550.0 207077.5 ;
      RECT  105670.0 206942.5 105740.0 207077.5 ;
      RECT  105480.0 207472.5 105550.0 207607.5 ;
      RECT  105860.0 207472.5 105930.0 207607.5 ;
      RECT  105470.0 206820.0 105540.0 207987.5 ;
      RECT  105805.0 206820.0 105875.0 207987.5 ;
      RECT  106175.0 206942.5 106252.5 207077.5 ;
      RECT  106377.5 206942.5 106580.0 207077.5 ;
      RECT  106175.0 207472.5 106252.5 207607.5 ;
      RECT  106510.0 207472.5 106632.5 207607.5 ;
      RECT  106185.0 206942.5 106255.0 207077.5 ;
      RECT  106375.0 206942.5 106445.0 207077.5 ;
      RECT  106185.0 207472.5 106255.0 207607.5 ;
      RECT  106565.0 207472.5 106635.0 207607.5 ;
      RECT  106175.0 206820.0 106245.0 207987.5 ;
      RECT  106510.0 206820.0 106580.0 207987.5 ;
      RECT  106880.0 206942.5 106957.5 207077.5 ;
      RECT  107082.5 206942.5 107285.0 207077.5 ;
      RECT  106880.0 207472.5 106957.5 207607.5 ;
      RECT  107215.0 207472.5 107337.5 207607.5 ;
      RECT  106890.0 206942.5 106960.0 207077.5 ;
      RECT  107080.0 206942.5 107150.0 207077.5 ;
      RECT  106890.0 207472.5 106960.0 207607.5 ;
      RECT  107270.0 207472.5 107340.0 207607.5 ;
      RECT  106880.0 206820.0 106950.0 207987.5 ;
      RECT  107215.0 206820.0 107285.0 207987.5 ;
      RECT  17345.0 206820.0 17415.0 207987.5 ;
      RECT  17680.0 206820.0 17750.0 207987.5 ;
      RECT  18050.0 206820.0 18120.0 207987.5 ;
      RECT  18385.0 206820.0 18455.0 207987.5 ;
      RECT  18755.0 206820.0 18825.0 207987.5 ;
      RECT  19090.0 206820.0 19160.0 207987.5 ;
      RECT  19460.0 206820.0 19530.0 207987.5 ;
      RECT  19795.0 206820.0 19865.0 207987.5 ;
      RECT  20165.0 206820.0 20235.0 207987.5 ;
      RECT  20500.0 206820.0 20570.0 207987.5 ;
      RECT  20870.0 206820.0 20940.0 207987.5 ;
      RECT  21205.0 206820.0 21275.0 207987.5 ;
      RECT  21575.0 206820.0 21645.0 207987.5 ;
      RECT  21910.0 206820.0 21980.0 207987.5 ;
      RECT  22280.0 206820.0 22350.0 207987.5 ;
      RECT  22615.0 206820.0 22685.0 207987.5 ;
      RECT  22985.0 206820.0 23055.0 207987.5 ;
      RECT  23320.0 206820.0 23390.0 207987.5 ;
      RECT  23690.0 206820.0 23760.0 207987.5 ;
      RECT  24025.0 206820.0 24095.0 207987.5 ;
      RECT  24395.0 206820.0 24465.0 207987.5 ;
      RECT  24730.0 206820.0 24800.0 207987.5 ;
      RECT  25100.0 206820.0 25170.0 207987.5 ;
      RECT  25435.0 206820.0 25505.0 207987.5 ;
      RECT  25805.0 206820.0 25875.0 207987.5 ;
      RECT  26140.0 206820.0 26210.0 207987.5 ;
      RECT  26510.0 206820.0 26580.0 207987.5 ;
      RECT  26845.0 206820.0 26915.0 207987.5 ;
      RECT  27215.0 206820.0 27285.0 207987.5 ;
      RECT  27550.0 206820.0 27620.0 207987.5 ;
      RECT  27920.0 206820.0 27990.0 207987.5 ;
      RECT  28255.0 206820.0 28325.0 207987.5 ;
      RECT  28625.0 206820.0 28695.0 207987.5 ;
      RECT  28960.0 206820.0 29030.0 207987.5 ;
      RECT  29330.0 206820.0 29400.0 207987.5 ;
      RECT  29665.0 206820.0 29735.0 207987.5 ;
      RECT  30035.0 206820.0 30105.0 207987.5 ;
      RECT  30370.0 206820.0 30440.0 207987.5 ;
      RECT  30740.0 206820.0 30810.0 207987.5 ;
      RECT  31075.0 206820.0 31145.0 207987.5 ;
      RECT  31445.0 206820.0 31515.0 207987.5 ;
      RECT  31780.0 206820.0 31850.0 207987.5 ;
      RECT  32150.0 206820.0 32220.0 207987.5 ;
      RECT  32485.0 206820.0 32555.0 207987.5 ;
      RECT  32855.0 206820.0 32925.0 207987.5 ;
      RECT  33190.0 206820.0 33260.0 207987.5 ;
      RECT  33560.0 206820.0 33630.0 207987.5 ;
      RECT  33895.0 206820.0 33965.0 207987.5 ;
      RECT  34265.0 206820.0 34335.0 207987.5 ;
      RECT  34600.0 206820.0 34670.0 207987.5 ;
      RECT  34970.0 206820.0 35040.0 207987.5 ;
      RECT  35305.0 206820.0 35375.0 207987.5 ;
      RECT  35675.0 206820.0 35745.0 207987.5 ;
      RECT  36010.0 206820.0 36080.0 207987.5 ;
      RECT  36380.0 206820.0 36450.0 207987.5 ;
      RECT  36715.0 206820.0 36785.0 207987.5 ;
      RECT  37085.0 206820.0 37155.0 207987.5 ;
      RECT  37420.0 206820.0 37490.0 207987.5 ;
      RECT  37790.0 206820.0 37860.0 207987.5 ;
      RECT  38125.0 206820.0 38195.0 207987.5 ;
      RECT  38495.0 206820.0 38565.0 207987.5 ;
      RECT  38830.0 206820.0 38900.0 207987.5 ;
      RECT  39200.0 206820.0 39270.0 207987.5 ;
      RECT  39535.0 206820.0 39605.0 207987.5 ;
      RECT  39905.0 206820.0 39975.0 207987.5 ;
      RECT  40240.0 206820.0 40310.0 207987.5 ;
      RECT  40610.0 206820.0 40680.0 207987.5 ;
      RECT  40945.0 206820.0 41015.0 207987.5 ;
      RECT  41315.0 206820.0 41385.0 207987.5 ;
      RECT  41650.0 206820.0 41720.0 207987.5 ;
      RECT  42020.0 206820.0 42090.0 207987.5 ;
      RECT  42355.0 206820.0 42425.0 207987.5 ;
      RECT  42725.0 206820.0 42795.0 207987.5 ;
      RECT  43060.0 206820.0 43130.0 207987.5 ;
      RECT  43430.0 206820.0 43500.0 207987.5 ;
      RECT  43765.0 206820.0 43835.0 207987.5 ;
      RECT  44135.0 206820.0 44205.0 207987.5 ;
      RECT  44470.0 206820.0 44540.0 207987.5 ;
      RECT  44840.0 206820.0 44910.0 207987.5 ;
      RECT  45175.0 206820.0 45245.0 207987.5 ;
      RECT  45545.0 206820.0 45615.0 207987.5 ;
      RECT  45880.0 206820.0 45950.0 207987.5 ;
      RECT  46250.0 206820.0 46320.0 207987.5 ;
      RECT  46585.0 206820.0 46655.0 207987.5 ;
      RECT  46955.0 206820.0 47025.0 207987.5 ;
      RECT  47290.0 206820.0 47360.0 207987.5 ;
      RECT  47660.0 206820.0 47730.0 207987.5 ;
      RECT  47995.0 206820.0 48065.0 207987.5 ;
      RECT  48365.0 206820.0 48435.0 207987.5 ;
      RECT  48700.0 206820.0 48770.0 207987.5 ;
      RECT  49070.0 206820.0 49140.0 207987.5 ;
      RECT  49405.0 206820.0 49475.0 207987.5 ;
      RECT  49775.0 206820.0 49845.0 207987.5 ;
      RECT  50110.0 206820.0 50180.0 207987.5 ;
      RECT  50480.0 206820.0 50550.0 207987.5 ;
      RECT  50815.0 206820.0 50885.0 207987.5 ;
      RECT  51185.0 206820.0 51255.0 207987.5 ;
      RECT  51520.0 206820.0 51590.0 207987.5 ;
      RECT  51890.0 206820.0 51960.0 207987.5 ;
      RECT  52225.0 206820.0 52295.0 207987.5 ;
      RECT  52595.0 206820.0 52665.0 207987.5 ;
      RECT  52930.0 206820.0 53000.0 207987.5 ;
      RECT  53300.0 206820.0 53370.0 207987.5 ;
      RECT  53635.0 206820.0 53705.0 207987.5 ;
      RECT  54005.0 206820.0 54075.0 207987.5 ;
      RECT  54340.0 206820.0 54410.0 207987.5 ;
      RECT  54710.0 206820.0 54780.0 207987.5 ;
      RECT  55045.0 206820.0 55115.0 207987.5 ;
      RECT  55415.0 206820.0 55485.0 207987.5 ;
      RECT  55750.0 206820.0 55820.0 207987.5 ;
      RECT  56120.0 206820.0 56190.0 207987.5 ;
      RECT  56455.0 206820.0 56525.0 207987.5 ;
      RECT  56825.0 206820.0 56895.0 207987.5 ;
      RECT  57160.0 206820.0 57230.0 207987.5 ;
      RECT  57530.0 206820.0 57600.0 207987.5 ;
      RECT  57865.0 206820.0 57935.0 207987.5 ;
      RECT  58235.0 206820.0 58305.0 207987.5 ;
      RECT  58570.0 206820.0 58640.0 207987.5 ;
      RECT  58940.0 206820.0 59010.0 207987.5 ;
      RECT  59275.0 206820.0 59345.0 207987.5 ;
      RECT  59645.0 206820.0 59715.0 207987.5 ;
      RECT  59980.0 206820.0 60050.0 207987.5 ;
      RECT  60350.0 206820.0 60420.0 207987.5 ;
      RECT  60685.0 206820.0 60755.0 207987.5 ;
      RECT  61055.0 206820.0 61125.0 207987.5 ;
      RECT  61390.0 206820.0 61460.0 207987.5 ;
      RECT  61760.0 206820.0 61830.0 207987.5 ;
      RECT  62095.0 206820.0 62165.0 207987.5 ;
      RECT  62465.0 206820.0 62535.0 207987.5 ;
      RECT  62800.0 206820.0 62870.0 207987.5 ;
      RECT  63170.0 206820.0 63240.0 207987.5 ;
      RECT  63505.0 206820.0 63575.0 207987.5 ;
      RECT  63875.0 206820.0 63945.0 207987.5 ;
      RECT  64210.0 206820.0 64280.0 207987.5 ;
      RECT  64580.0 206820.0 64650.0 207987.5 ;
      RECT  64915.0 206820.0 64985.0 207987.5 ;
      RECT  65285.0 206820.0 65355.0 207987.5 ;
      RECT  65620.0 206820.0 65690.0 207987.5 ;
      RECT  65990.0 206820.0 66060.0 207987.5 ;
      RECT  66325.0 206820.0 66395.0 207987.5 ;
      RECT  66695.0 206820.0 66765.0 207987.5 ;
      RECT  67030.0 206820.0 67100.0 207987.5 ;
      RECT  67400.0 206820.0 67470.0 207987.5 ;
      RECT  67735.0 206820.0 67805.0 207987.5 ;
      RECT  68105.0 206820.0 68175.0 207987.5 ;
      RECT  68440.0 206820.0 68510.0 207987.5 ;
      RECT  68810.0 206820.0 68880.0 207987.5 ;
      RECT  69145.0 206820.0 69215.0 207987.5 ;
      RECT  69515.0 206820.0 69585.0 207987.5 ;
      RECT  69850.0 206820.0 69920.0 207987.5 ;
      RECT  70220.0 206820.0 70290.0 207987.5 ;
      RECT  70555.0 206820.0 70625.0 207987.5 ;
      RECT  70925.0 206820.0 70995.0 207987.5 ;
      RECT  71260.0 206820.0 71330.0 207987.5 ;
      RECT  71630.0 206820.0 71700.0 207987.5 ;
      RECT  71965.0 206820.0 72035.0 207987.5 ;
      RECT  72335.0 206820.0 72405.0 207987.5 ;
      RECT  72670.0 206820.0 72740.0 207987.5 ;
      RECT  73040.0 206820.0 73110.0 207987.5 ;
      RECT  73375.0 206820.0 73445.0 207987.5 ;
      RECT  73745.0 206820.0 73815.0 207987.5 ;
      RECT  74080.0 206820.0 74150.0 207987.5 ;
      RECT  74450.0 206820.0 74520.0 207987.5 ;
      RECT  74785.0 206820.0 74855.0 207987.5 ;
      RECT  75155.0 206820.0 75225.0 207987.5 ;
      RECT  75490.0 206820.0 75560.0 207987.5 ;
      RECT  75860.0 206820.0 75930.0 207987.5 ;
      RECT  76195.0 206820.0 76265.0 207987.5 ;
      RECT  76565.0 206820.0 76635.0 207987.5 ;
      RECT  76900.0 206820.0 76970.0 207987.5 ;
      RECT  77270.0 206820.0 77340.0 207987.5 ;
      RECT  77605.0 206820.0 77675.0 207987.5 ;
      RECT  77975.0 206820.0 78045.0 207987.5 ;
      RECT  78310.0 206820.0 78380.0 207987.5 ;
      RECT  78680.0 206820.0 78750.0 207987.5 ;
      RECT  79015.0 206820.0 79085.0 207987.5 ;
      RECT  79385.0 206820.0 79455.0 207987.5 ;
      RECT  79720.0 206820.0 79790.0 207987.5 ;
      RECT  80090.0 206820.0 80160.0 207987.5 ;
      RECT  80425.0 206820.0 80495.0 207987.5 ;
      RECT  80795.0 206820.0 80865.0 207987.5 ;
      RECT  81130.0 206820.0 81200.0 207987.5 ;
      RECT  81500.0 206820.0 81570.0 207987.5 ;
      RECT  81835.0 206820.0 81905.0 207987.5 ;
      RECT  82205.0 206820.0 82275.0 207987.5 ;
      RECT  82540.0 206820.0 82610.0 207987.5 ;
      RECT  82910.0 206820.0 82980.0 207987.5 ;
      RECT  83245.0 206820.0 83315.0 207987.5 ;
      RECT  83615.0 206820.0 83685.0 207987.5 ;
      RECT  83950.0 206820.0 84020.0 207987.5 ;
      RECT  84320.0 206820.0 84390.0 207987.5 ;
      RECT  84655.0 206820.0 84725.0 207987.5 ;
      RECT  85025.0 206820.0 85095.0 207987.5 ;
      RECT  85360.0 206820.0 85430.0 207987.5 ;
      RECT  85730.0 206820.0 85800.0 207987.5 ;
      RECT  86065.0 206820.0 86135.0 207987.5 ;
      RECT  86435.0 206820.0 86505.0 207987.5 ;
      RECT  86770.0 206820.0 86840.0 207987.5 ;
      RECT  87140.0 206820.0 87210.0 207987.5 ;
      RECT  87475.0 206820.0 87545.0 207987.5 ;
      RECT  87845.0 206820.0 87915.0 207987.5 ;
      RECT  88180.0 206820.0 88250.0 207987.5 ;
      RECT  88550.0 206820.0 88620.0 207987.5 ;
      RECT  88885.0 206820.0 88955.0 207987.5 ;
      RECT  89255.0 206820.0 89325.0 207987.5 ;
      RECT  89590.0 206820.0 89660.0 207987.5 ;
      RECT  89960.0 206820.0 90030.0 207987.5 ;
      RECT  90295.0 206820.0 90365.0 207987.5 ;
      RECT  90665.0 206820.0 90735.0 207987.5 ;
      RECT  91000.0 206820.0 91070.0 207987.5 ;
      RECT  91370.0 206820.0 91440.0 207987.5 ;
      RECT  91705.0 206820.0 91775.0 207987.5 ;
      RECT  92075.0 206820.0 92145.0 207987.5 ;
      RECT  92410.0 206820.0 92480.0 207987.5 ;
      RECT  92780.0 206820.0 92850.0 207987.5 ;
      RECT  93115.0 206820.0 93185.0 207987.5 ;
      RECT  93485.0 206820.0 93555.0 207987.5 ;
      RECT  93820.0 206820.0 93890.0 207987.5 ;
      RECT  94190.0 206820.0 94260.0 207987.5 ;
      RECT  94525.0 206820.0 94595.0 207987.5 ;
      RECT  94895.0 206820.0 94965.0 207987.5 ;
      RECT  95230.0 206820.0 95300.0 207987.5 ;
      RECT  95600.0 206820.0 95670.0 207987.5 ;
      RECT  95935.0 206820.0 96005.0 207987.5 ;
      RECT  96305.0 206820.0 96375.0 207987.5 ;
      RECT  96640.0 206820.0 96710.0 207987.5 ;
      RECT  97010.0 206820.0 97080.0 207987.5 ;
      RECT  97345.0 206820.0 97415.0 207987.5 ;
      RECT  97715.0 206820.0 97785.0 207987.5 ;
      RECT  98050.0 206820.0 98120.0 207987.5 ;
      RECT  98420.0 206820.0 98490.0 207987.5 ;
      RECT  98755.0 206820.0 98825.0 207987.5 ;
      RECT  99125.0 206820.0 99195.0 207987.5 ;
      RECT  99460.0 206820.0 99530.0 207987.5 ;
      RECT  99830.0 206820.0 99900.0 207987.5 ;
      RECT  100165.0 206820.0 100235.0 207987.5 ;
      RECT  100535.0 206820.0 100605.0 207987.5 ;
      RECT  100870.0 206820.0 100940.0 207987.5 ;
      RECT  101240.0 206820.0 101310.0 207987.5 ;
      RECT  101575.0 206820.0 101645.0 207987.5 ;
      RECT  101945.0 206820.0 102015.0 207987.5 ;
      RECT  102280.0 206820.0 102350.0 207987.5 ;
      RECT  102650.0 206820.0 102720.0 207987.5 ;
      RECT  102985.0 206820.0 103055.0 207987.5 ;
      RECT  103355.0 206820.0 103425.0 207987.5 ;
      RECT  103690.0 206820.0 103760.0 207987.5 ;
      RECT  104060.0 206820.0 104130.0 207987.5 ;
      RECT  104395.0 206820.0 104465.0 207987.5 ;
      RECT  104765.0 206820.0 104835.0 207987.5 ;
      RECT  105100.0 206820.0 105170.0 207987.5 ;
      RECT  105470.0 206820.0 105540.0 207987.5 ;
      RECT  105805.0 206820.0 105875.0 207987.5 ;
      RECT  106175.0 206820.0 106245.0 207987.5 ;
      RECT  106510.0 206820.0 106580.0 207987.5 ;
      RECT  106880.0 206820.0 106950.0 207987.5 ;
      RECT  107215.0 206820.0 107285.0 207987.5 ;
      RECT  18050.0 31535.0 18120.0 32235.0 ;
      RECT  18385.0 31395.0 18455.0 32235.0 ;
      RECT  18755.0 31535.0 18825.0 32235.0 ;
      RECT  19090.0 31395.0 19160.0 32235.0 ;
      RECT  19460.0 31535.0 19530.0 32235.0 ;
      RECT  19795.0 31395.0 19865.0 32235.0 ;
      RECT  20870.0 31535.0 20940.0 32235.0 ;
      RECT  21205.0 31395.0 21275.0 32235.0 ;
      RECT  21575.0 31535.0 21645.0 32235.0 ;
      RECT  21910.0 31395.0 21980.0 32235.0 ;
      RECT  22280.0 31535.0 22350.0 32235.0 ;
      RECT  22615.0 31395.0 22685.0 32235.0 ;
      RECT  23690.0 31535.0 23760.0 32235.0 ;
      RECT  24025.0 31395.0 24095.0 32235.0 ;
      RECT  24395.0 31535.0 24465.0 32235.0 ;
      RECT  24730.0 31395.0 24800.0 32235.0 ;
      RECT  25100.0 31535.0 25170.0 32235.0 ;
      RECT  25435.0 31395.0 25505.0 32235.0 ;
      RECT  26510.0 31535.0 26580.0 32235.0 ;
      RECT  26845.0 31395.0 26915.0 32235.0 ;
      RECT  27215.0 31535.0 27285.0 32235.0 ;
      RECT  27550.0 31395.0 27620.0 32235.0 ;
      RECT  27920.0 31535.0 27990.0 32235.0 ;
      RECT  28255.0 31395.0 28325.0 32235.0 ;
      RECT  29330.0 31535.0 29400.0 32235.0 ;
      RECT  29665.0 31395.0 29735.0 32235.0 ;
      RECT  30035.0 31535.0 30105.0 32235.0 ;
      RECT  30370.0 31395.0 30440.0 32235.0 ;
      RECT  30740.0 31535.0 30810.0 32235.0 ;
      RECT  31075.0 31395.0 31145.0 32235.0 ;
      RECT  32150.0 31535.0 32220.0 32235.0 ;
      RECT  32485.0 31395.0 32555.0 32235.0 ;
      RECT  32855.0 31535.0 32925.0 32235.0 ;
      RECT  33190.0 31395.0 33260.0 32235.0 ;
      RECT  33560.0 31535.0 33630.0 32235.0 ;
      RECT  33895.0 31395.0 33965.0 32235.0 ;
      RECT  34970.0 31535.0 35040.0 32235.0 ;
      RECT  35305.0 31395.0 35375.0 32235.0 ;
      RECT  35675.0 31535.0 35745.0 32235.0 ;
      RECT  36010.0 31395.0 36080.0 32235.0 ;
      RECT  36380.0 31535.0 36450.0 32235.0 ;
      RECT  36715.0 31395.0 36785.0 32235.0 ;
      RECT  37790.0 31535.0 37860.0 32235.0 ;
      RECT  38125.0 31395.0 38195.0 32235.0 ;
      RECT  38495.0 31535.0 38565.0 32235.0 ;
      RECT  38830.0 31395.0 38900.0 32235.0 ;
      RECT  39200.0 31535.0 39270.0 32235.0 ;
      RECT  39535.0 31395.0 39605.0 32235.0 ;
      RECT  40610.0 31535.0 40680.0 32235.0 ;
      RECT  40945.0 31395.0 41015.0 32235.0 ;
      RECT  41315.0 31535.0 41385.0 32235.0 ;
      RECT  41650.0 31395.0 41720.0 32235.0 ;
      RECT  42020.0 31535.0 42090.0 32235.0 ;
      RECT  42355.0 31395.0 42425.0 32235.0 ;
      RECT  43430.0 31535.0 43500.0 32235.0 ;
      RECT  43765.0 31395.0 43835.0 32235.0 ;
      RECT  44135.0 31535.0 44205.0 32235.0 ;
      RECT  44470.0 31395.0 44540.0 32235.0 ;
      RECT  44840.0 31535.0 44910.0 32235.0 ;
      RECT  45175.0 31395.0 45245.0 32235.0 ;
      RECT  46250.0 31535.0 46320.0 32235.0 ;
      RECT  46585.0 31395.0 46655.0 32235.0 ;
      RECT  46955.0 31535.0 47025.0 32235.0 ;
      RECT  47290.0 31395.0 47360.0 32235.0 ;
      RECT  47660.0 31535.0 47730.0 32235.0 ;
      RECT  47995.0 31395.0 48065.0 32235.0 ;
      RECT  49070.0 31535.0 49140.0 32235.0 ;
      RECT  49405.0 31395.0 49475.0 32235.0 ;
      RECT  49775.0 31535.0 49845.0 32235.0 ;
      RECT  50110.0 31395.0 50180.0 32235.0 ;
      RECT  50480.0 31535.0 50550.0 32235.0 ;
      RECT  50815.0 31395.0 50885.0 32235.0 ;
      RECT  51890.0 31535.0 51960.0 32235.0 ;
      RECT  52225.0 31395.0 52295.0 32235.0 ;
      RECT  52595.0 31535.0 52665.0 32235.0 ;
      RECT  52930.0 31395.0 53000.0 32235.0 ;
      RECT  53300.0 31535.0 53370.0 32235.0 ;
      RECT  53635.0 31395.0 53705.0 32235.0 ;
      RECT  54710.0 31535.0 54780.0 32235.0 ;
      RECT  55045.0 31395.0 55115.0 32235.0 ;
      RECT  55415.0 31535.0 55485.0 32235.0 ;
      RECT  55750.0 31395.0 55820.0 32235.0 ;
      RECT  56120.0 31535.0 56190.0 32235.0 ;
      RECT  56455.0 31395.0 56525.0 32235.0 ;
      RECT  57530.0 31535.0 57600.0 32235.0 ;
      RECT  57865.0 31395.0 57935.0 32235.0 ;
      RECT  58235.0 31535.0 58305.0 32235.0 ;
      RECT  58570.0 31395.0 58640.0 32235.0 ;
      RECT  58940.0 31535.0 59010.0 32235.0 ;
      RECT  59275.0 31395.0 59345.0 32235.0 ;
      RECT  60350.0 31535.0 60420.0 32235.0 ;
      RECT  60685.0 31395.0 60755.0 32235.0 ;
      RECT  61055.0 31535.0 61125.0 32235.0 ;
      RECT  61390.0 31395.0 61460.0 32235.0 ;
      RECT  61760.0 31535.0 61830.0 32235.0 ;
      RECT  62095.0 31395.0 62165.0 32235.0 ;
      RECT  63170.0 31535.0 63240.0 32235.0 ;
      RECT  63505.0 31395.0 63575.0 32235.0 ;
      RECT  63875.0 31535.0 63945.0 32235.0 ;
      RECT  64210.0 31395.0 64280.0 32235.0 ;
      RECT  64580.0 31535.0 64650.0 32235.0 ;
      RECT  64915.0 31395.0 64985.0 32235.0 ;
      RECT  65990.0 31535.0 66060.0 32235.0 ;
      RECT  66325.0 31395.0 66395.0 32235.0 ;
      RECT  66695.0 31535.0 66765.0 32235.0 ;
      RECT  67030.0 31395.0 67100.0 32235.0 ;
      RECT  67400.0 31535.0 67470.0 32235.0 ;
      RECT  67735.0 31395.0 67805.0 32235.0 ;
      RECT  68810.0 31535.0 68880.0 32235.0 ;
      RECT  69145.0 31395.0 69215.0 32235.0 ;
      RECT  69515.0 31535.0 69585.0 32235.0 ;
      RECT  69850.0 31395.0 69920.0 32235.0 ;
      RECT  70220.0 31535.0 70290.0 32235.0 ;
      RECT  70555.0 31395.0 70625.0 32235.0 ;
      RECT  71630.0 31535.0 71700.0 32235.0 ;
      RECT  71965.0 31395.0 72035.0 32235.0 ;
      RECT  72335.0 31535.0 72405.0 32235.0 ;
      RECT  72670.0 31395.0 72740.0 32235.0 ;
      RECT  73040.0 31535.0 73110.0 32235.0 ;
      RECT  73375.0 31395.0 73445.0 32235.0 ;
      RECT  74450.0 31535.0 74520.0 32235.0 ;
      RECT  74785.0 31395.0 74855.0 32235.0 ;
      RECT  75155.0 31535.0 75225.0 32235.0 ;
      RECT  75490.0 31395.0 75560.0 32235.0 ;
      RECT  75860.0 31535.0 75930.0 32235.0 ;
      RECT  76195.0 31395.0 76265.0 32235.0 ;
      RECT  77270.0 31535.0 77340.0 32235.0 ;
      RECT  77605.0 31395.0 77675.0 32235.0 ;
      RECT  77975.0 31535.0 78045.0 32235.0 ;
      RECT  78310.0 31395.0 78380.0 32235.0 ;
      RECT  78680.0 31535.0 78750.0 32235.0 ;
      RECT  79015.0 31395.0 79085.0 32235.0 ;
      RECT  80090.0 31535.0 80160.0 32235.0 ;
      RECT  80425.0 31395.0 80495.0 32235.0 ;
      RECT  80795.0 31535.0 80865.0 32235.0 ;
      RECT  81130.0 31395.0 81200.0 32235.0 ;
      RECT  81500.0 31535.0 81570.0 32235.0 ;
      RECT  81835.0 31395.0 81905.0 32235.0 ;
      RECT  82910.0 31535.0 82980.0 32235.0 ;
      RECT  83245.0 31395.0 83315.0 32235.0 ;
      RECT  83615.0 31535.0 83685.0 32235.0 ;
      RECT  83950.0 31395.0 84020.0 32235.0 ;
      RECT  84320.0 31535.0 84390.0 32235.0 ;
      RECT  84655.0 31395.0 84725.0 32235.0 ;
      RECT  85730.0 31535.0 85800.0 32235.0 ;
      RECT  86065.0 31395.0 86135.0 32235.0 ;
      RECT  86435.0 31535.0 86505.0 32235.0 ;
      RECT  86770.0 31395.0 86840.0 32235.0 ;
      RECT  87140.0 31535.0 87210.0 32235.0 ;
      RECT  87475.0 31395.0 87545.0 32235.0 ;
      RECT  88550.0 31535.0 88620.0 32235.0 ;
      RECT  88885.0 31395.0 88955.0 32235.0 ;
      RECT  89255.0 31535.0 89325.0 32235.0 ;
      RECT  89590.0 31395.0 89660.0 32235.0 ;
      RECT  89960.0 31535.0 90030.0 32235.0 ;
      RECT  90295.0 31395.0 90365.0 32235.0 ;
      RECT  91370.0 31535.0 91440.0 32235.0 ;
      RECT  91705.0 31395.0 91775.0 32235.0 ;
      RECT  92075.0 31535.0 92145.0 32235.0 ;
      RECT  92410.0 31395.0 92480.0 32235.0 ;
      RECT  92780.0 31535.0 92850.0 32235.0 ;
      RECT  93115.0 31395.0 93185.0 32235.0 ;
      RECT  94190.0 31535.0 94260.0 32235.0 ;
      RECT  94525.0 31395.0 94595.0 32235.0 ;
      RECT  94895.0 31535.0 94965.0 32235.0 ;
      RECT  95230.0 31395.0 95300.0 32235.0 ;
      RECT  95600.0 31535.0 95670.0 32235.0 ;
      RECT  95935.0 31395.0 96005.0 32235.0 ;
      RECT  97010.0 31535.0 97080.0 32235.0 ;
      RECT  97345.0 31395.0 97415.0 32235.0 ;
      RECT  97715.0 31535.0 97785.0 32235.0 ;
      RECT  98050.0 31395.0 98120.0 32235.0 ;
      RECT  98420.0 31535.0 98490.0 32235.0 ;
      RECT  98755.0 31395.0 98825.0 32235.0 ;
      RECT  99830.0 31535.0 99900.0 32235.0 ;
      RECT  100165.0 31395.0 100235.0 32235.0 ;
      RECT  100535.0 31535.0 100605.0 32235.0 ;
      RECT  100870.0 31395.0 100940.0 32235.0 ;
      RECT  101240.0 31535.0 101310.0 32235.0 ;
      RECT  101575.0 31395.0 101645.0 32235.0 ;
      RECT  102650.0 31535.0 102720.0 32235.0 ;
      RECT  102985.0 31395.0 103055.0 32235.0 ;
      RECT  103355.0 31535.0 103425.0 32235.0 ;
      RECT  103690.0 31395.0 103760.0 32235.0 ;
      RECT  104060.0 31535.0 104130.0 32235.0 ;
      RECT  104395.0 31395.0 104465.0 32235.0 ;
      RECT  105470.0 31535.0 105540.0 32235.0 ;
      RECT  105805.0 31395.0 105875.0 32235.0 ;
      RECT  106175.0 31535.0 106245.0 32235.0 ;
      RECT  106510.0 31395.0 106580.0 32235.0 ;
      RECT  106880.0 31535.0 106950.0 32235.0 ;
      RECT  107215.0 31395.0 107285.0 32235.0 ;
      RECT  17345.0 32875.0 17415.0 32945.0 ;
      RECT  17417.5 32875.0 17487.5 32945.0 ;
      RECT  17345.0 32375.0 17415.0 32910.0 ;
      RECT  17380.0 32875.0 17452.5 32945.0 ;
      RECT  17417.5 32910.0 17487.5 33442.5 ;
      RECT  17680.0 33287.5 17750.0 33357.5 ;
      RECT  17607.5 33287.5 17677.5 33357.5 ;
      RECT  17680.0 33322.5 17750.0 33925.0 ;
      RECT  17642.5 33287.5 17715.0 33357.5 ;
      RECT  17607.5 32717.5 17677.5 33322.5 ;
      RECT  17345.0 33857.5 17415.0 33992.5 ;
      RECT  17680.0 32307.5 17750.0 32442.5 ;
      RECT  17417.5 33442.5 17487.5 33577.5 ;
      RECT  17607.5 32582.5 17677.5 32717.5 ;
      RECT  17865.0 32482.5 17935.0 32617.5 ;
      RECT  17345.0 33925.0 17415.0 34065.0 ;
      RECT  17680.0 33925.0 17750.0 34065.0 ;
      RECT  17345.0 32235.0 17415.0 32375.0 ;
      RECT  17680.0 32235.0 17750.0 32375.0 ;
      RECT  17160.0 32235.0 17230.0 34065.0 ;
      RECT  17865.0 32235.0 17935.0 34065.0 ;
      RECT  18050.0 32875.0 18120.0 32945.0 ;
      RECT  18122.5 32875.0 18192.5 32945.0 ;
      RECT  18050.0 32375.0 18120.0 32910.0 ;
      RECT  18085.0 32875.0 18157.5 32945.0 ;
      RECT  18122.5 32910.0 18192.5 33442.5 ;
      RECT  18385.0 33287.5 18455.0 33357.5 ;
      RECT  18312.5 33287.5 18382.5 33357.5 ;
      RECT  18385.0 33322.5 18455.0 33925.0 ;
      RECT  18347.5 33287.5 18420.0 33357.5 ;
      RECT  18312.5 32717.5 18382.5 33322.5 ;
      RECT  18050.0 33857.5 18120.0 33992.5 ;
      RECT  18385.0 32307.5 18455.0 32442.5 ;
      RECT  18122.5 33442.5 18192.5 33577.5 ;
      RECT  18312.5 32582.5 18382.5 32717.5 ;
      RECT  18570.0 32482.5 18640.0 32617.5 ;
      RECT  18050.0 33925.0 18120.0 34065.0 ;
      RECT  18385.0 33925.0 18455.0 34065.0 ;
      RECT  18050.0 32235.0 18120.0 32375.0 ;
      RECT  18385.0 32235.0 18455.0 32375.0 ;
      RECT  17865.0 32235.0 17935.0 34065.0 ;
      RECT  18570.0 32235.0 18640.0 34065.0 ;
      RECT  18755.0 32875.0 18825.0 32945.0 ;
      RECT  18827.5 32875.0 18897.5 32945.0 ;
      RECT  18755.0 32375.0 18825.0 32910.0 ;
      RECT  18790.0 32875.0 18862.5 32945.0 ;
      RECT  18827.5 32910.0 18897.5 33442.5 ;
      RECT  19090.0 33287.5 19160.0 33357.5 ;
      RECT  19017.5 33287.5 19087.5 33357.5 ;
      RECT  19090.0 33322.5 19160.0 33925.0 ;
      RECT  19052.5 33287.5 19125.0 33357.5 ;
      RECT  19017.5 32717.5 19087.5 33322.5 ;
      RECT  18755.0 33857.5 18825.0 33992.5 ;
      RECT  19090.0 32307.5 19160.0 32442.5 ;
      RECT  18827.5 33442.5 18897.5 33577.5 ;
      RECT  19017.5 32582.5 19087.5 32717.5 ;
      RECT  19275.0 32482.5 19345.0 32617.5 ;
      RECT  18755.0 33925.0 18825.0 34065.0 ;
      RECT  19090.0 33925.0 19160.0 34065.0 ;
      RECT  18755.0 32235.0 18825.0 32375.0 ;
      RECT  19090.0 32235.0 19160.0 32375.0 ;
      RECT  18570.0 32235.0 18640.0 34065.0 ;
      RECT  19275.0 32235.0 19345.0 34065.0 ;
      RECT  19460.0 32875.0 19530.0 32945.0 ;
      RECT  19532.5 32875.0 19602.5 32945.0 ;
      RECT  19460.0 32375.0 19530.0 32910.0 ;
      RECT  19495.0 32875.0 19567.5 32945.0 ;
      RECT  19532.5 32910.0 19602.5 33442.5 ;
      RECT  19795.0 33287.5 19865.0 33357.5 ;
      RECT  19722.5 33287.5 19792.5 33357.5 ;
      RECT  19795.0 33322.5 19865.0 33925.0 ;
      RECT  19757.5 33287.5 19830.0 33357.5 ;
      RECT  19722.5 32717.5 19792.5 33322.5 ;
      RECT  19460.0 33857.5 19530.0 33992.5 ;
      RECT  19795.0 32307.5 19865.0 32442.5 ;
      RECT  19532.5 33442.5 19602.5 33577.5 ;
      RECT  19722.5 32582.5 19792.5 32717.5 ;
      RECT  19980.0 32482.5 20050.0 32617.5 ;
      RECT  19460.0 33925.0 19530.0 34065.0 ;
      RECT  19795.0 33925.0 19865.0 34065.0 ;
      RECT  19460.0 32235.0 19530.0 32375.0 ;
      RECT  19795.0 32235.0 19865.0 32375.0 ;
      RECT  19275.0 32235.0 19345.0 34065.0 ;
      RECT  19980.0 32235.0 20050.0 34065.0 ;
      RECT  20165.0 32875.0 20235.0 32945.0 ;
      RECT  20237.5 32875.0 20307.5 32945.0 ;
      RECT  20165.0 32375.0 20235.0 32910.0 ;
      RECT  20200.0 32875.0 20272.5 32945.0 ;
      RECT  20237.5 32910.0 20307.5 33442.5 ;
      RECT  20500.0 33287.5 20570.0 33357.5 ;
      RECT  20427.5 33287.5 20497.5 33357.5 ;
      RECT  20500.0 33322.5 20570.0 33925.0 ;
      RECT  20462.5 33287.5 20535.0 33357.5 ;
      RECT  20427.5 32717.5 20497.5 33322.5 ;
      RECT  20165.0 33857.5 20235.0 33992.5 ;
      RECT  20500.0 32307.5 20570.0 32442.5 ;
      RECT  20237.5 33442.5 20307.5 33577.5 ;
      RECT  20427.5 32582.5 20497.5 32717.5 ;
      RECT  20685.0 32482.5 20755.0 32617.5 ;
      RECT  20165.0 33925.0 20235.0 34065.0 ;
      RECT  20500.0 33925.0 20570.0 34065.0 ;
      RECT  20165.0 32235.0 20235.0 32375.0 ;
      RECT  20500.0 32235.0 20570.0 32375.0 ;
      RECT  19980.0 32235.0 20050.0 34065.0 ;
      RECT  20685.0 32235.0 20755.0 34065.0 ;
      RECT  20870.0 32875.0 20940.0 32945.0 ;
      RECT  20942.5 32875.0 21012.5 32945.0 ;
      RECT  20870.0 32375.0 20940.0 32910.0 ;
      RECT  20905.0 32875.0 20977.5 32945.0 ;
      RECT  20942.5 32910.0 21012.5 33442.5 ;
      RECT  21205.0 33287.5 21275.0 33357.5 ;
      RECT  21132.5 33287.5 21202.5 33357.5 ;
      RECT  21205.0 33322.5 21275.0 33925.0 ;
      RECT  21167.5 33287.5 21240.0 33357.5 ;
      RECT  21132.5 32717.5 21202.5 33322.5 ;
      RECT  20870.0 33857.5 20940.0 33992.5 ;
      RECT  21205.0 32307.5 21275.0 32442.5 ;
      RECT  20942.5 33442.5 21012.5 33577.5 ;
      RECT  21132.5 32582.5 21202.5 32717.5 ;
      RECT  21390.0 32482.5 21460.0 32617.5 ;
      RECT  20870.0 33925.0 20940.0 34065.0 ;
      RECT  21205.0 33925.0 21275.0 34065.0 ;
      RECT  20870.0 32235.0 20940.0 32375.0 ;
      RECT  21205.0 32235.0 21275.0 32375.0 ;
      RECT  20685.0 32235.0 20755.0 34065.0 ;
      RECT  21390.0 32235.0 21460.0 34065.0 ;
      RECT  21575.0 32875.0 21645.0 32945.0 ;
      RECT  21647.5 32875.0 21717.5 32945.0 ;
      RECT  21575.0 32375.0 21645.0 32910.0 ;
      RECT  21610.0 32875.0 21682.5 32945.0 ;
      RECT  21647.5 32910.0 21717.5 33442.5 ;
      RECT  21910.0 33287.5 21980.0 33357.5 ;
      RECT  21837.5 33287.5 21907.5 33357.5 ;
      RECT  21910.0 33322.5 21980.0 33925.0 ;
      RECT  21872.5 33287.5 21945.0 33357.5 ;
      RECT  21837.5 32717.5 21907.5 33322.5 ;
      RECT  21575.0 33857.5 21645.0 33992.5 ;
      RECT  21910.0 32307.5 21980.0 32442.5 ;
      RECT  21647.5 33442.5 21717.5 33577.5 ;
      RECT  21837.5 32582.5 21907.5 32717.5 ;
      RECT  22095.0 32482.5 22165.0 32617.5 ;
      RECT  21575.0 33925.0 21645.0 34065.0 ;
      RECT  21910.0 33925.0 21980.0 34065.0 ;
      RECT  21575.0 32235.0 21645.0 32375.0 ;
      RECT  21910.0 32235.0 21980.0 32375.0 ;
      RECT  21390.0 32235.0 21460.0 34065.0 ;
      RECT  22095.0 32235.0 22165.0 34065.0 ;
      RECT  22280.0 32875.0 22350.0 32945.0 ;
      RECT  22352.5 32875.0 22422.5 32945.0 ;
      RECT  22280.0 32375.0 22350.0 32910.0 ;
      RECT  22315.0 32875.0 22387.5 32945.0 ;
      RECT  22352.5 32910.0 22422.5 33442.5 ;
      RECT  22615.0 33287.5 22685.0 33357.5 ;
      RECT  22542.5 33287.5 22612.5 33357.5 ;
      RECT  22615.0 33322.5 22685.0 33925.0 ;
      RECT  22577.5 33287.5 22650.0 33357.5 ;
      RECT  22542.5 32717.5 22612.5 33322.5 ;
      RECT  22280.0 33857.5 22350.0 33992.5 ;
      RECT  22615.0 32307.5 22685.0 32442.5 ;
      RECT  22352.5 33442.5 22422.5 33577.5 ;
      RECT  22542.5 32582.5 22612.5 32717.5 ;
      RECT  22800.0 32482.5 22870.0 32617.5 ;
      RECT  22280.0 33925.0 22350.0 34065.0 ;
      RECT  22615.0 33925.0 22685.0 34065.0 ;
      RECT  22280.0 32235.0 22350.0 32375.0 ;
      RECT  22615.0 32235.0 22685.0 32375.0 ;
      RECT  22095.0 32235.0 22165.0 34065.0 ;
      RECT  22800.0 32235.0 22870.0 34065.0 ;
      RECT  22985.0 32875.0 23055.0 32945.0 ;
      RECT  23057.5 32875.0 23127.5 32945.0 ;
      RECT  22985.0 32375.0 23055.0 32910.0 ;
      RECT  23020.0 32875.0 23092.5 32945.0 ;
      RECT  23057.5 32910.0 23127.5 33442.5 ;
      RECT  23320.0 33287.5 23390.0 33357.5 ;
      RECT  23247.5 33287.5 23317.5 33357.5 ;
      RECT  23320.0 33322.5 23390.0 33925.0 ;
      RECT  23282.5 33287.5 23355.0 33357.5 ;
      RECT  23247.5 32717.5 23317.5 33322.5 ;
      RECT  22985.0 33857.5 23055.0 33992.5 ;
      RECT  23320.0 32307.5 23390.0 32442.5 ;
      RECT  23057.5 33442.5 23127.5 33577.5 ;
      RECT  23247.5 32582.5 23317.5 32717.5 ;
      RECT  23505.0 32482.5 23575.0 32617.5 ;
      RECT  22985.0 33925.0 23055.0 34065.0 ;
      RECT  23320.0 33925.0 23390.0 34065.0 ;
      RECT  22985.0 32235.0 23055.0 32375.0 ;
      RECT  23320.0 32235.0 23390.0 32375.0 ;
      RECT  22800.0 32235.0 22870.0 34065.0 ;
      RECT  23505.0 32235.0 23575.0 34065.0 ;
      RECT  23690.0 32875.0 23760.0 32945.0 ;
      RECT  23762.5 32875.0 23832.5 32945.0 ;
      RECT  23690.0 32375.0 23760.0 32910.0 ;
      RECT  23725.0 32875.0 23797.5 32945.0 ;
      RECT  23762.5 32910.0 23832.5 33442.5 ;
      RECT  24025.0 33287.5 24095.0 33357.5 ;
      RECT  23952.5 33287.5 24022.5 33357.5 ;
      RECT  24025.0 33322.5 24095.0 33925.0 ;
      RECT  23987.5 33287.5 24060.0 33357.5 ;
      RECT  23952.5 32717.5 24022.5 33322.5 ;
      RECT  23690.0 33857.5 23760.0 33992.5 ;
      RECT  24025.0 32307.5 24095.0 32442.5 ;
      RECT  23762.5 33442.5 23832.5 33577.5 ;
      RECT  23952.5 32582.5 24022.5 32717.5 ;
      RECT  24210.0 32482.5 24280.0 32617.5 ;
      RECT  23690.0 33925.0 23760.0 34065.0 ;
      RECT  24025.0 33925.0 24095.0 34065.0 ;
      RECT  23690.0 32235.0 23760.0 32375.0 ;
      RECT  24025.0 32235.0 24095.0 32375.0 ;
      RECT  23505.0 32235.0 23575.0 34065.0 ;
      RECT  24210.0 32235.0 24280.0 34065.0 ;
      RECT  24395.0 32875.0 24465.0 32945.0 ;
      RECT  24467.5 32875.0 24537.5 32945.0 ;
      RECT  24395.0 32375.0 24465.0 32910.0 ;
      RECT  24430.0 32875.0 24502.5 32945.0 ;
      RECT  24467.5 32910.0 24537.5 33442.5 ;
      RECT  24730.0 33287.5 24800.0 33357.5 ;
      RECT  24657.5 33287.5 24727.5 33357.5 ;
      RECT  24730.0 33322.5 24800.0 33925.0 ;
      RECT  24692.5 33287.5 24765.0 33357.5 ;
      RECT  24657.5 32717.5 24727.5 33322.5 ;
      RECT  24395.0 33857.5 24465.0 33992.5 ;
      RECT  24730.0 32307.5 24800.0 32442.5 ;
      RECT  24467.5 33442.5 24537.5 33577.5 ;
      RECT  24657.5 32582.5 24727.5 32717.5 ;
      RECT  24915.0 32482.5 24985.0 32617.5 ;
      RECT  24395.0 33925.0 24465.0 34065.0 ;
      RECT  24730.0 33925.0 24800.0 34065.0 ;
      RECT  24395.0 32235.0 24465.0 32375.0 ;
      RECT  24730.0 32235.0 24800.0 32375.0 ;
      RECT  24210.0 32235.0 24280.0 34065.0 ;
      RECT  24915.0 32235.0 24985.0 34065.0 ;
      RECT  25100.0 32875.0 25170.0 32945.0 ;
      RECT  25172.5 32875.0 25242.5 32945.0 ;
      RECT  25100.0 32375.0 25170.0 32910.0 ;
      RECT  25135.0 32875.0 25207.5 32945.0 ;
      RECT  25172.5 32910.0 25242.5 33442.5 ;
      RECT  25435.0 33287.5 25505.0 33357.5 ;
      RECT  25362.5 33287.5 25432.5 33357.5 ;
      RECT  25435.0 33322.5 25505.0 33925.0 ;
      RECT  25397.5 33287.5 25470.0 33357.5 ;
      RECT  25362.5 32717.5 25432.5 33322.5 ;
      RECT  25100.0 33857.5 25170.0 33992.5 ;
      RECT  25435.0 32307.5 25505.0 32442.5 ;
      RECT  25172.5 33442.5 25242.5 33577.5 ;
      RECT  25362.5 32582.5 25432.5 32717.5 ;
      RECT  25620.0 32482.5 25690.0 32617.5 ;
      RECT  25100.0 33925.0 25170.0 34065.0 ;
      RECT  25435.0 33925.0 25505.0 34065.0 ;
      RECT  25100.0 32235.0 25170.0 32375.0 ;
      RECT  25435.0 32235.0 25505.0 32375.0 ;
      RECT  24915.0 32235.0 24985.0 34065.0 ;
      RECT  25620.0 32235.0 25690.0 34065.0 ;
      RECT  25805.0 32875.0 25875.0 32945.0 ;
      RECT  25877.5 32875.0 25947.5 32945.0 ;
      RECT  25805.0 32375.0 25875.0 32910.0 ;
      RECT  25840.0 32875.0 25912.5 32945.0 ;
      RECT  25877.5 32910.0 25947.5 33442.5 ;
      RECT  26140.0 33287.5 26210.0 33357.5 ;
      RECT  26067.5 33287.5 26137.5 33357.5 ;
      RECT  26140.0 33322.5 26210.0 33925.0 ;
      RECT  26102.5 33287.5 26175.0 33357.5 ;
      RECT  26067.5 32717.5 26137.5 33322.5 ;
      RECT  25805.0 33857.5 25875.0 33992.5 ;
      RECT  26140.0 32307.5 26210.0 32442.5 ;
      RECT  25877.5 33442.5 25947.5 33577.5 ;
      RECT  26067.5 32582.5 26137.5 32717.5 ;
      RECT  26325.0 32482.5 26395.0 32617.5 ;
      RECT  25805.0 33925.0 25875.0 34065.0 ;
      RECT  26140.0 33925.0 26210.0 34065.0 ;
      RECT  25805.0 32235.0 25875.0 32375.0 ;
      RECT  26140.0 32235.0 26210.0 32375.0 ;
      RECT  25620.0 32235.0 25690.0 34065.0 ;
      RECT  26325.0 32235.0 26395.0 34065.0 ;
      RECT  26510.0 32875.0 26580.0 32945.0 ;
      RECT  26582.5 32875.0 26652.5 32945.0 ;
      RECT  26510.0 32375.0 26580.0 32910.0 ;
      RECT  26545.0 32875.0 26617.5 32945.0 ;
      RECT  26582.5 32910.0 26652.5 33442.5 ;
      RECT  26845.0 33287.5 26915.0 33357.5 ;
      RECT  26772.5 33287.5 26842.5 33357.5 ;
      RECT  26845.0 33322.5 26915.0 33925.0 ;
      RECT  26807.5 33287.5 26880.0 33357.5 ;
      RECT  26772.5 32717.5 26842.5 33322.5 ;
      RECT  26510.0 33857.5 26580.0 33992.5 ;
      RECT  26845.0 32307.5 26915.0 32442.5 ;
      RECT  26582.5 33442.5 26652.5 33577.5 ;
      RECT  26772.5 32582.5 26842.5 32717.5 ;
      RECT  27030.0 32482.5 27100.0 32617.5 ;
      RECT  26510.0 33925.0 26580.0 34065.0 ;
      RECT  26845.0 33925.0 26915.0 34065.0 ;
      RECT  26510.0 32235.0 26580.0 32375.0 ;
      RECT  26845.0 32235.0 26915.0 32375.0 ;
      RECT  26325.0 32235.0 26395.0 34065.0 ;
      RECT  27030.0 32235.0 27100.0 34065.0 ;
      RECT  27215.0 32875.0 27285.0 32945.0 ;
      RECT  27287.5 32875.0 27357.5 32945.0 ;
      RECT  27215.0 32375.0 27285.0 32910.0 ;
      RECT  27250.0 32875.0 27322.5 32945.0 ;
      RECT  27287.5 32910.0 27357.5 33442.5 ;
      RECT  27550.0 33287.5 27620.0 33357.5 ;
      RECT  27477.5 33287.5 27547.5 33357.5 ;
      RECT  27550.0 33322.5 27620.0 33925.0 ;
      RECT  27512.5 33287.5 27585.0 33357.5 ;
      RECT  27477.5 32717.5 27547.5 33322.5 ;
      RECT  27215.0 33857.5 27285.0 33992.5 ;
      RECT  27550.0 32307.5 27620.0 32442.5 ;
      RECT  27287.5 33442.5 27357.5 33577.5 ;
      RECT  27477.5 32582.5 27547.5 32717.5 ;
      RECT  27735.0 32482.5 27805.0 32617.5 ;
      RECT  27215.0 33925.0 27285.0 34065.0 ;
      RECT  27550.0 33925.0 27620.0 34065.0 ;
      RECT  27215.0 32235.0 27285.0 32375.0 ;
      RECT  27550.0 32235.0 27620.0 32375.0 ;
      RECT  27030.0 32235.0 27100.0 34065.0 ;
      RECT  27735.0 32235.0 27805.0 34065.0 ;
      RECT  27920.0 32875.0 27990.0 32945.0 ;
      RECT  27992.5 32875.0 28062.5 32945.0 ;
      RECT  27920.0 32375.0 27990.0 32910.0 ;
      RECT  27955.0 32875.0 28027.5 32945.0 ;
      RECT  27992.5 32910.0 28062.5 33442.5 ;
      RECT  28255.0 33287.5 28325.0 33357.5 ;
      RECT  28182.5 33287.5 28252.5 33357.5 ;
      RECT  28255.0 33322.5 28325.0 33925.0 ;
      RECT  28217.5 33287.5 28290.0 33357.5 ;
      RECT  28182.5 32717.5 28252.5 33322.5 ;
      RECT  27920.0 33857.5 27990.0 33992.5 ;
      RECT  28255.0 32307.5 28325.0 32442.5 ;
      RECT  27992.5 33442.5 28062.5 33577.5 ;
      RECT  28182.5 32582.5 28252.5 32717.5 ;
      RECT  28440.0 32482.5 28510.0 32617.5 ;
      RECT  27920.0 33925.0 27990.0 34065.0 ;
      RECT  28255.0 33925.0 28325.0 34065.0 ;
      RECT  27920.0 32235.0 27990.0 32375.0 ;
      RECT  28255.0 32235.0 28325.0 32375.0 ;
      RECT  27735.0 32235.0 27805.0 34065.0 ;
      RECT  28440.0 32235.0 28510.0 34065.0 ;
      RECT  28625.0 32875.0 28695.0 32945.0 ;
      RECT  28697.5 32875.0 28767.5 32945.0 ;
      RECT  28625.0 32375.0 28695.0 32910.0 ;
      RECT  28660.0 32875.0 28732.5 32945.0 ;
      RECT  28697.5 32910.0 28767.5 33442.5 ;
      RECT  28960.0 33287.5 29030.0 33357.5 ;
      RECT  28887.5 33287.5 28957.5 33357.5 ;
      RECT  28960.0 33322.5 29030.0 33925.0 ;
      RECT  28922.5 33287.5 28995.0 33357.5 ;
      RECT  28887.5 32717.5 28957.5 33322.5 ;
      RECT  28625.0 33857.5 28695.0 33992.5 ;
      RECT  28960.0 32307.5 29030.0 32442.5 ;
      RECT  28697.5 33442.5 28767.5 33577.5 ;
      RECT  28887.5 32582.5 28957.5 32717.5 ;
      RECT  29145.0 32482.5 29215.0 32617.5 ;
      RECT  28625.0 33925.0 28695.0 34065.0 ;
      RECT  28960.0 33925.0 29030.0 34065.0 ;
      RECT  28625.0 32235.0 28695.0 32375.0 ;
      RECT  28960.0 32235.0 29030.0 32375.0 ;
      RECT  28440.0 32235.0 28510.0 34065.0 ;
      RECT  29145.0 32235.0 29215.0 34065.0 ;
      RECT  29330.0 32875.0 29400.0 32945.0 ;
      RECT  29402.5 32875.0 29472.5 32945.0 ;
      RECT  29330.0 32375.0 29400.0 32910.0 ;
      RECT  29365.0 32875.0 29437.5 32945.0 ;
      RECT  29402.5 32910.0 29472.5 33442.5 ;
      RECT  29665.0 33287.5 29735.0 33357.5 ;
      RECT  29592.5 33287.5 29662.5 33357.5 ;
      RECT  29665.0 33322.5 29735.0 33925.0 ;
      RECT  29627.5 33287.5 29700.0 33357.5 ;
      RECT  29592.5 32717.5 29662.5 33322.5 ;
      RECT  29330.0 33857.5 29400.0 33992.5 ;
      RECT  29665.0 32307.5 29735.0 32442.5 ;
      RECT  29402.5 33442.5 29472.5 33577.5 ;
      RECT  29592.5 32582.5 29662.5 32717.5 ;
      RECT  29850.0 32482.5 29920.0 32617.5 ;
      RECT  29330.0 33925.0 29400.0 34065.0 ;
      RECT  29665.0 33925.0 29735.0 34065.0 ;
      RECT  29330.0 32235.0 29400.0 32375.0 ;
      RECT  29665.0 32235.0 29735.0 32375.0 ;
      RECT  29145.0 32235.0 29215.0 34065.0 ;
      RECT  29850.0 32235.0 29920.0 34065.0 ;
      RECT  30035.0 32875.0 30105.0 32945.0 ;
      RECT  30107.5 32875.0 30177.5 32945.0 ;
      RECT  30035.0 32375.0 30105.0 32910.0 ;
      RECT  30070.0 32875.0 30142.5 32945.0 ;
      RECT  30107.5 32910.0 30177.5 33442.5 ;
      RECT  30370.0 33287.5 30440.0 33357.5 ;
      RECT  30297.5 33287.5 30367.5 33357.5 ;
      RECT  30370.0 33322.5 30440.0 33925.0 ;
      RECT  30332.5 33287.5 30405.0 33357.5 ;
      RECT  30297.5 32717.5 30367.5 33322.5 ;
      RECT  30035.0 33857.5 30105.0 33992.5 ;
      RECT  30370.0 32307.5 30440.0 32442.5 ;
      RECT  30107.5 33442.5 30177.5 33577.5 ;
      RECT  30297.5 32582.5 30367.5 32717.5 ;
      RECT  30555.0 32482.5 30625.0 32617.5 ;
      RECT  30035.0 33925.0 30105.0 34065.0 ;
      RECT  30370.0 33925.0 30440.0 34065.0 ;
      RECT  30035.0 32235.0 30105.0 32375.0 ;
      RECT  30370.0 32235.0 30440.0 32375.0 ;
      RECT  29850.0 32235.0 29920.0 34065.0 ;
      RECT  30555.0 32235.0 30625.0 34065.0 ;
      RECT  30740.0 32875.0 30810.0 32945.0 ;
      RECT  30812.5 32875.0 30882.5 32945.0 ;
      RECT  30740.0 32375.0 30810.0 32910.0 ;
      RECT  30775.0 32875.0 30847.5 32945.0 ;
      RECT  30812.5 32910.0 30882.5 33442.5 ;
      RECT  31075.0 33287.5 31145.0 33357.5 ;
      RECT  31002.5 33287.5 31072.5 33357.5 ;
      RECT  31075.0 33322.5 31145.0 33925.0 ;
      RECT  31037.5 33287.5 31110.0 33357.5 ;
      RECT  31002.5 32717.5 31072.5 33322.5 ;
      RECT  30740.0 33857.5 30810.0 33992.5 ;
      RECT  31075.0 32307.5 31145.0 32442.5 ;
      RECT  30812.5 33442.5 30882.5 33577.5 ;
      RECT  31002.5 32582.5 31072.5 32717.5 ;
      RECT  31260.0 32482.5 31330.0 32617.5 ;
      RECT  30740.0 33925.0 30810.0 34065.0 ;
      RECT  31075.0 33925.0 31145.0 34065.0 ;
      RECT  30740.0 32235.0 30810.0 32375.0 ;
      RECT  31075.0 32235.0 31145.0 32375.0 ;
      RECT  30555.0 32235.0 30625.0 34065.0 ;
      RECT  31260.0 32235.0 31330.0 34065.0 ;
      RECT  31445.0 32875.0 31515.0 32945.0 ;
      RECT  31517.5 32875.0 31587.5 32945.0 ;
      RECT  31445.0 32375.0 31515.0 32910.0 ;
      RECT  31480.0 32875.0 31552.5 32945.0 ;
      RECT  31517.5 32910.0 31587.5 33442.5 ;
      RECT  31780.0 33287.5 31850.0 33357.5 ;
      RECT  31707.5 33287.5 31777.5 33357.5 ;
      RECT  31780.0 33322.5 31850.0 33925.0 ;
      RECT  31742.5 33287.5 31815.0 33357.5 ;
      RECT  31707.5 32717.5 31777.5 33322.5 ;
      RECT  31445.0 33857.5 31515.0 33992.5 ;
      RECT  31780.0 32307.5 31850.0 32442.5 ;
      RECT  31517.5 33442.5 31587.5 33577.5 ;
      RECT  31707.5 32582.5 31777.5 32717.5 ;
      RECT  31965.0 32482.5 32035.0 32617.5 ;
      RECT  31445.0 33925.0 31515.0 34065.0 ;
      RECT  31780.0 33925.0 31850.0 34065.0 ;
      RECT  31445.0 32235.0 31515.0 32375.0 ;
      RECT  31780.0 32235.0 31850.0 32375.0 ;
      RECT  31260.0 32235.0 31330.0 34065.0 ;
      RECT  31965.0 32235.0 32035.0 34065.0 ;
      RECT  32150.0 32875.0 32220.0 32945.0 ;
      RECT  32222.5 32875.0 32292.5 32945.0 ;
      RECT  32150.0 32375.0 32220.0 32910.0 ;
      RECT  32185.0 32875.0 32257.5 32945.0 ;
      RECT  32222.5 32910.0 32292.5 33442.5 ;
      RECT  32485.0 33287.5 32555.0 33357.5 ;
      RECT  32412.5 33287.5 32482.5 33357.5 ;
      RECT  32485.0 33322.5 32555.0 33925.0 ;
      RECT  32447.5 33287.5 32520.0 33357.5 ;
      RECT  32412.5 32717.5 32482.5 33322.5 ;
      RECT  32150.0 33857.5 32220.0 33992.5 ;
      RECT  32485.0 32307.5 32555.0 32442.5 ;
      RECT  32222.5 33442.5 32292.5 33577.5 ;
      RECT  32412.5 32582.5 32482.5 32717.5 ;
      RECT  32670.0 32482.5 32740.0 32617.5 ;
      RECT  32150.0 33925.0 32220.0 34065.0 ;
      RECT  32485.0 33925.0 32555.0 34065.0 ;
      RECT  32150.0 32235.0 32220.0 32375.0 ;
      RECT  32485.0 32235.0 32555.0 32375.0 ;
      RECT  31965.0 32235.0 32035.0 34065.0 ;
      RECT  32670.0 32235.0 32740.0 34065.0 ;
      RECT  32855.0 32875.0 32925.0 32945.0 ;
      RECT  32927.5 32875.0 32997.5 32945.0 ;
      RECT  32855.0 32375.0 32925.0 32910.0 ;
      RECT  32890.0 32875.0 32962.5 32945.0 ;
      RECT  32927.5 32910.0 32997.5 33442.5 ;
      RECT  33190.0 33287.5 33260.0 33357.5 ;
      RECT  33117.5 33287.5 33187.5 33357.5 ;
      RECT  33190.0 33322.5 33260.0 33925.0 ;
      RECT  33152.5 33287.5 33225.0 33357.5 ;
      RECT  33117.5 32717.5 33187.5 33322.5 ;
      RECT  32855.0 33857.5 32925.0 33992.5 ;
      RECT  33190.0 32307.5 33260.0 32442.5 ;
      RECT  32927.5 33442.5 32997.5 33577.5 ;
      RECT  33117.5 32582.5 33187.5 32717.5 ;
      RECT  33375.0 32482.5 33445.0 32617.5 ;
      RECT  32855.0 33925.0 32925.0 34065.0 ;
      RECT  33190.0 33925.0 33260.0 34065.0 ;
      RECT  32855.0 32235.0 32925.0 32375.0 ;
      RECT  33190.0 32235.0 33260.0 32375.0 ;
      RECT  32670.0 32235.0 32740.0 34065.0 ;
      RECT  33375.0 32235.0 33445.0 34065.0 ;
      RECT  33560.0 32875.0 33630.0 32945.0 ;
      RECT  33632.5 32875.0 33702.5 32945.0 ;
      RECT  33560.0 32375.0 33630.0 32910.0 ;
      RECT  33595.0 32875.0 33667.5 32945.0 ;
      RECT  33632.5 32910.0 33702.5 33442.5 ;
      RECT  33895.0 33287.5 33965.0 33357.5 ;
      RECT  33822.5 33287.5 33892.5 33357.5 ;
      RECT  33895.0 33322.5 33965.0 33925.0 ;
      RECT  33857.5 33287.5 33930.0 33357.5 ;
      RECT  33822.5 32717.5 33892.5 33322.5 ;
      RECT  33560.0 33857.5 33630.0 33992.5 ;
      RECT  33895.0 32307.5 33965.0 32442.5 ;
      RECT  33632.5 33442.5 33702.5 33577.5 ;
      RECT  33822.5 32582.5 33892.5 32717.5 ;
      RECT  34080.0 32482.5 34150.0 32617.5 ;
      RECT  33560.0 33925.0 33630.0 34065.0 ;
      RECT  33895.0 33925.0 33965.0 34065.0 ;
      RECT  33560.0 32235.0 33630.0 32375.0 ;
      RECT  33895.0 32235.0 33965.0 32375.0 ;
      RECT  33375.0 32235.0 33445.0 34065.0 ;
      RECT  34080.0 32235.0 34150.0 34065.0 ;
      RECT  34265.0 32875.0 34335.0 32945.0 ;
      RECT  34337.5 32875.0 34407.5 32945.0 ;
      RECT  34265.0 32375.0 34335.0 32910.0 ;
      RECT  34300.0 32875.0 34372.5 32945.0 ;
      RECT  34337.5 32910.0 34407.5 33442.5 ;
      RECT  34600.0 33287.5 34670.0 33357.5 ;
      RECT  34527.5 33287.5 34597.5 33357.5 ;
      RECT  34600.0 33322.5 34670.0 33925.0 ;
      RECT  34562.5 33287.5 34635.0 33357.5 ;
      RECT  34527.5 32717.5 34597.5 33322.5 ;
      RECT  34265.0 33857.5 34335.0 33992.5 ;
      RECT  34600.0 32307.5 34670.0 32442.5 ;
      RECT  34337.5 33442.5 34407.5 33577.5 ;
      RECT  34527.5 32582.5 34597.5 32717.5 ;
      RECT  34785.0 32482.5 34855.0 32617.5 ;
      RECT  34265.0 33925.0 34335.0 34065.0 ;
      RECT  34600.0 33925.0 34670.0 34065.0 ;
      RECT  34265.0 32235.0 34335.0 32375.0 ;
      RECT  34600.0 32235.0 34670.0 32375.0 ;
      RECT  34080.0 32235.0 34150.0 34065.0 ;
      RECT  34785.0 32235.0 34855.0 34065.0 ;
      RECT  34970.0 32875.0 35040.0 32945.0 ;
      RECT  35042.5 32875.0 35112.5 32945.0 ;
      RECT  34970.0 32375.0 35040.0 32910.0 ;
      RECT  35005.0 32875.0 35077.5 32945.0 ;
      RECT  35042.5 32910.0 35112.5 33442.5 ;
      RECT  35305.0 33287.5 35375.0 33357.5 ;
      RECT  35232.5 33287.5 35302.5 33357.5 ;
      RECT  35305.0 33322.5 35375.0 33925.0 ;
      RECT  35267.5 33287.5 35340.0 33357.5 ;
      RECT  35232.5 32717.5 35302.5 33322.5 ;
      RECT  34970.0 33857.5 35040.0 33992.5 ;
      RECT  35305.0 32307.5 35375.0 32442.5 ;
      RECT  35042.5 33442.5 35112.5 33577.5 ;
      RECT  35232.5 32582.5 35302.5 32717.5 ;
      RECT  35490.0 32482.5 35560.0 32617.5 ;
      RECT  34970.0 33925.0 35040.0 34065.0 ;
      RECT  35305.0 33925.0 35375.0 34065.0 ;
      RECT  34970.0 32235.0 35040.0 32375.0 ;
      RECT  35305.0 32235.0 35375.0 32375.0 ;
      RECT  34785.0 32235.0 34855.0 34065.0 ;
      RECT  35490.0 32235.0 35560.0 34065.0 ;
      RECT  35675.0 32875.0 35745.0 32945.0 ;
      RECT  35747.5 32875.0 35817.5 32945.0 ;
      RECT  35675.0 32375.0 35745.0 32910.0 ;
      RECT  35710.0 32875.0 35782.5 32945.0 ;
      RECT  35747.5 32910.0 35817.5 33442.5 ;
      RECT  36010.0 33287.5 36080.0 33357.5 ;
      RECT  35937.5 33287.5 36007.5 33357.5 ;
      RECT  36010.0 33322.5 36080.0 33925.0 ;
      RECT  35972.5 33287.5 36045.0 33357.5 ;
      RECT  35937.5 32717.5 36007.5 33322.5 ;
      RECT  35675.0 33857.5 35745.0 33992.5 ;
      RECT  36010.0 32307.5 36080.0 32442.5 ;
      RECT  35747.5 33442.5 35817.5 33577.5 ;
      RECT  35937.5 32582.5 36007.5 32717.5 ;
      RECT  36195.0 32482.5 36265.0 32617.5 ;
      RECT  35675.0 33925.0 35745.0 34065.0 ;
      RECT  36010.0 33925.0 36080.0 34065.0 ;
      RECT  35675.0 32235.0 35745.0 32375.0 ;
      RECT  36010.0 32235.0 36080.0 32375.0 ;
      RECT  35490.0 32235.0 35560.0 34065.0 ;
      RECT  36195.0 32235.0 36265.0 34065.0 ;
      RECT  36380.0 32875.0 36450.0 32945.0 ;
      RECT  36452.5 32875.0 36522.5 32945.0 ;
      RECT  36380.0 32375.0 36450.0 32910.0 ;
      RECT  36415.0 32875.0 36487.5 32945.0 ;
      RECT  36452.5 32910.0 36522.5 33442.5 ;
      RECT  36715.0 33287.5 36785.0 33357.5 ;
      RECT  36642.5 33287.5 36712.5 33357.5 ;
      RECT  36715.0 33322.5 36785.0 33925.0 ;
      RECT  36677.5 33287.5 36750.0 33357.5 ;
      RECT  36642.5 32717.5 36712.5 33322.5 ;
      RECT  36380.0 33857.5 36450.0 33992.5 ;
      RECT  36715.0 32307.5 36785.0 32442.5 ;
      RECT  36452.5 33442.5 36522.5 33577.5 ;
      RECT  36642.5 32582.5 36712.5 32717.5 ;
      RECT  36900.0 32482.5 36970.0 32617.5 ;
      RECT  36380.0 33925.0 36450.0 34065.0 ;
      RECT  36715.0 33925.0 36785.0 34065.0 ;
      RECT  36380.0 32235.0 36450.0 32375.0 ;
      RECT  36715.0 32235.0 36785.0 32375.0 ;
      RECT  36195.0 32235.0 36265.0 34065.0 ;
      RECT  36900.0 32235.0 36970.0 34065.0 ;
      RECT  37085.0 32875.0 37155.0 32945.0 ;
      RECT  37157.5 32875.0 37227.5 32945.0 ;
      RECT  37085.0 32375.0 37155.0 32910.0 ;
      RECT  37120.0 32875.0 37192.5 32945.0 ;
      RECT  37157.5 32910.0 37227.5 33442.5 ;
      RECT  37420.0 33287.5 37490.0 33357.5 ;
      RECT  37347.5 33287.5 37417.5 33357.5 ;
      RECT  37420.0 33322.5 37490.0 33925.0 ;
      RECT  37382.5 33287.5 37455.0 33357.5 ;
      RECT  37347.5 32717.5 37417.5 33322.5 ;
      RECT  37085.0 33857.5 37155.0 33992.5 ;
      RECT  37420.0 32307.5 37490.0 32442.5 ;
      RECT  37157.5 33442.5 37227.5 33577.5 ;
      RECT  37347.5 32582.5 37417.5 32717.5 ;
      RECT  37605.0 32482.5 37675.0 32617.5 ;
      RECT  37085.0 33925.0 37155.0 34065.0 ;
      RECT  37420.0 33925.0 37490.0 34065.0 ;
      RECT  37085.0 32235.0 37155.0 32375.0 ;
      RECT  37420.0 32235.0 37490.0 32375.0 ;
      RECT  36900.0 32235.0 36970.0 34065.0 ;
      RECT  37605.0 32235.0 37675.0 34065.0 ;
      RECT  37790.0 32875.0 37860.0 32945.0 ;
      RECT  37862.5 32875.0 37932.5 32945.0 ;
      RECT  37790.0 32375.0 37860.0 32910.0 ;
      RECT  37825.0 32875.0 37897.5 32945.0 ;
      RECT  37862.5 32910.0 37932.5 33442.5 ;
      RECT  38125.0 33287.5 38195.0 33357.5 ;
      RECT  38052.5 33287.5 38122.5 33357.5 ;
      RECT  38125.0 33322.5 38195.0 33925.0 ;
      RECT  38087.5 33287.5 38160.0 33357.5 ;
      RECT  38052.5 32717.5 38122.5 33322.5 ;
      RECT  37790.0 33857.5 37860.0 33992.5 ;
      RECT  38125.0 32307.5 38195.0 32442.5 ;
      RECT  37862.5 33442.5 37932.5 33577.5 ;
      RECT  38052.5 32582.5 38122.5 32717.5 ;
      RECT  38310.0 32482.5 38380.0 32617.5 ;
      RECT  37790.0 33925.0 37860.0 34065.0 ;
      RECT  38125.0 33925.0 38195.0 34065.0 ;
      RECT  37790.0 32235.0 37860.0 32375.0 ;
      RECT  38125.0 32235.0 38195.0 32375.0 ;
      RECT  37605.0 32235.0 37675.0 34065.0 ;
      RECT  38310.0 32235.0 38380.0 34065.0 ;
      RECT  38495.0 32875.0 38565.0 32945.0 ;
      RECT  38567.5 32875.0 38637.5 32945.0 ;
      RECT  38495.0 32375.0 38565.0 32910.0 ;
      RECT  38530.0 32875.0 38602.5 32945.0 ;
      RECT  38567.5 32910.0 38637.5 33442.5 ;
      RECT  38830.0 33287.5 38900.0 33357.5 ;
      RECT  38757.5 33287.5 38827.5 33357.5 ;
      RECT  38830.0 33322.5 38900.0 33925.0 ;
      RECT  38792.5 33287.5 38865.0 33357.5 ;
      RECT  38757.5 32717.5 38827.5 33322.5 ;
      RECT  38495.0 33857.5 38565.0 33992.5 ;
      RECT  38830.0 32307.5 38900.0 32442.5 ;
      RECT  38567.5 33442.5 38637.5 33577.5 ;
      RECT  38757.5 32582.5 38827.5 32717.5 ;
      RECT  39015.0 32482.5 39085.0 32617.5 ;
      RECT  38495.0 33925.0 38565.0 34065.0 ;
      RECT  38830.0 33925.0 38900.0 34065.0 ;
      RECT  38495.0 32235.0 38565.0 32375.0 ;
      RECT  38830.0 32235.0 38900.0 32375.0 ;
      RECT  38310.0 32235.0 38380.0 34065.0 ;
      RECT  39015.0 32235.0 39085.0 34065.0 ;
      RECT  39200.0 32875.0 39270.0 32945.0 ;
      RECT  39272.5 32875.0 39342.5 32945.0 ;
      RECT  39200.0 32375.0 39270.0 32910.0 ;
      RECT  39235.0 32875.0 39307.5 32945.0 ;
      RECT  39272.5 32910.0 39342.5 33442.5 ;
      RECT  39535.0 33287.5 39605.0 33357.5 ;
      RECT  39462.5 33287.5 39532.5 33357.5 ;
      RECT  39535.0 33322.5 39605.0 33925.0 ;
      RECT  39497.5 33287.5 39570.0 33357.5 ;
      RECT  39462.5 32717.5 39532.5 33322.5 ;
      RECT  39200.0 33857.5 39270.0 33992.5 ;
      RECT  39535.0 32307.5 39605.0 32442.5 ;
      RECT  39272.5 33442.5 39342.5 33577.5 ;
      RECT  39462.5 32582.5 39532.5 32717.5 ;
      RECT  39720.0 32482.5 39790.0 32617.5 ;
      RECT  39200.0 33925.0 39270.0 34065.0 ;
      RECT  39535.0 33925.0 39605.0 34065.0 ;
      RECT  39200.0 32235.0 39270.0 32375.0 ;
      RECT  39535.0 32235.0 39605.0 32375.0 ;
      RECT  39015.0 32235.0 39085.0 34065.0 ;
      RECT  39720.0 32235.0 39790.0 34065.0 ;
      RECT  39905.0 32875.0 39975.0 32945.0 ;
      RECT  39977.5 32875.0 40047.5 32945.0 ;
      RECT  39905.0 32375.0 39975.0 32910.0 ;
      RECT  39940.0 32875.0 40012.5 32945.0 ;
      RECT  39977.5 32910.0 40047.5 33442.5 ;
      RECT  40240.0 33287.5 40310.0 33357.5 ;
      RECT  40167.5 33287.5 40237.5 33357.5 ;
      RECT  40240.0 33322.5 40310.0 33925.0 ;
      RECT  40202.5 33287.5 40275.0 33357.5 ;
      RECT  40167.5 32717.5 40237.5 33322.5 ;
      RECT  39905.0 33857.5 39975.0 33992.5 ;
      RECT  40240.0 32307.5 40310.0 32442.5 ;
      RECT  39977.5 33442.5 40047.5 33577.5 ;
      RECT  40167.5 32582.5 40237.5 32717.5 ;
      RECT  40425.0 32482.5 40495.0 32617.5 ;
      RECT  39905.0 33925.0 39975.0 34065.0 ;
      RECT  40240.0 33925.0 40310.0 34065.0 ;
      RECT  39905.0 32235.0 39975.0 32375.0 ;
      RECT  40240.0 32235.0 40310.0 32375.0 ;
      RECT  39720.0 32235.0 39790.0 34065.0 ;
      RECT  40425.0 32235.0 40495.0 34065.0 ;
      RECT  40610.0 32875.0 40680.0 32945.0 ;
      RECT  40682.5 32875.0 40752.5 32945.0 ;
      RECT  40610.0 32375.0 40680.0 32910.0 ;
      RECT  40645.0 32875.0 40717.5 32945.0 ;
      RECT  40682.5 32910.0 40752.5 33442.5 ;
      RECT  40945.0 33287.5 41015.0 33357.5 ;
      RECT  40872.5 33287.5 40942.5 33357.5 ;
      RECT  40945.0 33322.5 41015.0 33925.0 ;
      RECT  40907.5 33287.5 40980.0 33357.5 ;
      RECT  40872.5 32717.5 40942.5 33322.5 ;
      RECT  40610.0 33857.5 40680.0 33992.5 ;
      RECT  40945.0 32307.5 41015.0 32442.5 ;
      RECT  40682.5 33442.5 40752.5 33577.5 ;
      RECT  40872.5 32582.5 40942.5 32717.5 ;
      RECT  41130.0 32482.5 41200.0 32617.5 ;
      RECT  40610.0 33925.0 40680.0 34065.0 ;
      RECT  40945.0 33925.0 41015.0 34065.0 ;
      RECT  40610.0 32235.0 40680.0 32375.0 ;
      RECT  40945.0 32235.0 41015.0 32375.0 ;
      RECT  40425.0 32235.0 40495.0 34065.0 ;
      RECT  41130.0 32235.0 41200.0 34065.0 ;
      RECT  41315.0 32875.0 41385.0 32945.0 ;
      RECT  41387.5 32875.0 41457.5 32945.0 ;
      RECT  41315.0 32375.0 41385.0 32910.0 ;
      RECT  41350.0 32875.0 41422.5 32945.0 ;
      RECT  41387.5 32910.0 41457.5 33442.5 ;
      RECT  41650.0 33287.5 41720.0 33357.5 ;
      RECT  41577.5 33287.5 41647.5 33357.5 ;
      RECT  41650.0 33322.5 41720.0 33925.0 ;
      RECT  41612.5 33287.5 41685.0 33357.5 ;
      RECT  41577.5 32717.5 41647.5 33322.5 ;
      RECT  41315.0 33857.5 41385.0 33992.5 ;
      RECT  41650.0 32307.5 41720.0 32442.5 ;
      RECT  41387.5 33442.5 41457.5 33577.5 ;
      RECT  41577.5 32582.5 41647.5 32717.5 ;
      RECT  41835.0 32482.5 41905.0 32617.5 ;
      RECT  41315.0 33925.0 41385.0 34065.0 ;
      RECT  41650.0 33925.0 41720.0 34065.0 ;
      RECT  41315.0 32235.0 41385.0 32375.0 ;
      RECT  41650.0 32235.0 41720.0 32375.0 ;
      RECT  41130.0 32235.0 41200.0 34065.0 ;
      RECT  41835.0 32235.0 41905.0 34065.0 ;
      RECT  42020.0 32875.0 42090.0 32945.0 ;
      RECT  42092.5 32875.0 42162.5 32945.0 ;
      RECT  42020.0 32375.0 42090.0 32910.0 ;
      RECT  42055.0 32875.0 42127.5 32945.0 ;
      RECT  42092.5 32910.0 42162.5 33442.5 ;
      RECT  42355.0 33287.5 42425.0 33357.5 ;
      RECT  42282.5 33287.5 42352.5 33357.5 ;
      RECT  42355.0 33322.5 42425.0 33925.0 ;
      RECT  42317.5 33287.5 42390.0 33357.5 ;
      RECT  42282.5 32717.5 42352.5 33322.5 ;
      RECT  42020.0 33857.5 42090.0 33992.5 ;
      RECT  42355.0 32307.5 42425.0 32442.5 ;
      RECT  42092.5 33442.5 42162.5 33577.5 ;
      RECT  42282.5 32582.5 42352.5 32717.5 ;
      RECT  42540.0 32482.5 42610.0 32617.5 ;
      RECT  42020.0 33925.0 42090.0 34065.0 ;
      RECT  42355.0 33925.0 42425.0 34065.0 ;
      RECT  42020.0 32235.0 42090.0 32375.0 ;
      RECT  42355.0 32235.0 42425.0 32375.0 ;
      RECT  41835.0 32235.0 41905.0 34065.0 ;
      RECT  42540.0 32235.0 42610.0 34065.0 ;
      RECT  42725.0 32875.0 42795.0 32945.0 ;
      RECT  42797.5 32875.0 42867.5 32945.0 ;
      RECT  42725.0 32375.0 42795.0 32910.0 ;
      RECT  42760.0 32875.0 42832.5 32945.0 ;
      RECT  42797.5 32910.0 42867.5 33442.5 ;
      RECT  43060.0 33287.5 43130.0 33357.5 ;
      RECT  42987.5 33287.5 43057.5 33357.5 ;
      RECT  43060.0 33322.5 43130.0 33925.0 ;
      RECT  43022.5 33287.5 43095.0 33357.5 ;
      RECT  42987.5 32717.5 43057.5 33322.5 ;
      RECT  42725.0 33857.5 42795.0 33992.5 ;
      RECT  43060.0 32307.5 43130.0 32442.5 ;
      RECT  42797.5 33442.5 42867.5 33577.5 ;
      RECT  42987.5 32582.5 43057.5 32717.5 ;
      RECT  43245.0 32482.5 43315.0 32617.5 ;
      RECT  42725.0 33925.0 42795.0 34065.0 ;
      RECT  43060.0 33925.0 43130.0 34065.0 ;
      RECT  42725.0 32235.0 42795.0 32375.0 ;
      RECT  43060.0 32235.0 43130.0 32375.0 ;
      RECT  42540.0 32235.0 42610.0 34065.0 ;
      RECT  43245.0 32235.0 43315.0 34065.0 ;
      RECT  43430.0 32875.0 43500.0 32945.0 ;
      RECT  43502.5 32875.0 43572.5 32945.0 ;
      RECT  43430.0 32375.0 43500.0 32910.0 ;
      RECT  43465.0 32875.0 43537.5 32945.0 ;
      RECT  43502.5 32910.0 43572.5 33442.5 ;
      RECT  43765.0 33287.5 43835.0 33357.5 ;
      RECT  43692.5 33287.5 43762.5 33357.5 ;
      RECT  43765.0 33322.5 43835.0 33925.0 ;
      RECT  43727.5 33287.5 43800.0 33357.5 ;
      RECT  43692.5 32717.5 43762.5 33322.5 ;
      RECT  43430.0 33857.5 43500.0 33992.5 ;
      RECT  43765.0 32307.5 43835.0 32442.5 ;
      RECT  43502.5 33442.5 43572.5 33577.5 ;
      RECT  43692.5 32582.5 43762.5 32717.5 ;
      RECT  43950.0 32482.5 44020.0 32617.5 ;
      RECT  43430.0 33925.0 43500.0 34065.0 ;
      RECT  43765.0 33925.0 43835.0 34065.0 ;
      RECT  43430.0 32235.0 43500.0 32375.0 ;
      RECT  43765.0 32235.0 43835.0 32375.0 ;
      RECT  43245.0 32235.0 43315.0 34065.0 ;
      RECT  43950.0 32235.0 44020.0 34065.0 ;
      RECT  44135.0 32875.0 44205.0 32945.0 ;
      RECT  44207.5 32875.0 44277.5 32945.0 ;
      RECT  44135.0 32375.0 44205.0 32910.0 ;
      RECT  44170.0 32875.0 44242.5 32945.0 ;
      RECT  44207.5 32910.0 44277.5 33442.5 ;
      RECT  44470.0 33287.5 44540.0 33357.5 ;
      RECT  44397.5 33287.5 44467.5 33357.5 ;
      RECT  44470.0 33322.5 44540.0 33925.0 ;
      RECT  44432.5 33287.5 44505.0 33357.5 ;
      RECT  44397.5 32717.5 44467.5 33322.5 ;
      RECT  44135.0 33857.5 44205.0 33992.5 ;
      RECT  44470.0 32307.5 44540.0 32442.5 ;
      RECT  44207.5 33442.5 44277.5 33577.5 ;
      RECT  44397.5 32582.5 44467.5 32717.5 ;
      RECT  44655.0 32482.5 44725.0 32617.5 ;
      RECT  44135.0 33925.0 44205.0 34065.0 ;
      RECT  44470.0 33925.0 44540.0 34065.0 ;
      RECT  44135.0 32235.0 44205.0 32375.0 ;
      RECT  44470.0 32235.0 44540.0 32375.0 ;
      RECT  43950.0 32235.0 44020.0 34065.0 ;
      RECT  44655.0 32235.0 44725.0 34065.0 ;
      RECT  44840.0 32875.0 44910.0 32945.0 ;
      RECT  44912.5 32875.0 44982.5 32945.0 ;
      RECT  44840.0 32375.0 44910.0 32910.0 ;
      RECT  44875.0 32875.0 44947.5 32945.0 ;
      RECT  44912.5 32910.0 44982.5 33442.5 ;
      RECT  45175.0 33287.5 45245.0 33357.5 ;
      RECT  45102.5 33287.5 45172.5 33357.5 ;
      RECT  45175.0 33322.5 45245.0 33925.0 ;
      RECT  45137.5 33287.5 45210.0 33357.5 ;
      RECT  45102.5 32717.5 45172.5 33322.5 ;
      RECT  44840.0 33857.5 44910.0 33992.5 ;
      RECT  45175.0 32307.5 45245.0 32442.5 ;
      RECT  44912.5 33442.5 44982.5 33577.5 ;
      RECT  45102.5 32582.5 45172.5 32717.5 ;
      RECT  45360.0 32482.5 45430.0 32617.5 ;
      RECT  44840.0 33925.0 44910.0 34065.0 ;
      RECT  45175.0 33925.0 45245.0 34065.0 ;
      RECT  44840.0 32235.0 44910.0 32375.0 ;
      RECT  45175.0 32235.0 45245.0 32375.0 ;
      RECT  44655.0 32235.0 44725.0 34065.0 ;
      RECT  45360.0 32235.0 45430.0 34065.0 ;
      RECT  45545.0 32875.0 45615.0 32945.0 ;
      RECT  45617.5 32875.0 45687.5 32945.0 ;
      RECT  45545.0 32375.0 45615.0 32910.0 ;
      RECT  45580.0 32875.0 45652.5 32945.0 ;
      RECT  45617.5 32910.0 45687.5 33442.5 ;
      RECT  45880.0 33287.5 45950.0 33357.5 ;
      RECT  45807.5 33287.5 45877.5 33357.5 ;
      RECT  45880.0 33322.5 45950.0 33925.0 ;
      RECT  45842.5 33287.5 45915.0 33357.5 ;
      RECT  45807.5 32717.5 45877.5 33322.5 ;
      RECT  45545.0 33857.5 45615.0 33992.5 ;
      RECT  45880.0 32307.5 45950.0 32442.5 ;
      RECT  45617.5 33442.5 45687.5 33577.5 ;
      RECT  45807.5 32582.5 45877.5 32717.5 ;
      RECT  46065.0 32482.5 46135.0 32617.5 ;
      RECT  45545.0 33925.0 45615.0 34065.0 ;
      RECT  45880.0 33925.0 45950.0 34065.0 ;
      RECT  45545.0 32235.0 45615.0 32375.0 ;
      RECT  45880.0 32235.0 45950.0 32375.0 ;
      RECT  45360.0 32235.0 45430.0 34065.0 ;
      RECT  46065.0 32235.0 46135.0 34065.0 ;
      RECT  46250.0 32875.0 46320.0 32945.0 ;
      RECT  46322.5 32875.0 46392.5 32945.0 ;
      RECT  46250.0 32375.0 46320.0 32910.0 ;
      RECT  46285.0 32875.0 46357.5 32945.0 ;
      RECT  46322.5 32910.0 46392.5 33442.5 ;
      RECT  46585.0 33287.5 46655.0 33357.5 ;
      RECT  46512.5 33287.5 46582.5 33357.5 ;
      RECT  46585.0 33322.5 46655.0 33925.0 ;
      RECT  46547.5 33287.5 46620.0 33357.5 ;
      RECT  46512.5 32717.5 46582.5 33322.5 ;
      RECT  46250.0 33857.5 46320.0 33992.5 ;
      RECT  46585.0 32307.5 46655.0 32442.5 ;
      RECT  46322.5 33442.5 46392.5 33577.5 ;
      RECT  46512.5 32582.5 46582.5 32717.5 ;
      RECT  46770.0 32482.5 46840.0 32617.5 ;
      RECT  46250.0 33925.0 46320.0 34065.0 ;
      RECT  46585.0 33925.0 46655.0 34065.0 ;
      RECT  46250.0 32235.0 46320.0 32375.0 ;
      RECT  46585.0 32235.0 46655.0 32375.0 ;
      RECT  46065.0 32235.0 46135.0 34065.0 ;
      RECT  46770.0 32235.0 46840.0 34065.0 ;
      RECT  46955.0 32875.0 47025.0 32945.0 ;
      RECT  47027.5 32875.0 47097.5 32945.0 ;
      RECT  46955.0 32375.0 47025.0 32910.0 ;
      RECT  46990.0 32875.0 47062.5 32945.0 ;
      RECT  47027.5 32910.0 47097.5 33442.5 ;
      RECT  47290.0 33287.5 47360.0 33357.5 ;
      RECT  47217.5 33287.5 47287.5 33357.5 ;
      RECT  47290.0 33322.5 47360.0 33925.0 ;
      RECT  47252.5 33287.5 47325.0 33357.5 ;
      RECT  47217.5 32717.5 47287.5 33322.5 ;
      RECT  46955.0 33857.5 47025.0 33992.5 ;
      RECT  47290.0 32307.5 47360.0 32442.5 ;
      RECT  47027.5 33442.5 47097.5 33577.5 ;
      RECT  47217.5 32582.5 47287.5 32717.5 ;
      RECT  47475.0 32482.5 47545.0 32617.5 ;
      RECT  46955.0 33925.0 47025.0 34065.0 ;
      RECT  47290.0 33925.0 47360.0 34065.0 ;
      RECT  46955.0 32235.0 47025.0 32375.0 ;
      RECT  47290.0 32235.0 47360.0 32375.0 ;
      RECT  46770.0 32235.0 46840.0 34065.0 ;
      RECT  47475.0 32235.0 47545.0 34065.0 ;
      RECT  47660.0 32875.0 47730.0 32945.0 ;
      RECT  47732.5 32875.0 47802.5 32945.0 ;
      RECT  47660.0 32375.0 47730.0 32910.0 ;
      RECT  47695.0 32875.0 47767.5 32945.0 ;
      RECT  47732.5 32910.0 47802.5 33442.5 ;
      RECT  47995.0 33287.5 48065.0 33357.5 ;
      RECT  47922.5 33287.5 47992.5 33357.5 ;
      RECT  47995.0 33322.5 48065.0 33925.0 ;
      RECT  47957.5 33287.5 48030.0 33357.5 ;
      RECT  47922.5 32717.5 47992.5 33322.5 ;
      RECT  47660.0 33857.5 47730.0 33992.5 ;
      RECT  47995.0 32307.5 48065.0 32442.5 ;
      RECT  47732.5 33442.5 47802.5 33577.5 ;
      RECT  47922.5 32582.5 47992.5 32717.5 ;
      RECT  48180.0 32482.5 48250.0 32617.5 ;
      RECT  47660.0 33925.0 47730.0 34065.0 ;
      RECT  47995.0 33925.0 48065.0 34065.0 ;
      RECT  47660.0 32235.0 47730.0 32375.0 ;
      RECT  47995.0 32235.0 48065.0 32375.0 ;
      RECT  47475.0 32235.0 47545.0 34065.0 ;
      RECT  48180.0 32235.0 48250.0 34065.0 ;
      RECT  48365.0 32875.0 48435.0 32945.0 ;
      RECT  48437.5 32875.0 48507.5 32945.0 ;
      RECT  48365.0 32375.0 48435.0 32910.0 ;
      RECT  48400.0 32875.0 48472.5 32945.0 ;
      RECT  48437.5 32910.0 48507.5 33442.5 ;
      RECT  48700.0 33287.5 48770.0 33357.5 ;
      RECT  48627.5 33287.5 48697.5 33357.5 ;
      RECT  48700.0 33322.5 48770.0 33925.0 ;
      RECT  48662.5 33287.5 48735.0 33357.5 ;
      RECT  48627.5 32717.5 48697.5 33322.5 ;
      RECT  48365.0 33857.5 48435.0 33992.5 ;
      RECT  48700.0 32307.5 48770.0 32442.5 ;
      RECT  48437.5 33442.5 48507.5 33577.5 ;
      RECT  48627.5 32582.5 48697.5 32717.5 ;
      RECT  48885.0 32482.5 48955.0 32617.5 ;
      RECT  48365.0 33925.0 48435.0 34065.0 ;
      RECT  48700.0 33925.0 48770.0 34065.0 ;
      RECT  48365.0 32235.0 48435.0 32375.0 ;
      RECT  48700.0 32235.0 48770.0 32375.0 ;
      RECT  48180.0 32235.0 48250.0 34065.0 ;
      RECT  48885.0 32235.0 48955.0 34065.0 ;
      RECT  49070.0 32875.0 49140.0 32945.0 ;
      RECT  49142.5 32875.0 49212.5 32945.0 ;
      RECT  49070.0 32375.0 49140.0 32910.0 ;
      RECT  49105.0 32875.0 49177.5 32945.0 ;
      RECT  49142.5 32910.0 49212.5 33442.5 ;
      RECT  49405.0 33287.5 49475.0 33357.5 ;
      RECT  49332.5 33287.5 49402.5 33357.5 ;
      RECT  49405.0 33322.5 49475.0 33925.0 ;
      RECT  49367.5 33287.5 49440.0 33357.5 ;
      RECT  49332.5 32717.5 49402.5 33322.5 ;
      RECT  49070.0 33857.5 49140.0 33992.5 ;
      RECT  49405.0 32307.5 49475.0 32442.5 ;
      RECT  49142.5 33442.5 49212.5 33577.5 ;
      RECT  49332.5 32582.5 49402.5 32717.5 ;
      RECT  49590.0 32482.5 49660.0 32617.5 ;
      RECT  49070.0 33925.0 49140.0 34065.0 ;
      RECT  49405.0 33925.0 49475.0 34065.0 ;
      RECT  49070.0 32235.0 49140.0 32375.0 ;
      RECT  49405.0 32235.0 49475.0 32375.0 ;
      RECT  48885.0 32235.0 48955.0 34065.0 ;
      RECT  49590.0 32235.0 49660.0 34065.0 ;
      RECT  49775.0 32875.0 49845.0 32945.0 ;
      RECT  49847.5 32875.0 49917.5 32945.0 ;
      RECT  49775.0 32375.0 49845.0 32910.0 ;
      RECT  49810.0 32875.0 49882.5 32945.0 ;
      RECT  49847.5 32910.0 49917.5 33442.5 ;
      RECT  50110.0 33287.5 50180.0 33357.5 ;
      RECT  50037.5 33287.5 50107.5 33357.5 ;
      RECT  50110.0 33322.5 50180.0 33925.0 ;
      RECT  50072.5 33287.5 50145.0 33357.5 ;
      RECT  50037.5 32717.5 50107.5 33322.5 ;
      RECT  49775.0 33857.5 49845.0 33992.5 ;
      RECT  50110.0 32307.5 50180.0 32442.5 ;
      RECT  49847.5 33442.5 49917.5 33577.5 ;
      RECT  50037.5 32582.5 50107.5 32717.5 ;
      RECT  50295.0 32482.5 50365.0 32617.5 ;
      RECT  49775.0 33925.0 49845.0 34065.0 ;
      RECT  50110.0 33925.0 50180.0 34065.0 ;
      RECT  49775.0 32235.0 49845.0 32375.0 ;
      RECT  50110.0 32235.0 50180.0 32375.0 ;
      RECT  49590.0 32235.0 49660.0 34065.0 ;
      RECT  50295.0 32235.0 50365.0 34065.0 ;
      RECT  50480.0 32875.0 50550.0 32945.0 ;
      RECT  50552.5 32875.0 50622.5 32945.0 ;
      RECT  50480.0 32375.0 50550.0 32910.0 ;
      RECT  50515.0 32875.0 50587.5 32945.0 ;
      RECT  50552.5 32910.0 50622.5 33442.5 ;
      RECT  50815.0 33287.5 50885.0 33357.5 ;
      RECT  50742.5 33287.5 50812.5 33357.5 ;
      RECT  50815.0 33322.5 50885.0 33925.0 ;
      RECT  50777.5 33287.5 50850.0 33357.5 ;
      RECT  50742.5 32717.5 50812.5 33322.5 ;
      RECT  50480.0 33857.5 50550.0 33992.5 ;
      RECT  50815.0 32307.5 50885.0 32442.5 ;
      RECT  50552.5 33442.5 50622.5 33577.5 ;
      RECT  50742.5 32582.5 50812.5 32717.5 ;
      RECT  51000.0 32482.5 51070.0 32617.5 ;
      RECT  50480.0 33925.0 50550.0 34065.0 ;
      RECT  50815.0 33925.0 50885.0 34065.0 ;
      RECT  50480.0 32235.0 50550.0 32375.0 ;
      RECT  50815.0 32235.0 50885.0 32375.0 ;
      RECT  50295.0 32235.0 50365.0 34065.0 ;
      RECT  51000.0 32235.0 51070.0 34065.0 ;
      RECT  51185.0 32875.0 51255.0 32945.0 ;
      RECT  51257.5 32875.0 51327.5 32945.0 ;
      RECT  51185.0 32375.0 51255.0 32910.0 ;
      RECT  51220.0 32875.0 51292.5 32945.0 ;
      RECT  51257.5 32910.0 51327.5 33442.5 ;
      RECT  51520.0 33287.5 51590.0 33357.5 ;
      RECT  51447.5 33287.5 51517.5 33357.5 ;
      RECT  51520.0 33322.5 51590.0 33925.0 ;
      RECT  51482.5 33287.5 51555.0 33357.5 ;
      RECT  51447.5 32717.5 51517.5 33322.5 ;
      RECT  51185.0 33857.5 51255.0 33992.5 ;
      RECT  51520.0 32307.5 51590.0 32442.5 ;
      RECT  51257.5 33442.5 51327.5 33577.5 ;
      RECT  51447.5 32582.5 51517.5 32717.5 ;
      RECT  51705.0 32482.5 51775.0 32617.5 ;
      RECT  51185.0 33925.0 51255.0 34065.0 ;
      RECT  51520.0 33925.0 51590.0 34065.0 ;
      RECT  51185.0 32235.0 51255.0 32375.0 ;
      RECT  51520.0 32235.0 51590.0 32375.0 ;
      RECT  51000.0 32235.0 51070.0 34065.0 ;
      RECT  51705.0 32235.0 51775.0 34065.0 ;
      RECT  51890.0 32875.0 51960.0 32945.0 ;
      RECT  51962.5 32875.0 52032.5 32945.0 ;
      RECT  51890.0 32375.0 51960.0 32910.0 ;
      RECT  51925.0 32875.0 51997.5 32945.0 ;
      RECT  51962.5 32910.0 52032.5 33442.5 ;
      RECT  52225.0 33287.5 52295.0 33357.5 ;
      RECT  52152.5 33287.5 52222.5 33357.5 ;
      RECT  52225.0 33322.5 52295.0 33925.0 ;
      RECT  52187.5 33287.5 52260.0 33357.5 ;
      RECT  52152.5 32717.5 52222.5 33322.5 ;
      RECT  51890.0 33857.5 51960.0 33992.5 ;
      RECT  52225.0 32307.5 52295.0 32442.5 ;
      RECT  51962.5 33442.5 52032.5 33577.5 ;
      RECT  52152.5 32582.5 52222.5 32717.5 ;
      RECT  52410.0 32482.5 52480.0 32617.5 ;
      RECT  51890.0 33925.0 51960.0 34065.0 ;
      RECT  52225.0 33925.0 52295.0 34065.0 ;
      RECT  51890.0 32235.0 51960.0 32375.0 ;
      RECT  52225.0 32235.0 52295.0 32375.0 ;
      RECT  51705.0 32235.0 51775.0 34065.0 ;
      RECT  52410.0 32235.0 52480.0 34065.0 ;
      RECT  52595.0 32875.0 52665.0 32945.0 ;
      RECT  52667.5 32875.0 52737.5 32945.0 ;
      RECT  52595.0 32375.0 52665.0 32910.0 ;
      RECT  52630.0 32875.0 52702.5 32945.0 ;
      RECT  52667.5 32910.0 52737.5 33442.5 ;
      RECT  52930.0 33287.5 53000.0 33357.5 ;
      RECT  52857.5 33287.5 52927.5 33357.5 ;
      RECT  52930.0 33322.5 53000.0 33925.0 ;
      RECT  52892.5 33287.5 52965.0 33357.5 ;
      RECT  52857.5 32717.5 52927.5 33322.5 ;
      RECT  52595.0 33857.5 52665.0 33992.5 ;
      RECT  52930.0 32307.5 53000.0 32442.5 ;
      RECT  52667.5 33442.5 52737.5 33577.5 ;
      RECT  52857.5 32582.5 52927.5 32717.5 ;
      RECT  53115.0 32482.5 53185.0 32617.5 ;
      RECT  52595.0 33925.0 52665.0 34065.0 ;
      RECT  52930.0 33925.0 53000.0 34065.0 ;
      RECT  52595.0 32235.0 52665.0 32375.0 ;
      RECT  52930.0 32235.0 53000.0 32375.0 ;
      RECT  52410.0 32235.0 52480.0 34065.0 ;
      RECT  53115.0 32235.0 53185.0 34065.0 ;
      RECT  53300.0 32875.0 53370.0 32945.0 ;
      RECT  53372.5 32875.0 53442.5 32945.0 ;
      RECT  53300.0 32375.0 53370.0 32910.0 ;
      RECT  53335.0 32875.0 53407.5 32945.0 ;
      RECT  53372.5 32910.0 53442.5 33442.5 ;
      RECT  53635.0 33287.5 53705.0 33357.5 ;
      RECT  53562.5 33287.5 53632.5 33357.5 ;
      RECT  53635.0 33322.5 53705.0 33925.0 ;
      RECT  53597.5 33287.5 53670.0 33357.5 ;
      RECT  53562.5 32717.5 53632.5 33322.5 ;
      RECT  53300.0 33857.5 53370.0 33992.5 ;
      RECT  53635.0 32307.5 53705.0 32442.5 ;
      RECT  53372.5 33442.5 53442.5 33577.5 ;
      RECT  53562.5 32582.5 53632.5 32717.5 ;
      RECT  53820.0 32482.5 53890.0 32617.5 ;
      RECT  53300.0 33925.0 53370.0 34065.0 ;
      RECT  53635.0 33925.0 53705.0 34065.0 ;
      RECT  53300.0 32235.0 53370.0 32375.0 ;
      RECT  53635.0 32235.0 53705.0 32375.0 ;
      RECT  53115.0 32235.0 53185.0 34065.0 ;
      RECT  53820.0 32235.0 53890.0 34065.0 ;
      RECT  54005.0 32875.0 54075.0 32945.0 ;
      RECT  54077.5 32875.0 54147.5 32945.0 ;
      RECT  54005.0 32375.0 54075.0 32910.0 ;
      RECT  54040.0 32875.0 54112.5 32945.0 ;
      RECT  54077.5 32910.0 54147.5 33442.5 ;
      RECT  54340.0 33287.5 54410.0 33357.5 ;
      RECT  54267.5 33287.5 54337.5 33357.5 ;
      RECT  54340.0 33322.5 54410.0 33925.0 ;
      RECT  54302.5 33287.5 54375.0 33357.5 ;
      RECT  54267.5 32717.5 54337.5 33322.5 ;
      RECT  54005.0 33857.5 54075.0 33992.5 ;
      RECT  54340.0 32307.5 54410.0 32442.5 ;
      RECT  54077.5 33442.5 54147.5 33577.5 ;
      RECT  54267.5 32582.5 54337.5 32717.5 ;
      RECT  54525.0 32482.5 54595.0 32617.5 ;
      RECT  54005.0 33925.0 54075.0 34065.0 ;
      RECT  54340.0 33925.0 54410.0 34065.0 ;
      RECT  54005.0 32235.0 54075.0 32375.0 ;
      RECT  54340.0 32235.0 54410.0 32375.0 ;
      RECT  53820.0 32235.0 53890.0 34065.0 ;
      RECT  54525.0 32235.0 54595.0 34065.0 ;
      RECT  54710.0 32875.0 54780.0 32945.0 ;
      RECT  54782.5 32875.0 54852.5 32945.0 ;
      RECT  54710.0 32375.0 54780.0 32910.0 ;
      RECT  54745.0 32875.0 54817.5 32945.0 ;
      RECT  54782.5 32910.0 54852.5 33442.5 ;
      RECT  55045.0 33287.5 55115.0 33357.5 ;
      RECT  54972.5 33287.5 55042.5 33357.5 ;
      RECT  55045.0 33322.5 55115.0 33925.0 ;
      RECT  55007.5 33287.5 55080.0 33357.5 ;
      RECT  54972.5 32717.5 55042.5 33322.5 ;
      RECT  54710.0 33857.5 54780.0 33992.5 ;
      RECT  55045.0 32307.5 55115.0 32442.5 ;
      RECT  54782.5 33442.5 54852.5 33577.5 ;
      RECT  54972.5 32582.5 55042.5 32717.5 ;
      RECT  55230.0 32482.5 55300.0 32617.5 ;
      RECT  54710.0 33925.0 54780.0 34065.0 ;
      RECT  55045.0 33925.0 55115.0 34065.0 ;
      RECT  54710.0 32235.0 54780.0 32375.0 ;
      RECT  55045.0 32235.0 55115.0 32375.0 ;
      RECT  54525.0 32235.0 54595.0 34065.0 ;
      RECT  55230.0 32235.0 55300.0 34065.0 ;
      RECT  55415.0 32875.0 55485.0 32945.0 ;
      RECT  55487.5 32875.0 55557.5 32945.0 ;
      RECT  55415.0 32375.0 55485.0 32910.0 ;
      RECT  55450.0 32875.0 55522.5 32945.0 ;
      RECT  55487.5 32910.0 55557.5 33442.5 ;
      RECT  55750.0 33287.5 55820.0 33357.5 ;
      RECT  55677.5 33287.5 55747.5 33357.5 ;
      RECT  55750.0 33322.5 55820.0 33925.0 ;
      RECT  55712.5 33287.5 55785.0 33357.5 ;
      RECT  55677.5 32717.5 55747.5 33322.5 ;
      RECT  55415.0 33857.5 55485.0 33992.5 ;
      RECT  55750.0 32307.5 55820.0 32442.5 ;
      RECT  55487.5 33442.5 55557.5 33577.5 ;
      RECT  55677.5 32582.5 55747.5 32717.5 ;
      RECT  55935.0 32482.5 56005.0 32617.5 ;
      RECT  55415.0 33925.0 55485.0 34065.0 ;
      RECT  55750.0 33925.0 55820.0 34065.0 ;
      RECT  55415.0 32235.0 55485.0 32375.0 ;
      RECT  55750.0 32235.0 55820.0 32375.0 ;
      RECT  55230.0 32235.0 55300.0 34065.0 ;
      RECT  55935.0 32235.0 56005.0 34065.0 ;
      RECT  56120.0 32875.0 56190.0 32945.0 ;
      RECT  56192.5 32875.0 56262.5 32945.0 ;
      RECT  56120.0 32375.0 56190.0 32910.0 ;
      RECT  56155.0 32875.0 56227.5 32945.0 ;
      RECT  56192.5 32910.0 56262.5 33442.5 ;
      RECT  56455.0 33287.5 56525.0 33357.5 ;
      RECT  56382.5 33287.5 56452.5 33357.5 ;
      RECT  56455.0 33322.5 56525.0 33925.0 ;
      RECT  56417.5 33287.5 56490.0 33357.5 ;
      RECT  56382.5 32717.5 56452.5 33322.5 ;
      RECT  56120.0 33857.5 56190.0 33992.5 ;
      RECT  56455.0 32307.5 56525.0 32442.5 ;
      RECT  56192.5 33442.5 56262.5 33577.5 ;
      RECT  56382.5 32582.5 56452.5 32717.5 ;
      RECT  56640.0 32482.5 56710.0 32617.5 ;
      RECT  56120.0 33925.0 56190.0 34065.0 ;
      RECT  56455.0 33925.0 56525.0 34065.0 ;
      RECT  56120.0 32235.0 56190.0 32375.0 ;
      RECT  56455.0 32235.0 56525.0 32375.0 ;
      RECT  55935.0 32235.0 56005.0 34065.0 ;
      RECT  56640.0 32235.0 56710.0 34065.0 ;
      RECT  56825.0 32875.0 56895.0 32945.0 ;
      RECT  56897.5 32875.0 56967.5 32945.0 ;
      RECT  56825.0 32375.0 56895.0 32910.0 ;
      RECT  56860.0 32875.0 56932.5 32945.0 ;
      RECT  56897.5 32910.0 56967.5 33442.5 ;
      RECT  57160.0 33287.5 57230.0 33357.5 ;
      RECT  57087.5 33287.5 57157.5 33357.5 ;
      RECT  57160.0 33322.5 57230.0 33925.0 ;
      RECT  57122.5 33287.5 57195.0 33357.5 ;
      RECT  57087.5 32717.5 57157.5 33322.5 ;
      RECT  56825.0 33857.5 56895.0 33992.5 ;
      RECT  57160.0 32307.5 57230.0 32442.5 ;
      RECT  56897.5 33442.5 56967.5 33577.5 ;
      RECT  57087.5 32582.5 57157.5 32717.5 ;
      RECT  57345.0 32482.5 57415.0 32617.5 ;
      RECT  56825.0 33925.0 56895.0 34065.0 ;
      RECT  57160.0 33925.0 57230.0 34065.0 ;
      RECT  56825.0 32235.0 56895.0 32375.0 ;
      RECT  57160.0 32235.0 57230.0 32375.0 ;
      RECT  56640.0 32235.0 56710.0 34065.0 ;
      RECT  57345.0 32235.0 57415.0 34065.0 ;
      RECT  57530.0 32875.0 57600.0 32945.0 ;
      RECT  57602.5 32875.0 57672.5 32945.0 ;
      RECT  57530.0 32375.0 57600.0 32910.0 ;
      RECT  57565.0 32875.0 57637.5 32945.0 ;
      RECT  57602.5 32910.0 57672.5 33442.5 ;
      RECT  57865.0 33287.5 57935.0 33357.5 ;
      RECT  57792.5 33287.5 57862.5 33357.5 ;
      RECT  57865.0 33322.5 57935.0 33925.0 ;
      RECT  57827.5 33287.5 57900.0 33357.5 ;
      RECT  57792.5 32717.5 57862.5 33322.5 ;
      RECT  57530.0 33857.5 57600.0 33992.5 ;
      RECT  57865.0 32307.5 57935.0 32442.5 ;
      RECT  57602.5 33442.5 57672.5 33577.5 ;
      RECT  57792.5 32582.5 57862.5 32717.5 ;
      RECT  58050.0 32482.5 58120.0 32617.5 ;
      RECT  57530.0 33925.0 57600.0 34065.0 ;
      RECT  57865.0 33925.0 57935.0 34065.0 ;
      RECT  57530.0 32235.0 57600.0 32375.0 ;
      RECT  57865.0 32235.0 57935.0 32375.0 ;
      RECT  57345.0 32235.0 57415.0 34065.0 ;
      RECT  58050.0 32235.0 58120.0 34065.0 ;
      RECT  58235.0 32875.0 58305.0 32945.0 ;
      RECT  58307.5 32875.0 58377.5 32945.0 ;
      RECT  58235.0 32375.0 58305.0 32910.0 ;
      RECT  58270.0 32875.0 58342.5 32945.0 ;
      RECT  58307.5 32910.0 58377.5 33442.5 ;
      RECT  58570.0 33287.5 58640.0 33357.5 ;
      RECT  58497.5 33287.5 58567.5 33357.5 ;
      RECT  58570.0 33322.5 58640.0 33925.0 ;
      RECT  58532.5 33287.5 58605.0 33357.5 ;
      RECT  58497.5 32717.5 58567.5 33322.5 ;
      RECT  58235.0 33857.5 58305.0 33992.5 ;
      RECT  58570.0 32307.5 58640.0 32442.5 ;
      RECT  58307.5 33442.5 58377.5 33577.5 ;
      RECT  58497.5 32582.5 58567.5 32717.5 ;
      RECT  58755.0 32482.5 58825.0 32617.5 ;
      RECT  58235.0 33925.0 58305.0 34065.0 ;
      RECT  58570.0 33925.0 58640.0 34065.0 ;
      RECT  58235.0 32235.0 58305.0 32375.0 ;
      RECT  58570.0 32235.0 58640.0 32375.0 ;
      RECT  58050.0 32235.0 58120.0 34065.0 ;
      RECT  58755.0 32235.0 58825.0 34065.0 ;
      RECT  58940.0 32875.0 59010.0 32945.0 ;
      RECT  59012.5 32875.0 59082.5 32945.0 ;
      RECT  58940.0 32375.0 59010.0 32910.0 ;
      RECT  58975.0 32875.0 59047.5 32945.0 ;
      RECT  59012.5 32910.0 59082.5 33442.5 ;
      RECT  59275.0 33287.5 59345.0 33357.5 ;
      RECT  59202.5 33287.5 59272.5 33357.5 ;
      RECT  59275.0 33322.5 59345.0 33925.0 ;
      RECT  59237.5 33287.5 59310.0 33357.5 ;
      RECT  59202.5 32717.5 59272.5 33322.5 ;
      RECT  58940.0 33857.5 59010.0 33992.5 ;
      RECT  59275.0 32307.5 59345.0 32442.5 ;
      RECT  59012.5 33442.5 59082.5 33577.5 ;
      RECT  59202.5 32582.5 59272.5 32717.5 ;
      RECT  59460.0 32482.5 59530.0 32617.5 ;
      RECT  58940.0 33925.0 59010.0 34065.0 ;
      RECT  59275.0 33925.0 59345.0 34065.0 ;
      RECT  58940.0 32235.0 59010.0 32375.0 ;
      RECT  59275.0 32235.0 59345.0 32375.0 ;
      RECT  58755.0 32235.0 58825.0 34065.0 ;
      RECT  59460.0 32235.0 59530.0 34065.0 ;
      RECT  59645.0 32875.0 59715.0 32945.0 ;
      RECT  59717.5 32875.0 59787.5 32945.0 ;
      RECT  59645.0 32375.0 59715.0 32910.0 ;
      RECT  59680.0 32875.0 59752.5 32945.0 ;
      RECT  59717.5 32910.0 59787.5 33442.5 ;
      RECT  59980.0 33287.5 60050.0 33357.5 ;
      RECT  59907.5 33287.5 59977.5 33357.5 ;
      RECT  59980.0 33322.5 60050.0 33925.0 ;
      RECT  59942.5 33287.5 60015.0 33357.5 ;
      RECT  59907.5 32717.5 59977.5 33322.5 ;
      RECT  59645.0 33857.5 59715.0 33992.5 ;
      RECT  59980.0 32307.5 60050.0 32442.5 ;
      RECT  59717.5 33442.5 59787.5 33577.5 ;
      RECT  59907.5 32582.5 59977.5 32717.5 ;
      RECT  60165.0 32482.5 60235.0 32617.5 ;
      RECT  59645.0 33925.0 59715.0 34065.0 ;
      RECT  59980.0 33925.0 60050.0 34065.0 ;
      RECT  59645.0 32235.0 59715.0 32375.0 ;
      RECT  59980.0 32235.0 60050.0 32375.0 ;
      RECT  59460.0 32235.0 59530.0 34065.0 ;
      RECT  60165.0 32235.0 60235.0 34065.0 ;
      RECT  60350.0 32875.0 60420.0 32945.0 ;
      RECT  60422.5 32875.0 60492.5 32945.0 ;
      RECT  60350.0 32375.0 60420.0 32910.0 ;
      RECT  60385.0 32875.0 60457.5 32945.0 ;
      RECT  60422.5 32910.0 60492.5 33442.5 ;
      RECT  60685.0 33287.5 60755.0 33357.5 ;
      RECT  60612.5 33287.5 60682.5 33357.5 ;
      RECT  60685.0 33322.5 60755.0 33925.0 ;
      RECT  60647.5 33287.5 60720.0 33357.5 ;
      RECT  60612.5 32717.5 60682.5 33322.5 ;
      RECT  60350.0 33857.5 60420.0 33992.5 ;
      RECT  60685.0 32307.5 60755.0 32442.5 ;
      RECT  60422.5 33442.5 60492.5 33577.5 ;
      RECT  60612.5 32582.5 60682.5 32717.5 ;
      RECT  60870.0 32482.5 60940.0 32617.5 ;
      RECT  60350.0 33925.0 60420.0 34065.0 ;
      RECT  60685.0 33925.0 60755.0 34065.0 ;
      RECT  60350.0 32235.0 60420.0 32375.0 ;
      RECT  60685.0 32235.0 60755.0 32375.0 ;
      RECT  60165.0 32235.0 60235.0 34065.0 ;
      RECT  60870.0 32235.0 60940.0 34065.0 ;
      RECT  61055.0 32875.0 61125.0 32945.0 ;
      RECT  61127.5 32875.0 61197.5 32945.0 ;
      RECT  61055.0 32375.0 61125.0 32910.0 ;
      RECT  61090.0 32875.0 61162.5 32945.0 ;
      RECT  61127.5 32910.0 61197.5 33442.5 ;
      RECT  61390.0 33287.5 61460.0 33357.5 ;
      RECT  61317.5 33287.5 61387.5 33357.5 ;
      RECT  61390.0 33322.5 61460.0 33925.0 ;
      RECT  61352.5 33287.5 61425.0 33357.5 ;
      RECT  61317.5 32717.5 61387.5 33322.5 ;
      RECT  61055.0 33857.5 61125.0 33992.5 ;
      RECT  61390.0 32307.5 61460.0 32442.5 ;
      RECT  61127.5 33442.5 61197.5 33577.5 ;
      RECT  61317.5 32582.5 61387.5 32717.5 ;
      RECT  61575.0 32482.5 61645.0 32617.5 ;
      RECT  61055.0 33925.0 61125.0 34065.0 ;
      RECT  61390.0 33925.0 61460.0 34065.0 ;
      RECT  61055.0 32235.0 61125.0 32375.0 ;
      RECT  61390.0 32235.0 61460.0 32375.0 ;
      RECT  60870.0 32235.0 60940.0 34065.0 ;
      RECT  61575.0 32235.0 61645.0 34065.0 ;
      RECT  61760.0 32875.0 61830.0 32945.0 ;
      RECT  61832.5 32875.0 61902.5 32945.0 ;
      RECT  61760.0 32375.0 61830.0 32910.0 ;
      RECT  61795.0 32875.0 61867.5 32945.0 ;
      RECT  61832.5 32910.0 61902.5 33442.5 ;
      RECT  62095.0 33287.5 62165.0 33357.5 ;
      RECT  62022.5 33287.5 62092.5 33357.5 ;
      RECT  62095.0 33322.5 62165.0 33925.0 ;
      RECT  62057.5 33287.5 62130.0 33357.5 ;
      RECT  62022.5 32717.5 62092.5 33322.5 ;
      RECT  61760.0 33857.5 61830.0 33992.5 ;
      RECT  62095.0 32307.5 62165.0 32442.5 ;
      RECT  61832.5 33442.5 61902.5 33577.5 ;
      RECT  62022.5 32582.5 62092.5 32717.5 ;
      RECT  62280.0 32482.5 62350.0 32617.5 ;
      RECT  61760.0 33925.0 61830.0 34065.0 ;
      RECT  62095.0 33925.0 62165.0 34065.0 ;
      RECT  61760.0 32235.0 61830.0 32375.0 ;
      RECT  62095.0 32235.0 62165.0 32375.0 ;
      RECT  61575.0 32235.0 61645.0 34065.0 ;
      RECT  62280.0 32235.0 62350.0 34065.0 ;
      RECT  62465.0 32875.0 62535.0 32945.0 ;
      RECT  62537.5 32875.0 62607.5 32945.0 ;
      RECT  62465.0 32375.0 62535.0 32910.0 ;
      RECT  62500.0 32875.0 62572.5 32945.0 ;
      RECT  62537.5 32910.0 62607.5 33442.5 ;
      RECT  62800.0 33287.5 62870.0 33357.5 ;
      RECT  62727.5 33287.5 62797.5 33357.5 ;
      RECT  62800.0 33322.5 62870.0 33925.0 ;
      RECT  62762.5 33287.5 62835.0 33357.5 ;
      RECT  62727.5 32717.5 62797.5 33322.5 ;
      RECT  62465.0 33857.5 62535.0 33992.5 ;
      RECT  62800.0 32307.5 62870.0 32442.5 ;
      RECT  62537.5 33442.5 62607.5 33577.5 ;
      RECT  62727.5 32582.5 62797.5 32717.5 ;
      RECT  62985.0 32482.5 63055.0 32617.5 ;
      RECT  62465.0 33925.0 62535.0 34065.0 ;
      RECT  62800.0 33925.0 62870.0 34065.0 ;
      RECT  62465.0 32235.0 62535.0 32375.0 ;
      RECT  62800.0 32235.0 62870.0 32375.0 ;
      RECT  62280.0 32235.0 62350.0 34065.0 ;
      RECT  62985.0 32235.0 63055.0 34065.0 ;
      RECT  63170.0 32875.0 63240.0 32945.0 ;
      RECT  63242.5 32875.0 63312.5 32945.0 ;
      RECT  63170.0 32375.0 63240.0 32910.0 ;
      RECT  63205.0 32875.0 63277.5 32945.0 ;
      RECT  63242.5 32910.0 63312.5 33442.5 ;
      RECT  63505.0 33287.5 63575.0 33357.5 ;
      RECT  63432.5 33287.5 63502.5 33357.5 ;
      RECT  63505.0 33322.5 63575.0 33925.0 ;
      RECT  63467.5 33287.5 63540.0 33357.5 ;
      RECT  63432.5 32717.5 63502.5 33322.5 ;
      RECT  63170.0 33857.5 63240.0 33992.5 ;
      RECT  63505.0 32307.5 63575.0 32442.5 ;
      RECT  63242.5 33442.5 63312.5 33577.5 ;
      RECT  63432.5 32582.5 63502.5 32717.5 ;
      RECT  63690.0 32482.5 63760.0 32617.5 ;
      RECT  63170.0 33925.0 63240.0 34065.0 ;
      RECT  63505.0 33925.0 63575.0 34065.0 ;
      RECT  63170.0 32235.0 63240.0 32375.0 ;
      RECT  63505.0 32235.0 63575.0 32375.0 ;
      RECT  62985.0 32235.0 63055.0 34065.0 ;
      RECT  63690.0 32235.0 63760.0 34065.0 ;
      RECT  63875.0 32875.0 63945.0 32945.0 ;
      RECT  63947.5 32875.0 64017.5 32945.0 ;
      RECT  63875.0 32375.0 63945.0 32910.0 ;
      RECT  63910.0 32875.0 63982.5 32945.0 ;
      RECT  63947.5 32910.0 64017.5 33442.5 ;
      RECT  64210.0 33287.5 64280.0 33357.5 ;
      RECT  64137.5 33287.5 64207.5 33357.5 ;
      RECT  64210.0 33322.5 64280.0 33925.0 ;
      RECT  64172.5 33287.5 64245.0 33357.5 ;
      RECT  64137.5 32717.5 64207.5 33322.5 ;
      RECT  63875.0 33857.5 63945.0 33992.5 ;
      RECT  64210.0 32307.5 64280.0 32442.5 ;
      RECT  63947.5 33442.5 64017.5 33577.5 ;
      RECT  64137.5 32582.5 64207.5 32717.5 ;
      RECT  64395.0 32482.5 64465.0 32617.5 ;
      RECT  63875.0 33925.0 63945.0 34065.0 ;
      RECT  64210.0 33925.0 64280.0 34065.0 ;
      RECT  63875.0 32235.0 63945.0 32375.0 ;
      RECT  64210.0 32235.0 64280.0 32375.0 ;
      RECT  63690.0 32235.0 63760.0 34065.0 ;
      RECT  64395.0 32235.0 64465.0 34065.0 ;
      RECT  64580.0 32875.0 64650.0 32945.0 ;
      RECT  64652.5 32875.0 64722.5 32945.0 ;
      RECT  64580.0 32375.0 64650.0 32910.0 ;
      RECT  64615.0 32875.0 64687.5 32945.0 ;
      RECT  64652.5 32910.0 64722.5 33442.5 ;
      RECT  64915.0 33287.5 64985.0 33357.5 ;
      RECT  64842.5 33287.5 64912.5 33357.5 ;
      RECT  64915.0 33322.5 64985.0 33925.0 ;
      RECT  64877.5 33287.5 64950.0 33357.5 ;
      RECT  64842.5 32717.5 64912.5 33322.5 ;
      RECT  64580.0 33857.5 64650.0 33992.5 ;
      RECT  64915.0 32307.5 64985.0 32442.5 ;
      RECT  64652.5 33442.5 64722.5 33577.5 ;
      RECT  64842.5 32582.5 64912.5 32717.5 ;
      RECT  65100.0 32482.5 65170.0 32617.5 ;
      RECT  64580.0 33925.0 64650.0 34065.0 ;
      RECT  64915.0 33925.0 64985.0 34065.0 ;
      RECT  64580.0 32235.0 64650.0 32375.0 ;
      RECT  64915.0 32235.0 64985.0 32375.0 ;
      RECT  64395.0 32235.0 64465.0 34065.0 ;
      RECT  65100.0 32235.0 65170.0 34065.0 ;
      RECT  65285.0 32875.0 65355.0 32945.0 ;
      RECT  65357.5 32875.0 65427.5 32945.0 ;
      RECT  65285.0 32375.0 65355.0 32910.0 ;
      RECT  65320.0 32875.0 65392.5 32945.0 ;
      RECT  65357.5 32910.0 65427.5 33442.5 ;
      RECT  65620.0 33287.5 65690.0 33357.5 ;
      RECT  65547.5 33287.5 65617.5 33357.5 ;
      RECT  65620.0 33322.5 65690.0 33925.0 ;
      RECT  65582.5 33287.5 65655.0 33357.5 ;
      RECT  65547.5 32717.5 65617.5 33322.5 ;
      RECT  65285.0 33857.5 65355.0 33992.5 ;
      RECT  65620.0 32307.5 65690.0 32442.5 ;
      RECT  65357.5 33442.5 65427.5 33577.5 ;
      RECT  65547.5 32582.5 65617.5 32717.5 ;
      RECT  65805.0 32482.5 65875.0 32617.5 ;
      RECT  65285.0 33925.0 65355.0 34065.0 ;
      RECT  65620.0 33925.0 65690.0 34065.0 ;
      RECT  65285.0 32235.0 65355.0 32375.0 ;
      RECT  65620.0 32235.0 65690.0 32375.0 ;
      RECT  65100.0 32235.0 65170.0 34065.0 ;
      RECT  65805.0 32235.0 65875.0 34065.0 ;
      RECT  65990.0 32875.0 66060.0 32945.0 ;
      RECT  66062.5 32875.0 66132.5 32945.0 ;
      RECT  65990.0 32375.0 66060.0 32910.0 ;
      RECT  66025.0 32875.0 66097.5 32945.0 ;
      RECT  66062.5 32910.0 66132.5 33442.5 ;
      RECT  66325.0 33287.5 66395.0 33357.5 ;
      RECT  66252.5 33287.5 66322.5 33357.5 ;
      RECT  66325.0 33322.5 66395.0 33925.0 ;
      RECT  66287.5 33287.5 66360.0 33357.5 ;
      RECT  66252.5 32717.5 66322.5 33322.5 ;
      RECT  65990.0 33857.5 66060.0 33992.5 ;
      RECT  66325.0 32307.5 66395.0 32442.5 ;
      RECT  66062.5 33442.5 66132.5 33577.5 ;
      RECT  66252.5 32582.5 66322.5 32717.5 ;
      RECT  66510.0 32482.5 66580.0 32617.5 ;
      RECT  65990.0 33925.0 66060.0 34065.0 ;
      RECT  66325.0 33925.0 66395.0 34065.0 ;
      RECT  65990.0 32235.0 66060.0 32375.0 ;
      RECT  66325.0 32235.0 66395.0 32375.0 ;
      RECT  65805.0 32235.0 65875.0 34065.0 ;
      RECT  66510.0 32235.0 66580.0 34065.0 ;
      RECT  66695.0 32875.0 66765.0 32945.0 ;
      RECT  66767.5 32875.0 66837.5 32945.0 ;
      RECT  66695.0 32375.0 66765.0 32910.0 ;
      RECT  66730.0 32875.0 66802.5 32945.0 ;
      RECT  66767.5 32910.0 66837.5 33442.5 ;
      RECT  67030.0 33287.5 67100.0 33357.5 ;
      RECT  66957.5 33287.5 67027.5 33357.5 ;
      RECT  67030.0 33322.5 67100.0 33925.0 ;
      RECT  66992.5 33287.5 67065.0 33357.5 ;
      RECT  66957.5 32717.5 67027.5 33322.5 ;
      RECT  66695.0 33857.5 66765.0 33992.5 ;
      RECT  67030.0 32307.5 67100.0 32442.5 ;
      RECT  66767.5 33442.5 66837.5 33577.5 ;
      RECT  66957.5 32582.5 67027.5 32717.5 ;
      RECT  67215.0 32482.5 67285.0 32617.5 ;
      RECT  66695.0 33925.0 66765.0 34065.0 ;
      RECT  67030.0 33925.0 67100.0 34065.0 ;
      RECT  66695.0 32235.0 66765.0 32375.0 ;
      RECT  67030.0 32235.0 67100.0 32375.0 ;
      RECT  66510.0 32235.0 66580.0 34065.0 ;
      RECT  67215.0 32235.0 67285.0 34065.0 ;
      RECT  67400.0 32875.0 67470.0 32945.0 ;
      RECT  67472.5 32875.0 67542.5 32945.0 ;
      RECT  67400.0 32375.0 67470.0 32910.0 ;
      RECT  67435.0 32875.0 67507.5 32945.0 ;
      RECT  67472.5 32910.0 67542.5 33442.5 ;
      RECT  67735.0 33287.5 67805.0 33357.5 ;
      RECT  67662.5 33287.5 67732.5 33357.5 ;
      RECT  67735.0 33322.5 67805.0 33925.0 ;
      RECT  67697.5 33287.5 67770.0 33357.5 ;
      RECT  67662.5 32717.5 67732.5 33322.5 ;
      RECT  67400.0 33857.5 67470.0 33992.5 ;
      RECT  67735.0 32307.5 67805.0 32442.5 ;
      RECT  67472.5 33442.5 67542.5 33577.5 ;
      RECT  67662.5 32582.5 67732.5 32717.5 ;
      RECT  67920.0 32482.5 67990.0 32617.5 ;
      RECT  67400.0 33925.0 67470.0 34065.0 ;
      RECT  67735.0 33925.0 67805.0 34065.0 ;
      RECT  67400.0 32235.0 67470.0 32375.0 ;
      RECT  67735.0 32235.0 67805.0 32375.0 ;
      RECT  67215.0 32235.0 67285.0 34065.0 ;
      RECT  67920.0 32235.0 67990.0 34065.0 ;
      RECT  68105.0 32875.0 68175.0 32945.0 ;
      RECT  68177.5 32875.0 68247.5 32945.0 ;
      RECT  68105.0 32375.0 68175.0 32910.0 ;
      RECT  68140.0 32875.0 68212.5 32945.0 ;
      RECT  68177.5 32910.0 68247.5 33442.5 ;
      RECT  68440.0 33287.5 68510.0 33357.5 ;
      RECT  68367.5 33287.5 68437.5 33357.5 ;
      RECT  68440.0 33322.5 68510.0 33925.0 ;
      RECT  68402.5 33287.5 68475.0 33357.5 ;
      RECT  68367.5 32717.5 68437.5 33322.5 ;
      RECT  68105.0 33857.5 68175.0 33992.5 ;
      RECT  68440.0 32307.5 68510.0 32442.5 ;
      RECT  68177.5 33442.5 68247.5 33577.5 ;
      RECT  68367.5 32582.5 68437.5 32717.5 ;
      RECT  68625.0 32482.5 68695.0 32617.5 ;
      RECT  68105.0 33925.0 68175.0 34065.0 ;
      RECT  68440.0 33925.0 68510.0 34065.0 ;
      RECT  68105.0 32235.0 68175.0 32375.0 ;
      RECT  68440.0 32235.0 68510.0 32375.0 ;
      RECT  67920.0 32235.0 67990.0 34065.0 ;
      RECT  68625.0 32235.0 68695.0 34065.0 ;
      RECT  68810.0 32875.0 68880.0 32945.0 ;
      RECT  68882.5 32875.0 68952.5 32945.0 ;
      RECT  68810.0 32375.0 68880.0 32910.0 ;
      RECT  68845.0 32875.0 68917.5 32945.0 ;
      RECT  68882.5 32910.0 68952.5 33442.5 ;
      RECT  69145.0 33287.5 69215.0 33357.5 ;
      RECT  69072.5 33287.5 69142.5 33357.5 ;
      RECT  69145.0 33322.5 69215.0 33925.0 ;
      RECT  69107.5 33287.5 69180.0 33357.5 ;
      RECT  69072.5 32717.5 69142.5 33322.5 ;
      RECT  68810.0 33857.5 68880.0 33992.5 ;
      RECT  69145.0 32307.5 69215.0 32442.5 ;
      RECT  68882.5 33442.5 68952.5 33577.5 ;
      RECT  69072.5 32582.5 69142.5 32717.5 ;
      RECT  69330.0 32482.5 69400.0 32617.5 ;
      RECT  68810.0 33925.0 68880.0 34065.0 ;
      RECT  69145.0 33925.0 69215.0 34065.0 ;
      RECT  68810.0 32235.0 68880.0 32375.0 ;
      RECT  69145.0 32235.0 69215.0 32375.0 ;
      RECT  68625.0 32235.0 68695.0 34065.0 ;
      RECT  69330.0 32235.0 69400.0 34065.0 ;
      RECT  69515.0 32875.0 69585.0 32945.0 ;
      RECT  69587.5 32875.0 69657.5 32945.0 ;
      RECT  69515.0 32375.0 69585.0 32910.0 ;
      RECT  69550.0 32875.0 69622.5 32945.0 ;
      RECT  69587.5 32910.0 69657.5 33442.5 ;
      RECT  69850.0 33287.5 69920.0 33357.5 ;
      RECT  69777.5 33287.5 69847.5 33357.5 ;
      RECT  69850.0 33322.5 69920.0 33925.0 ;
      RECT  69812.5 33287.5 69885.0 33357.5 ;
      RECT  69777.5 32717.5 69847.5 33322.5 ;
      RECT  69515.0 33857.5 69585.0 33992.5 ;
      RECT  69850.0 32307.5 69920.0 32442.5 ;
      RECT  69587.5 33442.5 69657.5 33577.5 ;
      RECT  69777.5 32582.5 69847.5 32717.5 ;
      RECT  70035.0 32482.5 70105.0 32617.5 ;
      RECT  69515.0 33925.0 69585.0 34065.0 ;
      RECT  69850.0 33925.0 69920.0 34065.0 ;
      RECT  69515.0 32235.0 69585.0 32375.0 ;
      RECT  69850.0 32235.0 69920.0 32375.0 ;
      RECT  69330.0 32235.0 69400.0 34065.0 ;
      RECT  70035.0 32235.0 70105.0 34065.0 ;
      RECT  70220.0 32875.0 70290.0 32945.0 ;
      RECT  70292.5 32875.0 70362.5 32945.0 ;
      RECT  70220.0 32375.0 70290.0 32910.0 ;
      RECT  70255.0 32875.0 70327.5 32945.0 ;
      RECT  70292.5 32910.0 70362.5 33442.5 ;
      RECT  70555.0 33287.5 70625.0 33357.5 ;
      RECT  70482.5 33287.5 70552.5 33357.5 ;
      RECT  70555.0 33322.5 70625.0 33925.0 ;
      RECT  70517.5 33287.5 70590.0 33357.5 ;
      RECT  70482.5 32717.5 70552.5 33322.5 ;
      RECT  70220.0 33857.5 70290.0 33992.5 ;
      RECT  70555.0 32307.5 70625.0 32442.5 ;
      RECT  70292.5 33442.5 70362.5 33577.5 ;
      RECT  70482.5 32582.5 70552.5 32717.5 ;
      RECT  70740.0 32482.5 70810.0 32617.5 ;
      RECT  70220.0 33925.0 70290.0 34065.0 ;
      RECT  70555.0 33925.0 70625.0 34065.0 ;
      RECT  70220.0 32235.0 70290.0 32375.0 ;
      RECT  70555.0 32235.0 70625.0 32375.0 ;
      RECT  70035.0 32235.0 70105.0 34065.0 ;
      RECT  70740.0 32235.0 70810.0 34065.0 ;
      RECT  70925.0 32875.0 70995.0 32945.0 ;
      RECT  70997.5 32875.0 71067.5 32945.0 ;
      RECT  70925.0 32375.0 70995.0 32910.0 ;
      RECT  70960.0 32875.0 71032.5 32945.0 ;
      RECT  70997.5 32910.0 71067.5 33442.5 ;
      RECT  71260.0 33287.5 71330.0 33357.5 ;
      RECT  71187.5 33287.5 71257.5 33357.5 ;
      RECT  71260.0 33322.5 71330.0 33925.0 ;
      RECT  71222.5 33287.5 71295.0 33357.5 ;
      RECT  71187.5 32717.5 71257.5 33322.5 ;
      RECT  70925.0 33857.5 70995.0 33992.5 ;
      RECT  71260.0 32307.5 71330.0 32442.5 ;
      RECT  70997.5 33442.5 71067.5 33577.5 ;
      RECT  71187.5 32582.5 71257.5 32717.5 ;
      RECT  71445.0 32482.5 71515.0 32617.5 ;
      RECT  70925.0 33925.0 70995.0 34065.0 ;
      RECT  71260.0 33925.0 71330.0 34065.0 ;
      RECT  70925.0 32235.0 70995.0 32375.0 ;
      RECT  71260.0 32235.0 71330.0 32375.0 ;
      RECT  70740.0 32235.0 70810.0 34065.0 ;
      RECT  71445.0 32235.0 71515.0 34065.0 ;
      RECT  71630.0 32875.0 71700.0 32945.0 ;
      RECT  71702.5 32875.0 71772.5 32945.0 ;
      RECT  71630.0 32375.0 71700.0 32910.0 ;
      RECT  71665.0 32875.0 71737.5 32945.0 ;
      RECT  71702.5 32910.0 71772.5 33442.5 ;
      RECT  71965.0 33287.5 72035.0 33357.5 ;
      RECT  71892.5 33287.5 71962.5 33357.5 ;
      RECT  71965.0 33322.5 72035.0 33925.0 ;
      RECT  71927.5 33287.5 72000.0 33357.5 ;
      RECT  71892.5 32717.5 71962.5 33322.5 ;
      RECT  71630.0 33857.5 71700.0 33992.5 ;
      RECT  71965.0 32307.5 72035.0 32442.5 ;
      RECT  71702.5 33442.5 71772.5 33577.5 ;
      RECT  71892.5 32582.5 71962.5 32717.5 ;
      RECT  72150.0 32482.5 72220.0 32617.5 ;
      RECT  71630.0 33925.0 71700.0 34065.0 ;
      RECT  71965.0 33925.0 72035.0 34065.0 ;
      RECT  71630.0 32235.0 71700.0 32375.0 ;
      RECT  71965.0 32235.0 72035.0 32375.0 ;
      RECT  71445.0 32235.0 71515.0 34065.0 ;
      RECT  72150.0 32235.0 72220.0 34065.0 ;
      RECT  72335.0 32875.0 72405.0 32945.0 ;
      RECT  72407.5 32875.0 72477.5 32945.0 ;
      RECT  72335.0 32375.0 72405.0 32910.0 ;
      RECT  72370.0 32875.0 72442.5 32945.0 ;
      RECT  72407.5 32910.0 72477.5 33442.5 ;
      RECT  72670.0 33287.5 72740.0 33357.5 ;
      RECT  72597.5 33287.5 72667.5 33357.5 ;
      RECT  72670.0 33322.5 72740.0 33925.0 ;
      RECT  72632.5 33287.5 72705.0 33357.5 ;
      RECT  72597.5 32717.5 72667.5 33322.5 ;
      RECT  72335.0 33857.5 72405.0 33992.5 ;
      RECT  72670.0 32307.5 72740.0 32442.5 ;
      RECT  72407.5 33442.5 72477.5 33577.5 ;
      RECT  72597.5 32582.5 72667.5 32717.5 ;
      RECT  72855.0 32482.5 72925.0 32617.5 ;
      RECT  72335.0 33925.0 72405.0 34065.0 ;
      RECT  72670.0 33925.0 72740.0 34065.0 ;
      RECT  72335.0 32235.0 72405.0 32375.0 ;
      RECT  72670.0 32235.0 72740.0 32375.0 ;
      RECT  72150.0 32235.0 72220.0 34065.0 ;
      RECT  72855.0 32235.0 72925.0 34065.0 ;
      RECT  73040.0 32875.0 73110.0 32945.0 ;
      RECT  73112.5 32875.0 73182.5 32945.0 ;
      RECT  73040.0 32375.0 73110.0 32910.0 ;
      RECT  73075.0 32875.0 73147.5 32945.0 ;
      RECT  73112.5 32910.0 73182.5 33442.5 ;
      RECT  73375.0 33287.5 73445.0 33357.5 ;
      RECT  73302.5 33287.5 73372.5 33357.5 ;
      RECT  73375.0 33322.5 73445.0 33925.0 ;
      RECT  73337.5 33287.5 73410.0 33357.5 ;
      RECT  73302.5 32717.5 73372.5 33322.5 ;
      RECT  73040.0 33857.5 73110.0 33992.5 ;
      RECT  73375.0 32307.5 73445.0 32442.5 ;
      RECT  73112.5 33442.5 73182.5 33577.5 ;
      RECT  73302.5 32582.5 73372.5 32717.5 ;
      RECT  73560.0 32482.5 73630.0 32617.5 ;
      RECT  73040.0 33925.0 73110.0 34065.0 ;
      RECT  73375.0 33925.0 73445.0 34065.0 ;
      RECT  73040.0 32235.0 73110.0 32375.0 ;
      RECT  73375.0 32235.0 73445.0 32375.0 ;
      RECT  72855.0 32235.0 72925.0 34065.0 ;
      RECT  73560.0 32235.0 73630.0 34065.0 ;
      RECT  73745.0 32875.0 73815.0 32945.0 ;
      RECT  73817.5 32875.0 73887.5 32945.0 ;
      RECT  73745.0 32375.0 73815.0 32910.0 ;
      RECT  73780.0 32875.0 73852.5 32945.0 ;
      RECT  73817.5 32910.0 73887.5 33442.5 ;
      RECT  74080.0 33287.5 74150.0 33357.5 ;
      RECT  74007.5 33287.5 74077.5 33357.5 ;
      RECT  74080.0 33322.5 74150.0 33925.0 ;
      RECT  74042.5 33287.5 74115.0 33357.5 ;
      RECT  74007.5 32717.5 74077.5 33322.5 ;
      RECT  73745.0 33857.5 73815.0 33992.5 ;
      RECT  74080.0 32307.5 74150.0 32442.5 ;
      RECT  73817.5 33442.5 73887.5 33577.5 ;
      RECT  74007.5 32582.5 74077.5 32717.5 ;
      RECT  74265.0 32482.5 74335.0 32617.5 ;
      RECT  73745.0 33925.0 73815.0 34065.0 ;
      RECT  74080.0 33925.0 74150.0 34065.0 ;
      RECT  73745.0 32235.0 73815.0 32375.0 ;
      RECT  74080.0 32235.0 74150.0 32375.0 ;
      RECT  73560.0 32235.0 73630.0 34065.0 ;
      RECT  74265.0 32235.0 74335.0 34065.0 ;
      RECT  74450.0 32875.0 74520.0 32945.0 ;
      RECT  74522.5 32875.0 74592.5 32945.0 ;
      RECT  74450.0 32375.0 74520.0 32910.0 ;
      RECT  74485.0 32875.0 74557.5 32945.0 ;
      RECT  74522.5 32910.0 74592.5 33442.5 ;
      RECT  74785.0 33287.5 74855.0 33357.5 ;
      RECT  74712.5 33287.5 74782.5 33357.5 ;
      RECT  74785.0 33322.5 74855.0 33925.0 ;
      RECT  74747.5 33287.5 74820.0 33357.5 ;
      RECT  74712.5 32717.5 74782.5 33322.5 ;
      RECT  74450.0 33857.5 74520.0 33992.5 ;
      RECT  74785.0 32307.5 74855.0 32442.5 ;
      RECT  74522.5 33442.5 74592.5 33577.5 ;
      RECT  74712.5 32582.5 74782.5 32717.5 ;
      RECT  74970.0 32482.5 75040.0 32617.5 ;
      RECT  74450.0 33925.0 74520.0 34065.0 ;
      RECT  74785.0 33925.0 74855.0 34065.0 ;
      RECT  74450.0 32235.0 74520.0 32375.0 ;
      RECT  74785.0 32235.0 74855.0 32375.0 ;
      RECT  74265.0 32235.0 74335.0 34065.0 ;
      RECT  74970.0 32235.0 75040.0 34065.0 ;
      RECT  75155.0 32875.0 75225.0 32945.0 ;
      RECT  75227.5 32875.0 75297.5 32945.0 ;
      RECT  75155.0 32375.0 75225.0 32910.0 ;
      RECT  75190.0 32875.0 75262.5 32945.0 ;
      RECT  75227.5 32910.0 75297.5 33442.5 ;
      RECT  75490.0 33287.5 75560.0 33357.5 ;
      RECT  75417.5 33287.5 75487.5 33357.5 ;
      RECT  75490.0 33322.5 75560.0 33925.0 ;
      RECT  75452.5 33287.5 75525.0 33357.5 ;
      RECT  75417.5 32717.5 75487.5 33322.5 ;
      RECT  75155.0 33857.5 75225.0 33992.5 ;
      RECT  75490.0 32307.5 75560.0 32442.5 ;
      RECT  75227.5 33442.5 75297.5 33577.5 ;
      RECT  75417.5 32582.5 75487.5 32717.5 ;
      RECT  75675.0 32482.5 75745.0 32617.5 ;
      RECT  75155.0 33925.0 75225.0 34065.0 ;
      RECT  75490.0 33925.0 75560.0 34065.0 ;
      RECT  75155.0 32235.0 75225.0 32375.0 ;
      RECT  75490.0 32235.0 75560.0 32375.0 ;
      RECT  74970.0 32235.0 75040.0 34065.0 ;
      RECT  75675.0 32235.0 75745.0 34065.0 ;
      RECT  75860.0 32875.0 75930.0 32945.0 ;
      RECT  75932.5 32875.0 76002.5 32945.0 ;
      RECT  75860.0 32375.0 75930.0 32910.0 ;
      RECT  75895.0 32875.0 75967.5 32945.0 ;
      RECT  75932.5 32910.0 76002.5 33442.5 ;
      RECT  76195.0 33287.5 76265.0 33357.5 ;
      RECT  76122.5 33287.5 76192.5 33357.5 ;
      RECT  76195.0 33322.5 76265.0 33925.0 ;
      RECT  76157.5 33287.5 76230.0 33357.5 ;
      RECT  76122.5 32717.5 76192.5 33322.5 ;
      RECT  75860.0 33857.5 75930.0 33992.5 ;
      RECT  76195.0 32307.5 76265.0 32442.5 ;
      RECT  75932.5 33442.5 76002.5 33577.5 ;
      RECT  76122.5 32582.5 76192.5 32717.5 ;
      RECT  76380.0 32482.5 76450.0 32617.5 ;
      RECT  75860.0 33925.0 75930.0 34065.0 ;
      RECT  76195.0 33925.0 76265.0 34065.0 ;
      RECT  75860.0 32235.0 75930.0 32375.0 ;
      RECT  76195.0 32235.0 76265.0 32375.0 ;
      RECT  75675.0 32235.0 75745.0 34065.0 ;
      RECT  76380.0 32235.0 76450.0 34065.0 ;
      RECT  76565.0 32875.0 76635.0 32945.0 ;
      RECT  76637.5 32875.0 76707.5 32945.0 ;
      RECT  76565.0 32375.0 76635.0 32910.0 ;
      RECT  76600.0 32875.0 76672.5 32945.0 ;
      RECT  76637.5 32910.0 76707.5 33442.5 ;
      RECT  76900.0 33287.5 76970.0 33357.5 ;
      RECT  76827.5 33287.5 76897.5 33357.5 ;
      RECT  76900.0 33322.5 76970.0 33925.0 ;
      RECT  76862.5 33287.5 76935.0 33357.5 ;
      RECT  76827.5 32717.5 76897.5 33322.5 ;
      RECT  76565.0 33857.5 76635.0 33992.5 ;
      RECT  76900.0 32307.5 76970.0 32442.5 ;
      RECT  76637.5 33442.5 76707.5 33577.5 ;
      RECT  76827.5 32582.5 76897.5 32717.5 ;
      RECT  77085.0 32482.5 77155.0 32617.5 ;
      RECT  76565.0 33925.0 76635.0 34065.0 ;
      RECT  76900.0 33925.0 76970.0 34065.0 ;
      RECT  76565.0 32235.0 76635.0 32375.0 ;
      RECT  76900.0 32235.0 76970.0 32375.0 ;
      RECT  76380.0 32235.0 76450.0 34065.0 ;
      RECT  77085.0 32235.0 77155.0 34065.0 ;
      RECT  77270.0 32875.0 77340.0 32945.0 ;
      RECT  77342.5 32875.0 77412.5 32945.0 ;
      RECT  77270.0 32375.0 77340.0 32910.0 ;
      RECT  77305.0 32875.0 77377.5 32945.0 ;
      RECT  77342.5 32910.0 77412.5 33442.5 ;
      RECT  77605.0 33287.5 77675.0 33357.5 ;
      RECT  77532.5 33287.5 77602.5 33357.5 ;
      RECT  77605.0 33322.5 77675.0 33925.0 ;
      RECT  77567.5 33287.5 77640.0 33357.5 ;
      RECT  77532.5 32717.5 77602.5 33322.5 ;
      RECT  77270.0 33857.5 77340.0 33992.5 ;
      RECT  77605.0 32307.5 77675.0 32442.5 ;
      RECT  77342.5 33442.5 77412.5 33577.5 ;
      RECT  77532.5 32582.5 77602.5 32717.5 ;
      RECT  77790.0 32482.5 77860.0 32617.5 ;
      RECT  77270.0 33925.0 77340.0 34065.0 ;
      RECT  77605.0 33925.0 77675.0 34065.0 ;
      RECT  77270.0 32235.0 77340.0 32375.0 ;
      RECT  77605.0 32235.0 77675.0 32375.0 ;
      RECT  77085.0 32235.0 77155.0 34065.0 ;
      RECT  77790.0 32235.0 77860.0 34065.0 ;
      RECT  77975.0 32875.0 78045.0 32945.0 ;
      RECT  78047.5 32875.0 78117.5 32945.0 ;
      RECT  77975.0 32375.0 78045.0 32910.0 ;
      RECT  78010.0 32875.0 78082.5 32945.0 ;
      RECT  78047.5 32910.0 78117.5 33442.5 ;
      RECT  78310.0 33287.5 78380.0 33357.5 ;
      RECT  78237.5 33287.5 78307.5 33357.5 ;
      RECT  78310.0 33322.5 78380.0 33925.0 ;
      RECT  78272.5 33287.5 78345.0 33357.5 ;
      RECT  78237.5 32717.5 78307.5 33322.5 ;
      RECT  77975.0 33857.5 78045.0 33992.5 ;
      RECT  78310.0 32307.5 78380.0 32442.5 ;
      RECT  78047.5 33442.5 78117.5 33577.5 ;
      RECT  78237.5 32582.5 78307.5 32717.5 ;
      RECT  78495.0 32482.5 78565.0 32617.5 ;
      RECT  77975.0 33925.0 78045.0 34065.0 ;
      RECT  78310.0 33925.0 78380.0 34065.0 ;
      RECT  77975.0 32235.0 78045.0 32375.0 ;
      RECT  78310.0 32235.0 78380.0 32375.0 ;
      RECT  77790.0 32235.0 77860.0 34065.0 ;
      RECT  78495.0 32235.0 78565.0 34065.0 ;
      RECT  78680.0 32875.0 78750.0 32945.0 ;
      RECT  78752.5 32875.0 78822.5 32945.0 ;
      RECT  78680.0 32375.0 78750.0 32910.0 ;
      RECT  78715.0 32875.0 78787.5 32945.0 ;
      RECT  78752.5 32910.0 78822.5 33442.5 ;
      RECT  79015.0 33287.5 79085.0 33357.5 ;
      RECT  78942.5 33287.5 79012.5 33357.5 ;
      RECT  79015.0 33322.5 79085.0 33925.0 ;
      RECT  78977.5 33287.5 79050.0 33357.5 ;
      RECT  78942.5 32717.5 79012.5 33322.5 ;
      RECT  78680.0 33857.5 78750.0 33992.5 ;
      RECT  79015.0 32307.5 79085.0 32442.5 ;
      RECT  78752.5 33442.5 78822.5 33577.5 ;
      RECT  78942.5 32582.5 79012.5 32717.5 ;
      RECT  79200.0 32482.5 79270.0 32617.5 ;
      RECT  78680.0 33925.0 78750.0 34065.0 ;
      RECT  79015.0 33925.0 79085.0 34065.0 ;
      RECT  78680.0 32235.0 78750.0 32375.0 ;
      RECT  79015.0 32235.0 79085.0 32375.0 ;
      RECT  78495.0 32235.0 78565.0 34065.0 ;
      RECT  79200.0 32235.0 79270.0 34065.0 ;
      RECT  79385.0 32875.0 79455.0 32945.0 ;
      RECT  79457.5 32875.0 79527.5 32945.0 ;
      RECT  79385.0 32375.0 79455.0 32910.0 ;
      RECT  79420.0 32875.0 79492.5 32945.0 ;
      RECT  79457.5 32910.0 79527.5 33442.5 ;
      RECT  79720.0 33287.5 79790.0 33357.5 ;
      RECT  79647.5 33287.5 79717.5 33357.5 ;
      RECT  79720.0 33322.5 79790.0 33925.0 ;
      RECT  79682.5 33287.5 79755.0 33357.5 ;
      RECT  79647.5 32717.5 79717.5 33322.5 ;
      RECT  79385.0 33857.5 79455.0 33992.5 ;
      RECT  79720.0 32307.5 79790.0 32442.5 ;
      RECT  79457.5 33442.5 79527.5 33577.5 ;
      RECT  79647.5 32582.5 79717.5 32717.5 ;
      RECT  79905.0 32482.5 79975.0 32617.5 ;
      RECT  79385.0 33925.0 79455.0 34065.0 ;
      RECT  79720.0 33925.0 79790.0 34065.0 ;
      RECT  79385.0 32235.0 79455.0 32375.0 ;
      RECT  79720.0 32235.0 79790.0 32375.0 ;
      RECT  79200.0 32235.0 79270.0 34065.0 ;
      RECT  79905.0 32235.0 79975.0 34065.0 ;
      RECT  80090.0 32875.0 80160.0 32945.0 ;
      RECT  80162.5 32875.0 80232.5 32945.0 ;
      RECT  80090.0 32375.0 80160.0 32910.0 ;
      RECT  80125.0 32875.0 80197.5 32945.0 ;
      RECT  80162.5 32910.0 80232.5 33442.5 ;
      RECT  80425.0 33287.5 80495.0 33357.5 ;
      RECT  80352.5 33287.5 80422.5 33357.5 ;
      RECT  80425.0 33322.5 80495.0 33925.0 ;
      RECT  80387.5 33287.5 80460.0 33357.5 ;
      RECT  80352.5 32717.5 80422.5 33322.5 ;
      RECT  80090.0 33857.5 80160.0 33992.5 ;
      RECT  80425.0 32307.5 80495.0 32442.5 ;
      RECT  80162.5 33442.5 80232.5 33577.5 ;
      RECT  80352.5 32582.5 80422.5 32717.5 ;
      RECT  80610.0 32482.5 80680.0 32617.5 ;
      RECT  80090.0 33925.0 80160.0 34065.0 ;
      RECT  80425.0 33925.0 80495.0 34065.0 ;
      RECT  80090.0 32235.0 80160.0 32375.0 ;
      RECT  80425.0 32235.0 80495.0 32375.0 ;
      RECT  79905.0 32235.0 79975.0 34065.0 ;
      RECT  80610.0 32235.0 80680.0 34065.0 ;
      RECT  80795.0 32875.0 80865.0 32945.0 ;
      RECT  80867.5 32875.0 80937.5 32945.0 ;
      RECT  80795.0 32375.0 80865.0 32910.0 ;
      RECT  80830.0 32875.0 80902.5 32945.0 ;
      RECT  80867.5 32910.0 80937.5 33442.5 ;
      RECT  81130.0 33287.5 81200.0 33357.5 ;
      RECT  81057.5 33287.5 81127.5 33357.5 ;
      RECT  81130.0 33322.5 81200.0 33925.0 ;
      RECT  81092.5 33287.5 81165.0 33357.5 ;
      RECT  81057.5 32717.5 81127.5 33322.5 ;
      RECT  80795.0 33857.5 80865.0 33992.5 ;
      RECT  81130.0 32307.5 81200.0 32442.5 ;
      RECT  80867.5 33442.5 80937.5 33577.5 ;
      RECT  81057.5 32582.5 81127.5 32717.5 ;
      RECT  81315.0 32482.5 81385.0 32617.5 ;
      RECT  80795.0 33925.0 80865.0 34065.0 ;
      RECT  81130.0 33925.0 81200.0 34065.0 ;
      RECT  80795.0 32235.0 80865.0 32375.0 ;
      RECT  81130.0 32235.0 81200.0 32375.0 ;
      RECT  80610.0 32235.0 80680.0 34065.0 ;
      RECT  81315.0 32235.0 81385.0 34065.0 ;
      RECT  81500.0 32875.0 81570.0 32945.0 ;
      RECT  81572.5 32875.0 81642.5 32945.0 ;
      RECT  81500.0 32375.0 81570.0 32910.0 ;
      RECT  81535.0 32875.0 81607.5 32945.0 ;
      RECT  81572.5 32910.0 81642.5 33442.5 ;
      RECT  81835.0 33287.5 81905.0 33357.5 ;
      RECT  81762.5 33287.5 81832.5 33357.5 ;
      RECT  81835.0 33322.5 81905.0 33925.0 ;
      RECT  81797.5 33287.5 81870.0 33357.5 ;
      RECT  81762.5 32717.5 81832.5 33322.5 ;
      RECT  81500.0 33857.5 81570.0 33992.5 ;
      RECT  81835.0 32307.5 81905.0 32442.5 ;
      RECT  81572.5 33442.5 81642.5 33577.5 ;
      RECT  81762.5 32582.5 81832.5 32717.5 ;
      RECT  82020.0 32482.5 82090.0 32617.5 ;
      RECT  81500.0 33925.0 81570.0 34065.0 ;
      RECT  81835.0 33925.0 81905.0 34065.0 ;
      RECT  81500.0 32235.0 81570.0 32375.0 ;
      RECT  81835.0 32235.0 81905.0 32375.0 ;
      RECT  81315.0 32235.0 81385.0 34065.0 ;
      RECT  82020.0 32235.0 82090.0 34065.0 ;
      RECT  82205.0 32875.0 82275.0 32945.0 ;
      RECT  82277.5 32875.0 82347.5 32945.0 ;
      RECT  82205.0 32375.0 82275.0 32910.0 ;
      RECT  82240.0 32875.0 82312.5 32945.0 ;
      RECT  82277.5 32910.0 82347.5 33442.5 ;
      RECT  82540.0 33287.5 82610.0 33357.5 ;
      RECT  82467.5 33287.5 82537.5 33357.5 ;
      RECT  82540.0 33322.5 82610.0 33925.0 ;
      RECT  82502.5 33287.5 82575.0 33357.5 ;
      RECT  82467.5 32717.5 82537.5 33322.5 ;
      RECT  82205.0 33857.5 82275.0 33992.5 ;
      RECT  82540.0 32307.5 82610.0 32442.5 ;
      RECT  82277.5 33442.5 82347.5 33577.5 ;
      RECT  82467.5 32582.5 82537.5 32717.5 ;
      RECT  82725.0 32482.5 82795.0 32617.5 ;
      RECT  82205.0 33925.0 82275.0 34065.0 ;
      RECT  82540.0 33925.0 82610.0 34065.0 ;
      RECT  82205.0 32235.0 82275.0 32375.0 ;
      RECT  82540.0 32235.0 82610.0 32375.0 ;
      RECT  82020.0 32235.0 82090.0 34065.0 ;
      RECT  82725.0 32235.0 82795.0 34065.0 ;
      RECT  82910.0 32875.0 82980.0 32945.0 ;
      RECT  82982.5 32875.0 83052.5 32945.0 ;
      RECT  82910.0 32375.0 82980.0 32910.0 ;
      RECT  82945.0 32875.0 83017.5 32945.0 ;
      RECT  82982.5 32910.0 83052.5 33442.5 ;
      RECT  83245.0 33287.5 83315.0 33357.5 ;
      RECT  83172.5 33287.5 83242.5 33357.5 ;
      RECT  83245.0 33322.5 83315.0 33925.0 ;
      RECT  83207.5 33287.5 83280.0 33357.5 ;
      RECT  83172.5 32717.5 83242.5 33322.5 ;
      RECT  82910.0 33857.5 82980.0 33992.5 ;
      RECT  83245.0 32307.5 83315.0 32442.5 ;
      RECT  82982.5 33442.5 83052.5 33577.5 ;
      RECT  83172.5 32582.5 83242.5 32717.5 ;
      RECT  83430.0 32482.5 83500.0 32617.5 ;
      RECT  82910.0 33925.0 82980.0 34065.0 ;
      RECT  83245.0 33925.0 83315.0 34065.0 ;
      RECT  82910.0 32235.0 82980.0 32375.0 ;
      RECT  83245.0 32235.0 83315.0 32375.0 ;
      RECT  82725.0 32235.0 82795.0 34065.0 ;
      RECT  83430.0 32235.0 83500.0 34065.0 ;
      RECT  83615.0 32875.0 83685.0 32945.0 ;
      RECT  83687.5 32875.0 83757.5 32945.0 ;
      RECT  83615.0 32375.0 83685.0 32910.0 ;
      RECT  83650.0 32875.0 83722.5 32945.0 ;
      RECT  83687.5 32910.0 83757.5 33442.5 ;
      RECT  83950.0 33287.5 84020.0 33357.5 ;
      RECT  83877.5 33287.5 83947.5 33357.5 ;
      RECT  83950.0 33322.5 84020.0 33925.0 ;
      RECT  83912.5 33287.5 83985.0 33357.5 ;
      RECT  83877.5 32717.5 83947.5 33322.5 ;
      RECT  83615.0 33857.5 83685.0 33992.5 ;
      RECT  83950.0 32307.5 84020.0 32442.5 ;
      RECT  83687.5 33442.5 83757.5 33577.5 ;
      RECT  83877.5 32582.5 83947.5 32717.5 ;
      RECT  84135.0 32482.5 84205.0 32617.5 ;
      RECT  83615.0 33925.0 83685.0 34065.0 ;
      RECT  83950.0 33925.0 84020.0 34065.0 ;
      RECT  83615.0 32235.0 83685.0 32375.0 ;
      RECT  83950.0 32235.0 84020.0 32375.0 ;
      RECT  83430.0 32235.0 83500.0 34065.0 ;
      RECT  84135.0 32235.0 84205.0 34065.0 ;
      RECT  84320.0 32875.0 84390.0 32945.0 ;
      RECT  84392.5 32875.0 84462.5 32945.0 ;
      RECT  84320.0 32375.0 84390.0 32910.0 ;
      RECT  84355.0 32875.0 84427.5 32945.0 ;
      RECT  84392.5 32910.0 84462.5 33442.5 ;
      RECT  84655.0 33287.5 84725.0 33357.5 ;
      RECT  84582.5 33287.5 84652.5 33357.5 ;
      RECT  84655.0 33322.5 84725.0 33925.0 ;
      RECT  84617.5 33287.5 84690.0 33357.5 ;
      RECT  84582.5 32717.5 84652.5 33322.5 ;
      RECT  84320.0 33857.5 84390.0 33992.5 ;
      RECT  84655.0 32307.5 84725.0 32442.5 ;
      RECT  84392.5 33442.5 84462.5 33577.5 ;
      RECT  84582.5 32582.5 84652.5 32717.5 ;
      RECT  84840.0 32482.5 84910.0 32617.5 ;
      RECT  84320.0 33925.0 84390.0 34065.0 ;
      RECT  84655.0 33925.0 84725.0 34065.0 ;
      RECT  84320.0 32235.0 84390.0 32375.0 ;
      RECT  84655.0 32235.0 84725.0 32375.0 ;
      RECT  84135.0 32235.0 84205.0 34065.0 ;
      RECT  84840.0 32235.0 84910.0 34065.0 ;
      RECT  85025.0 32875.0 85095.0 32945.0 ;
      RECT  85097.5 32875.0 85167.5 32945.0 ;
      RECT  85025.0 32375.0 85095.0 32910.0 ;
      RECT  85060.0 32875.0 85132.5 32945.0 ;
      RECT  85097.5 32910.0 85167.5 33442.5 ;
      RECT  85360.0 33287.5 85430.0 33357.5 ;
      RECT  85287.5 33287.5 85357.5 33357.5 ;
      RECT  85360.0 33322.5 85430.0 33925.0 ;
      RECT  85322.5 33287.5 85395.0 33357.5 ;
      RECT  85287.5 32717.5 85357.5 33322.5 ;
      RECT  85025.0 33857.5 85095.0 33992.5 ;
      RECT  85360.0 32307.5 85430.0 32442.5 ;
      RECT  85097.5 33442.5 85167.5 33577.5 ;
      RECT  85287.5 32582.5 85357.5 32717.5 ;
      RECT  85545.0 32482.5 85615.0 32617.5 ;
      RECT  85025.0 33925.0 85095.0 34065.0 ;
      RECT  85360.0 33925.0 85430.0 34065.0 ;
      RECT  85025.0 32235.0 85095.0 32375.0 ;
      RECT  85360.0 32235.0 85430.0 32375.0 ;
      RECT  84840.0 32235.0 84910.0 34065.0 ;
      RECT  85545.0 32235.0 85615.0 34065.0 ;
      RECT  85730.0 32875.0 85800.0 32945.0 ;
      RECT  85802.5 32875.0 85872.5 32945.0 ;
      RECT  85730.0 32375.0 85800.0 32910.0 ;
      RECT  85765.0 32875.0 85837.5 32945.0 ;
      RECT  85802.5 32910.0 85872.5 33442.5 ;
      RECT  86065.0 33287.5 86135.0 33357.5 ;
      RECT  85992.5 33287.5 86062.5 33357.5 ;
      RECT  86065.0 33322.5 86135.0 33925.0 ;
      RECT  86027.5 33287.5 86100.0 33357.5 ;
      RECT  85992.5 32717.5 86062.5 33322.5 ;
      RECT  85730.0 33857.5 85800.0 33992.5 ;
      RECT  86065.0 32307.5 86135.0 32442.5 ;
      RECT  85802.5 33442.5 85872.5 33577.5 ;
      RECT  85992.5 32582.5 86062.5 32717.5 ;
      RECT  86250.0 32482.5 86320.0 32617.5 ;
      RECT  85730.0 33925.0 85800.0 34065.0 ;
      RECT  86065.0 33925.0 86135.0 34065.0 ;
      RECT  85730.0 32235.0 85800.0 32375.0 ;
      RECT  86065.0 32235.0 86135.0 32375.0 ;
      RECT  85545.0 32235.0 85615.0 34065.0 ;
      RECT  86250.0 32235.0 86320.0 34065.0 ;
      RECT  86435.0 32875.0 86505.0 32945.0 ;
      RECT  86507.5 32875.0 86577.5 32945.0 ;
      RECT  86435.0 32375.0 86505.0 32910.0 ;
      RECT  86470.0 32875.0 86542.5 32945.0 ;
      RECT  86507.5 32910.0 86577.5 33442.5 ;
      RECT  86770.0 33287.5 86840.0 33357.5 ;
      RECT  86697.5 33287.5 86767.5 33357.5 ;
      RECT  86770.0 33322.5 86840.0 33925.0 ;
      RECT  86732.5 33287.5 86805.0 33357.5 ;
      RECT  86697.5 32717.5 86767.5 33322.5 ;
      RECT  86435.0 33857.5 86505.0 33992.5 ;
      RECT  86770.0 32307.5 86840.0 32442.5 ;
      RECT  86507.5 33442.5 86577.5 33577.5 ;
      RECT  86697.5 32582.5 86767.5 32717.5 ;
      RECT  86955.0 32482.5 87025.0 32617.5 ;
      RECT  86435.0 33925.0 86505.0 34065.0 ;
      RECT  86770.0 33925.0 86840.0 34065.0 ;
      RECT  86435.0 32235.0 86505.0 32375.0 ;
      RECT  86770.0 32235.0 86840.0 32375.0 ;
      RECT  86250.0 32235.0 86320.0 34065.0 ;
      RECT  86955.0 32235.0 87025.0 34065.0 ;
      RECT  87140.0 32875.0 87210.0 32945.0 ;
      RECT  87212.5 32875.0 87282.5 32945.0 ;
      RECT  87140.0 32375.0 87210.0 32910.0 ;
      RECT  87175.0 32875.0 87247.5 32945.0 ;
      RECT  87212.5 32910.0 87282.5 33442.5 ;
      RECT  87475.0 33287.5 87545.0 33357.5 ;
      RECT  87402.5 33287.5 87472.5 33357.5 ;
      RECT  87475.0 33322.5 87545.0 33925.0 ;
      RECT  87437.5 33287.5 87510.0 33357.5 ;
      RECT  87402.5 32717.5 87472.5 33322.5 ;
      RECT  87140.0 33857.5 87210.0 33992.5 ;
      RECT  87475.0 32307.5 87545.0 32442.5 ;
      RECT  87212.5 33442.5 87282.5 33577.5 ;
      RECT  87402.5 32582.5 87472.5 32717.5 ;
      RECT  87660.0 32482.5 87730.0 32617.5 ;
      RECT  87140.0 33925.0 87210.0 34065.0 ;
      RECT  87475.0 33925.0 87545.0 34065.0 ;
      RECT  87140.0 32235.0 87210.0 32375.0 ;
      RECT  87475.0 32235.0 87545.0 32375.0 ;
      RECT  86955.0 32235.0 87025.0 34065.0 ;
      RECT  87660.0 32235.0 87730.0 34065.0 ;
      RECT  87845.0 32875.0 87915.0 32945.0 ;
      RECT  87917.5 32875.0 87987.5 32945.0 ;
      RECT  87845.0 32375.0 87915.0 32910.0 ;
      RECT  87880.0 32875.0 87952.5 32945.0 ;
      RECT  87917.5 32910.0 87987.5 33442.5 ;
      RECT  88180.0 33287.5 88250.0 33357.5 ;
      RECT  88107.5 33287.5 88177.5 33357.5 ;
      RECT  88180.0 33322.5 88250.0 33925.0 ;
      RECT  88142.5 33287.5 88215.0 33357.5 ;
      RECT  88107.5 32717.5 88177.5 33322.5 ;
      RECT  87845.0 33857.5 87915.0 33992.5 ;
      RECT  88180.0 32307.5 88250.0 32442.5 ;
      RECT  87917.5 33442.5 87987.5 33577.5 ;
      RECT  88107.5 32582.5 88177.5 32717.5 ;
      RECT  88365.0 32482.5 88435.0 32617.5 ;
      RECT  87845.0 33925.0 87915.0 34065.0 ;
      RECT  88180.0 33925.0 88250.0 34065.0 ;
      RECT  87845.0 32235.0 87915.0 32375.0 ;
      RECT  88180.0 32235.0 88250.0 32375.0 ;
      RECT  87660.0 32235.0 87730.0 34065.0 ;
      RECT  88365.0 32235.0 88435.0 34065.0 ;
      RECT  88550.0 32875.0 88620.0 32945.0 ;
      RECT  88622.5 32875.0 88692.5 32945.0 ;
      RECT  88550.0 32375.0 88620.0 32910.0 ;
      RECT  88585.0 32875.0 88657.5 32945.0 ;
      RECT  88622.5 32910.0 88692.5 33442.5 ;
      RECT  88885.0 33287.5 88955.0 33357.5 ;
      RECT  88812.5 33287.5 88882.5 33357.5 ;
      RECT  88885.0 33322.5 88955.0 33925.0 ;
      RECT  88847.5 33287.5 88920.0 33357.5 ;
      RECT  88812.5 32717.5 88882.5 33322.5 ;
      RECT  88550.0 33857.5 88620.0 33992.5 ;
      RECT  88885.0 32307.5 88955.0 32442.5 ;
      RECT  88622.5 33442.5 88692.5 33577.5 ;
      RECT  88812.5 32582.5 88882.5 32717.5 ;
      RECT  89070.0 32482.5 89140.0 32617.5 ;
      RECT  88550.0 33925.0 88620.0 34065.0 ;
      RECT  88885.0 33925.0 88955.0 34065.0 ;
      RECT  88550.0 32235.0 88620.0 32375.0 ;
      RECT  88885.0 32235.0 88955.0 32375.0 ;
      RECT  88365.0 32235.0 88435.0 34065.0 ;
      RECT  89070.0 32235.0 89140.0 34065.0 ;
      RECT  89255.0 32875.0 89325.0 32945.0 ;
      RECT  89327.5 32875.0 89397.5 32945.0 ;
      RECT  89255.0 32375.0 89325.0 32910.0 ;
      RECT  89290.0 32875.0 89362.5 32945.0 ;
      RECT  89327.5 32910.0 89397.5 33442.5 ;
      RECT  89590.0 33287.5 89660.0 33357.5 ;
      RECT  89517.5 33287.5 89587.5 33357.5 ;
      RECT  89590.0 33322.5 89660.0 33925.0 ;
      RECT  89552.5 33287.5 89625.0 33357.5 ;
      RECT  89517.5 32717.5 89587.5 33322.5 ;
      RECT  89255.0 33857.5 89325.0 33992.5 ;
      RECT  89590.0 32307.5 89660.0 32442.5 ;
      RECT  89327.5 33442.5 89397.5 33577.5 ;
      RECT  89517.5 32582.5 89587.5 32717.5 ;
      RECT  89775.0 32482.5 89845.0 32617.5 ;
      RECT  89255.0 33925.0 89325.0 34065.0 ;
      RECT  89590.0 33925.0 89660.0 34065.0 ;
      RECT  89255.0 32235.0 89325.0 32375.0 ;
      RECT  89590.0 32235.0 89660.0 32375.0 ;
      RECT  89070.0 32235.0 89140.0 34065.0 ;
      RECT  89775.0 32235.0 89845.0 34065.0 ;
      RECT  89960.0 32875.0 90030.0 32945.0 ;
      RECT  90032.5 32875.0 90102.5 32945.0 ;
      RECT  89960.0 32375.0 90030.0 32910.0 ;
      RECT  89995.0 32875.0 90067.5 32945.0 ;
      RECT  90032.5 32910.0 90102.5 33442.5 ;
      RECT  90295.0 33287.5 90365.0 33357.5 ;
      RECT  90222.5 33287.5 90292.5 33357.5 ;
      RECT  90295.0 33322.5 90365.0 33925.0 ;
      RECT  90257.5 33287.5 90330.0 33357.5 ;
      RECT  90222.5 32717.5 90292.5 33322.5 ;
      RECT  89960.0 33857.5 90030.0 33992.5 ;
      RECT  90295.0 32307.5 90365.0 32442.5 ;
      RECT  90032.5 33442.5 90102.5 33577.5 ;
      RECT  90222.5 32582.5 90292.5 32717.5 ;
      RECT  90480.0 32482.5 90550.0 32617.5 ;
      RECT  89960.0 33925.0 90030.0 34065.0 ;
      RECT  90295.0 33925.0 90365.0 34065.0 ;
      RECT  89960.0 32235.0 90030.0 32375.0 ;
      RECT  90295.0 32235.0 90365.0 32375.0 ;
      RECT  89775.0 32235.0 89845.0 34065.0 ;
      RECT  90480.0 32235.0 90550.0 34065.0 ;
      RECT  90665.0 32875.0 90735.0 32945.0 ;
      RECT  90737.5 32875.0 90807.5 32945.0 ;
      RECT  90665.0 32375.0 90735.0 32910.0 ;
      RECT  90700.0 32875.0 90772.5 32945.0 ;
      RECT  90737.5 32910.0 90807.5 33442.5 ;
      RECT  91000.0 33287.5 91070.0 33357.5 ;
      RECT  90927.5 33287.5 90997.5 33357.5 ;
      RECT  91000.0 33322.5 91070.0 33925.0 ;
      RECT  90962.5 33287.5 91035.0 33357.5 ;
      RECT  90927.5 32717.5 90997.5 33322.5 ;
      RECT  90665.0 33857.5 90735.0 33992.5 ;
      RECT  91000.0 32307.5 91070.0 32442.5 ;
      RECT  90737.5 33442.5 90807.5 33577.5 ;
      RECT  90927.5 32582.5 90997.5 32717.5 ;
      RECT  91185.0 32482.5 91255.0 32617.5 ;
      RECT  90665.0 33925.0 90735.0 34065.0 ;
      RECT  91000.0 33925.0 91070.0 34065.0 ;
      RECT  90665.0 32235.0 90735.0 32375.0 ;
      RECT  91000.0 32235.0 91070.0 32375.0 ;
      RECT  90480.0 32235.0 90550.0 34065.0 ;
      RECT  91185.0 32235.0 91255.0 34065.0 ;
      RECT  91370.0 32875.0 91440.0 32945.0 ;
      RECT  91442.5 32875.0 91512.5 32945.0 ;
      RECT  91370.0 32375.0 91440.0 32910.0 ;
      RECT  91405.0 32875.0 91477.5 32945.0 ;
      RECT  91442.5 32910.0 91512.5 33442.5 ;
      RECT  91705.0 33287.5 91775.0 33357.5 ;
      RECT  91632.5 33287.5 91702.5 33357.5 ;
      RECT  91705.0 33322.5 91775.0 33925.0 ;
      RECT  91667.5 33287.5 91740.0 33357.5 ;
      RECT  91632.5 32717.5 91702.5 33322.5 ;
      RECT  91370.0 33857.5 91440.0 33992.5 ;
      RECT  91705.0 32307.5 91775.0 32442.5 ;
      RECT  91442.5 33442.5 91512.5 33577.5 ;
      RECT  91632.5 32582.5 91702.5 32717.5 ;
      RECT  91890.0 32482.5 91960.0 32617.5 ;
      RECT  91370.0 33925.0 91440.0 34065.0 ;
      RECT  91705.0 33925.0 91775.0 34065.0 ;
      RECT  91370.0 32235.0 91440.0 32375.0 ;
      RECT  91705.0 32235.0 91775.0 32375.0 ;
      RECT  91185.0 32235.0 91255.0 34065.0 ;
      RECT  91890.0 32235.0 91960.0 34065.0 ;
      RECT  92075.0 32875.0 92145.0 32945.0 ;
      RECT  92147.5 32875.0 92217.5 32945.0 ;
      RECT  92075.0 32375.0 92145.0 32910.0 ;
      RECT  92110.0 32875.0 92182.5 32945.0 ;
      RECT  92147.5 32910.0 92217.5 33442.5 ;
      RECT  92410.0 33287.5 92480.0 33357.5 ;
      RECT  92337.5 33287.5 92407.5 33357.5 ;
      RECT  92410.0 33322.5 92480.0 33925.0 ;
      RECT  92372.5 33287.5 92445.0 33357.5 ;
      RECT  92337.5 32717.5 92407.5 33322.5 ;
      RECT  92075.0 33857.5 92145.0 33992.5 ;
      RECT  92410.0 32307.5 92480.0 32442.5 ;
      RECT  92147.5 33442.5 92217.5 33577.5 ;
      RECT  92337.5 32582.5 92407.5 32717.5 ;
      RECT  92595.0 32482.5 92665.0 32617.5 ;
      RECT  92075.0 33925.0 92145.0 34065.0 ;
      RECT  92410.0 33925.0 92480.0 34065.0 ;
      RECT  92075.0 32235.0 92145.0 32375.0 ;
      RECT  92410.0 32235.0 92480.0 32375.0 ;
      RECT  91890.0 32235.0 91960.0 34065.0 ;
      RECT  92595.0 32235.0 92665.0 34065.0 ;
      RECT  92780.0 32875.0 92850.0 32945.0 ;
      RECT  92852.5 32875.0 92922.5 32945.0 ;
      RECT  92780.0 32375.0 92850.0 32910.0 ;
      RECT  92815.0 32875.0 92887.5 32945.0 ;
      RECT  92852.5 32910.0 92922.5 33442.5 ;
      RECT  93115.0 33287.5 93185.0 33357.5 ;
      RECT  93042.5 33287.5 93112.5 33357.5 ;
      RECT  93115.0 33322.5 93185.0 33925.0 ;
      RECT  93077.5 33287.5 93150.0 33357.5 ;
      RECT  93042.5 32717.5 93112.5 33322.5 ;
      RECT  92780.0 33857.5 92850.0 33992.5 ;
      RECT  93115.0 32307.5 93185.0 32442.5 ;
      RECT  92852.5 33442.5 92922.5 33577.5 ;
      RECT  93042.5 32582.5 93112.5 32717.5 ;
      RECT  93300.0 32482.5 93370.0 32617.5 ;
      RECT  92780.0 33925.0 92850.0 34065.0 ;
      RECT  93115.0 33925.0 93185.0 34065.0 ;
      RECT  92780.0 32235.0 92850.0 32375.0 ;
      RECT  93115.0 32235.0 93185.0 32375.0 ;
      RECT  92595.0 32235.0 92665.0 34065.0 ;
      RECT  93300.0 32235.0 93370.0 34065.0 ;
      RECT  93485.0 32875.0 93555.0 32945.0 ;
      RECT  93557.5 32875.0 93627.5 32945.0 ;
      RECT  93485.0 32375.0 93555.0 32910.0 ;
      RECT  93520.0 32875.0 93592.5 32945.0 ;
      RECT  93557.5 32910.0 93627.5 33442.5 ;
      RECT  93820.0 33287.5 93890.0 33357.5 ;
      RECT  93747.5 33287.5 93817.5 33357.5 ;
      RECT  93820.0 33322.5 93890.0 33925.0 ;
      RECT  93782.5 33287.5 93855.0 33357.5 ;
      RECT  93747.5 32717.5 93817.5 33322.5 ;
      RECT  93485.0 33857.5 93555.0 33992.5 ;
      RECT  93820.0 32307.5 93890.0 32442.5 ;
      RECT  93557.5 33442.5 93627.5 33577.5 ;
      RECT  93747.5 32582.5 93817.5 32717.5 ;
      RECT  94005.0 32482.5 94075.0 32617.5 ;
      RECT  93485.0 33925.0 93555.0 34065.0 ;
      RECT  93820.0 33925.0 93890.0 34065.0 ;
      RECT  93485.0 32235.0 93555.0 32375.0 ;
      RECT  93820.0 32235.0 93890.0 32375.0 ;
      RECT  93300.0 32235.0 93370.0 34065.0 ;
      RECT  94005.0 32235.0 94075.0 34065.0 ;
      RECT  94190.0 32875.0 94260.0 32945.0 ;
      RECT  94262.5 32875.0 94332.5 32945.0 ;
      RECT  94190.0 32375.0 94260.0 32910.0 ;
      RECT  94225.0 32875.0 94297.5 32945.0 ;
      RECT  94262.5 32910.0 94332.5 33442.5 ;
      RECT  94525.0 33287.5 94595.0 33357.5 ;
      RECT  94452.5 33287.5 94522.5 33357.5 ;
      RECT  94525.0 33322.5 94595.0 33925.0 ;
      RECT  94487.5 33287.5 94560.0 33357.5 ;
      RECT  94452.5 32717.5 94522.5 33322.5 ;
      RECT  94190.0 33857.5 94260.0 33992.5 ;
      RECT  94525.0 32307.5 94595.0 32442.5 ;
      RECT  94262.5 33442.5 94332.5 33577.5 ;
      RECT  94452.5 32582.5 94522.5 32717.5 ;
      RECT  94710.0 32482.5 94780.0 32617.5 ;
      RECT  94190.0 33925.0 94260.0 34065.0 ;
      RECT  94525.0 33925.0 94595.0 34065.0 ;
      RECT  94190.0 32235.0 94260.0 32375.0 ;
      RECT  94525.0 32235.0 94595.0 32375.0 ;
      RECT  94005.0 32235.0 94075.0 34065.0 ;
      RECT  94710.0 32235.0 94780.0 34065.0 ;
      RECT  94895.0 32875.0 94965.0 32945.0 ;
      RECT  94967.5 32875.0 95037.5 32945.0 ;
      RECT  94895.0 32375.0 94965.0 32910.0 ;
      RECT  94930.0 32875.0 95002.5 32945.0 ;
      RECT  94967.5 32910.0 95037.5 33442.5 ;
      RECT  95230.0 33287.5 95300.0 33357.5 ;
      RECT  95157.5 33287.5 95227.5 33357.5 ;
      RECT  95230.0 33322.5 95300.0 33925.0 ;
      RECT  95192.5 33287.5 95265.0 33357.5 ;
      RECT  95157.5 32717.5 95227.5 33322.5 ;
      RECT  94895.0 33857.5 94965.0 33992.5 ;
      RECT  95230.0 32307.5 95300.0 32442.5 ;
      RECT  94967.5 33442.5 95037.5 33577.5 ;
      RECT  95157.5 32582.5 95227.5 32717.5 ;
      RECT  95415.0 32482.5 95485.0 32617.5 ;
      RECT  94895.0 33925.0 94965.0 34065.0 ;
      RECT  95230.0 33925.0 95300.0 34065.0 ;
      RECT  94895.0 32235.0 94965.0 32375.0 ;
      RECT  95230.0 32235.0 95300.0 32375.0 ;
      RECT  94710.0 32235.0 94780.0 34065.0 ;
      RECT  95415.0 32235.0 95485.0 34065.0 ;
      RECT  95600.0 32875.0 95670.0 32945.0 ;
      RECT  95672.5 32875.0 95742.5 32945.0 ;
      RECT  95600.0 32375.0 95670.0 32910.0 ;
      RECT  95635.0 32875.0 95707.5 32945.0 ;
      RECT  95672.5 32910.0 95742.5 33442.5 ;
      RECT  95935.0 33287.5 96005.0 33357.5 ;
      RECT  95862.5 33287.5 95932.5 33357.5 ;
      RECT  95935.0 33322.5 96005.0 33925.0 ;
      RECT  95897.5 33287.5 95970.0 33357.5 ;
      RECT  95862.5 32717.5 95932.5 33322.5 ;
      RECT  95600.0 33857.5 95670.0 33992.5 ;
      RECT  95935.0 32307.5 96005.0 32442.5 ;
      RECT  95672.5 33442.5 95742.5 33577.5 ;
      RECT  95862.5 32582.5 95932.5 32717.5 ;
      RECT  96120.0 32482.5 96190.0 32617.5 ;
      RECT  95600.0 33925.0 95670.0 34065.0 ;
      RECT  95935.0 33925.0 96005.0 34065.0 ;
      RECT  95600.0 32235.0 95670.0 32375.0 ;
      RECT  95935.0 32235.0 96005.0 32375.0 ;
      RECT  95415.0 32235.0 95485.0 34065.0 ;
      RECT  96120.0 32235.0 96190.0 34065.0 ;
      RECT  96305.0 32875.0 96375.0 32945.0 ;
      RECT  96377.5 32875.0 96447.5 32945.0 ;
      RECT  96305.0 32375.0 96375.0 32910.0 ;
      RECT  96340.0 32875.0 96412.5 32945.0 ;
      RECT  96377.5 32910.0 96447.5 33442.5 ;
      RECT  96640.0 33287.5 96710.0 33357.5 ;
      RECT  96567.5 33287.5 96637.5 33357.5 ;
      RECT  96640.0 33322.5 96710.0 33925.0 ;
      RECT  96602.5 33287.5 96675.0 33357.5 ;
      RECT  96567.5 32717.5 96637.5 33322.5 ;
      RECT  96305.0 33857.5 96375.0 33992.5 ;
      RECT  96640.0 32307.5 96710.0 32442.5 ;
      RECT  96377.5 33442.5 96447.5 33577.5 ;
      RECT  96567.5 32582.5 96637.5 32717.5 ;
      RECT  96825.0 32482.5 96895.0 32617.5 ;
      RECT  96305.0 33925.0 96375.0 34065.0 ;
      RECT  96640.0 33925.0 96710.0 34065.0 ;
      RECT  96305.0 32235.0 96375.0 32375.0 ;
      RECT  96640.0 32235.0 96710.0 32375.0 ;
      RECT  96120.0 32235.0 96190.0 34065.0 ;
      RECT  96825.0 32235.0 96895.0 34065.0 ;
      RECT  97010.0 32875.0 97080.0 32945.0 ;
      RECT  97082.5 32875.0 97152.5 32945.0 ;
      RECT  97010.0 32375.0 97080.0 32910.0 ;
      RECT  97045.0 32875.0 97117.5 32945.0 ;
      RECT  97082.5 32910.0 97152.5 33442.5 ;
      RECT  97345.0 33287.5 97415.0 33357.5 ;
      RECT  97272.5 33287.5 97342.5 33357.5 ;
      RECT  97345.0 33322.5 97415.0 33925.0 ;
      RECT  97307.5 33287.5 97380.0 33357.5 ;
      RECT  97272.5 32717.5 97342.5 33322.5 ;
      RECT  97010.0 33857.5 97080.0 33992.5 ;
      RECT  97345.0 32307.5 97415.0 32442.5 ;
      RECT  97082.5 33442.5 97152.5 33577.5 ;
      RECT  97272.5 32582.5 97342.5 32717.5 ;
      RECT  97530.0 32482.5 97600.0 32617.5 ;
      RECT  97010.0 33925.0 97080.0 34065.0 ;
      RECT  97345.0 33925.0 97415.0 34065.0 ;
      RECT  97010.0 32235.0 97080.0 32375.0 ;
      RECT  97345.0 32235.0 97415.0 32375.0 ;
      RECT  96825.0 32235.0 96895.0 34065.0 ;
      RECT  97530.0 32235.0 97600.0 34065.0 ;
      RECT  97715.0 32875.0 97785.0 32945.0 ;
      RECT  97787.5 32875.0 97857.5 32945.0 ;
      RECT  97715.0 32375.0 97785.0 32910.0 ;
      RECT  97750.0 32875.0 97822.5 32945.0 ;
      RECT  97787.5 32910.0 97857.5 33442.5 ;
      RECT  98050.0 33287.5 98120.0 33357.5 ;
      RECT  97977.5 33287.5 98047.5 33357.5 ;
      RECT  98050.0 33322.5 98120.0 33925.0 ;
      RECT  98012.5 33287.5 98085.0 33357.5 ;
      RECT  97977.5 32717.5 98047.5 33322.5 ;
      RECT  97715.0 33857.5 97785.0 33992.5 ;
      RECT  98050.0 32307.5 98120.0 32442.5 ;
      RECT  97787.5 33442.5 97857.5 33577.5 ;
      RECT  97977.5 32582.5 98047.5 32717.5 ;
      RECT  98235.0 32482.5 98305.0 32617.5 ;
      RECT  97715.0 33925.0 97785.0 34065.0 ;
      RECT  98050.0 33925.0 98120.0 34065.0 ;
      RECT  97715.0 32235.0 97785.0 32375.0 ;
      RECT  98050.0 32235.0 98120.0 32375.0 ;
      RECT  97530.0 32235.0 97600.0 34065.0 ;
      RECT  98235.0 32235.0 98305.0 34065.0 ;
      RECT  98420.0 32875.0 98490.0 32945.0 ;
      RECT  98492.5 32875.0 98562.5 32945.0 ;
      RECT  98420.0 32375.0 98490.0 32910.0 ;
      RECT  98455.0 32875.0 98527.5 32945.0 ;
      RECT  98492.5 32910.0 98562.5 33442.5 ;
      RECT  98755.0 33287.5 98825.0 33357.5 ;
      RECT  98682.5 33287.5 98752.5 33357.5 ;
      RECT  98755.0 33322.5 98825.0 33925.0 ;
      RECT  98717.5 33287.5 98790.0 33357.5 ;
      RECT  98682.5 32717.5 98752.5 33322.5 ;
      RECT  98420.0 33857.5 98490.0 33992.5 ;
      RECT  98755.0 32307.5 98825.0 32442.5 ;
      RECT  98492.5 33442.5 98562.5 33577.5 ;
      RECT  98682.5 32582.5 98752.5 32717.5 ;
      RECT  98940.0 32482.5 99010.0 32617.5 ;
      RECT  98420.0 33925.0 98490.0 34065.0 ;
      RECT  98755.0 33925.0 98825.0 34065.0 ;
      RECT  98420.0 32235.0 98490.0 32375.0 ;
      RECT  98755.0 32235.0 98825.0 32375.0 ;
      RECT  98235.0 32235.0 98305.0 34065.0 ;
      RECT  98940.0 32235.0 99010.0 34065.0 ;
      RECT  99125.0 32875.0 99195.0 32945.0 ;
      RECT  99197.5 32875.0 99267.5 32945.0 ;
      RECT  99125.0 32375.0 99195.0 32910.0 ;
      RECT  99160.0 32875.0 99232.5 32945.0 ;
      RECT  99197.5 32910.0 99267.5 33442.5 ;
      RECT  99460.0 33287.5 99530.0 33357.5 ;
      RECT  99387.5 33287.5 99457.5 33357.5 ;
      RECT  99460.0 33322.5 99530.0 33925.0 ;
      RECT  99422.5 33287.5 99495.0 33357.5 ;
      RECT  99387.5 32717.5 99457.5 33322.5 ;
      RECT  99125.0 33857.5 99195.0 33992.5 ;
      RECT  99460.0 32307.5 99530.0 32442.5 ;
      RECT  99197.5 33442.5 99267.5 33577.5 ;
      RECT  99387.5 32582.5 99457.5 32717.5 ;
      RECT  99645.0 32482.5 99715.0 32617.5 ;
      RECT  99125.0 33925.0 99195.0 34065.0 ;
      RECT  99460.0 33925.0 99530.0 34065.0 ;
      RECT  99125.0 32235.0 99195.0 32375.0 ;
      RECT  99460.0 32235.0 99530.0 32375.0 ;
      RECT  98940.0 32235.0 99010.0 34065.0 ;
      RECT  99645.0 32235.0 99715.0 34065.0 ;
      RECT  99830.0 32875.0 99900.0 32945.0 ;
      RECT  99902.5 32875.0 99972.5 32945.0 ;
      RECT  99830.0 32375.0 99900.0 32910.0 ;
      RECT  99865.0 32875.0 99937.5 32945.0 ;
      RECT  99902.5 32910.0 99972.5 33442.5 ;
      RECT  100165.0 33287.5 100235.0 33357.5 ;
      RECT  100092.5 33287.5 100162.5 33357.5 ;
      RECT  100165.0 33322.5 100235.0 33925.0 ;
      RECT  100127.5 33287.5 100200.0 33357.5 ;
      RECT  100092.5 32717.5 100162.5 33322.5 ;
      RECT  99830.0 33857.5 99900.0 33992.5 ;
      RECT  100165.0 32307.5 100235.0 32442.5 ;
      RECT  99902.5 33442.5 99972.5 33577.5 ;
      RECT  100092.5 32582.5 100162.5 32717.5 ;
      RECT  100350.0 32482.5 100420.0 32617.5 ;
      RECT  99830.0 33925.0 99900.0 34065.0 ;
      RECT  100165.0 33925.0 100235.0 34065.0 ;
      RECT  99830.0 32235.0 99900.0 32375.0 ;
      RECT  100165.0 32235.0 100235.0 32375.0 ;
      RECT  99645.0 32235.0 99715.0 34065.0 ;
      RECT  100350.0 32235.0 100420.0 34065.0 ;
      RECT  100535.0 32875.0 100605.0 32945.0 ;
      RECT  100607.5 32875.0 100677.5 32945.0 ;
      RECT  100535.0 32375.0 100605.0 32910.0 ;
      RECT  100570.0 32875.0 100642.5 32945.0 ;
      RECT  100607.5 32910.0 100677.5 33442.5 ;
      RECT  100870.0 33287.5 100940.0 33357.5 ;
      RECT  100797.5 33287.5 100867.5 33357.5 ;
      RECT  100870.0 33322.5 100940.0 33925.0 ;
      RECT  100832.5 33287.5 100905.0 33357.5 ;
      RECT  100797.5 32717.5 100867.5 33322.5 ;
      RECT  100535.0 33857.5 100605.0 33992.5 ;
      RECT  100870.0 32307.5 100940.0 32442.5 ;
      RECT  100607.5 33442.5 100677.5 33577.5 ;
      RECT  100797.5 32582.5 100867.5 32717.5 ;
      RECT  101055.0 32482.5 101125.0 32617.5 ;
      RECT  100535.0 33925.0 100605.0 34065.0 ;
      RECT  100870.0 33925.0 100940.0 34065.0 ;
      RECT  100535.0 32235.0 100605.0 32375.0 ;
      RECT  100870.0 32235.0 100940.0 32375.0 ;
      RECT  100350.0 32235.0 100420.0 34065.0 ;
      RECT  101055.0 32235.0 101125.0 34065.0 ;
      RECT  101240.0 32875.0 101310.0 32945.0 ;
      RECT  101312.5 32875.0 101382.5 32945.0 ;
      RECT  101240.0 32375.0 101310.0 32910.0 ;
      RECT  101275.0 32875.0 101347.5 32945.0 ;
      RECT  101312.5 32910.0 101382.5 33442.5 ;
      RECT  101575.0 33287.5 101645.0 33357.5 ;
      RECT  101502.5 33287.5 101572.5 33357.5 ;
      RECT  101575.0 33322.5 101645.0 33925.0 ;
      RECT  101537.5 33287.5 101610.0 33357.5 ;
      RECT  101502.5 32717.5 101572.5 33322.5 ;
      RECT  101240.0 33857.5 101310.0 33992.5 ;
      RECT  101575.0 32307.5 101645.0 32442.5 ;
      RECT  101312.5 33442.5 101382.5 33577.5 ;
      RECT  101502.5 32582.5 101572.5 32717.5 ;
      RECT  101760.0 32482.5 101830.0 32617.5 ;
      RECT  101240.0 33925.0 101310.0 34065.0 ;
      RECT  101575.0 33925.0 101645.0 34065.0 ;
      RECT  101240.0 32235.0 101310.0 32375.0 ;
      RECT  101575.0 32235.0 101645.0 32375.0 ;
      RECT  101055.0 32235.0 101125.0 34065.0 ;
      RECT  101760.0 32235.0 101830.0 34065.0 ;
      RECT  101945.0 32875.0 102015.0 32945.0 ;
      RECT  102017.5 32875.0 102087.5 32945.0 ;
      RECT  101945.0 32375.0 102015.0 32910.0 ;
      RECT  101980.0 32875.0 102052.5 32945.0 ;
      RECT  102017.5 32910.0 102087.5 33442.5 ;
      RECT  102280.0 33287.5 102350.0 33357.5 ;
      RECT  102207.5 33287.5 102277.5 33357.5 ;
      RECT  102280.0 33322.5 102350.0 33925.0 ;
      RECT  102242.5 33287.5 102315.0 33357.5 ;
      RECT  102207.5 32717.5 102277.5 33322.5 ;
      RECT  101945.0 33857.5 102015.0 33992.5 ;
      RECT  102280.0 32307.5 102350.0 32442.5 ;
      RECT  102017.5 33442.5 102087.5 33577.5 ;
      RECT  102207.5 32582.5 102277.5 32717.5 ;
      RECT  102465.0 32482.5 102535.0 32617.5 ;
      RECT  101945.0 33925.0 102015.0 34065.0 ;
      RECT  102280.0 33925.0 102350.0 34065.0 ;
      RECT  101945.0 32235.0 102015.0 32375.0 ;
      RECT  102280.0 32235.0 102350.0 32375.0 ;
      RECT  101760.0 32235.0 101830.0 34065.0 ;
      RECT  102465.0 32235.0 102535.0 34065.0 ;
      RECT  102650.0 32875.0 102720.0 32945.0 ;
      RECT  102722.5 32875.0 102792.5 32945.0 ;
      RECT  102650.0 32375.0 102720.0 32910.0 ;
      RECT  102685.0 32875.0 102757.5 32945.0 ;
      RECT  102722.5 32910.0 102792.5 33442.5 ;
      RECT  102985.0 33287.5 103055.0 33357.5 ;
      RECT  102912.5 33287.5 102982.5 33357.5 ;
      RECT  102985.0 33322.5 103055.0 33925.0 ;
      RECT  102947.5 33287.5 103020.0 33357.5 ;
      RECT  102912.5 32717.5 102982.5 33322.5 ;
      RECT  102650.0 33857.5 102720.0 33992.5 ;
      RECT  102985.0 32307.5 103055.0 32442.5 ;
      RECT  102722.5 33442.5 102792.5 33577.5 ;
      RECT  102912.5 32582.5 102982.5 32717.5 ;
      RECT  103170.0 32482.5 103240.0 32617.5 ;
      RECT  102650.0 33925.0 102720.0 34065.0 ;
      RECT  102985.0 33925.0 103055.0 34065.0 ;
      RECT  102650.0 32235.0 102720.0 32375.0 ;
      RECT  102985.0 32235.0 103055.0 32375.0 ;
      RECT  102465.0 32235.0 102535.0 34065.0 ;
      RECT  103170.0 32235.0 103240.0 34065.0 ;
      RECT  103355.0 32875.0 103425.0 32945.0 ;
      RECT  103427.5 32875.0 103497.5 32945.0 ;
      RECT  103355.0 32375.0 103425.0 32910.0 ;
      RECT  103390.0 32875.0 103462.5 32945.0 ;
      RECT  103427.5 32910.0 103497.5 33442.5 ;
      RECT  103690.0 33287.5 103760.0 33357.5 ;
      RECT  103617.5 33287.5 103687.5 33357.5 ;
      RECT  103690.0 33322.5 103760.0 33925.0 ;
      RECT  103652.5 33287.5 103725.0 33357.5 ;
      RECT  103617.5 32717.5 103687.5 33322.5 ;
      RECT  103355.0 33857.5 103425.0 33992.5 ;
      RECT  103690.0 32307.5 103760.0 32442.5 ;
      RECT  103427.5 33442.5 103497.5 33577.5 ;
      RECT  103617.5 32582.5 103687.5 32717.5 ;
      RECT  103875.0 32482.5 103945.0 32617.5 ;
      RECT  103355.0 33925.0 103425.0 34065.0 ;
      RECT  103690.0 33925.0 103760.0 34065.0 ;
      RECT  103355.0 32235.0 103425.0 32375.0 ;
      RECT  103690.0 32235.0 103760.0 32375.0 ;
      RECT  103170.0 32235.0 103240.0 34065.0 ;
      RECT  103875.0 32235.0 103945.0 34065.0 ;
      RECT  104060.0 32875.0 104130.0 32945.0 ;
      RECT  104132.5 32875.0 104202.5 32945.0 ;
      RECT  104060.0 32375.0 104130.0 32910.0 ;
      RECT  104095.0 32875.0 104167.5 32945.0 ;
      RECT  104132.5 32910.0 104202.5 33442.5 ;
      RECT  104395.0 33287.5 104465.0 33357.5 ;
      RECT  104322.5 33287.5 104392.5 33357.5 ;
      RECT  104395.0 33322.5 104465.0 33925.0 ;
      RECT  104357.5 33287.5 104430.0 33357.5 ;
      RECT  104322.5 32717.5 104392.5 33322.5 ;
      RECT  104060.0 33857.5 104130.0 33992.5 ;
      RECT  104395.0 32307.5 104465.0 32442.5 ;
      RECT  104132.5 33442.5 104202.5 33577.5 ;
      RECT  104322.5 32582.5 104392.5 32717.5 ;
      RECT  104580.0 32482.5 104650.0 32617.5 ;
      RECT  104060.0 33925.0 104130.0 34065.0 ;
      RECT  104395.0 33925.0 104465.0 34065.0 ;
      RECT  104060.0 32235.0 104130.0 32375.0 ;
      RECT  104395.0 32235.0 104465.0 32375.0 ;
      RECT  103875.0 32235.0 103945.0 34065.0 ;
      RECT  104580.0 32235.0 104650.0 34065.0 ;
      RECT  104765.0 32875.0 104835.0 32945.0 ;
      RECT  104837.5 32875.0 104907.5 32945.0 ;
      RECT  104765.0 32375.0 104835.0 32910.0 ;
      RECT  104800.0 32875.0 104872.5 32945.0 ;
      RECT  104837.5 32910.0 104907.5 33442.5 ;
      RECT  105100.0 33287.5 105170.0 33357.5 ;
      RECT  105027.5 33287.5 105097.5 33357.5 ;
      RECT  105100.0 33322.5 105170.0 33925.0 ;
      RECT  105062.5 33287.5 105135.0 33357.5 ;
      RECT  105027.5 32717.5 105097.5 33322.5 ;
      RECT  104765.0 33857.5 104835.0 33992.5 ;
      RECT  105100.0 32307.5 105170.0 32442.5 ;
      RECT  104837.5 33442.5 104907.5 33577.5 ;
      RECT  105027.5 32582.5 105097.5 32717.5 ;
      RECT  105285.0 32482.5 105355.0 32617.5 ;
      RECT  104765.0 33925.0 104835.0 34065.0 ;
      RECT  105100.0 33925.0 105170.0 34065.0 ;
      RECT  104765.0 32235.0 104835.0 32375.0 ;
      RECT  105100.0 32235.0 105170.0 32375.0 ;
      RECT  104580.0 32235.0 104650.0 34065.0 ;
      RECT  105285.0 32235.0 105355.0 34065.0 ;
      RECT  105470.0 32875.0 105540.0 32945.0 ;
      RECT  105542.5 32875.0 105612.5 32945.0 ;
      RECT  105470.0 32375.0 105540.0 32910.0 ;
      RECT  105505.0 32875.0 105577.5 32945.0 ;
      RECT  105542.5 32910.0 105612.5 33442.5 ;
      RECT  105805.0 33287.5 105875.0 33357.5 ;
      RECT  105732.5 33287.5 105802.5 33357.5 ;
      RECT  105805.0 33322.5 105875.0 33925.0 ;
      RECT  105767.5 33287.5 105840.0 33357.5 ;
      RECT  105732.5 32717.5 105802.5 33322.5 ;
      RECT  105470.0 33857.5 105540.0 33992.5 ;
      RECT  105805.0 32307.5 105875.0 32442.5 ;
      RECT  105542.5 33442.5 105612.5 33577.5 ;
      RECT  105732.5 32582.5 105802.5 32717.5 ;
      RECT  105990.0 32482.5 106060.0 32617.5 ;
      RECT  105470.0 33925.0 105540.0 34065.0 ;
      RECT  105805.0 33925.0 105875.0 34065.0 ;
      RECT  105470.0 32235.0 105540.0 32375.0 ;
      RECT  105805.0 32235.0 105875.0 32375.0 ;
      RECT  105285.0 32235.0 105355.0 34065.0 ;
      RECT  105990.0 32235.0 106060.0 34065.0 ;
      RECT  106175.0 32875.0 106245.0 32945.0 ;
      RECT  106247.5 32875.0 106317.5 32945.0 ;
      RECT  106175.0 32375.0 106245.0 32910.0 ;
      RECT  106210.0 32875.0 106282.5 32945.0 ;
      RECT  106247.5 32910.0 106317.5 33442.5 ;
      RECT  106510.0 33287.5 106580.0 33357.5 ;
      RECT  106437.5 33287.5 106507.5 33357.5 ;
      RECT  106510.0 33322.5 106580.0 33925.0 ;
      RECT  106472.5 33287.5 106545.0 33357.5 ;
      RECT  106437.5 32717.5 106507.5 33322.5 ;
      RECT  106175.0 33857.5 106245.0 33992.5 ;
      RECT  106510.0 32307.5 106580.0 32442.5 ;
      RECT  106247.5 33442.5 106317.5 33577.5 ;
      RECT  106437.5 32582.5 106507.5 32717.5 ;
      RECT  106695.0 32482.5 106765.0 32617.5 ;
      RECT  106175.0 33925.0 106245.0 34065.0 ;
      RECT  106510.0 33925.0 106580.0 34065.0 ;
      RECT  106175.0 32235.0 106245.0 32375.0 ;
      RECT  106510.0 32235.0 106580.0 32375.0 ;
      RECT  105990.0 32235.0 106060.0 34065.0 ;
      RECT  106695.0 32235.0 106765.0 34065.0 ;
      RECT  106880.0 32875.0 106950.0 32945.0 ;
      RECT  106952.5 32875.0 107022.5 32945.0 ;
      RECT  106880.0 32375.0 106950.0 32910.0 ;
      RECT  106915.0 32875.0 106987.5 32945.0 ;
      RECT  106952.5 32910.0 107022.5 33442.5 ;
      RECT  107215.0 33287.5 107285.0 33357.5 ;
      RECT  107142.5 33287.5 107212.5 33357.5 ;
      RECT  107215.0 33322.5 107285.0 33925.0 ;
      RECT  107177.5 33287.5 107250.0 33357.5 ;
      RECT  107142.5 32717.5 107212.5 33322.5 ;
      RECT  106880.0 33857.5 106950.0 33992.5 ;
      RECT  107215.0 32307.5 107285.0 32442.5 ;
      RECT  106952.5 33442.5 107022.5 33577.5 ;
      RECT  107142.5 32582.5 107212.5 32717.5 ;
      RECT  107400.0 32482.5 107470.0 32617.5 ;
      RECT  106880.0 33925.0 106950.0 34065.0 ;
      RECT  107215.0 33925.0 107285.0 34065.0 ;
      RECT  106880.0 32235.0 106950.0 32375.0 ;
      RECT  107215.0 32235.0 107285.0 32375.0 ;
      RECT  106695.0 32235.0 106765.0 34065.0 ;
      RECT  107400.0 32235.0 107470.0 34065.0 ;
      RECT  17480.0 31535.0 17345.0 31605.0 ;
      RECT  17680.0 31395.0 17545.0 31465.0 ;
      RECT  18185.0 31535.0 18050.0 31605.0 ;
      RECT  18385.0 31395.0 18250.0 31465.0 ;
      RECT  18890.0 31535.0 18755.0 31605.0 ;
      RECT  19090.0 31395.0 18955.0 31465.0 ;
      RECT  19595.0 31535.0 19460.0 31605.0 ;
      RECT  19795.0 31395.0 19660.0 31465.0 ;
      RECT  20300.0 31535.0 20165.0 31605.0 ;
      RECT  20500.0 31395.0 20365.0 31465.0 ;
      RECT  21005.0 31535.0 20870.0 31605.0 ;
      RECT  21205.0 31395.0 21070.0 31465.0 ;
      RECT  21710.0 31535.0 21575.0 31605.0 ;
      RECT  21910.0 31395.0 21775.0 31465.0 ;
      RECT  22415.0 31535.0 22280.0 31605.0 ;
      RECT  22615.0 31395.0 22480.0 31465.0 ;
      RECT  23120.0 31535.0 22985.0 31605.0 ;
      RECT  23320.0 31395.0 23185.0 31465.0 ;
      RECT  23825.0 31535.0 23690.0 31605.0 ;
      RECT  24025.0 31395.0 23890.0 31465.0 ;
      RECT  24530.0 31535.0 24395.0 31605.0 ;
      RECT  24730.0 31395.0 24595.0 31465.0 ;
      RECT  25235.0 31535.0 25100.0 31605.0 ;
      RECT  25435.0 31395.0 25300.0 31465.0 ;
      RECT  25940.0 31535.0 25805.0 31605.0 ;
      RECT  26140.0 31395.0 26005.0 31465.0 ;
      RECT  26645.0 31535.0 26510.0 31605.0 ;
      RECT  26845.0 31395.0 26710.0 31465.0 ;
      RECT  27350.0 31535.0 27215.0 31605.0 ;
      RECT  27550.0 31395.0 27415.0 31465.0 ;
      RECT  28055.0 31535.0 27920.0 31605.0 ;
      RECT  28255.0 31395.0 28120.0 31465.0 ;
      RECT  28760.0 31535.0 28625.0 31605.0 ;
      RECT  28960.0 31395.0 28825.0 31465.0 ;
      RECT  29465.0 31535.0 29330.0 31605.0 ;
      RECT  29665.0 31395.0 29530.0 31465.0 ;
      RECT  30170.0 31535.0 30035.0 31605.0 ;
      RECT  30370.0 31395.0 30235.0 31465.0 ;
      RECT  30875.0 31535.0 30740.0 31605.0 ;
      RECT  31075.0 31395.0 30940.0 31465.0 ;
      RECT  31580.0 31535.0 31445.0 31605.0 ;
      RECT  31780.0 31395.0 31645.0 31465.0 ;
      RECT  32285.0 31535.0 32150.0 31605.0 ;
      RECT  32485.0 31395.0 32350.0 31465.0 ;
      RECT  32990.0 31535.0 32855.0 31605.0 ;
      RECT  33190.0 31395.0 33055.0 31465.0 ;
      RECT  33695.0 31535.0 33560.0 31605.0 ;
      RECT  33895.0 31395.0 33760.0 31465.0 ;
      RECT  34400.0 31535.0 34265.0 31605.0 ;
      RECT  34600.0 31395.0 34465.0 31465.0 ;
      RECT  35105.0 31535.0 34970.0 31605.0 ;
      RECT  35305.0 31395.0 35170.0 31465.0 ;
      RECT  35810.0 31535.0 35675.0 31605.0 ;
      RECT  36010.0 31395.0 35875.0 31465.0 ;
      RECT  36515.0 31535.0 36380.0 31605.0 ;
      RECT  36715.0 31395.0 36580.0 31465.0 ;
      RECT  37220.0 31535.0 37085.0 31605.0 ;
      RECT  37420.0 31395.0 37285.0 31465.0 ;
      RECT  37925.0 31535.0 37790.0 31605.0 ;
      RECT  38125.0 31395.0 37990.0 31465.0 ;
      RECT  38630.0 31535.0 38495.0 31605.0 ;
      RECT  38830.0 31395.0 38695.0 31465.0 ;
      RECT  39335.0 31535.0 39200.0 31605.0 ;
      RECT  39535.0 31395.0 39400.0 31465.0 ;
      RECT  40040.0 31535.0 39905.0 31605.0 ;
      RECT  40240.0 31395.0 40105.0 31465.0 ;
      RECT  40745.0 31535.0 40610.0 31605.0 ;
      RECT  40945.0 31395.0 40810.0 31465.0 ;
      RECT  41450.0 31535.0 41315.0 31605.0 ;
      RECT  41650.0 31395.0 41515.0 31465.0 ;
      RECT  42155.0 31535.0 42020.0 31605.0 ;
      RECT  42355.0 31395.0 42220.0 31465.0 ;
      RECT  42860.0 31535.0 42725.0 31605.0 ;
      RECT  43060.0 31395.0 42925.0 31465.0 ;
      RECT  43565.0 31535.0 43430.0 31605.0 ;
      RECT  43765.0 31395.0 43630.0 31465.0 ;
      RECT  44270.0 31535.0 44135.0 31605.0 ;
      RECT  44470.0 31395.0 44335.0 31465.0 ;
      RECT  44975.0 31535.0 44840.0 31605.0 ;
      RECT  45175.0 31395.0 45040.0 31465.0 ;
      RECT  45680.0 31535.0 45545.0 31605.0 ;
      RECT  45880.0 31395.0 45745.0 31465.0 ;
      RECT  46385.0 31535.0 46250.0 31605.0 ;
      RECT  46585.0 31395.0 46450.0 31465.0 ;
      RECT  47090.0 31535.0 46955.0 31605.0 ;
      RECT  47290.0 31395.0 47155.0 31465.0 ;
      RECT  47795.0 31535.0 47660.0 31605.0 ;
      RECT  47995.0 31395.0 47860.0 31465.0 ;
      RECT  48500.0 31535.0 48365.0 31605.0 ;
      RECT  48700.0 31395.0 48565.0 31465.0 ;
      RECT  49205.0 31535.0 49070.0 31605.0 ;
      RECT  49405.0 31395.0 49270.0 31465.0 ;
      RECT  49910.0 31535.0 49775.0 31605.0 ;
      RECT  50110.0 31395.0 49975.0 31465.0 ;
      RECT  50615.0 31535.0 50480.0 31605.0 ;
      RECT  50815.0 31395.0 50680.0 31465.0 ;
      RECT  51320.0 31535.0 51185.0 31605.0 ;
      RECT  51520.0 31395.0 51385.0 31465.0 ;
      RECT  52025.0 31535.0 51890.0 31605.0 ;
      RECT  52225.0 31395.0 52090.0 31465.0 ;
      RECT  52730.0 31535.0 52595.0 31605.0 ;
      RECT  52930.0 31395.0 52795.0 31465.0 ;
      RECT  53435.0 31535.0 53300.0 31605.0 ;
      RECT  53635.0 31395.0 53500.0 31465.0 ;
      RECT  54140.0 31535.0 54005.0 31605.0 ;
      RECT  54340.0 31395.0 54205.0 31465.0 ;
      RECT  54845.0 31535.0 54710.0 31605.0 ;
      RECT  55045.0 31395.0 54910.0 31465.0 ;
      RECT  55550.0 31535.0 55415.0 31605.0 ;
      RECT  55750.0 31395.0 55615.0 31465.0 ;
      RECT  56255.0 31535.0 56120.0 31605.0 ;
      RECT  56455.0 31395.0 56320.0 31465.0 ;
      RECT  56960.0 31535.0 56825.0 31605.0 ;
      RECT  57160.0 31395.0 57025.0 31465.0 ;
      RECT  57665.0 31535.0 57530.0 31605.0 ;
      RECT  57865.0 31395.0 57730.0 31465.0 ;
      RECT  58370.0 31535.0 58235.0 31605.0 ;
      RECT  58570.0 31395.0 58435.0 31465.0 ;
      RECT  59075.0 31535.0 58940.0 31605.0 ;
      RECT  59275.0 31395.0 59140.0 31465.0 ;
      RECT  59780.0 31535.0 59645.0 31605.0 ;
      RECT  59980.0 31395.0 59845.0 31465.0 ;
      RECT  60485.0 31535.0 60350.0 31605.0 ;
      RECT  60685.0 31395.0 60550.0 31465.0 ;
      RECT  61190.0 31535.0 61055.0 31605.0 ;
      RECT  61390.0 31395.0 61255.0 31465.0 ;
      RECT  61895.0 31535.0 61760.0 31605.0 ;
      RECT  62095.0 31395.0 61960.0 31465.0 ;
      RECT  62600.0 31535.0 62465.0 31605.0 ;
      RECT  62800.0 31395.0 62665.0 31465.0 ;
      RECT  63305.0 31535.0 63170.0 31605.0 ;
      RECT  63505.0 31395.0 63370.0 31465.0 ;
      RECT  64010.0 31535.0 63875.0 31605.0 ;
      RECT  64210.0 31395.0 64075.0 31465.0 ;
      RECT  64715.0 31535.0 64580.0 31605.0 ;
      RECT  64915.0 31395.0 64780.0 31465.0 ;
      RECT  65420.0 31535.0 65285.0 31605.0 ;
      RECT  65620.0 31395.0 65485.0 31465.0 ;
      RECT  66125.0 31535.0 65990.0 31605.0 ;
      RECT  66325.0 31395.0 66190.0 31465.0 ;
      RECT  66830.0 31535.0 66695.0 31605.0 ;
      RECT  67030.0 31395.0 66895.0 31465.0 ;
      RECT  67535.0 31535.0 67400.0 31605.0 ;
      RECT  67735.0 31395.0 67600.0 31465.0 ;
      RECT  68240.0 31535.0 68105.0 31605.0 ;
      RECT  68440.0 31395.0 68305.0 31465.0 ;
      RECT  68945.0 31535.0 68810.0 31605.0 ;
      RECT  69145.0 31395.0 69010.0 31465.0 ;
      RECT  69650.0 31535.0 69515.0 31605.0 ;
      RECT  69850.0 31395.0 69715.0 31465.0 ;
      RECT  70355.0 31535.0 70220.0 31605.0 ;
      RECT  70555.0 31395.0 70420.0 31465.0 ;
      RECT  71060.0 31535.0 70925.0 31605.0 ;
      RECT  71260.0 31395.0 71125.0 31465.0 ;
      RECT  71765.0 31535.0 71630.0 31605.0 ;
      RECT  71965.0 31395.0 71830.0 31465.0 ;
      RECT  72470.0 31535.0 72335.0 31605.0 ;
      RECT  72670.0 31395.0 72535.0 31465.0 ;
      RECT  73175.0 31535.0 73040.0 31605.0 ;
      RECT  73375.0 31395.0 73240.0 31465.0 ;
      RECT  73880.0 31535.0 73745.0 31605.0 ;
      RECT  74080.0 31395.0 73945.0 31465.0 ;
      RECT  74585.0 31535.0 74450.0 31605.0 ;
      RECT  74785.0 31395.0 74650.0 31465.0 ;
      RECT  75290.0 31535.0 75155.0 31605.0 ;
      RECT  75490.0 31395.0 75355.0 31465.0 ;
      RECT  75995.0 31535.0 75860.0 31605.0 ;
      RECT  76195.0 31395.0 76060.0 31465.0 ;
      RECT  76700.0 31535.0 76565.0 31605.0 ;
      RECT  76900.0 31395.0 76765.0 31465.0 ;
      RECT  77405.0 31535.0 77270.0 31605.0 ;
      RECT  77605.0 31395.0 77470.0 31465.0 ;
      RECT  78110.0 31535.0 77975.0 31605.0 ;
      RECT  78310.0 31395.0 78175.0 31465.0 ;
      RECT  78815.0 31535.0 78680.0 31605.0 ;
      RECT  79015.0 31395.0 78880.0 31465.0 ;
      RECT  79520.0 31535.0 79385.0 31605.0 ;
      RECT  79720.0 31395.0 79585.0 31465.0 ;
      RECT  80225.0 31535.0 80090.0 31605.0 ;
      RECT  80425.0 31395.0 80290.0 31465.0 ;
      RECT  80930.0 31535.0 80795.0 31605.0 ;
      RECT  81130.0 31395.0 80995.0 31465.0 ;
      RECT  81635.0 31535.0 81500.0 31605.0 ;
      RECT  81835.0 31395.0 81700.0 31465.0 ;
      RECT  82340.0 31535.0 82205.0 31605.0 ;
      RECT  82540.0 31395.0 82405.0 31465.0 ;
      RECT  83045.0 31535.0 82910.0 31605.0 ;
      RECT  83245.0 31395.0 83110.0 31465.0 ;
      RECT  83750.0 31535.0 83615.0 31605.0 ;
      RECT  83950.0 31395.0 83815.0 31465.0 ;
      RECT  84455.0 31535.0 84320.0 31605.0 ;
      RECT  84655.0 31395.0 84520.0 31465.0 ;
      RECT  85160.0 31535.0 85025.0 31605.0 ;
      RECT  85360.0 31395.0 85225.0 31465.0 ;
      RECT  85865.0 31535.0 85730.0 31605.0 ;
      RECT  86065.0 31395.0 85930.0 31465.0 ;
      RECT  86570.0 31535.0 86435.0 31605.0 ;
      RECT  86770.0 31395.0 86635.0 31465.0 ;
      RECT  87275.0 31535.0 87140.0 31605.0 ;
      RECT  87475.0 31395.0 87340.0 31465.0 ;
      RECT  87980.0 31535.0 87845.0 31605.0 ;
      RECT  88180.0 31395.0 88045.0 31465.0 ;
      RECT  88685.0 31535.0 88550.0 31605.0 ;
      RECT  88885.0 31395.0 88750.0 31465.0 ;
      RECT  89390.0 31535.0 89255.0 31605.0 ;
      RECT  89590.0 31395.0 89455.0 31465.0 ;
      RECT  90095.0 31535.0 89960.0 31605.0 ;
      RECT  90295.0 31395.0 90160.0 31465.0 ;
      RECT  90800.0 31535.0 90665.0 31605.0 ;
      RECT  91000.0 31395.0 90865.0 31465.0 ;
      RECT  91505.0 31535.0 91370.0 31605.0 ;
      RECT  91705.0 31395.0 91570.0 31465.0 ;
      RECT  92210.0 31535.0 92075.0 31605.0 ;
      RECT  92410.0 31395.0 92275.0 31465.0 ;
      RECT  92915.0 31535.0 92780.0 31605.0 ;
      RECT  93115.0 31395.0 92980.0 31465.0 ;
      RECT  93620.0 31535.0 93485.0 31605.0 ;
      RECT  93820.0 31395.0 93685.0 31465.0 ;
      RECT  94325.0 31535.0 94190.0 31605.0 ;
      RECT  94525.0 31395.0 94390.0 31465.0 ;
      RECT  95030.0 31535.0 94895.0 31605.0 ;
      RECT  95230.0 31395.0 95095.0 31465.0 ;
      RECT  95735.0 31535.0 95600.0 31605.0 ;
      RECT  95935.0 31395.0 95800.0 31465.0 ;
      RECT  96440.0 31535.0 96305.0 31605.0 ;
      RECT  96640.0 31395.0 96505.0 31465.0 ;
      RECT  97145.0 31535.0 97010.0 31605.0 ;
      RECT  97345.0 31395.0 97210.0 31465.0 ;
      RECT  97850.0 31535.0 97715.0 31605.0 ;
      RECT  98050.0 31395.0 97915.0 31465.0 ;
      RECT  98555.0 31535.0 98420.0 31605.0 ;
      RECT  98755.0 31395.0 98620.0 31465.0 ;
      RECT  99260.0 31535.0 99125.0 31605.0 ;
      RECT  99460.0 31395.0 99325.0 31465.0 ;
      RECT  99965.0 31535.0 99830.0 31605.0 ;
      RECT  100165.0 31395.0 100030.0 31465.0 ;
      RECT  100670.0 31535.0 100535.0 31605.0 ;
      RECT  100870.0 31395.0 100735.0 31465.0 ;
      RECT  101375.0 31535.0 101240.0 31605.0 ;
      RECT  101575.0 31395.0 101440.0 31465.0 ;
      RECT  102080.0 31535.0 101945.0 31605.0 ;
      RECT  102280.0 31395.0 102145.0 31465.0 ;
      RECT  102785.0 31535.0 102650.0 31605.0 ;
      RECT  102985.0 31395.0 102850.0 31465.0 ;
      RECT  103490.0 31535.0 103355.0 31605.0 ;
      RECT  103690.0 31395.0 103555.0 31465.0 ;
      RECT  104195.0 31535.0 104060.0 31605.0 ;
      RECT  104395.0 31395.0 104260.0 31465.0 ;
      RECT  104900.0 31535.0 104765.0 31605.0 ;
      RECT  105100.0 31395.0 104965.0 31465.0 ;
      RECT  105605.0 31535.0 105470.0 31605.0 ;
      RECT  105805.0 31395.0 105670.0 31465.0 ;
      RECT  106310.0 31535.0 106175.0 31605.0 ;
      RECT  106510.0 31395.0 106375.0 31465.0 ;
      RECT  107015.0 31535.0 106880.0 31605.0 ;
      RECT  107215.0 31395.0 107080.0 31465.0 ;
      RECT  17345.0 33925.0 17415.0 34065.0 ;
      RECT  17680.0 33925.0 17750.0 34065.0 ;
      RECT  18050.0 33925.0 18120.0 34065.0 ;
      RECT  18385.0 33925.0 18455.0 34065.0 ;
      RECT  18755.0 33925.0 18825.0 34065.0 ;
      RECT  19090.0 33925.0 19160.0 34065.0 ;
      RECT  19460.0 33925.0 19530.0 34065.0 ;
      RECT  19795.0 33925.0 19865.0 34065.0 ;
      RECT  20165.0 33925.0 20235.0 34065.0 ;
      RECT  20500.0 33925.0 20570.0 34065.0 ;
      RECT  20870.0 33925.0 20940.0 34065.0 ;
      RECT  21205.0 33925.0 21275.0 34065.0 ;
      RECT  21575.0 33925.0 21645.0 34065.0 ;
      RECT  21910.0 33925.0 21980.0 34065.0 ;
      RECT  22280.0 33925.0 22350.0 34065.0 ;
      RECT  22615.0 33925.0 22685.0 34065.0 ;
      RECT  22985.0 33925.0 23055.0 34065.0 ;
      RECT  23320.0 33925.0 23390.0 34065.0 ;
      RECT  23690.0 33925.0 23760.0 34065.0 ;
      RECT  24025.0 33925.0 24095.0 34065.0 ;
      RECT  24395.0 33925.0 24465.0 34065.0 ;
      RECT  24730.0 33925.0 24800.0 34065.0 ;
      RECT  25100.0 33925.0 25170.0 34065.0 ;
      RECT  25435.0 33925.0 25505.0 34065.0 ;
      RECT  25805.0 33925.0 25875.0 34065.0 ;
      RECT  26140.0 33925.0 26210.0 34065.0 ;
      RECT  26510.0 33925.0 26580.0 34065.0 ;
      RECT  26845.0 33925.0 26915.0 34065.0 ;
      RECT  27215.0 33925.0 27285.0 34065.0 ;
      RECT  27550.0 33925.0 27620.0 34065.0 ;
      RECT  27920.0 33925.0 27990.0 34065.0 ;
      RECT  28255.0 33925.0 28325.0 34065.0 ;
      RECT  28625.0 33925.0 28695.0 34065.0 ;
      RECT  28960.0 33925.0 29030.0 34065.0 ;
      RECT  29330.0 33925.0 29400.0 34065.0 ;
      RECT  29665.0 33925.0 29735.0 34065.0 ;
      RECT  30035.0 33925.0 30105.0 34065.0 ;
      RECT  30370.0 33925.0 30440.0 34065.0 ;
      RECT  30740.0 33925.0 30810.0 34065.0 ;
      RECT  31075.0 33925.0 31145.0 34065.0 ;
      RECT  31445.0 33925.0 31515.0 34065.0 ;
      RECT  31780.0 33925.0 31850.0 34065.0 ;
      RECT  32150.0 33925.0 32220.0 34065.0 ;
      RECT  32485.0 33925.0 32555.0 34065.0 ;
      RECT  32855.0 33925.0 32925.0 34065.0 ;
      RECT  33190.0 33925.0 33260.0 34065.0 ;
      RECT  33560.0 33925.0 33630.0 34065.0 ;
      RECT  33895.0 33925.0 33965.0 34065.0 ;
      RECT  34265.0 33925.0 34335.0 34065.0 ;
      RECT  34600.0 33925.0 34670.0 34065.0 ;
      RECT  34970.0 33925.0 35040.0 34065.0 ;
      RECT  35305.0 33925.0 35375.0 34065.0 ;
      RECT  35675.0 33925.0 35745.0 34065.0 ;
      RECT  36010.0 33925.0 36080.0 34065.0 ;
      RECT  36380.0 33925.0 36450.0 34065.0 ;
      RECT  36715.0 33925.0 36785.0 34065.0 ;
      RECT  37085.0 33925.0 37155.0 34065.0 ;
      RECT  37420.0 33925.0 37490.0 34065.0 ;
      RECT  37790.0 33925.0 37860.0 34065.0 ;
      RECT  38125.0 33925.0 38195.0 34065.0 ;
      RECT  38495.0 33925.0 38565.0 34065.0 ;
      RECT  38830.0 33925.0 38900.0 34065.0 ;
      RECT  39200.0 33925.0 39270.0 34065.0 ;
      RECT  39535.0 33925.0 39605.0 34065.0 ;
      RECT  39905.0 33925.0 39975.0 34065.0 ;
      RECT  40240.0 33925.0 40310.0 34065.0 ;
      RECT  40610.0 33925.0 40680.0 34065.0 ;
      RECT  40945.0 33925.0 41015.0 34065.0 ;
      RECT  41315.0 33925.0 41385.0 34065.0 ;
      RECT  41650.0 33925.0 41720.0 34065.0 ;
      RECT  42020.0 33925.0 42090.0 34065.0 ;
      RECT  42355.0 33925.0 42425.0 34065.0 ;
      RECT  42725.0 33925.0 42795.0 34065.0 ;
      RECT  43060.0 33925.0 43130.0 34065.0 ;
      RECT  43430.0 33925.0 43500.0 34065.0 ;
      RECT  43765.0 33925.0 43835.0 34065.0 ;
      RECT  44135.0 33925.0 44205.0 34065.0 ;
      RECT  44470.0 33925.0 44540.0 34065.0 ;
      RECT  44840.0 33925.0 44910.0 34065.0 ;
      RECT  45175.0 33925.0 45245.0 34065.0 ;
      RECT  45545.0 33925.0 45615.0 34065.0 ;
      RECT  45880.0 33925.0 45950.0 34065.0 ;
      RECT  46250.0 33925.0 46320.0 34065.0 ;
      RECT  46585.0 33925.0 46655.0 34065.0 ;
      RECT  46955.0 33925.0 47025.0 34065.0 ;
      RECT  47290.0 33925.0 47360.0 34065.0 ;
      RECT  47660.0 33925.0 47730.0 34065.0 ;
      RECT  47995.0 33925.0 48065.0 34065.0 ;
      RECT  48365.0 33925.0 48435.0 34065.0 ;
      RECT  48700.0 33925.0 48770.0 34065.0 ;
      RECT  49070.0 33925.0 49140.0 34065.0 ;
      RECT  49405.0 33925.0 49475.0 34065.0 ;
      RECT  49775.0 33925.0 49845.0 34065.0 ;
      RECT  50110.0 33925.0 50180.0 34065.0 ;
      RECT  50480.0 33925.0 50550.0 34065.0 ;
      RECT  50815.0 33925.0 50885.0 34065.0 ;
      RECT  51185.0 33925.0 51255.0 34065.0 ;
      RECT  51520.0 33925.0 51590.0 34065.0 ;
      RECT  51890.0 33925.0 51960.0 34065.0 ;
      RECT  52225.0 33925.0 52295.0 34065.0 ;
      RECT  52595.0 33925.0 52665.0 34065.0 ;
      RECT  52930.0 33925.0 53000.0 34065.0 ;
      RECT  53300.0 33925.0 53370.0 34065.0 ;
      RECT  53635.0 33925.0 53705.0 34065.0 ;
      RECT  54005.0 33925.0 54075.0 34065.0 ;
      RECT  54340.0 33925.0 54410.0 34065.0 ;
      RECT  54710.0 33925.0 54780.0 34065.0 ;
      RECT  55045.0 33925.0 55115.0 34065.0 ;
      RECT  55415.0 33925.0 55485.0 34065.0 ;
      RECT  55750.0 33925.0 55820.0 34065.0 ;
      RECT  56120.0 33925.0 56190.0 34065.0 ;
      RECT  56455.0 33925.0 56525.0 34065.0 ;
      RECT  56825.0 33925.0 56895.0 34065.0 ;
      RECT  57160.0 33925.0 57230.0 34065.0 ;
      RECT  57530.0 33925.0 57600.0 34065.0 ;
      RECT  57865.0 33925.0 57935.0 34065.0 ;
      RECT  58235.0 33925.0 58305.0 34065.0 ;
      RECT  58570.0 33925.0 58640.0 34065.0 ;
      RECT  58940.0 33925.0 59010.0 34065.0 ;
      RECT  59275.0 33925.0 59345.0 34065.0 ;
      RECT  59645.0 33925.0 59715.0 34065.0 ;
      RECT  59980.0 33925.0 60050.0 34065.0 ;
      RECT  60350.0 33925.0 60420.0 34065.0 ;
      RECT  60685.0 33925.0 60755.0 34065.0 ;
      RECT  61055.0 33925.0 61125.0 34065.0 ;
      RECT  61390.0 33925.0 61460.0 34065.0 ;
      RECT  61760.0 33925.0 61830.0 34065.0 ;
      RECT  62095.0 33925.0 62165.0 34065.0 ;
      RECT  62465.0 33925.0 62535.0 34065.0 ;
      RECT  62800.0 33925.0 62870.0 34065.0 ;
      RECT  63170.0 33925.0 63240.0 34065.0 ;
      RECT  63505.0 33925.0 63575.0 34065.0 ;
      RECT  63875.0 33925.0 63945.0 34065.0 ;
      RECT  64210.0 33925.0 64280.0 34065.0 ;
      RECT  64580.0 33925.0 64650.0 34065.0 ;
      RECT  64915.0 33925.0 64985.0 34065.0 ;
      RECT  65285.0 33925.0 65355.0 34065.0 ;
      RECT  65620.0 33925.0 65690.0 34065.0 ;
      RECT  65990.0 33925.0 66060.0 34065.0 ;
      RECT  66325.0 33925.0 66395.0 34065.0 ;
      RECT  66695.0 33925.0 66765.0 34065.0 ;
      RECT  67030.0 33925.0 67100.0 34065.0 ;
      RECT  67400.0 33925.0 67470.0 34065.0 ;
      RECT  67735.0 33925.0 67805.0 34065.0 ;
      RECT  68105.0 33925.0 68175.0 34065.0 ;
      RECT  68440.0 33925.0 68510.0 34065.0 ;
      RECT  68810.0 33925.0 68880.0 34065.0 ;
      RECT  69145.0 33925.0 69215.0 34065.0 ;
      RECT  69515.0 33925.0 69585.0 34065.0 ;
      RECT  69850.0 33925.0 69920.0 34065.0 ;
      RECT  70220.0 33925.0 70290.0 34065.0 ;
      RECT  70555.0 33925.0 70625.0 34065.0 ;
      RECT  70925.0 33925.0 70995.0 34065.0 ;
      RECT  71260.0 33925.0 71330.0 34065.0 ;
      RECT  71630.0 33925.0 71700.0 34065.0 ;
      RECT  71965.0 33925.0 72035.0 34065.0 ;
      RECT  72335.0 33925.0 72405.0 34065.0 ;
      RECT  72670.0 33925.0 72740.0 34065.0 ;
      RECT  73040.0 33925.0 73110.0 34065.0 ;
      RECT  73375.0 33925.0 73445.0 34065.0 ;
      RECT  73745.0 33925.0 73815.0 34065.0 ;
      RECT  74080.0 33925.0 74150.0 34065.0 ;
      RECT  74450.0 33925.0 74520.0 34065.0 ;
      RECT  74785.0 33925.0 74855.0 34065.0 ;
      RECT  75155.0 33925.0 75225.0 34065.0 ;
      RECT  75490.0 33925.0 75560.0 34065.0 ;
      RECT  75860.0 33925.0 75930.0 34065.0 ;
      RECT  76195.0 33925.0 76265.0 34065.0 ;
      RECT  76565.0 33925.0 76635.0 34065.0 ;
      RECT  76900.0 33925.0 76970.0 34065.0 ;
      RECT  77270.0 33925.0 77340.0 34065.0 ;
      RECT  77605.0 33925.0 77675.0 34065.0 ;
      RECT  77975.0 33925.0 78045.0 34065.0 ;
      RECT  78310.0 33925.0 78380.0 34065.0 ;
      RECT  78680.0 33925.0 78750.0 34065.0 ;
      RECT  79015.0 33925.0 79085.0 34065.0 ;
      RECT  79385.0 33925.0 79455.0 34065.0 ;
      RECT  79720.0 33925.0 79790.0 34065.0 ;
      RECT  80090.0 33925.0 80160.0 34065.0 ;
      RECT  80425.0 33925.0 80495.0 34065.0 ;
      RECT  80795.0 33925.0 80865.0 34065.0 ;
      RECT  81130.0 33925.0 81200.0 34065.0 ;
      RECT  81500.0 33925.0 81570.0 34065.0 ;
      RECT  81835.0 33925.0 81905.0 34065.0 ;
      RECT  82205.0 33925.0 82275.0 34065.0 ;
      RECT  82540.0 33925.0 82610.0 34065.0 ;
      RECT  82910.0 33925.0 82980.0 34065.0 ;
      RECT  83245.0 33925.0 83315.0 34065.0 ;
      RECT  83615.0 33925.0 83685.0 34065.0 ;
      RECT  83950.0 33925.0 84020.0 34065.0 ;
      RECT  84320.0 33925.0 84390.0 34065.0 ;
      RECT  84655.0 33925.0 84725.0 34065.0 ;
      RECT  85025.0 33925.0 85095.0 34065.0 ;
      RECT  85360.0 33925.0 85430.0 34065.0 ;
      RECT  85730.0 33925.0 85800.0 34065.0 ;
      RECT  86065.0 33925.0 86135.0 34065.0 ;
      RECT  86435.0 33925.0 86505.0 34065.0 ;
      RECT  86770.0 33925.0 86840.0 34065.0 ;
      RECT  87140.0 33925.0 87210.0 34065.0 ;
      RECT  87475.0 33925.0 87545.0 34065.0 ;
      RECT  87845.0 33925.0 87915.0 34065.0 ;
      RECT  88180.0 33925.0 88250.0 34065.0 ;
      RECT  88550.0 33925.0 88620.0 34065.0 ;
      RECT  88885.0 33925.0 88955.0 34065.0 ;
      RECT  89255.0 33925.0 89325.0 34065.0 ;
      RECT  89590.0 33925.0 89660.0 34065.0 ;
      RECT  89960.0 33925.0 90030.0 34065.0 ;
      RECT  90295.0 33925.0 90365.0 34065.0 ;
      RECT  90665.0 33925.0 90735.0 34065.0 ;
      RECT  91000.0 33925.0 91070.0 34065.0 ;
      RECT  91370.0 33925.0 91440.0 34065.0 ;
      RECT  91705.0 33925.0 91775.0 34065.0 ;
      RECT  92075.0 33925.0 92145.0 34065.0 ;
      RECT  92410.0 33925.0 92480.0 34065.0 ;
      RECT  92780.0 33925.0 92850.0 34065.0 ;
      RECT  93115.0 33925.0 93185.0 34065.0 ;
      RECT  93485.0 33925.0 93555.0 34065.0 ;
      RECT  93820.0 33925.0 93890.0 34065.0 ;
      RECT  94190.0 33925.0 94260.0 34065.0 ;
      RECT  94525.0 33925.0 94595.0 34065.0 ;
      RECT  94895.0 33925.0 94965.0 34065.0 ;
      RECT  95230.0 33925.0 95300.0 34065.0 ;
      RECT  95600.0 33925.0 95670.0 34065.0 ;
      RECT  95935.0 33925.0 96005.0 34065.0 ;
      RECT  96305.0 33925.0 96375.0 34065.0 ;
      RECT  96640.0 33925.0 96710.0 34065.0 ;
      RECT  97010.0 33925.0 97080.0 34065.0 ;
      RECT  97345.0 33925.0 97415.0 34065.0 ;
      RECT  97715.0 33925.0 97785.0 34065.0 ;
      RECT  98050.0 33925.0 98120.0 34065.0 ;
      RECT  98420.0 33925.0 98490.0 34065.0 ;
      RECT  98755.0 33925.0 98825.0 34065.0 ;
      RECT  99125.0 33925.0 99195.0 34065.0 ;
      RECT  99460.0 33925.0 99530.0 34065.0 ;
      RECT  99830.0 33925.0 99900.0 34065.0 ;
      RECT  100165.0 33925.0 100235.0 34065.0 ;
      RECT  100535.0 33925.0 100605.0 34065.0 ;
      RECT  100870.0 33925.0 100940.0 34065.0 ;
      RECT  101240.0 33925.0 101310.0 34065.0 ;
      RECT  101575.0 33925.0 101645.0 34065.0 ;
      RECT  101945.0 33925.0 102015.0 34065.0 ;
      RECT  102280.0 33925.0 102350.0 34065.0 ;
      RECT  102650.0 33925.0 102720.0 34065.0 ;
      RECT  102985.0 33925.0 103055.0 34065.0 ;
      RECT  103355.0 33925.0 103425.0 34065.0 ;
      RECT  103690.0 33925.0 103760.0 34065.0 ;
      RECT  104060.0 33925.0 104130.0 34065.0 ;
      RECT  104395.0 33925.0 104465.0 34065.0 ;
      RECT  104765.0 33925.0 104835.0 34065.0 ;
      RECT  105100.0 33925.0 105170.0 34065.0 ;
      RECT  105470.0 33925.0 105540.0 34065.0 ;
      RECT  105805.0 33925.0 105875.0 34065.0 ;
      RECT  106175.0 33925.0 106245.0 34065.0 ;
      RECT  106510.0 33925.0 106580.0 34065.0 ;
      RECT  106880.0 33925.0 106950.0 34065.0 ;
      RECT  107215.0 33925.0 107285.0 34065.0 ;
      RECT  17345.0 31255.0 17415.0 32235.0 ;
      RECT  17680.0 31255.0 17750.0 32235.0 ;
      RECT  20165.0 31255.0 20235.0 32235.0 ;
      RECT  20500.0 31255.0 20570.0 32235.0 ;
      RECT  22985.0 31255.0 23055.0 32235.0 ;
      RECT  23320.0 31255.0 23390.0 32235.0 ;
      RECT  25805.0 31255.0 25875.0 32235.0 ;
      RECT  26140.0 31255.0 26210.0 32235.0 ;
      RECT  28625.0 31255.0 28695.0 32235.0 ;
      RECT  28960.0 31255.0 29030.0 32235.0 ;
      RECT  31445.0 31255.0 31515.0 32235.0 ;
      RECT  31780.0 31255.0 31850.0 32235.0 ;
      RECT  34265.0 31255.0 34335.0 32235.0 ;
      RECT  34600.0 31255.0 34670.0 32235.0 ;
      RECT  37085.0 31255.0 37155.0 32235.0 ;
      RECT  37420.0 31255.0 37490.0 32235.0 ;
      RECT  39905.0 31255.0 39975.0 32235.0 ;
      RECT  40240.0 31255.0 40310.0 32235.0 ;
      RECT  42725.0 31255.0 42795.0 32235.0 ;
      RECT  43060.0 31255.0 43130.0 32235.0 ;
      RECT  45545.0 31255.0 45615.0 32235.0 ;
      RECT  45880.0 31255.0 45950.0 32235.0 ;
      RECT  48365.0 31255.0 48435.0 32235.0 ;
      RECT  48700.0 31255.0 48770.0 32235.0 ;
      RECT  51185.0 31255.0 51255.0 32235.0 ;
      RECT  51520.0 31255.0 51590.0 32235.0 ;
      RECT  54005.0 31255.0 54075.0 32235.0 ;
      RECT  54340.0 31255.0 54410.0 32235.0 ;
      RECT  56825.0 31255.0 56895.0 32235.0 ;
      RECT  57160.0 31255.0 57230.0 32235.0 ;
      RECT  59645.0 31255.0 59715.0 32235.0 ;
      RECT  59980.0 31255.0 60050.0 32235.0 ;
      RECT  62465.0 31255.0 62535.0 32235.0 ;
      RECT  62800.0 31255.0 62870.0 32235.0 ;
      RECT  65285.0 31255.0 65355.0 32235.0 ;
      RECT  65620.0 31255.0 65690.0 32235.0 ;
      RECT  68105.0 31255.0 68175.0 32235.0 ;
      RECT  68440.0 31255.0 68510.0 32235.0 ;
      RECT  70925.0 31255.0 70995.0 32235.0 ;
      RECT  71260.0 31255.0 71330.0 32235.0 ;
      RECT  73745.0 31255.0 73815.0 32235.0 ;
      RECT  74080.0 31255.0 74150.0 32235.0 ;
      RECT  76565.0 31255.0 76635.0 32235.0 ;
      RECT  76900.0 31255.0 76970.0 32235.0 ;
      RECT  79385.0 31255.0 79455.0 32235.0 ;
      RECT  79720.0 31255.0 79790.0 32235.0 ;
      RECT  82205.0 31255.0 82275.0 32235.0 ;
      RECT  82540.0 31255.0 82610.0 32235.0 ;
      RECT  85025.0 31255.0 85095.0 32235.0 ;
      RECT  85360.0 31255.0 85430.0 32235.0 ;
      RECT  87845.0 31255.0 87915.0 32235.0 ;
      RECT  88180.0 31255.0 88250.0 32235.0 ;
      RECT  90665.0 31255.0 90735.0 32235.0 ;
      RECT  91000.0 31255.0 91070.0 32235.0 ;
      RECT  93485.0 31255.0 93555.0 32235.0 ;
      RECT  93820.0 31255.0 93890.0 32235.0 ;
      RECT  96305.0 31255.0 96375.0 32235.0 ;
      RECT  96640.0 31255.0 96710.0 32235.0 ;
      RECT  99125.0 31255.0 99195.0 32235.0 ;
      RECT  99460.0 31255.0 99530.0 32235.0 ;
      RECT  101945.0 31255.0 102015.0 32235.0 ;
      RECT  102280.0 31255.0 102350.0 32235.0 ;
      RECT  104765.0 31255.0 104835.0 32235.0 ;
      RECT  105100.0 31255.0 105170.0 32235.0 ;
      RECT  17160.0 31255.0 17230.0 34065.0 ;
      RECT  17865.0 31255.0 17935.0 34065.0 ;
      RECT  18570.0 31255.0 18640.0 34065.0 ;
      RECT  19275.0 31255.0 19345.0 34065.0 ;
      RECT  19980.0 31255.0 20050.0 34065.0 ;
      RECT  20685.0 31255.0 20755.0 34065.0 ;
      RECT  21390.0 31255.0 21460.0 34065.0 ;
      RECT  22095.0 31255.0 22165.0 34065.0 ;
      RECT  22800.0 31255.0 22870.0 34065.0 ;
      RECT  23505.0 31255.0 23575.0 34065.0 ;
      RECT  24210.0 31255.0 24280.0 34065.0 ;
      RECT  24915.0 31255.0 24985.0 34065.0 ;
      RECT  25620.0 31255.0 25690.0 34065.0 ;
      RECT  26325.0 31255.0 26395.0 34065.0 ;
      RECT  27030.0 31255.0 27100.0 34065.0 ;
      RECT  27735.0 31255.0 27805.0 34065.0 ;
      RECT  28440.0 31255.0 28510.0 34065.0 ;
      RECT  29145.0 31255.0 29215.0 34065.0 ;
      RECT  29850.0 31255.0 29920.0 34065.0 ;
      RECT  30555.0 31255.0 30625.0 34065.0 ;
      RECT  31260.0 31255.0 31330.0 34065.0 ;
      RECT  31965.0 31255.0 32035.0 34065.0 ;
      RECT  32670.0 31255.0 32740.0 34065.0 ;
      RECT  33375.0 31255.0 33445.0 34065.0 ;
      RECT  34080.0 31255.0 34150.0 34065.0 ;
      RECT  34785.0 31255.0 34855.0 34065.0 ;
      RECT  35490.0 31255.0 35560.0 34065.0 ;
      RECT  36195.0 31255.0 36265.0 34065.0 ;
      RECT  36900.0 31255.0 36970.0 34065.0 ;
      RECT  37605.0 31255.0 37675.0 34065.0 ;
      RECT  38310.0 31255.0 38380.0 34065.0 ;
      RECT  39015.0 31255.0 39085.0 34065.0 ;
      RECT  39720.0 31255.0 39790.0 34065.0 ;
      RECT  40425.0 31255.0 40495.0 34065.0 ;
      RECT  41130.0 31255.0 41200.0 34065.0 ;
      RECT  41835.0 31255.0 41905.0 34065.0 ;
      RECT  42540.0 31255.0 42610.0 34065.0 ;
      RECT  43245.0 31255.0 43315.0 34065.0 ;
      RECT  43950.0 31255.0 44020.0 34065.0 ;
      RECT  44655.0 31255.0 44725.0 34065.0 ;
      RECT  45360.0 31255.0 45430.0 34065.0 ;
      RECT  46065.0 31255.0 46135.0 34065.0 ;
      RECT  46770.0 31255.0 46840.0 34065.0 ;
      RECT  47475.0 31255.0 47545.0 34065.0 ;
      RECT  48180.0 31255.0 48250.0 34065.0 ;
      RECT  48885.0 31255.0 48955.0 34065.0 ;
      RECT  49590.0 31255.0 49660.0 34065.0 ;
      RECT  50295.0 31255.0 50365.0 34065.0 ;
      RECT  51000.0 31255.0 51070.0 34065.0 ;
      RECT  51705.0 31255.0 51775.0 34065.0 ;
      RECT  52410.0 31255.0 52480.0 34065.0 ;
      RECT  53115.0 31255.0 53185.0 34065.0 ;
      RECT  53820.0 31255.0 53890.0 34065.0 ;
      RECT  54525.0 31255.0 54595.0 34065.0 ;
      RECT  55230.0 31255.0 55300.0 34065.0 ;
      RECT  55935.0 31255.0 56005.0 34065.0 ;
      RECT  56640.0 31255.0 56710.0 34065.0 ;
      RECT  57345.0 31255.0 57415.0 34065.0 ;
      RECT  58050.0 31255.0 58120.0 34065.0 ;
      RECT  58755.0 31255.0 58825.0 34065.0 ;
      RECT  59460.0 31255.0 59530.0 34065.0 ;
      RECT  60165.0 31255.0 60235.0 34065.0 ;
      RECT  60870.0 31255.0 60940.0 34065.0 ;
      RECT  61575.0 31255.0 61645.0 34065.0 ;
      RECT  62280.0 31255.0 62350.0 34065.0 ;
      RECT  62985.0 31255.0 63055.0 34065.0 ;
      RECT  63690.0 31255.0 63760.0 34065.0 ;
      RECT  64395.0 31255.0 64465.0 34065.0 ;
      RECT  65100.0 31255.0 65170.0 34065.0 ;
      RECT  65805.0 31255.0 65875.0 34065.0 ;
      RECT  66510.0 31255.0 66580.0 34065.0 ;
      RECT  67215.0 31255.0 67285.0 34065.0 ;
      RECT  67920.0 31255.0 67990.0 34065.0 ;
      RECT  68625.0 31255.0 68695.0 34065.0 ;
      RECT  69330.0 31255.0 69400.0 34065.0 ;
      RECT  70035.0 31255.0 70105.0 34065.0 ;
      RECT  70740.0 31255.0 70810.0 34065.0 ;
      RECT  71445.0 31255.0 71515.0 34065.0 ;
      RECT  72150.0 31255.0 72220.0 34065.0 ;
      RECT  72855.0 31255.0 72925.0 34065.0 ;
      RECT  73560.0 31255.0 73630.0 34065.0 ;
      RECT  74265.0 31255.0 74335.0 34065.0 ;
      RECT  74970.0 31255.0 75040.0 34065.0 ;
      RECT  75675.0 31255.0 75745.0 34065.0 ;
      RECT  76380.0 31255.0 76450.0 34065.0 ;
      RECT  77085.0 31255.0 77155.0 34065.0 ;
      RECT  77790.0 31255.0 77860.0 34065.0 ;
      RECT  78495.0 31255.0 78565.0 34065.0 ;
      RECT  79200.0 31255.0 79270.0 34065.0 ;
      RECT  79905.0 31255.0 79975.0 34065.0 ;
      RECT  80610.0 31255.0 80680.0 34065.0 ;
      RECT  81315.0 31255.0 81385.0 34065.0 ;
      RECT  82020.0 31255.0 82090.0 34065.0 ;
      RECT  82725.0 31255.0 82795.0 34065.0 ;
      RECT  83430.0 31255.0 83500.0 34065.0 ;
      RECT  84135.0 31255.0 84205.0 34065.0 ;
      RECT  84840.0 31255.0 84910.0 34065.0 ;
      RECT  85545.0 31255.0 85615.0 34065.0 ;
      RECT  86250.0 31255.0 86320.0 34065.0 ;
      RECT  86955.0 31255.0 87025.0 34065.0 ;
      RECT  87660.0 31255.0 87730.0 34065.0 ;
      RECT  88365.0 31255.0 88435.0 34065.0 ;
      RECT  89070.0 31255.0 89140.0 34065.0 ;
      RECT  89775.0 31255.0 89845.0 34065.0 ;
      RECT  90480.0 31255.0 90550.0 34065.0 ;
      RECT  91185.0 31255.0 91255.0 34065.0 ;
      RECT  91890.0 31255.0 91960.0 34065.0 ;
      RECT  92595.0 31255.0 92665.0 34065.0 ;
      RECT  93300.0 31255.0 93370.0 34065.0 ;
      RECT  94005.0 31255.0 94075.0 34065.0 ;
      RECT  94710.0 31255.0 94780.0 34065.0 ;
      RECT  95415.0 31255.0 95485.0 34065.0 ;
      RECT  96120.0 31255.0 96190.0 34065.0 ;
      RECT  96825.0 31255.0 96895.0 34065.0 ;
      RECT  97530.0 31255.0 97600.0 34065.0 ;
      RECT  98235.0 31255.0 98305.0 34065.0 ;
      RECT  98940.0 31255.0 99010.0 34065.0 ;
      RECT  99645.0 31255.0 99715.0 34065.0 ;
      RECT  100350.0 31255.0 100420.0 34065.0 ;
      RECT  101055.0 31255.0 101125.0 34065.0 ;
      RECT  101760.0 31255.0 101830.0 34065.0 ;
      RECT  102465.0 31255.0 102535.0 34065.0 ;
      RECT  103170.0 31255.0 103240.0 34065.0 ;
      RECT  103875.0 31255.0 103945.0 34065.0 ;
      RECT  104580.0 31255.0 104650.0 34065.0 ;
      RECT  105285.0 31255.0 105355.0 34065.0 ;
      RECT  105990.0 31255.0 106060.0 34065.0 ;
      RECT  106695.0 31255.0 106765.0 34065.0 ;
      RECT  9895.0 35.0 9965.0 5275.0 ;
      RECT  10170.0 35.0 10240.0 5275.0 ;
      RECT  9345.0 35.0 9415.0 5275.0 ;
      RECT  9620.0 35.0 9690.0 5275.0 ;
      RECT  10700.0 640.0 10770.0 710.0 ;
      RECT  10890.0 640.0 10960.0 710.0 ;
      RECT  10700.0 675.0 10770.0 1037.5 ;
      RECT  10735.0 640.0 10925.0 710.0 ;
      RECT  10890.0 332.5 10960.0 675.0 ;
      RECT  10700.0 1037.5 10770.0 1172.5 ;
      RECT  10890.0 197.5 10960.0 332.5 ;
      RECT  10992.5 640.0 10857.5 710.0 ;
      RECT  10700.0 2120.0 10770.0 2050.0 ;
      RECT  10890.0 2120.0 10960.0 2050.0 ;
      RECT  10700.0 2085.0 10770.0 1722.5 ;
      RECT  10735.0 2120.0 10925.0 2050.0 ;
      RECT  10890.0 2427.5 10960.0 2085.0 ;
      RECT  10700.0 1722.5 10770.0 1587.5 ;
      RECT  10890.0 2562.5 10960.0 2427.5 ;
      RECT  10992.5 2120.0 10857.5 2050.0 ;
      RECT  10700.0 3330.0 10770.0 3400.0 ;
      RECT  10890.0 3330.0 10960.0 3400.0 ;
      RECT  10700.0 3365.0 10770.0 3727.5 ;
      RECT  10735.0 3330.0 10925.0 3400.0 ;
      RECT  10890.0 3022.5 10960.0 3365.0 ;
      RECT  10700.0 3727.5 10770.0 3862.5 ;
      RECT  10890.0 2887.5 10960.0 3022.5 ;
      RECT  10992.5 3330.0 10857.5 3400.0 ;
      RECT  10700.0 4810.0 10770.0 4740.0 ;
      RECT  10890.0 4810.0 10960.0 4740.0 ;
      RECT  10700.0 4775.0 10770.0 4412.5 ;
      RECT  10735.0 4810.0 10925.0 4740.0 ;
      RECT  10890.0 5117.5 10960.0 4775.0 ;
      RECT  10700.0 4412.5 10770.0 4277.5 ;
      RECT  10890.0 5252.5 10960.0 5117.5 ;
      RECT  10992.5 4810.0 10857.5 4740.0 ;
      RECT  9447.5 1150.0 9312.5 1220.0 ;
      RECT  8062.5 627.5 7927.5 697.5 ;
      RECT  9722.5 2495.0 9587.5 2565.0 ;
      RECT  8337.5 2062.5 8202.5 2132.5 ;
      RECT  8062.5 2825.0 7927.5 2895.0 ;
      RECT  9997.5 2825.0 9862.5 2895.0 ;
      RECT  8337.5 4170.0 8202.5 4240.0 ;
      RECT  10272.5 4170.0 10137.5 4240.0 ;
      RECT  9447.5 640.0 9312.5 710.0 ;
      RECT  9722.5 425.0 9587.5 495.0 ;
      RECT  9997.5 2050.0 9862.5 2120.0 ;
      RECT  9722.5 2265.0 9587.5 2335.0 ;
      RECT  9447.5 3330.0 9312.5 3400.0 ;
      RECT  10272.5 3115.0 10137.5 3185.0 ;
      RECT  9997.5 4740.0 9862.5 4810.0 ;
      RECT  10272.5 4955.0 10137.5 5025.0 ;
      RECT  7960.0 35.0 8030.0 5275.0 ;
      RECT  8235.0 35.0 8305.0 5275.0 ;
      RECT  17195.0 26370.0 17900.0 31255.0 ;
      RECT  20015.0 26370.0 20720.0 31255.0 ;
      RECT  22835.0 26370.0 23540.0 31255.0 ;
      RECT  25655.0 26370.0 26360.0 31255.0 ;
      RECT  28475.0 26370.0 29180.0 31255.0 ;
      RECT  31295.0 26370.0 32000.0 31255.0 ;
      RECT  34115.0 26370.0 34820.0 31255.0 ;
      RECT  36935.0 26370.0 37640.0 31255.0 ;
      RECT  39755.0 26370.0 40460.0 31255.0 ;
      RECT  42575.0 26370.0 43280.0 31255.0 ;
      RECT  45395.0 26370.0 46100.0 31255.0 ;
      RECT  48215.0 26370.0 48920.0 31255.0 ;
      RECT  51035.0 26370.0 51740.0 31255.0 ;
      RECT  53855.0 26370.0 54560.0 31255.0 ;
      RECT  56675.0 26370.0 57380.0 31255.0 ;
      RECT  59495.0 26370.0 60200.0 31255.0 ;
      RECT  62315.0 26370.0 63020.0 31255.0 ;
      RECT  65135.0 26370.0 65840.0 31255.0 ;
      RECT  67955.0 26370.0 68660.0 31255.0 ;
      RECT  70775.0 26370.0 71480.0 31255.0 ;
      RECT  73595.0 26370.0 74300.0 31255.0 ;
      RECT  76415.0 26370.0 77120.0 31255.0 ;
      RECT  79235.0 26370.0 79940.0 31255.0 ;
      RECT  82055.0 26370.0 82760.0 31255.0 ;
      RECT  84875.0 26370.0 85580.0 31255.0 ;
      RECT  87695.0 26370.0 88400.0 31255.0 ;
      RECT  90515.0 26370.0 91220.0 31255.0 ;
      RECT  93335.0 26370.0 94040.0 31255.0 ;
      RECT  96155.0 26370.0 96860.0 31255.0 ;
      RECT  98975.0 26370.0 99680.0 31255.0 ;
      RECT  101795.0 26370.0 102500.0 31255.0 ;
      RECT  104615.0 26370.0 105320.0 31255.0 ;
      RECT  17345.0 26370.0 17415.0 31255.0 ;
      RECT  17680.0 26370.0 17750.0 30455.0 ;
      RECT  20165.0 26370.0 20235.0 31255.0 ;
      RECT  20500.0 26370.0 20570.0 30455.0 ;
      RECT  22985.0 26370.0 23055.0 31255.0 ;
      RECT  23320.0 26370.0 23390.0 30455.0 ;
      RECT  25805.0 26370.0 25875.0 31255.0 ;
      RECT  26140.0 26370.0 26210.0 30455.0 ;
      RECT  28625.0 26370.0 28695.0 31255.0 ;
      RECT  28960.0 26370.0 29030.0 30455.0 ;
      RECT  31445.0 26370.0 31515.0 31255.0 ;
      RECT  31780.0 26370.0 31850.0 30455.0 ;
      RECT  34265.0 26370.0 34335.0 31255.0 ;
      RECT  34600.0 26370.0 34670.0 30455.0 ;
      RECT  37085.0 26370.0 37155.0 31255.0 ;
      RECT  37420.0 26370.0 37490.0 30455.0 ;
      RECT  39905.0 26370.0 39975.0 31255.0 ;
      RECT  40240.0 26370.0 40310.0 30455.0 ;
      RECT  42725.0 26370.0 42795.0 31255.0 ;
      RECT  43060.0 26370.0 43130.0 30455.0 ;
      RECT  45545.0 26370.0 45615.0 31255.0 ;
      RECT  45880.0 26370.0 45950.0 30455.0 ;
      RECT  48365.0 26370.0 48435.0 31255.0 ;
      RECT  48700.0 26370.0 48770.0 30455.0 ;
      RECT  51185.0 26370.0 51255.0 31255.0 ;
      RECT  51520.0 26370.0 51590.0 30455.0 ;
      RECT  54005.0 26370.0 54075.0 31255.0 ;
      RECT  54340.0 26370.0 54410.0 30455.0 ;
      RECT  56825.0 26370.0 56895.0 31255.0 ;
      RECT  57160.0 26370.0 57230.0 30455.0 ;
      RECT  59645.0 26370.0 59715.0 31255.0 ;
      RECT  59980.0 26370.0 60050.0 30455.0 ;
      RECT  62465.0 26370.0 62535.0 31255.0 ;
      RECT  62800.0 26370.0 62870.0 30455.0 ;
      RECT  65285.0 26370.0 65355.0 31255.0 ;
      RECT  65620.0 26370.0 65690.0 30455.0 ;
      RECT  68105.0 26370.0 68175.0 31255.0 ;
      RECT  68440.0 26370.0 68510.0 30455.0 ;
      RECT  70925.0 26370.0 70995.0 31255.0 ;
      RECT  71260.0 26370.0 71330.0 30455.0 ;
      RECT  73745.0 26370.0 73815.0 31255.0 ;
      RECT  74080.0 26370.0 74150.0 30455.0 ;
      RECT  76565.0 26370.0 76635.0 31255.0 ;
      RECT  76900.0 26370.0 76970.0 30455.0 ;
      RECT  79385.0 26370.0 79455.0 31255.0 ;
      RECT  79720.0 26370.0 79790.0 30455.0 ;
      RECT  82205.0 26370.0 82275.0 31255.0 ;
      RECT  82540.0 26370.0 82610.0 30455.0 ;
      RECT  85025.0 26370.0 85095.0 31255.0 ;
      RECT  85360.0 26370.0 85430.0 30455.0 ;
      RECT  87845.0 26370.0 87915.0 31255.0 ;
      RECT  88180.0 26370.0 88250.0 30455.0 ;
      RECT  90665.0 26370.0 90735.0 31255.0 ;
      RECT  91000.0 26370.0 91070.0 30455.0 ;
      RECT  93485.0 26370.0 93555.0 31255.0 ;
      RECT  93820.0 26370.0 93890.0 30455.0 ;
      RECT  96305.0 26370.0 96375.0 31255.0 ;
      RECT  96640.0 26370.0 96710.0 30455.0 ;
      RECT  99125.0 26370.0 99195.0 31255.0 ;
      RECT  99460.0 26370.0 99530.0 30455.0 ;
      RECT  101945.0 26370.0 102015.0 31255.0 ;
      RECT  102280.0 26370.0 102350.0 30455.0 ;
      RECT  104765.0 26370.0 104835.0 31255.0 ;
      RECT  105100.0 26370.0 105170.0 30455.0 ;
      RECT  17195.0 22195.0 17900.0 26370.0 ;
      RECT  20015.0 22195.0 20720.0 26370.0 ;
      RECT  22835.0 22195.0 23540.0 26370.0 ;
      RECT  25655.0 22195.0 26360.0 26370.0 ;
      RECT  28475.0 22195.0 29180.0 26370.0 ;
      RECT  31295.0 22195.0 32000.0 26370.0 ;
      RECT  34115.0 22195.0 34820.0 26370.0 ;
      RECT  36935.0 22195.0 37640.0 26370.0 ;
      RECT  39755.0 22195.0 40460.0 26370.0 ;
      RECT  42575.0 22195.0 43280.0 26370.0 ;
      RECT  45395.0 22195.0 46100.0 26370.0 ;
      RECT  48215.0 22195.0 48920.0 26370.0 ;
      RECT  51035.0 22195.0 51740.0 26370.0 ;
      RECT  53855.0 22195.0 54560.0 26370.0 ;
      RECT  56675.0 22195.0 57380.0 26370.0 ;
      RECT  59495.0 22195.0 60200.0 26370.0 ;
      RECT  62315.0 22195.0 63020.0 26370.0 ;
      RECT  65135.0 22195.0 65840.0 26370.0 ;
      RECT  67955.0 22195.0 68660.0 26370.0 ;
      RECT  70775.0 22195.0 71480.0 26370.0 ;
      RECT  73595.0 22195.0 74300.0 26370.0 ;
      RECT  76415.0 22195.0 77120.0 26370.0 ;
      RECT  79235.0 22195.0 79940.0 26370.0 ;
      RECT  82055.0 22195.0 82760.0 26370.0 ;
      RECT  84875.0 22195.0 85580.0 26370.0 ;
      RECT  87695.0 22195.0 88400.0 26370.0 ;
      RECT  90515.0 22195.0 91220.0 26370.0 ;
      RECT  93335.0 22195.0 94040.0 26370.0 ;
      RECT  96155.0 22195.0 96860.0 26370.0 ;
      RECT  98975.0 22195.0 99680.0 26370.0 ;
      RECT  101795.0 22195.0 102500.0 26370.0 ;
      RECT  104615.0 22195.0 105320.0 26370.0 ;
      RECT  17512.5 22195.0 17582.5 22335.0 ;
      RECT  20332.5 22195.0 20402.5 22335.0 ;
      RECT  23152.5 22195.0 23222.5 22335.0 ;
      RECT  25972.5 22195.0 26042.5 22335.0 ;
      RECT  28792.5 22195.0 28862.5 22335.0 ;
      RECT  31612.5 22195.0 31682.5 22335.0 ;
      RECT  34432.5 22195.0 34502.5 22335.0 ;
      RECT  37252.5 22195.0 37322.5 22335.0 ;
      RECT  40072.5 22195.0 40142.5 22335.0 ;
      RECT  42892.5 22195.0 42962.5 22335.0 ;
      RECT  45712.5 22195.0 45782.5 22335.0 ;
      RECT  48532.5 22195.0 48602.5 22335.0 ;
      RECT  51352.5 22195.0 51422.5 22335.0 ;
      RECT  54172.5 22195.0 54242.5 22335.0 ;
      RECT  56992.5 22195.0 57062.5 22335.0 ;
      RECT  59812.5 22195.0 59882.5 22335.0 ;
      RECT  62632.5 22195.0 62702.5 22335.0 ;
      RECT  65452.5 22195.0 65522.5 22335.0 ;
      RECT  68272.5 22195.0 68342.5 22335.0 ;
      RECT  71092.5 22195.0 71162.5 22335.0 ;
      RECT  73912.5 22195.0 73982.5 22335.0 ;
      RECT  76732.5 22195.0 76802.5 22335.0 ;
      RECT  79552.5 22195.0 79622.5 22335.0 ;
      RECT  82372.5 22195.0 82442.5 22335.0 ;
      RECT  85192.5 22195.0 85262.5 22335.0 ;
      RECT  88012.5 22195.0 88082.5 22335.0 ;
      RECT  90832.5 22195.0 90902.5 22335.0 ;
      RECT  93652.5 22195.0 93722.5 22335.0 ;
      RECT  96472.5 22195.0 96542.5 22335.0 ;
      RECT  99292.5 22195.0 99362.5 22335.0 ;
      RECT  102112.5 22195.0 102182.5 22335.0 ;
      RECT  104932.5 22195.0 105002.5 22335.0 ;
      RECT  17345.0 26070.0 17415.0 26370.0 ;
      RECT  17680.0 23930.0 17750.0 26370.0 ;
      RECT  20165.0 26070.0 20235.0 26370.0 ;
      RECT  20500.0 23930.0 20570.0 26370.0 ;
      RECT  22985.0 26070.0 23055.0 26370.0 ;
      RECT  23320.0 23930.0 23390.0 26370.0 ;
      RECT  25805.0 26070.0 25875.0 26370.0 ;
      RECT  26140.0 23930.0 26210.0 26370.0 ;
      RECT  28625.0 26070.0 28695.0 26370.0 ;
      RECT  28960.0 23930.0 29030.0 26370.0 ;
      RECT  31445.0 26070.0 31515.0 26370.0 ;
      RECT  31780.0 23930.0 31850.0 26370.0 ;
      RECT  34265.0 26070.0 34335.0 26370.0 ;
      RECT  34600.0 23930.0 34670.0 26370.0 ;
      RECT  37085.0 26070.0 37155.0 26370.0 ;
      RECT  37420.0 23930.0 37490.0 26370.0 ;
      RECT  39905.0 26070.0 39975.0 26370.0 ;
      RECT  40240.0 23930.0 40310.0 26370.0 ;
      RECT  42725.0 26070.0 42795.0 26370.0 ;
      RECT  43060.0 23930.0 43130.0 26370.0 ;
      RECT  45545.0 26070.0 45615.0 26370.0 ;
      RECT  45880.0 23930.0 45950.0 26370.0 ;
      RECT  48365.0 26070.0 48435.0 26370.0 ;
      RECT  48700.0 23930.0 48770.0 26370.0 ;
      RECT  51185.0 26070.0 51255.0 26370.0 ;
      RECT  51520.0 23930.0 51590.0 26370.0 ;
      RECT  54005.0 26070.0 54075.0 26370.0 ;
      RECT  54340.0 23930.0 54410.0 26370.0 ;
      RECT  56825.0 26070.0 56895.0 26370.0 ;
      RECT  57160.0 23930.0 57230.0 26370.0 ;
      RECT  59645.0 26070.0 59715.0 26370.0 ;
      RECT  59980.0 23930.0 60050.0 26370.0 ;
      RECT  62465.0 26070.0 62535.0 26370.0 ;
      RECT  62800.0 23930.0 62870.0 26370.0 ;
      RECT  65285.0 26070.0 65355.0 26370.0 ;
      RECT  65620.0 23930.0 65690.0 26370.0 ;
      RECT  68105.0 26070.0 68175.0 26370.0 ;
      RECT  68440.0 23930.0 68510.0 26370.0 ;
      RECT  70925.0 26070.0 70995.0 26370.0 ;
      RECT  71260.0 23930.0 71330.0 26370.0 ;
      RECT  73745.0 26070.0 73815.0 26370.0 ;
      RECT  74080.0 23930.0 74150.0 26370.0 ;
      RECT  76565.0 26070.0 76635.0 26370.0 ;
      RECT  76900.0 23930.0 76970.0 26370.0 ;
      RECT  79385.0 26070.0 79455.0 26370.0 ;
      RECT  79720.0 23930.0 79790.0 26370.0 ;
      RECT  82205.0 26070.0 82275.0 26370.0 ;
      RECT  82540.0 23930.0 82610.0 26370.0 ;
      RECT  85025.0 26070.0 85095.0 26370.0 ;
      RECT  85360.0 23930.0 85430.0 26370.0 ;
      RECT  87845.0 26070.0 87915.0 26370.0 ;
      RECT  88180.0 23930.0 88250.0 26370.0 ;
      RECT  90665.0 26070.0 90735.0 26370.0 ;
      RECT  91000.0 23930.0 91070.0 26370.0 ;
      RECT  93485.0 26070.0 93555.0 26370.0 ;
      RECT  93820.0 23930.0 93890.0 26370.0 ;
      RECT  96305.0 26070.0 96375.0 26370.0 ;
      RECT  96640.0 23930.0 96710.0 26370.0 ;
      RECT  99125.0 26070.0 99195.0 26370.0 ;
      RECT  99460.0 23930.0 99530.0 26370.0 ;
      RECT  101945.0 26070.0 102015.0 26370.0 ;
      RECT  102280.0 23930.0 102350.0 26370.0 ;
      RECT  104765.0 26070.0 104835.0 26370.0 ;
      RECT  105100.0 23930.0 105170.0 26370.0 ;
      RECT  17195.0 15755.0 17900.0 22195.0 ;
      RECT  20015.0 15755.0 20720.0 22195.0 ;
      RECT  22835.0 15755.0 23540.0 22195.0 ;
      RECT  25655.0 15755.0 26360.0 22195.0 ;
      RECT  28475.0 15755.0 29180.0 22195.0 ;
      RECT  31295.0 15755.0 32000.0 22195.0 ;
      RECT  34115.0 15755.0 34820.0 22195.0 ;
      RECT  36935.0 15755.0 37640.0 22195.0 ;
      RECT  39755.0 15755.0 40460.0 22195.0 ;
      RECT  42575.0 15755.0 43280.0 22195.0 ;
      RECT  45395.0 15755.0 46100.0 22195.0 ;
      RECT  48215.0 15755.0 48920.0 22195.0 ;
      RECT  51035.0 15755.0 51740.0 22195.0 ;
      RECT  53855.0 15755.0 54560.0 22195.0 ;
      RECT  56675.0 15755.0 57380.0 22195.0 ;
      RECT  59495.0 15755.0 60200.0 22195.0 ;
      RECT  62315.0 15755.0 63020.0 22195.0 ;
      RECT  65135.0 15755.0 65840.0 22195.0 ;
      RECT  67955.0 15755.0 68660.0 22195.0 ;
      RECT  70775.0 15755.0 71480.0 22195.0 ;
      RECT  73595.0 15755.0 74300.0 22195.0 ;
      RECT  76415.0 15755.0 77120.0 22195.0 ;
      RECT  79235.0 15755.0 79940.0 22195.0 ;
      RECT  82055.0 15755.0 82760.0 22195.0 ;
      RECT  84875.0 15755.0 85580.0 22195.0 ;
      RECT  87695.0 15755.0 88400.0 22195.0 ;
      RECT  90515.0 15755.0 91220.0 22195.0 ;
      RECT  93335.0 15755.0 94040.0 22195.0 ;
      RECT  96155.0 15755.0 96860.0 22195.0 ;
      RECT  98975.0 15755.0 99680.0 22195.0 ;
      RECT  101795.0 15755.0 102500.0 22195.0 ;
      RECT  104615.0 15755.0 105320.0 22195.0 ;
      RECT  17512.5 15755.0 17582.5 15900.0 ;
      RECT  20332.5 15755.0 20402.5 15900.0 ;
      RECT  23152.5 15755.0 23222.5 15900.0 ;
      RECT  25972.5 15755.0 26042.5 15900.0 ;
      RECT  28792.5 15755.0 28862.5 15900.0 ;
      RECT  31612.5 15755.0 31682.5 15900.0 ;
      RECT  34432.5 15755.0 34502.5 15900.0 ;
      RECT  37252.5 15755.0 37322.5 15900.0 ;
      RECT  40072.5 15755.0 40142.5 15900.0 ;
      RECT  42892.5 15755.0 42962.5 15900.0 ;
      RECT  45712.5 15755.0 45782.5 15900.0 ;
      RECT  48532.5 15755.0 48602.5 15900.0 ;
      RECT  51352.5 15755.0 51422.5 15900.0 ;
      RECT  54172.5 15755.0 54242.5 15900.0 ;
      RECT  56992.5 15755.0 57062.5 15900.0 ;
      RECT  59812.5 15755.0 59882.5 15900.0 ;
      RECT  62632.5 15755.0 62702.5 15900.0 ;
      RECT  65452.5 15755.0 65522.5 15900.0 ;
      RECT  68272.5 15755.0 68342.5 15900.0 ;
      RECT  71092.5 15755.0 71162.5 15900.0 ;
      RECT  73912.5 15755.0 73982.5 15900.0 ;
      RECT  76732.5 15755.0 76802.5 15900.0 ;
      RECT  79552.5 15755.0 79622.5 15900.0 ;
      RECT  82372.5 15755.0 82442.5 15900.0 ;
      RECT  85192.5 15755.0 85262.5 15900.0 ;
      RECT  88012.5 15755.0 88082.5 15900.0 ;
      RECT  90832.5 15755.0 90902.5 15900.0 ;
      RECT  93652.5 15755.0 93722.5 15900.0 ;
      RECT  96472.5 15755.0 96542.5 15900.0 ;
      RECT  99292.5 15755.0 99362.5 15900.0 ;
      RECT  102112.5 15755.0 102182.5 15900.0 ;
      RECT  104932.5 15755.0 105002.5 15900.0 ;
      RECT  17512.5 21925.0 17582.5 22195.0 ;
      RECT  17357.5 21507.5 17427.5 22195.0 ;
      RECT  20332.5 21925.0 20402.5 22195.0 ;
      RECT  20177.5 21507.5 20247.5 22195.0 ;
      RECT  23152.5 21925.0 23222.5 22195.0 ;
      RECT  22997.5 21507.5 23067.5 22195.0 ;
      RECT  25972.5 21925.0 26042.5 22195.0 ;
      RECT  25817.5 21507.5 25887.5 22195.0 ;
      RECT  28792.5 21925.0 28862.5 22195.0 ;
      RECT  28637.5 21507.5 28707.5 22195.0 ;
      RECT  31612.5 21925.0 31682.5 22195.0 ;
      RECT  31457.5 21507.5 31527.5 22195.0 ;
      RECT  34432.5 21925.0 34502.5 22195.0 ;
      RECT  34277.5 21507.5 34347.5 22195.0 ;
      RECT  37252.5 21925.0 37322.5 22195.0 ;
      RECT  37097.5 21507.5 37167.5 22195.0 ;
      RECT  40072.5 21925.0 40142.5 22195.0 ;
      RECT  39917.5 21507.5 39987.5 22195.0 ;
      RECT  42892.5 21925.0 42962.5 22195.0 ;
      RECT  42737.5 21507.5 42807.5 22195.0 ;
      RECT  45712.5 21925.0 45782.5 22195.0 ;
      RECT  45557.5 21507.5 45627.5 22195.0 ;
      RECT  48532.5 21925.0 48602.5 22195.0 ;
      RECT  48377.5 21507.5 48447.5 22195.0 ;
      RECT  51352.5 21925.0 51422.5 22195.0 ;
      RECT  51197.5 21507.5 51267.5 22195.0 ;
      RECT  54172.5 21925.0 54242.5 22195.0 ;
      RECT  54017.5 21507.5 54087.5 22195.0 ;
      RECT  56992.5 21925.0 57062.5 22195.0 ;
      RECT  56837.5 21507.5 56907.5 22195.0 ;
      RECT  59812.5 21925.0 59882.5 22195.0 ;
      RECT  59657.5 21507.5 59727.5 22195.0 ;
      RECT  62632.5 21925.0 62702.5 22195.0 ;
      RECT  62477.5 21507.5 62547.5 22195.0 ;
      RECT  65452.5 21925.0 65522.5 22195.0 ;
      RECT  65297.5 21507.5 65367.5 22195.0 ;
      RECT  68272.5 21925.0 68342.5 22195.0 ;
      RECT  68117.5 21507.5 68187.5 22195.0 ;
      RECT  71092.5 21925.0 71162.5 22195.0 ;
      RECT  70937.5 21507.5 71007.5 22195.0 ;
      RECT  73912.5 21925.0 73982.5 22195.0 ;
      RECT  73757.5 21507.5 73827.5 22195.0 ;
      RECT  76732.5 21925.0 76802.5 22195.0 ;
      RECT  76577.5 21507.5 76647.5 22195.0 ;
      RECT  79552.5 21925.0 79622.5 22195.0 ;
      RECT  79397.5 21507.5 79467.5 22195.0 ;
      RECT  82372.5 21925.0 82442.5 22195.0 ;
      RECT  82217.5 21507.5 82287.5 22195.0 ;
      RECT  85192.5 21925.0 85262.5 22195.0 ;
      RECT  85037.5 21507.5 85107.5 22195.0 ;
      RECT  88012.5 21925.0 88082.5 22195.0 ;
      RECT  87857.5 21507.5 87927.5 22195.0 ;
      RECT  90832.5 21925.0 90902.5 22195.0 ;
      RECT  90677.5 21507.5 90747.5 22195.0 ;
      RECT  93652.5 21925.0 93722.5 22195.0 ;
      RECT  93497.5 21507.5 93567.5 22195.0 ;
      RECT  96472.5 21925.0 96542.5 22195.0 ;
      RECT  96317.5 21507.5 96387.5 22195.0 ;
      RECT  99292.5 21925.0 99362.5 22195.0 ;
      RECT  99137.5 21507.5 99207.5 22195.0 ;
      RECT  102112.5 21925.0 102182.5 22195.0 ;
      RECT  101957.5 21507.5 102027.5 22195.0 ;
      RECT  104932.5 21925.0 105002.5 22195.0 ;
      RECT  104777.5 21507.5 104847.5 22195.0 ;
      RECT  17160.0 15755.0 17230.0 22195.0 ;
      RECT  17865.0 15755.0 17935.0 22195.0 ;
      RECT  19980.0 15755.0 20050.0 22195.0 ;
      RECT  20685.0 15755.0 20755.0 22195.0 ;
      RECT  22800.0 15755.0 22870.0 22195.0 ;
      RECT  23505.0 15755.0 23575.0 22195.0 ;
      RECT  25620.0 15755.0 25690.0 22195.0 ;
      RECT  26325.0 15755.0 26395.0 22195.0 ;
      RECT  28440.0 15755.0 28510.0 22195.0 ;
      RECT  29145.0 15755.0 29215.0 22195.0 ;
      RECT  31260.0 15755.0 31330.0 22195.0 ;
      RECT  31965.0 15755.0 32035.0 22195.0 ;
      RECT  34080.0 15755.0 34150.0 22195.0 ;
      RECT  34785.0 15755.0 34855.0 22195.0 ;
      RECT  36900.0 15755.0 36970.0 22195.0 ;
      RECT  37605.0 15755.0 37675.0 22195.0 ;
      RECT  39720.0 15755.0 39790.0 22195.0 ;
      RECT  40425.0 15755.0 40495.0 22195.0 ;
      RECT  42540.0 15755.0 42610.0 22195.0 ;
      RECT  43245.0 15755.0 43315.0 22195.0 ;
      RECT  45360.0 15755.0 45430.0 22195.0 ;
      RECT  46065.0 15755.0 46135.0 22195.0 ;
      RECT  48180.0 15755.0 48250.0 22195.0 ;
      RECT  48885.0 15755.0 48955.0 22195.0 ;
      RECT  51000.0 15755.0 51070.0 22195.0 ;
      RECT  51705.0 15755.0 51775.0 22195.0 ;
      RECT  53820.0 15755.0 53890.0 22195.0 ;
      RECT  54525.0 15755.0 54595.0 22195.0 ;
      RECT  56640.0 15755.0 56710.0 22195.0 ;
      RECT  57345.0 15755.0 57415.0 22195.0 ;
      RECT  59460.0 15755.0 59530.0 22195.0 ;
      RECT  60165.0 15755.0 60235.0 22195.0 ;
      RECT  62280.0 15755.0 62350.0 22195.0 ;
      RECT  62985.0 15755.0 63055.0 22195.0 ;
      RECT  65100.0 15755.0 65170.0 22195.0 ;
      RECT  65805.0 15755.0 65875.0 22195.0 ;
      RECT  67920.0 15755.0 67990.0 22195.0 ;
      RECT  68625.0 15755.0 68695.0 22195.0 ;
      RECT  70740.0 15755.0 70810.0 22195.0 ;
      RECT  71445.0 15755.0 71515.0 22195.0 ;
      RECT  73560.0 15755.0 73630.0 22195.0 ;
      RECT  74265.0 15755.0 74335.0 22195.0 ;
      RECT  76380.0 15755.0 76450.0 22195.0 ;
      RECT  77085.0 15755.0 77155.0 22195.0 ;
      RECT  79200.0 15755.0 79270.0 22195.0 ;
      RECT  79905.0 15755.0 79975.0 22195.0 ;
      RECT  82020.0 15755.0 82090.0 22195.0 ;
      RECT  82725.0 15755.0 82795.0 22195.0 ;
      RECT  84840.0 15755.0 84910.0 22195.0 ;
      RECT  85545.0 15755.0 85615.0 22195.0 ;
      RECT  87660.0 15755.0 87730.0 22195.0 ;
      RECT  88365.0 15755.0 88435.0 22195.0 ;
      RECT  90480.0 15755.0 90550.0 22195.0 ;
      RECT  91185.0 15755.0 91255.0 22195.0 ;
      RECT  93300.0 15755.0 93370.0 22195.0 ;
      RECT  94005.0 15755.0 94075.0 22195.0 ;
      RECT  96120.0 15755.0 96190.0 22195.0 ;
      RECT  96825.0 15755.0 96895.0 22195.0 ;
      RECT  98940.0 15755.0 99010.0 22195.0 ;
      RECT  99645.0 15755.0 99715.0 22195.0 ;
      RECT  101760.0 15755.0 101830.0 22195.0 ;
      RECT  102465.0 15755.0 102535.0 22195.0 ;
      RECT  104580.0 15755.0 104650.0 22195.0 ;
      RECT  105285.0 15755.0 105355.0 22195.0 ;
      RECT  17195.0 15755.0 17900.0 12780.0 ;
      RECT  20015.0 15755.0 20720.0 12780.0 ;
      RECT  22835.0 15755.0 23540.0 12780.0 ;
      RECT  25655.0 15755.0 26360.0 12780.0 ;
      RECT  28475.0 15755.0 29180.0 12780.0 ;
      RECT  31295.0 15755.0 32000.0 12780.0 ;
      RECT  34115.0 15755.0 34820.0 12780.0 ;
      RECT  36935.0 15755.0 37640.0 12780.0 ;
      RECT  39755.0 15755.0 40460.0 12780.0 ;
      RECT  42575.0 15755.0 43280.0 12780.0 ;
      RECT  45395.0 15755.0 46100.0 12780.0 ;
      RECT  48215.0 15755.0 48920.0 12780.0 ;
      RECT  51035.0 15755.0 51740.0 12780.0 ;
      RECT  53855.0 15755.0 54560.0 12780.0 ;
      RECT  56675.0 15755.0 57380.0 12780.0 ;
      RECT  59495.0 15755.0 60200.0 12780.0 ;
      RECT  62315.0 15755.0 63020.0 12780.0 ;
      RECT  65135.0 15755.0 65840.0 12780.0 ;
      RECT  67955.0 15755.0 68660.0 12780.0 ;
      RECT  70775.0 15755.0 71480.0 12780.0 ;
      RECT  73595.0 15755.0 74300.0 12780.0 ;
      RECT  76415.0 15755.0 77120.0 12780.0 ;
      RECT  79235.0 15755.0 79940.0 12780.0 ;
      RECT  82055.0 15755.0 82760.0 12780.0 ;
      RECT  84875.0 15755.0 85580.0 12780.0 ;
      RECT  87695.0 15755.0 88400.0 12780.0 ;
      RECT  90515.0 15755.0 91220.0 12780.0 ;
      RECT  93335.0 15755.0 94040.0 12780.0 ;
      RECT  96155.0 15755.0 96860.0 12780.0 ;
      RECT  98975.0 15755.0 99680.0 12780.0 ;
      RECT  101795.0 15755.0 102500.0 12780.0 ;
      RECT  104615.0 15755.0 105320.0 12780.0 ;
      RECT  17512.5 13020.0 17582.5 12780.0 ;
      RECT  20332.5 13020.0 20402.5 12780.0 ;
      RECT  23152.5 13020.0 23222.5 12780.0 ;
      RECT  25972.5 13020.0 26042.5 12780.0 ;
      RECT  28792.5 13020.0 28862.5 12780.0 ;
      RECT  31612.5 13020.0 31682.5 12780.0 ;
      RECT  34432.5 13020.0 34502.5 12780.0 ;
      RECT  37252.5 13020.0 37322.5 12780.0 ;
      RECT  40072.5 13020.0 40142.5 12780.0 ;
      RECT  42892.5 13020.0 42962.5 12780.0 ;
      RECT  45712.5 13020.0 45782.5 12780.0 ;
      RECT  48532.5 13020.0 48602.5 12780.0 ;
      RECT  51352.5 13020.0 51422.5 12780.0 ;
      RECT  54172.5 13020.0 54242.5 12780.0 ;
      RECT  56992.5 13020.0 57062.5 12780.0 ;
      RECT  59812.5 13020.0 59882.5 12780.0 ;
      RECT  62632.5 13020.0 62702.5 12780.0 ;
      RECT  65452.5 13020.0 65522.5 12780.0 ;
      RECT  68272.5 13020.0 68342.5 12780.0 ;
      RECT  71092.5 13020.0 71162.5 12780.0 ;
      RECT  73912.5 13020.0 73982.5 12780.0 ;
      RECT  76732.5 13020.0 76802.5 12780.0 ;
      RECT  79552.5 13020.0 79622.5 12780.0 ;
      RECT  82372.5 13020.0 82442.5 12780.0 ;
      RECT  85192.5 13020.0 85262.5 12780.0 ;
      RECT  88012.5 13020.0 88082.5 12780.0 ;
      RECT  90832.5 13020.0 90902.5 12780.0 ;
      RECT  93652.5 13020.0 93722.5 12780.0 ;
      RECT  96472.5 13020.0 96542.5 12780.0 ;
      RECT  99292.5 13020.0 99362.5 12780.0 ;
      RECT  102112.5 13020.0 102182.5 12780.0 ;
      RECT  104932.5 13020.0 105002.5 12780.0 ;
      RECT  17512.5 15755.0 17582.5 15405.0 ;
      RECT  20332.5 15755.0 20402.5 15405.0 ;
      RECT  23152.5 15755.0 23222.5 15405.0 ;
      RECT  25972.5 15755.0 26042.5 15405.0 ;
      RECT  28792.5 15755.0 28862.5 15405.0 ;
      RECT  31612.5 15755.0 31682.5 15405.0 ;
      RECT  34432.5 15755.0 34502.5 15405.0 ;
      RECT  37252.5 15755.0 37322.5 15405.0 ;
      RECT  40072.5 15755.0 40142.5 15405.0 ;
      RECT  42892.5 15755.0 42962.5 15405.0 ;
      RECT  45712.5 15755.0 45782.5 15405.0 ;
      RECT  48532.5 15755.0 48602.5 15405.0 ;
      RECT  51352.5 15755.0 51422.5 15405.0 ;
      RECT  54172.5 15755.0 54242.5 15405.0 ;
      RECT  56992.5 15755.0 57062.5 15405.0 ;
      RECT  59812.5 15755.0 59882.5 15405.0 ;
      RECT  62632.5 15755.0 62702.5 15405.0 ;
      RECT  65452.5 15755.0 65522.5 15405.0 ;
      RECT  68272.5 15755.0 68342.5 15405.0 ;
      RECT  71092.5 15755.0 71162.5 15405.0 ;
      RECT  73912.5 15755.0 73982.5 15405.0 ;
      RECT  76732.5 15755.0 76802.5 15405.0 ;
      RECT  79552.5 15755.0 79622.5 15405.0 ;
      RECT  82372.5 15755.0 82442.5 15405.0 ;
      RECT  85192.5 15755.0 85262.5 15405.0 ;
      RECT  88012.5 15755.0 88082.5 15405.0 ;
      RECT  90832.5 15755.0 90902.5 15405.0 ;
      RECT  93652.5 15755.0 93722.5 15405.0 ;
      RECT  96472.5 15755.0 96542.5 15405.0 ;
      RECT  99292.5 15755.0 99362.5 15405.0 ;
      RECT  102112.5 15755.0 102182.5 15405.0 ;
      RECT  104932.5 15755.0 105002.5 15405.0 ;
      RECT  4655.0 12580.0 4725.0 206260.0 ;
      RECT  4830.0 12580.0 4900.0 206260.0 ;
      RECT  5005.0 12580.0 5075.0 206260.0 ;
      RECT  5180.0 12580.0 5250.0 206260.0 ;
      RECT  5355.0 12580.0 5425.0 206260.0 ;
      RECT  5530.0 12580.0 5600.0 206260.0 ;
      RECT  5705.0 12580.0 5775.0 206260.0 ;
      RECT  5880.0 12580.0 5950.0 206260.0 ;
      RECT  6055.0 12580.0 6125.0 206260.0 ;
      RECT  6230.0 12580.0 6300.0 206260.0 ;
      RECT  6405.0 12580.0 6475.0 206260.0 ;
      RECT  6580.0 12580.0 6650.0 206260.0 ;
      RECT  6755.0 12580.0 6825.0 206260.0 ;
      RECT  6930.0 12580.0 7000.0 206260.0 ;
      RECT  7105.0 12580.0 7175.0 206260.0 ;
      RECT  7280.0 12580.0 7350.0 206260.0 ;
      RECT  9485.0 12580.0 9415.0 17820.0 ;
      RECT  9210.0 12580.0 9140.0 17820.0 ;
      RECT  10035.0 12580.0 9965.0 17820.0 ;
      RECT  9760.0 12580.0 9690.0 17820.0 ;
      RECT  8680.0 13185.0 8610.0 13255.0 ;
      RECT  8490.0 13185.0 8420.0 13255.0 ;
      RECT  8680.0 13220.0 8610.0 13582.5 ;
      RECT  8645.0 13185.0 8455.0 13255.0 ;
      RECT  8490.0 12877.5 8420.0 13220.0 ;
      RECT  8680.0 13582.5 8610.0 13717.5 ;
      RECT  8490.0 12742.5 8420.0 12877.5 ;
      RECT  8387.5 13185.0 8522.5 13255.0 ;
      RECT  8680.0 14665.0 8610.0 14595.0 ;
      RECT  8490.0 14665.0 8420.0 14595.0 ;
      RECT  8680.0 14630.0 8610.0 14267.5 ;
      RECT  8645.0 14665.0 8455.0 14595.0 ;
      RECT  8490.0 14972.5 8420.0 14630.0 ;
      RECT  8680.0 14267.5 8610.0 14132.5 ;
      RECT  8490.0 15107.5 8420.0 14972.5 ;
      RECT  8387.5 14665.0 8522.5 14595.0 ;
      RECT  8680.0 15875.0 8610.0 15945.0 ;
      RECT  8490.0 15875.0 8420.0 15945.0 ;
      RECT  8680.0 15910.0 8610.0 16272.5 ;
      RECT  8645.0 15875.0 8455.0 15945.0 ;
      RECT  8490.0 15567.5 8420.0 15910.0 ;
      RECT  8680.0 16272.5 8610.0 16407.5 ;
      RECT  8490.0 15432.5 8420.0 15567.5 ;
      RECT  8387.5 15875.0 8522.5 15945.0 ;
      RECT  8680.0 17355.0 8610.0 17285.0 ;
      RECT  8490.0 17355.0 8420.0 17285.0 ;
      RECT  8680.0 17320.0 8610.0 16957.5 ;
      RECT  8645.0 17355.0 8455.0 17285.0 ;
      RECT  8490.0 17662.5 8420.0 17320.0 ;
      RECT  8680.0 16957.5 8610.0 16822.5 ;
      RECT  8490.0 17797.5 8420.0 17662.5 ;
      RECT  8387.5 17355.0 8522.5 17285.0 ;
      RECT  9932.5 13695.0 10067.5 13765.0 ;
      RECT  11317.5 13172.5 11452.5 13242.5 ;
      RECT  9657.5 15040.0 9792.5 15110.0 ;
      RECT  11042.5 14607.5 11177.5 14677.5 ;
      RECT  11317.5 15370.0 11452.5 15440.0 ;
      RECT  9382.5 15370.0 9517.5 15440.0 ;
      RECT  11042.5 16715.0 11177.5 16785.0 ;
      RECT  9107.5 16715.0 9242.5 16785.0 ;
      RECT  9932.5 13185.0 10067.5 13255.0 ;
      RECT  9657.5 12970.0 9792.5 13040.0 ;
      RECT  9382.5 14595.0 9517.5 14665.0 ;
      RECT  9657.5 14810.0 9792.5 14880.0 ;
      RECT  9932.5 15875.0 10067.5 15945.0 ;
      RECT  9107.5 15660.0 9242.5 15730.0 ;
      RECT  9382.5 17285.0 9517.5 17355.0 ;
      RECT  9107.5 17500.0 9242.5 17570.0 ;
      RECT  11420.0 12580.0 11350.0 17820.0 ;
      RECT  11145.0 12580.0 11075.0 17820.0 ;
      RECT  9485.0 17960.0 9415.0 23200.0 ;
      RECT  9210.0 17960.0 9140.0 23200.0 ;
      RECT  10035.0 17960.0 9965.0 23200.0 ;
      RECT  9760.0 17960.0 9690.0 23200.0 ;
      RECT  8680.0 18565.0 8610.0 18635.0 ;
      RECT  8490.0 18565.0 8420.0 18635.0 ;
      RECT  8680.0 18600.0 8610.0 18962.5 ;
      RECT  8645.0 18565.0 8455.0 18635.0 ;
      RECT  8490.0 18257.5 8420.0 18600.0 ;
      RECT  8680.0 18962.5 8610.0 19097.5 ;
      RECT  8490.0 18122.5 8420.0 18257.5 ;
      RECT  8387.5 18565.0 8522.5 18635.0 ;
      RECT  8680.0 20045.0 8610.0 19975.0 ;
      RECT  8490.0 20045.0 8420.0 19975.0 ;
      RECT  8680.0 20010.0 8610.0 19647.5 ;
      RECT  8645.0 20045.0 8455.0 19975.0 ;
      RECT  8490.0 20352.5 8420.0 20010.0 ;
      RECT  8680.0 19647.5 8610.0 19512.5 ;
      RECT  8490.0 20487.5 8420.0 20352.5 ;
      RECT  8387.5 20045.0 8522.5 19975.0 ;
      RECT  8680.0 21255.0 8610.0 21325.0 ;
      RECT  8490.0 21255.0 8420.0 21325.0 ;
      RECT  8680.0 21290.0 8610.0 21652.5 ;
      RECT  8645.0 21255.0 8455.0 21325.0 ;
      RECT  8490.0 20947.5 8420.0 21290.0 ;
      RECT  8680.0 21652.5 8610.0 21787.5 ;
      RECT  8490.0 20812.5 8420.0 20947.5 ;
      RECT  8387.5 21255.0 8522.5 21325.0 ;
      RECT  8680.0 22735.0 8610.0 22665.0 ;
      RECT  8490.0 22735.0 8420.0 22665.0 ;
      RECT  8680.0 22700.0 8610.0 22337.5 ;
      RECT  8645.0 22735.0 8455.0 22665.0 ;
      RECT  8490.0 23042.5 8420.0 22700.0 ;
      RECT  8680.0 22337.5 8610.0 22202.5 ;
      RECT  8490.0 23177.5 8420.0 23042.5 ;
      RECT  8387.5 22735.0 8522.5 22665.0 ;
      RECT  9932.5 19075.0 10067.5 19145.0 ;
      RECT  11317.5 18552.5 11452.5 18622.5 ;
      RECT  9657.5 20420.0 9792.5 20490.0 ;
      RECT  11042.5 19987.5 11177.5 20057.5 ;
      RECT  11317.5 20750.0 11452.5 20820.0 ;
      RECT  9382.5 20750.0 9517.5 20820.0 ;
      RECT  11042.5 22095.0 11177.5 22165.0 ;
      RECT  9107.5 22095.0 9242.5 22165.0 ;
      RECT  9932.5 18565.0 10067.5 18635.0 ;
      RECT  9657.5 18350.0 9792.5 18420.0 ;
      RECT  9382.5 19975.0 9517.5 20045.0 ;
      RECT  9657.5 20190.0 9792.5 20260.0 ;
      RECT  9932.5 21255.0 10067.5 21325.0 ;
      RECT  9107.5 21040.0 9242.5 21110.0 ;
      RECT  9382.5 22665.0 9517.5 22735.0 ;
      RECT  9107.5 22880.0 9242.5 22950.0 ;
      RECT  11420.0 17960.0 11350.0 23200.0 ;
      RECT  11145.0 17960.0 11075.0 23200.0 ;
      RECT  10125.0 23340.0 10055.0 33960.0 ;
      RECT  9850.0 23340.0 9780.0 33960.0 ;
      RECT  9575.0 23340.0 9505.0 33960.0 ;
      RECT  10675.0 23340.0 10605.0 33960.0 ;
      RECT  10400.0 23340.0 10330.0 33960.0 ;
      RECT  9300.0 23340.0 9230.0 33960.0 ;
      RECT  8390.0 23637.5 8320.0 24342.5 ;
      RECT  8770.0 23992.5 8700.0 24062.5 ;
      RECT  8390.0 23992.5 8320.0 24062.5 ;
      RECT  8770.0 24027.5 8700.0 24342.5 ;
      RECT  8735.0 23992.5 8355.0 24062.5 ;
      RECT  8390.0 23637.5 8320.0 24027.5 ;
      RECT  8770.0 24342.5 8700.0 24477.5 ;
      RECT  8390.0 24342.5 8320.0 24477.5 ;
      RECT  8390.0 23502.5 8320.0 23637.5 ;
      RECT  8390.0 23960.0 8320.0 24095.0 ;
      RECT  8390.0 25732.5 8320.0 25027.5 ;
      RECT  8770.0 25377.5 8700.0 25307.5 ;
      RECT  8390.0 25377.5 8320.0 25307.5 ;
      RECT  8770.0 25342.5 8700.0 25027.5 ;
      RECT  8735.0 25377.5 8355.0 25307.5 ;
      RECT  8390.0 25732.5 8320.0 25342.5 ;
      RECT  8770.0 25027.5 8700.0 24892.5 ;
      RECT  8390.0 25027.5 8320.0 24892.5 ;
      RECT  8390.0 25867.5 8320.0 25732.5 ;
      RECT  8390.0 25410.0 8320.0 25275.0 ;
      RECT  8390.0 26327.5 8320.0 27032.5 ;
      RECT  8770.0 26682.5 8700.0 26752.5 ;
      RECT  8390.0 26682.5 8320.0 26752.5 ;
      RECT  8770.0 26717.5 8700.0 27032.5 ;
      RECT  8735.0 26682.5 8355.0 26752.5 ;
      RECT  8390.0 26327.5 8320.0 26717.5 ;
      RECT  8770.0 27032.5 8700.0 27167.5 ;
      RECT  8390.0 27032.5 8320.0 27167.5 ;
      RECT  8390.0 26192.5 8320.0 26327.5 ;
      RECT  8390.0 26650.0 8320.0 26785.0 ;
      RECT  8390.0 28422.5 8320.0 27717.5 ;
      RECT  8770.0 28067.5 8700.0 27997.5 ;
      RECT  8390.0 28067.5 8320.0 27997.5 ;
      RECT  8770.0 28032.5 8700.0 27717.5 ;
      RECT  8735.0 28067.5 8355.0 27997.5 ;
      RECT  8390.0 28422.5 8320.0 28032.5 ;
      RECT  8770.0 27717.5 8700.0 27582.5 ;
      RECT  8390.0 27717.5 8320.0 27582.5 ;
      RECT  8390.0 28557.5 8320.0 28422.5 ;
      RECT  8390.0 28100.0 8320.0 27965.0 ;
      RECT  8390.0 29017.5 8320.0 29722.5 ;
      RECT  8770.0 29372.5 8700.0 29442.5 ;
      RECT  8390.0 29372.5 8320.0 29442.5 ;
      RECT  8770.0 29407.5 8700.0 29722.5 ;
      RECT  8735.0 29372.5 8355.0 29442.5 ;
      RECT  8390.0 29017.5 8320.0 29407.5 ;
      RECT  8770.0 29722.5 8700.0 29857.5 ;
      RECT  8390.0 29722.5 8320.0 29857.5 ;
      RECT  8390.0 28882.5 8320.0 29017.5 ;
      RECT  8390.0 29340.0 8320.0 29475.0 ;
      RECT  8390.0 31112.5 8320.0 30407.5 ;
      RECT  8770.0 30757.5 8700.0 30687.5 ;
      RECT  8390.0 30757.5 8320.0 30687.5 ;
      RECT  8770.0 30722.5 8700.0 30407.5 ;
      RECT  8735.0 30757.5 8355.0 30687.5 ;
      RECT  8390.0 31112.5 8320.0 30722.5 ;
      RECT  8770.0 30407.5 8700.0 30272.5 ;
      RECT  8390.0 30407.5 8320.0 30272.5 ;
      RECT  8390.0 31247.5 8320.0 31112.5 ;
      RECT  8390.0 30790.0 8320.0 30655.0 ;
      RECT  8390.0 31707.5 8320.0 32412.5 ;
      RECT  8770.0 32062.5 8700.0 32132.5 ;
      RECT  8390.0 32062.5 8320.0 32132.5 ;
      RECT  8770.0 32097.5 8700.0 32412.5 ;
      RECT  8735.0 32062.5 8355.0 32132.5 ;
      RECT  8390.0 31707.5 8320.0 32097.5 ;
      RECT  8770.0 32412.5 8700.0 32547.5 ;
      RECT  8390.0 32412.5 8320.0 32547.5 ;
      RECT  8390.0 31572.5 8320.0 31707.5 ;
      RECT  8390.0 32030.0 8320.0 32165.0 ;
      RECT  8390.0 33802.5 8320.0 33097.5 ;
      RECT  8770.0 33447.5 8700.0 33377.5 ;
      RECT  8390.0 33447.5 8320.0 33377.5 ;
      RECT  8770.0 33412.5 8700.0 33097.5 ;
      RECT  8735.0 33447.5 8355.0 33377.5 ;
      RECT  8390.0 33802.5 8320.0 33412.5 ;
      RECT  8770.0 33097.5 8700.0 32962.5 ;
      RECT  8390.0 33097.5 8320.0 32962.5 ;
      RECT  8390.0 33937.5 8320.0 33802.5 ;
      RECT  8390.0 33480.0 8320.0 33345.0 ;
      RECT  10572.5 24455.0 10707.5 24525.0 ;
      RECT  12232.5 23932.5 12367.5 24002.5 ;
      RECT  10297.5 25800.0 10432.5 25870.0 ;
      RECT  11957.5 25367.5 12092.5 25437.5 ;
      RECT  10022.5 27145.0 10157.5 27215.0 ;
      RECT  11682.5 26622.5 11817.5 26692.5 ;
      RECT  12232.5 27475.0 12367.5 27545.0 ;
      RECT  9747.5 27475.0 9882.5 27545.0 ;
      RECT  11957.5 28820.0 12092.5 28890.0 ;
      RECT  9472.5 28820.0 9607.5 28890.0 ;
      RECT  11682.5 30165.0 11817.5 30235.0 ;
      RECT  9197.5 30165.0 9332.5 30235.0 ;
      RECT  10572.5 23992.5 10707.5 24062.5 ;
      RECT  10297.5 23852.5 10432.5 23922.5 ;
      RECT  10022.5 23712.5 10157.5 23782.5 ;
      RECT  9747.5 25307.5 9882.5 25377.5 ;
      RECT  10297.5 25447.5 10432.5 25517.5 ;
      RECT  10022.5 25587.5 10157.5 25657.5 ;
      RECT  10572.5 26682.5 10707.5 26752.5 ;
      RECT  9472.5 26542.5 9607.5 26612.5 ;
      RECT  10022.5 26402.5 10157.5 26472.5 ;
      RECT  9747.5 27997.5 9882.5 28067.5 ;
      RECT  9472.5 28137.5 9607.5 28207.5 ;
      RECT  10022.5 28277.5 10157.5 28347.5 ;
      RECT  10572.5 29372.5 10707.5 29442.5 ;
      RECT  10297.5 29232.5 10432.5 29302.5 ;
      RECT  9197.5 29092.5 9332.5 29162.5 ;
      RECT  9747.5 30687.5 9882.5 30757.5 ;
      RECT  10297.5 30827.5 10432.5 30897.5 ;
      RECT  9197.5 30967.5 9332.5 31037.5 ;
      RECT  10572.5 32062.5 10707.5 32132.5 ;
      RECT  9472.5 31922.5 9607.5 31992.5 ;
      RECT  9197.5 31782.5 9332.5 31852.5 ;
      RECT  9747.5 33377.5 9882.5 33447.5 ;
      RECT  9472.5 33517.5 9607.5 33587.5 ;
      RECT  9197.5 33657.5 9332.5 33727.5 ;
      RECT  12335.0 23340.0 12265.0 33960.0 ;
      RECT  12060.0 23340.0 11990.0 33960.0 ;
      RECT  11785.0 23340.0 11715.0 33960.0 ;
      RECT  8090.0 34397.5 8160.0 35102.5 ;
      RECT  7710.0 34752.5 7780.0 34822.5 ;
      RECT  8090.0 34752.5 8160.0 34822.5 ;
      RECT  7710.0 34787.5 7780.0 35102.5 ;
      RECT  7745.0 34752.5 8125.0 34822.5 ;
      RECT  8090.0 34397.5 8160.0 34787.5 ;
      RECT  7710.0 35102.5 7780.0 35237.5 ;
      RECT  8090.0 35102.5 8160.0 35237.5 ;
      RECT  8090.0 34262.5 8160.0 34397.5 ;
      RECT  8090.0 34720.0 8160.0 34855.0 ;
      RECT  8090.0 36492.5 8160.0 35787.5 ;
      RECT  7710.0 36137.5 7780.0 36067.5 ;
      RECT  8090.0 36137.5 8160.0 36067.5 ;
      RECT  7710.0 36102.5 7780.0 35787.5 ;
      RECT  7745.0 36137.5 8125.0 36067.5 ;
      RECT  8090.0 36492.5 8160.0 36102.5 ;
      RECT  7710.0 35787.5 7780.0 35652.5 ;
      RECT  8090.0 35787.5 8160.0 35652.5 ;
      RECT  8090.0 36627.5 8160.0 36492.5 ;
      RECT  8090.0 36170.0 8160.0 36035.0 ;
      RECT  8090.0 37087.5 8160.0 37792.5 ;
      RECT  7710.0 37442.5 7780.0 37512.5 ;
      RECT  8090.0 37442.5 8160.0 37512.5 ;
      RECT  7710.0 37477.5 7780.0 37792.5 ;
      RECT  7745.0 37442.5 8125.0 37512.5 ;
      RECT  8090.0 37087.5 8160.0 37477.5 ;
      RECT  7710.0 37792.5 7780.0 37927.5 ;
      RECT  8090.0 37792.5 8160.0 37927.5 ;
      RECT  8090.0 36952.5 8160.0 37087.5 ;
      RECT  8090.0 37410.0 8160.0 37545.0 ;
      RECT  8090.0 39182.5 8160.0 38477.5 ;
      RECT  7710.0 38827.5 7780.0 38757.5 ;
      RECT  8090.0 38827.5 8160.0 38757.5 ;
      RECT  7710.0 38792.5 7780.0 38477.5 ;
      RECT  7745.0 38827.5 8125.0 38757.5 ;
      RECT  8090.0 39182.5 8160.0 38792.5 ;
      RECT  7710.0 38477.5 7780.0 38342.5 ;
      RECT  8090.0 38477.5 8160.0 38342.5 ;
      RECT  8090.0 39317.5 8160.0 39182.5 ;
      RECT  8090.0 38860.0 8160.0 38725.0 ;
      RECT  8090.0 39777.5 8160.0 40482.5 ;
      RECT  7710.0 40132.5 7780.0 40202.5 ;
      RECT  8090.0 40132.5 8160.0 40202.5 ;
      RECT  7710.0 40167.5 7780.0 40482.5 ;
      RECT  7745.0 40132.5 8125.0 40202.5 ;
      RECT  8090.0 39777.5 8160.0 40167.5 ;
      RECT  7710.0 40482.5 7780.0 40617.5 ;
      RECT  8090.0 40482.5 8160.0 40617.5 ;
      RECT  8090.0 39642.5 8160.0 39777.5 ;
      RECT  8090.0 40100.0 8160.0 40235.0 ;
      RECT  8090.0 41872.5 8160.0 41167.5 ;
      RECT  7710.0 41517.5 7780.0 41447.5 ;
      RECT  8090.0 41517.5 8160.0 41447.5 ;
      RECT  7710.0 41482.5 7780.0 41167.5 ;
      RECT  7745.0 41517.5 8125.0 41447.5 ;
      RECT  8090.0 41872.5 8160.0 41482.5 ;
      RECT  7710.0 41167.5 7780.0 41032.5 ;
      RECT  8090.0 41167.5 8160.0 41032.5 ;
      RECT  8090.0 42007.5 8160.0 41872.5 ;
      RECT  8090.0 41550.0 8160.0 41415.0 ;
      RECT  8090.0 42467.5 8160.0 43172.5 ;
      RECT  7710.0 42822.5 7780.0 42892.5 ;
      RECT  8090.0 42822.5 8160.0 42892.5 ;
      RECT  7710.0 42857.5 7780.0 43172.5 ;
      RECT  7745.0 42822.5 8125.0 42892.5 ;
      RECT  8090.0 42467.5 8160.0 42857.5 ;
      RECT  7710.0 43172.5 7780.0 43307.5 ;
      RECT  8090.0 43172.5 8160.0 43307.5 ;
      RECT  8090.0 42332.5 8160.0 42467.5 ;
      RECT  8090.0 42790.0 8160.0 42925.0 ;
      RECT  8090.0 44562.5 8160.0 43857.5 ;
      RECT  7710.0 44207.5 7780.0 44137.5 ;
      RECT  8090.0 44207.5 8160.0 44137.5 ;
      RECT  7710.0 44172.5 7780.0 43857.5 ;
      RECT  7745.0 44207.5 8125.0 44137.5 ;
      RECT  8090.0 44562.5 8160.0 44172.5 ;
      RECT  7710.0 43857.5 7780.0 43722.5 ;
      RECT  8090.0 43857.5 8160.0 43722.5 ;
      RECT  8090.0 44697.5 8160.0 44562.5 ;
      RECT  8090.0 44240.0 8160.0 44105.0 ;
      RECT  8090.0 45157.5 8160.0 45862.5 ;
      RECT  7710.0 45512.5 7780.0 45582.5 ;
      RECT  8090.0 45512.5 8160.0 45582.5 ;
      RECT  7710.0 45547.5 7780.0 45862.5 ;
      RECT  7745.0 45512.5 8125.0 45582.5 ;
      RECT  8090.0 45157.5 8160.0 45547.5 ;
      RECT  7710.0 45862.5 7780.0 45997.5 ;
      RECT  8090.0 45862.5 8160.0 45997.5 ;
      RECT  8090.0 45022.5 8160.0 45157.5 ;
      RECT  8090.0 45480.0 8160.0 45615.0 ;
      RECT  8090.0 47252.5 8160.0 46547.5 ;
      RECT  7710.0 46897.5 7780.0 46827.5 ;
      RECT  8090.0 46897.5 8160.0 46827.5 ;
      RECT  7710.0 46862.5 7780.0 46547.5 ;
      RECT  7745.0 46897.5 8125.0 46827.5 ;
      RECT  8090.0 47252.5 8160.0 46862.5 ;
      RECT  7710.0 46547.5 7780.0 46412.5 ;
      RECT  8090.0 46547.5 8160.0 46412.5 ;
      RECT  8090.0 47387.5 8160.0 47252.5 ;
      RECT  8090.0 46930.0 8160.0 46795.0 ;
      RECT  8090.0 47847.5 8160.0 48552.5 ;
      RECT  7710.0 48202.5 7780.0 48272.5 ;
      RECT  8090.0 48202.5 8160.0 48272.5 ;
      RECT  7710.0 48237.5 7780.0 48552.5 ;
      RECT  7745.0 48202.5 8125.0 48272.5 ;
      RECT  8090.0 47847.5 8160.0 48237.5 ;
      RECT  7710.0 48552.5 7780.0 48687.5 ;
      RECT  8090.0 48552.5 8160.0 48687.5 ;
      RECT  8090.0 47712.5 8160.0 47847.5 ;
      RECT  8090.0 48170.0 8160.0 48305.0 ;
      RECT  8090.0 49942.5 8160.0 49237.5 ;
      RECT  7710.0 49587.5 7780.0 49517.5 ;
      RECT  8090.0 49587.5 8160.0 49517.5 ;
      RECT  7710.0 49552.5 7780.0 49237.5 ;
      RECT  7745.0 49587.5 8125.0 49517.5 ;
      RECT  8090.0 49942.5 8160.0 49552.5 ;
      RECT  7710.0 49237.5 7780.0 49102.5 ;
      RECT  8090.0 49237.5 8160.0 49102.5 ;
      RECT  8090.0 50077.5 8160.0 49942.5 ;
      RECT  8090.0 49620.0 8160.0 49485.0 ;
      RECT  8090.0 50537.5 8160.0 51242.5 ;
      RECT  7710.0 50892.5 7780.0 50962.5 ;
      RECT  8090.0 50892.5 8160.0 50962.5 ;
      RECT  7710.0 50927.5 7780.0 51242.5 ;
      RECT  7745.0 50892.5 8125.0 50962.5 ;
      RECT  8090.0 50537.5 8160.0 50927.5 ;
      RECT  7710.0 51242.5 7780.0 51377.5 ;
      RECT  8090.0 51242.5 8160.0 51377.5 ;
      RECT  8090.0 50402.5 8160.0 50537.5 ;
      RECT  8090.0 50860.0 8160.0 50995.0 ;
      RECT  8090.0 52632.5 8160.0 51927.5 ;
      RECT  7710.0 52277.5 7780.0 52207.5 ;
      RECT  8090.0 52277.5 8160.0 52207.5 ;
      RECT  7710.0 52242.5 7780.0 51927.5 ;
      RECT  7745.0 52277.5 8125.0 52207.5 ;
      RECT  8090.0 52632.5 8160.0 52242.5 ;
      RECT  7710.0 51927.5 7780.0 51792.5 ;
      RECT  8090.0 51927.5 8160.0 51792.5 ;
      RECT  8090.0 52767.5 8160.0 52632.5 ;
      RECT  8090.0 52310.0 8160.0 52175.0 ;
      RECT  8090.0 53227.5 8160.0 53932.5 ;
      RECT  7710.0 53582.5 7780.0 53652.5 ;
      RECT  8090.0 53582.5 8160.0 53652.5 ;
      RECT  7710.0 53617.5 7780.0 53932.5 ;
      RECT  7745.0 53582.5 8125.0 53652.5 ;
      RECT  8090.0 53227.5 8160.0 53617.5 ;
      RECT  7710.0 53932.5 7780.0 54067.5 ;
      RECT  8090.0 53932.5 8160.0 54067.5 ;
      RECT  8090.0 53092.5 8160.0 53227.5 ;
      RECT  8090.0 53550.0 8160.0 53685.0 ;
      RECT  8090.0 55322.5 8160.0 54617.5 ;
      RECT  7710.0 54967.5 7780.0 54897.5 ;
      RECT  8090.0 54967.5 8160.0 54897.5 ;
      RECT  7710.0 54932.5 7780.0 54617.5 ;
      RECT  7745.0 54967.5 8125.0 54897.5 ;
      RECT  8090.0 55322.5 8160.0 54932.5 ;
      RECT  7710.0 54617.5 7780.0 54482.5 ;
      RECT  8090.0 54617.5 8160.0 54482.5 ;
      RECT  8090.0 55457.5 8160.0 55322.5 ;
      RECT  8090.0 55000.0 8160.0 54865.0 ;
      RECT  8090.0 55917.5 8160.0 56622.5 ;
      RECT  7710.0 56272.5 7780.0 56342.5 ;
      RECT  8090.0 56272.5 8160.0 56342.5 ;
      RECT  7710.0 56307.5 7780.0 56622.5 ;
      RECT  7745.0 56272.5 8125.0 56342.5 ;
      RECT  8090.0 55917.5 8160.0 56307.5 ;
      RECT  7710.0 56622.5 7780.0 56757.5 ;
      RECT  8090.0 56622.5 8160.0 56757.5 ;
      RECT  8090.0 55782.5 8160.0 55917.5 ;
      RECT  8090.0 56240.0 8160.0 56375.0 ;
      RECT  8090.0 58012.5 8160.0 57307.5 ;
      RECT  7710.0 57657.5 7780.0 57587.5 ;
      RECT  8090.0 57657.5 8160.0 57587.5 ;
      RECT  7710.0 57622.5 7780.0 57307.5 ;
      RECT  7745.0 57657.5 8125.0 57587.5 ;
      RECT  8090.0 58012.5 8160.0 57622.5 ;
      RECT  7710.0 57307.5 7780.0 57172.5 ;
      RECT  8090.0 57307.5 8160.0 57172.5 ;
      RECT  8090.0 58147.5 8160.0 58012.5 ;
      RECT  8090.0 57690.0 8160.0 57555.0 ;
      RECT  8090.0 58607.5 8160.0 59312.5 ;
      RECT  7710.0 58962.5 7780.0 59032.5 ;
      RECT  8090.0 58962.5 8160.0 59032.5 ;
      RECT  7710.0 58997.5 7780.0 59312.5 ;
      RECT  7745.0 58962.5 8125.0 59032.5 ;
      RECT  8090.0 58607.5 8160.0 58997.5 ;
      RECT  7710.0 59312.5 7780.0 59447.5 ;
      RECT  8090.0 59312.5 8160.0 59447.5 ;
      RECT  8090.0 58472.5 8160.0 58607.5 ;
      RECT  8090.0 58930.0 8160.0 59065.0 ;
      RECT  8090.0 60702.5 8160.0 59997.5 ;
      RECT  7710.0 60347.5 7780.0 60277.5 ;
      RECT  8090.0 60347.5 8160.0 60277.5 ;
      RECT  7710.0 60312.5 7780.0 59997.5 ;
      RECT  7745.0 60347.5 8125.0 60277.5 ;
      RECT  8090.0 60702.5 8160.0 60312.5 ;
      RECT  7710.0 59997.5 7780.0 59862.5 ;
      RECT  8090.0 59997.5 8160.0 59862.5 ;
      RECT  8090.0 60837.5 8160.0 60702.5 ;
      RECT  8090.0 60380.0 8160.0 60245.0 ;
      RECT  8090.0 61297.5 8160.0 62002.5 ;
      RECT  7710.0 61652.5 7780.0 61722.5 ;
      RECT  8090.0 61652.5 8160.0 61722.5 ;
      RECT  7710.0 61687.5 7780.0 62002.5 ;
      RECT  7745.0 61652.5 8125.0 61722.5 ;
      RECT  8090.0 61297.5 8160.0 61687.5 ;
      RECT  7710.0 62002.5 7780.0 62137.5 ;
      RECT  8090.0 62002.5 8160.0 62137.5 ;
      RECT  8090.0 61162.5 8160.0 61297.5 ;
      RECT  8090.0 61620.0 8160.0 61755.0 ;
      RECT  8090.0 63392.5 8160.0 62687.5 ;
      RECT  7710.0 63037.5 7780.0 62967.5 ;
      RECT  8090.0 63037.5 8160.0 62967.5 ;
      RECT  7710.0 63002.5 7780.0 62687.5 ;
      RECT  7745.0 63037.5 8125.0 62967.5 ;
      RECT  8090.0 63392.5 8160.0 63002.5 ;
      RECT  7710.0 62687.5 7780.0 62552.5 ;
      RECT  8090.0 62687.5 8160.0 62552.5 ;
      RECT  8090.0 63527.5 8160.0 63392.5 ;
      RECT  8090.0 63070.0 8160.0 62935.0 ;
      RECT  8090.0 63987.5 8160.0 64692.5 ;
      RECT  7710.0 64342.5 7780.0 64412.5 ;
      RECT  8090.0 64342.5 8160.0 64412.5 ;
      RECT  7710.0 64377.5 7780.0 64692.5 ;
      RECT  7745.0 64342.5 8125.0 64412.5 ;
      RECT  8090.0 63987.5 8160.0 64377.5 ;
      RECT  7710.0 64692.5 7780.0 64827.5 ;
      RECT  8090.0 64692.5 8160.0 64827.5 ;
      RECT  8090.0 63852.5 8160.0 63987.5 ;
      RECT  8090.0 64310.0 8160.0 64445.0 ;
      RECT  8090.0 66082.5 8160.0 65377.5 ;
      RECT  7710.0 65727.5 7780.0 65657.5 ;
      RECT  8090.0 65727.5 8160.0 65657.5 ;
      RECT  7710.0 65692.5 7780.0 65377.5 ;
      RECT  7745.0 65727.5 8125.0 65657.5 ;
      RECT  8090.0 66082.5 8160.0 65692.5 ;
      RECT  7710.0 65377.5 7780.0 65242.5 ;
      RECT  8090.0 65377.5 8160.0 65242.5 ;
      RECT  8090.0 66217.5 8160.0 66082.5 ;
      RECT  8090.0 65760.0 8160.0 65625.0 ;
      RECT  8090.0 66677.5 8160.0 67382.5 ;
      RECT  7710.0 67032.5 7780.0 67102.5 ;
      RECT  8090.0 67032.5 8160.0 67102.5 ;
      RECT  7710.0 67067.5 7780.0 67382.5 ;
      RECT  7745.0 67032.5 8125.0 67102.5 ;
      RECT  8090.0 66677.5 8160.0 67067.5 ;
      RECT  7710.0 67382.5 7780.0 67517.5 ;
      RECT  8090.0 67382.5 8160.0 67517.5 ;
      RECT  8090.0 66542.5 8160.0 66677.5 ;
      RECT  8090.0 67000.0 8160.0 67135.0 ;
      RECT  8090.0 68772.5 8160.0 68067.5 ;
      RECT  7710.0 68417.5 7780.0 68347.5 ;
      RECT  8090.0 68417.5 8160.0 68347.5 ;
      RECT  7710.0 68382.5 7780.0 68067.5 ;
      RECT  7745.0 68417.5 8125.0 68347.5 ;
      RECT  8090.0 68772.5 8160.0 68382.5 ;
      RECT  7710.0 68067.5 7780.0 67932.5 ;
      RECT  8090.0 68067.5 8160.0 67932.5 ;
      RECT  8090.0 68907.5 8160.0 68772.5 ;
      RECT  8090.0 68450.0 8160.0 68315.0 ;
      RECT  8090.0 69367.5 8160.0 70072.5 ;
      RECT  7710.0 69722.5 7780.0 69792.5 ;
      RECT  8090.0 69722.5 8160.0 69792.5 ;
      RECT  7710.0 69757.5 7780.0 70072.5 ;
      RECT  7745.0 69722.5 8125.0 69792.5 ;
      RECT  8090.0 69367.5 8160.0 69757.5 ;
      RECT  7710.0 70072.5 7780.0 70207.5 ;
      RECT  8090.0 70072.5 8160.0 70207.5 ;
      RECT  8090.0 69232.5 8160.0 69367.5 ;
      RECT  8090.0 69690.0 8160.0 69825.0 ;
      RECT  8090.0 71462.5 8160.0 70757.5 ;
      RECT  7710.0 71107.5 7780.0 71037.5 ;
      RECT  8090.0 71107.5 8160.0 71037.5 ;
      RECT  7710.0 71072.5 7780.0 70757.5 ;
      RECT  7745.0 71107.5 8125.0 71037.5 ;
      RECT  8090.0 71462.5 8160.0 71072.5 ;
      RECT  7710.0 70757.5 7780.0 70622.5 ;
      RECT  8090.0 70757.5 8160.0 70622.5 ;
      RECT  8090.0 71597.5 8160.0 71462.5 ;
      RECT  8090.0 71140.0 8160.0 71005.0 ;
      RECT  8090.0 72057.5 8160.0 72762.5 ;
      RECT  7710.0 72412.5 7780.0 72482.5 ;
      RECT  8090.0 72412.5 8160.0 72482.5 ;
      RECT  7710.0 72447.5 7780.0 72762.5 ;
      RECT  7745.0 72412.5 8125.0 72482.5 ;
      RECT  8090.0 72057.5 8160.0 72447.5 ;
      RECT  7710.0 72762.5 7780.0 72897.5 ;
      RECT  8090.0 72762.5 8160.0 72897.5 ;
      RECT  8090.0 71922.5 8160.0 72057.5 ;
      RECT  8090.0 72380.0 8160.0 72515.0 ;
      RECT  8090.0 74152.5 8160.0 73447.5 ;
      RECT  7710.0 73797.5 7780.0 73727.5 ;
      RECT  8090.0 73797.5 8160.0 73727.5 ;
      RECT  7710.0 73762.5 7780.0 73447.5 ;
      RECT  7745.0 73797.5 8125.0 73727.5 ;
      RECT  8090.0 74152.5 8160.0 73762.5 ;
      RECT  7710.0 73447.5 7780.0 73312.5 ;
      RECT  8090.0 73447.5 8160.0 73312.5 ;
      RECT  8090.0 74287.5 8160.0 74152.5 ;
      RECT  8090.0 73830.0 8160.0 73695.0 ;
      RECT  8090.0 74747.5 8160.0 75452.5 ;
      RECT  7710.0 75102.5 7780.0 75172.5 ;
      RECT  8090.0 75102.5 8160.0 75172.5 ;
      RECT  7710.0 75137.5 7780.0 75452.5 ;
      RECT  7745.0 75102.5 8125.0 75172.5 ;
      RECT  8090.0 74747.5 8160.0 75137.5 ;
      RECT  7710.0 75452.5 7780.0 75587.5 ;
      RECT  8090.0 75452.5 8160.0 75587.5 ;
      RECT  8090.0 74612.5 8160.0 74747.5 ;
      RECT  8090.0 75070.0 8160.0 75205.0 ;
      RECT  8090.0 76842.5 8160.0 76137.5 ;
      RECT  7710.0 76487.5 7780.0 76417.5 ;
      RECT  8090.0 76487.5 8160.0 76417.5 ;
      RECT  7710.0 76452.5 7780.0 76137.5 ;
      RECT  7745.0 76487.5 8125.0 76417.5 ;
      RECT  8090.0 76842.5 8160.0 76452.5 ;
      RECT  7710.0 76137.5 7780.0 76002.5 ;
      RECT  8090.0 76137.5 8160.0 76002.5 ;
      RECT  8090.0 76977.5 8160.0 76842.5 ;
      RECT  8090.0 76520.0 8160.0 76385.0 ;
      RECT  8090.0 77437.5 8160.0 78142.5 ;
      RECT  7710.0 77792.5 7780.0 77862.5 ;
      RECT  8090.0 77792.5 8160.0 77862.5 ;
      RECT  7710.0 77827.5 7780.0 78142.5 ;
      RECT  7745.0 77792.5 8125.0 77862.5 ;
      RECT  8090.0 77437.5 8160.0 77827.5 ;
      RECT  7710.0 78142.5 7780.0 78277.5 ;
      RECT  8090.0 78142.5 8160.0 78277.5 ;
      RECT  8090.0 77302.5 8160.0 77437.5 ;
      RECT  8090.0 77760.0 8160.0 77895.0 ;
      RECT  8090.0 79532.5 8160.0 78827.5 ;
      RECT  7710.0 79177.5 7780.0 79107.5 ;
      RECT  8090.0 79177.5 8160.0 79107.5 ;
      RECT  7710.0 79142.5 7780.0 78827.5 ;
      RECT  7745.0 79177.5 8125.0 79107.5 ;
      RECT  8090.0 79532.5 8160.0 79142.5 ;
      RECT  7710.0 78827.5 7780.0 78692.5 ;
      RECT  8090.0 78827.5 8160.0 78692.5 ;
      RECT  8090.0 79667.5 8160.0 79532.5 ;
      RECT  8090.0 79210.0 8160.0 79075.0 ;
      RECT  8090.0 80127.5 8160.0 80832.5 ;
      RECT  7710.0 80482.5 7780.0 80552.5 ;
      RECT  8090.0 80482.5 8160.0 80552.5 ;
      RECT  7710.0 80517.5 7780.0 80832.5 ;
      RECT  7745.0 80482.5 8125.0 80552.5 ;
      RECT  8090.0 80127.5 8160.0 80517.5 ;
      RECT  7710.0 80832.5 7780.0 80967.5 ;
      RECT  8090.0 80832.5 8160.0 80967.5 ;
      RECT  8090.0 79992.5 8160.0 80127.5 ;
      RECT  8090.0 80450.0 8160.0 80585.0 ;
      RECT  8090.0 82222.5 8160.0 81517.5 ;
      RECT  7710.0 81867.5 7780.0 81797.5 ;
      RECT  8090.0 81867.5 8160.0 81797.5 ;
      RECT  7710.0 81832.5 7780.0 81517.5 ;
      RECT  7745.0 81867.5 8125.0 81797.5 ;
      RECT  8090.0 82222.5 8160.0 81832.5 ;
      RECT  7710.0 81517.5 7780.0 81382.5 ;
      RECT  8090.0 81517.5 8160.0 81382.5 ;
      RECT  8090.0 82357.5 8160.0 82222.5 ;
      RECT  8090.0 81900.0 8160.0 81765.0 ;
      RECT  8090.0 82817.5 8160.0 83522.5 ;
      RECT  7710.0 83172.5 7780.0 83242.5 ;
      RECT  8090.0 83172.5 8160.0 83242.5 ;
      RECT  7710.0 83207.5 7780.0 83522.5 ;
      RECT  7745.0 83172.5 8125.0 83242.5 ;
      RECT  8090.0 82817.5 8160.0 83207.5 ;
      RECT  7710.0 83522.5 7780.0 83657.5 ;
      RECT  8090.0 83522.5 8160.0 83657.5 ;
      RECT  8090.0 82682.5 8160.0 82817.5 ;
      RECT  8090.0 83140.0 8160.0 83275.0 ;
      RECT  8090.0 84912.5 8160.0 84207.5 ;
      RECT  7710.0 84557.5 7780.0 84487.5 ;
      RECT  8090.0 84557.5 8160.0 84487.5 ;
      RECT  7710.0 84522.5 7780.0 84207.5 ;
      RECT  7745.0 84557.5 8125.0 84487.5 ;
      RECT  8090.0 84912.5 8160.0 84522.5 ;
      RECT  7710.0 84207.5 7780.0 84072.5 ;
      RECT  8090.0 84207.5 8160.0 84072.5 ;
      RECT  8090.0 85047.5 8160.0 84912.5 ;
      RECT  8090.0 84590.0 8160.0 84455.0 ;
      RECT  8090.0 85507.5 8160.0 86212.5 ;
      RECT  7710.0 85862.5 7780.0 85932.5 ;
      RECT  8090.0 85862.5 8160.0 85932.5 ;
      RECT  7710.0 85897.5 7780.0 86212.5 ;
      RECT  7745.0 85862.5 8125.0 85932.5 ;
      RECT  8090.0 85507.5 8160.0 85897.5 ;
      RECT  7710.0 86212.5 7780.0 86347.5 ;
      RECT  8090.0 86212.5 8160.0 86347.5 ;
      RECT  8090.0 85372.5 8160.0 85507.5 ;
      RECT  8090.0 85830.0 8160.0 85965.0 ;
      RECT  8090.0 87602.5 8160.0 86897.5 ;
      RECT  7710.0 87247.5 7780.0 87177.5 ;
      RECT  8090.0 87247.5 8160.0 87177.5 ;
      RECT  7710.0 87212.5 7780.0 86897.5 ;
      RECT  7745.0 87247.5 8125.0 87177.5 ;
      RECT  8090.0 87602.5 8160.0 87212.5 ;
      RECT  7710.0 86897.5 7780.0 86762.5 ;
      RECT  8090.0 86897.5 8160.0 86762.5 ;
      RECT  8090.0 87737.5 8160.0 87602.5 ;
      RECT  8090.0 87280.0 8160.0 87145.0 ;
      RECT  8090.0 88197.5 8160.0 88902.5 ;
      RECT  7710.0 88552.5 7780.0 88622.5 ;
      RECT  8090.0 88552.5 8160.0 88622.5 ;
      RECT  7710.0 88587.5 7780.0 88902.5 ;
      RECT  7745.0 88552.5 8125.0 88622.5 ;
      RECT  8090.0 88197.5 8160.0 88587.5 ;
      RECT  7710.0 88902.5 7780.0 89037.5 ;
      RECT  8090.0 88902.5 8160.0 89037.5 ;
      RECT  8090.0 88062.5 8160.0 88197.5 ;
      RECT  8090.0 88520.0 8160.0 88655.0 ;
      RECT  8090.0 90292.5 8160.0 89587.5 ;
      RECT  7710.0 89937.5 7780.0 89867.5 ;
      RECT  8090.0 89937.5 8160.0 89867.5 ;
      RECT  7710.0 89902.5 7780.0 89587.5 ;
      RECT  7745.0 89937.5 8125.0 89867.5 ;
      RECT  8090.0 90292.5 8160.0 89902.5 ;
      RECT  7710.0 89587.5 7780.0 89452.5 ;
      RECT  8090.0 89587.5 8160.0 89452.5 ;
      RECT  8090.0 90427.5 8160.0 90292.5 ;
      RECT  8090.0 89970.0 8160.0 89835.0 ;
      RECT  8090.0 90887.5 8160.0 91592.5 ;
      RECT  7710.0 91242.5 7780.0 91312.5 ;
      RECT  8090.0 91242.5 8160.0 91312.5 ;
      RECT  7710.0 91277.5 7780.0 91592.5 ;
      RECT  7745.0 91242.5 8125.0 91312.5 ;
      RECT  8090.0 90887.5 8160.0 91277.5 ;
      RECT  7710.0 91592.5 7780.0 91727.5 ;
      RECT  8090.0 91592.5 8160.0 91727.5 ;
      RECT  8090.0 90752.5 8160.0 90887.5 ;
      RECT  8090.0 91210.0 8160.0 91345.0 ;
      RECT  8090.0 92982.5 8160.0 92277.5 ;
      RECT  7710.0 92627.5 7780.0 92557.5 ;
      RECT  8090.0 92627.5 8160.0 92557.5 ;
      RECT  7710.0 92592.5 7780.0 92277.5 ;
      RECT  7745.0 92627.5 8125.0 92557.5 ;
      RECT  8090.0 92982.5 8160.0 92592.5 ;
      RECT  7710.0 92277.5 7780.0 92142.5 ;
      RECT  8090.0 92277.5 8160.0 92142.5 ;
      RECT  8090.0 93117.5 8160.0 92982.5 ;
      RECT  8090.0 92660.0 8160.0 92525.0 ;
      RECT  8090.0 93577.5 8160.0 94282.5 ;
      RECT  7710.0 93932.5 7780.0 94002.5 ;
      RECT  8090.0 93932.5 8160.0 94002.5 ;
      RECT  7710.0 93967.5 7780.0 94282.5 ;
      RECT  7745.0 93932.5 8125.0 94002.5 ;
      RECT  8090.0 93577.5 8160.0 93967.5 ;
      RECT  7710.0 94282.5 7780.0 94417.5 ;
      RECT  8090.0 94282.5 8160.0 94417.5 ;
      RECT  8090.0 93442.5 8160.0 93577.5 ;
      RECT  8090.0 93900.0 8160.0 94035.0 ;
      RECT  8090.0 95672.5 8160.0 94967.5 ;
      RECT  7710.0 95317.5 7780.0 95247.5 ;
      RECT  8090.0 95317.5 8160.0 95247.5 ;
      RECT  7710.0 95282.5 7780.0 94967.5 ;
      RECT  7745.0 95317.5 8125.0 95247.5 ;
      RECT  8090.0 95672.5 8160.0 95282.5 ;
      RECT  7710.0 94967.5 7780.0 94832.5 ;
      RECT  8090.0 94967.5 8160.0 94832.5 ;
      RECT  8090.0 95807.5 8160.0 95672.5 ;
      RECT  8090.0 95350.0 8160.0 95215.0 ;
      RECT  8090.0 96267.5 8160.0 96972.5 ;
      RECT  7710.0 96622.5 7780.0 96692.5 ;
      RECT  8090.0 96622.5 8160.0 96692.5 ;
      RECT  7710.0 96657.5 7780.0 96972.5 ;
      RECT  7745.0 96622.5 8125.0 96692.5 ;
      RECT  8090.0 96267.5 8160.0 96657.5 ;
      RECT  7710.0 96972.5 7780.0 97107.5 ;
      RECT  8090.0 96972.5 8160.0 97107.5 ;
      RECT  8090.0 96132.5 8160.0 96267.5 ;
      RECT  8090.0 96590.0 8160.0 96725.0 ;
      RECT  8090.0 98362.5 8160.0 97657.5 ;
      RECT  7710.0 98007.5 7780.0 97937.5 ;
      RECT  8090.0 98007.5 8160.0 97937.5 ;
      RECT  7710.0 97972.5 7780.0 97657.5 ;
      RECT  7745.0 98007.5 8125.0 97937.5 ;
      RECT  8090.0 98362.5 8160.0 97972.5 ;
      RECT  7710.0 97657.5 7780.0 97522.5 ;
      RECT  8090.0 97657.5 8160.0 97522.5 ;
      RECT  8090.0 98497.5 8160.0 98362.5 ;
      RECT  8090.0 98040.0 8160.0 97905.0 ;
      RECT  8090.0 98957.5 8160.0 99662.5 ;
      RECT  7710.0 99312.5 7780.0 99382.5 ;
      RECT  8090.0 99312.5 8160.0 99382.5 ;
      RECT  7710.0 99347.5 7780.0 99662.5 ;
      RECT  7745.0 99312.5 8125.0 99382.5 ;
      RECT  8090.0 98957.5 8160.0 99347.5 ;
      RECT  7710.0 99662.5 7780.0 99797.5 ;
      RECT  8090.0 99662.5 8160.0 99797.5 ;
      RECT  8090.0 98822.5 8160.0 98957.5 ;
      RECT  8090.0 99280.0 8160.0 99415.0 ;
      RECT  8090.0 101052.5 8160.0 100347.5 ;
      RECT  7710.0 100697.5 7780.0 100627.5 ;
      RECT  8090.0 100697.5 8160.0 100627.5 ;
      RECT  7710.0 100662.5 7780.0 100347.5 ;
      RECT  7745.0 100697.5 8125.0 100627.5 ;
      RECT  8090.0 101052.5 8160.0 100662.5 ;
      RECT  7710.0 100347.5 7780.0 100212.5 ;
      RECT  8090.0 100347.5 8160.0 100212.5 ;
      RECT  8090.0 101187.5 8160.0 101052.5 ;
      RECT  8090.0 100730.0 8160.0 100595.0 ;
      RECT  8090.0 101647.5 8160.0 102352.5 ;
      RECT  7710.0 102002.5 7780.0 102072.5 ;
      RECT  8090.0 102002.5 8160.0 102072.5 ;
      RECT  7710.0 102037.5 7780.0 102352.5 ;
      RECT  7745.0 102002.5 8125.0 102072.5 ;
      RECT  8090.0 101647.5 8160.0 102037.5 ;
      RECT  7710.0 102352.5 7780.0 102487.5 ;
      RECT  8090.0 102352.5 8160.0 102487.5 ;
      RECT  8090.0 101512.5 8160.0 101647.5 ;
      RECT  8090.0 101970.0 8160.0 102105.0 ;
      RECT  8090.0 103742.5 8160.0 103037.5 ;
      RECT  7710.0 103387.5 7780.0 103317.5 ;
      RECT  8090.0 103387.5 8160.0 103317.5 ;
      RECT  7710.0 103352.5 7780.0 103037.5 ;
      RECT  7745.0 103387.5 8125.0 103317.5 ;
      RECT  8090.0 103742.5 8160.0 103352.5 ;
      RECT  7710.0 103037.5 7780.0 102902.5 ;
      RECT  8090.0 103037.5 8160.0 102902.5 ;
      RECT  8090.0 103877.5 8160.0 103742.5 ;
      RECT  8090.0 103420.0 8160.0 103285.0 ;
      RECT  8090.0 104337.5 8160.0 105042.5 ;
      RECT  7710.0 104692.5 7780.0 104762.5 ;
      RECT  8090.0 104692.5 8160.0 104762.5 ;
      RECT  7710.0 104727.5 7780.0 105042.5 ;
      RECT  7745.0 104692.5 8125.0 104762.5 ;
      RECT  8090.0 104337.5 8160.0 104727.5 ;
      RECT  7710.0 105042.5 7780.0 105177.5 ;
      RECT  8090.0 105042.5 8160.0 105177.5 ;
      RECT  8090.0 104202.5 8160.0 104337.5 ;
      RECT  8090.0 104660.0 8160.0 104795.0 ;
      RECT  8090.0 106432.5 8160.0 105727.5 ;
      RECT  7710.0 106077.5 7780.0 106007.5 ;
      RECT  8090.0 106077.5 8160.0 106007.5 ;
      RECT  7710.0 106042.5 7780.0 105727.5 ;
      RECT  7745.0 106077.5 8125.0 106007.5 ;
      RECT  8090.0 106432.5 8160.0 106042.5 ;
      RECT  7710.0 105727.5 7780.0 105592.5 ;
      RECT  8090.0 105727.5 8160.0 105592.5 ;
      RECT  8090.0 106567.5 8160.0 106432.5 ;
      RECT  8090.0 106110.0 8160.0 105975.0 ;
      RECT  8090.0 107027.5 8160.0 107732.5 ;
      RECT  7710.0 107382.5 7780.0 107452.5 ;
      RECT  8090.0 107382.5 8160.0 107452.5 ;
      RECT  7710.0 107417.5 7780.0 107732.5 ;
      RECT  7745.0 107382.5 8125.0 107452.5 ;
      RECT  8090.0 107027.5 8160.0 107417.5 ;
      RECT  7710.0 107732.5 7780.0 107867.5 ;
      RECT  8090.0 107732.5 8160.0 107867.5 ;
      RECT  8090.0 106892.5 8160.0 107027.5 ;
      RECT  8090.0 107350.0 8160.0 107485.0 ;
      RECT  8090.0 109122.5 8160.0 108417.5 ;
      RECT  7710.0 108767.5 7780.0 108697.5 ;
      RECT  8090.0 108767.5 8160.0 108697.5 ;
      RECT  7710.0 108732.5 7780.0 108417.5 ;
      RECT  7745.0 108767.5 8125.0 108697.5 ;
      RECT  8090.0 109122.5 8160.0 108732.5 ;
      RECT  7710.0 108417.5 7780.0 108282.5 ;
      RECT  8090.0 108417.5 8160.0 108282.5 ;
      RECT  8090.0 109257.5 8160.0 109122.5 ;
      RECT  8090.0 108800.0 8160.0 108665.0 ;
      RECT  8090.0 109717.5 8160.0 110422.5 ;
      RECT  7710.0 110072.5 7780.0 110142.5 ;
      RECT  8090.0 110072.5 8160.0 110142.5 ;
      RECT  7710.0 110107.5 7780.0 110422.5 ;
      RECT  7745.0 110072.5 8125.0 110142.5 ;
      RECT  8090.0 109717.5 8160.0 110107.5 ;
      RECT  7710.0 110422.5 7780.0 110557.5 ;
      RECT  8090.0 110422.5 8160.0 110557.5 ;
      RECT  8090.0 109582.5 8160.0 109717.5 ;
      RECT  8090.0 110040.0 8160.0 110175.0 ;
      RECT  8090.0 111812.5 8160.0 111107.5 ;
      RECT  7710.0 111457.5 7780.0 111387.5 ;
      RECT  8090.0 111457.5 8160.0 111387.5 ;
      RECT  7710.0 111422.5 7780.0 111107.5 ;
      RECT  7745.0 111457.5 8125.0 111387.5 ;
      RECT  8090.0 111812.5 8160.0 111422.5 ;
      RECT  7710.0 111107.5 7780.0 110972.5 ;
      RECT  8090.0 111107.5 8160.0 110972.5 ;
      RECT  8090.0 111947.5 8160.0 111812.5 ;
      RECT  8090.0 111490.0 8160.0 111355.0 ;
      RECT  8090.0 112407.5 8160.0 113112.5 ;
      RECT  7710.0 112762.5 7780.0 112832.5 ;
      RECT  8090.0 112762.5 8160.0 112832.5 ;
      RECT  7710.0 112797.5 7780.0 113112.5 ;
      RECT  7745.0 112762.5 8125.0 112832.5 ;
      RECT  8090.0 112407.5 8160.0 112797.5 ;
      RECT  7710.0 113112.5 7780.0 113247.5 ;
      RECT  8090.0 113112.5 8160.0 113247.5 ;
      RECT  8090.0 112272.5 8160.0 112407.5 ;
      RECT  8090.0 112730.0 8160.0 112865.0 ;
      RECT  8090.0 114502.5 8160.0 113797.5 ;
      RECT  7710.0 114147.5 7780.0 114077.5 ;
      RECT  8090.0 114147.5 8160.0 114077.5 ;
      RECT  7710.0 114112.5 7780.0 113797.5 ;
      RECT  7745.0 114147.5 8125.0 114077.5 ;
      RECT  8090.0 114502.5 8160.0 114112.5 ;
      RECT  7710.0 113797.5 7780.0 113662.5 ;
      RECT  8090.0 113797.5 8160.0 113662.5 ;
      RECT  8090.0 114637.5 8160.0 114502.5 ;
      RECT  8090.0 114180.0 8160.0 114045.0 ;
      RECT  8090.0 115097.5 8160.0 115802.5 ;
      RECT  7710.0 115452.5 7780.0 115522.5 ;
      RECT  8090.0 115452.5 8160.0 115522.5 ;
      RECT  7710.0 115487.5 7780.0 115802.5 ;
      RECT  7745.0 115452.5 8125.0 115522.5 ;
      RECT  8090.0 115097.5 8160.0 115487.5 ;
      RECT  7710.0 115802.5 7780.0 115937.5 ;
      RECT  8090.0 115802.5 8160.0 115937.5 ;
      RECT  8090.0 114962.5 8160.0 115097.5 ;
      RECT  8090.0 115420.0 8160.0 115555.0 ;
      RECT  8090.0 117192.5 8160.0 116487.5 ;
      RECT  7710.0 116837.5 7780.0 116767.5 ;
      RECT  8090.0 116837.5 8160.0 116767.5 ;
      RECT  7710.0 116802.5 7780.0 116487.5 ;
      RECT  7745.0 116837.5 8125.0 116767.5 ;
      RECT  8090.0 117192.5 8160.0 116802.5 ;
      RECT  7710.0 116487.5 7780.0 116352.5 ;
      RECT  8090.0 116487.5 8160.0 116352.5 ;
      RECT  8090.0 117327.5 8160.0 117192.5 ;
      RECT  8090.0 116870.0 8160.0 116735.0 ;
      RECT  8090.0 117787.5 8160.0 118492.5 ;
      RECT  7710.0 118142.5 7780.0 118212.5 ;
      RECT  8090.0 118142.5 8160.0 118212.5 ;
      RECT  7710.0 118177.5 7780.0 118492.5 ;
      RECT  7745.0 118142.5 8125.0 118212.5 ;
      RECT  8090.0 117787.5 8160.0 118177.5 ;
      RECT  7710.0 118492.5 7780.0 118627.5 ;
      RECT  8090.0 118492.5 8160.0 118627.5 ;
      RECT  8090.0 117652.5 8160.0 117787.5 ;
      RECT  8090.0 118110.0 8160.0 118245.0 ;
      RECT  8090.0 119882.5 8160.0 119177.5 ;
      RECT  7710.0 119527.5 7780.0 119457.5 ;
      RECT  8090.0 119527.5 8160.0 119457.5 ;
      RECT  7710.0 119492.5 7780.0 119177.5 ;
      RECT  7745.0 119527.5 8125.0 119457.5 ;
      RECT  8090.0 119882.5 8160.0 119492.5 ;
      RECT  7710.0 119177.5 7780.0 119042.5 ;
      RECT  8090.0 119177.5 8160.0 119042.5 ;
      RECT  8090.0 120017.5 8160.0 119882.5 ;
      RECT  8090.0 119560.0 8160.0 119425.0 ;
      RECT  8090.0 120477.5 8160.0 121182.5 ;
      RECT  7710.0 120832.5 7780.0 120902.5 ;
      RECT  8090.0 120832.5 8160.0 120902.5 ;
      RECT  7710.0 120867.5 7780.0 121182.5 ;
      RECT  7745.0 120832.5 8125.0 120902.5 ;
      RECT  8090.0 120477.5 8160.0 120867.5 ;
      RECT  7710.0 121182.5 7780.0 121317.5 ;
      RECT  8090.0 121182.5 8160.0 121317.5 ;
      RECT  8090.0 120342.5 8160.0 120477.5 ;
      RECT  8090.0 120800.0 8160.0 120935.0 ;
      RECT  8090.0 122572.5 8160.0 121867.5 ;
      RECT  7710.0 122217.5 7780.0 122147.5 ;
      RECT  8090.0 122217.5 8160.0 122147.5 ;
      RECT  7710.0 122182.5 7780.0 121867.5 ;
      RECT  7745.0 122217.5 8125.0 122147.5 ;
      RECT  8090.0 122572.5 8160.0 122182.5 ;
      RECT  7710.0 121867.5 7780.0 121732.5 ;
      RECT  8090.0 121867.5 8160.0 121732.5 ;
      RECT  8090.0 122707.5 8160.0 122572.5 ;
      RECT  8090.0 122250.0 8160.0 122115.0 ;
      RECT  8090.0 123167.5 8160.0 123872.5 ;
      RECT  7710.0 123522.5 7780.0 123592.5 ;
      RECT  8090.0 123522.5 8160.0 123592.5 ;
      RECT  7710.0 123557.5 7780.0 123872.5 ;
      RECT  7745.0 123522.5 8125.0 123592.5 ;
      RECT  8090.0 123167.5 8160.0 123557.5 ;
      RECT  7710.0 123872.5 7780.0 124007.5 ;
      RECT  8090.0 123872.5 8160.0 124007.5 ;
      RECT  8090.0 123032.5 8160.0 123167.5 ;
      RECT  8090.0 123490.0 8160.0 123625.0 ;
      RECT  8090.0 125262.5 8160.0 124557.5 ;
      RECT  7710.0 124907.5 7780.0 124837.5 ;
      RECT  8090.0 124907.5 8160.0 124837.5 ;
      RECT  7710.0 124872.5 7780.0 124557.5 ;
      RECT  7745.0 124907.5 8125.0 124837.5 ;
      RECT  8090.0 125262.5 8160.0 124872.5 ;
      RECT  7710.0 124557.5 7780.0 124422.5 ;
      RECT  8090.0 124557.5 8160.0 124422.5 ;
      RECT  8090.0 125397.5 8160.0 125262.5 ;
      RECT  8090.0 124940.0 8160.0 124805.0 ;
      RECT  8090.0 125857.5 8160.0 126562.5 ;
      RECT  7710.0 126212.5 7780.0 126282.5 ;
      RECT  8090.0 126212.5 8160.0 126282.5 ;
      RECT  7710.0 126247.5 7780.0 126562.5 ;
      RECT  7745.0 126212.5 8125.0 126282.5 ;
      RECT  8090.0 125857.5 8160.0 126247.5 ;
      RECT  7710.0 126562.5 7780.0 126697.5 ;
      RECT  8090.0 126562.5 8160.0 126697.5 ;
      RECT  8090.0 125722.5 8160.0 125857.5 ;
      RECT  8090.0 126180.0 8160.0 126315.0 ;
      RECT  8090.0 127952.5 8160.0 127247.5 ;
      RECT  7710.0 127597.5 7780.0 127527.5 ;
      RECT  8090.0 127597.5 8160.0 127527.5 ;
      RECT  7710.0 127562.5 7780.0 127247.5 ;
      RECT  7745.0 127597.5 8125.0 127527.5 ;
      RECT  8090.0 127952.5 8160.0 127562.5 ;
      RECT  7710.0 127247.5 7780.0 127112.5 ;
      RECT  8090.0 127247.5 8160.0 127112.5 ;
      RECT  8090.0 128087.5 8160.0 127952.5 ;
      RECT  8090.0 127630.0 8160.0 127495.0 ;
      RECT  8090.0 128547.5 8160.0 129252.5 ;
      RECT  7710.0 128902.5 7780.0 128972.5 ;
      RECT  8090.0 128902.5 8160.0 128972.5 ;
      RECT  7710.0 128937.5 7780.0 129252.5 ;
      RECT  7745.0 128902.5 8125.0 128972.5 ;
      RECT  8090.0 128547.5 8160.0 128937.5 ;
      RECT  7710.0 129252.5 7780.0 129387.5 ;
      RECT  8090.0 129252.5 8160.0 129387.5 ;
      RECT  8090.0 128412.5 8160.0 128547.5 ;
      RECT  8090.0 128870.0 8160.0 129005.0 ;
      RECT  8090.0 130642.5 8160.0 129937.5 ;
      RECT  7710.0 130287.5 7780.0 130217.5 ;
      RECT  8090.0 130287.5 8160.0 130217.5 ;
      RECT  7710.0 130252.5 7780.0 129937.5 ;
      RECT  7745.0 130287.5 8125.0 130217.5 ;
      RECT  8090.0 130642.5 8160.0 130252.5 ;
      RECT  7710.0 129937.5 7780.0 129802.5 ;
      RECT  8090.0 129937.5 8160.0 129802.5 ;
      RECT  8090.0 130777.5 8160.0 130642.5 ;
      RECT  8090.0 130320.0 8160.0 130185.0 ;
      RECT  8090.0 131237.5 8160.0 131942.5 ;
      RECT  7710.0 131592.5 7780.0 131662.5 ;
      RECT  8090.0 131592.5 8160.0 131662.5 ;
      RECT  7710.0 131627.5 7780.0 131942.5 ;
      RECT  7745.0 131592.5 8125.0 131662.5 ;
      RECT  8090.0 131237.5 8160.0 131627.5 ;
      RECT  7710.0 131942.5 7780.0 132077.5 ;
      RECT  8090.0 131942.5 8160.0 132077.5 ;
      RECT  8090.0 131102.5 8160.0 131237.5 ;
      RECT  8090.0 131560.0 8160.0 131695.0 ;
      RECT  8090.0 133332.5 8160.0 132627.5 ;
      RECT  7710.0 132977.5 7780.0 132907.5 ;
      RECT  8090.0 132977.5 8160.0 132907.5 ;
      RECT  7710.0 132942.5 7780.0 132627.5 ;
      RECT  7745.0 132977.5 8125.0 132907.5 ;
      RECT  8090.0 133332.5 8160.0 132942.5 ;
      RECT  7710.0 132627.5 7780.0 132492.5 ;
      RECT  8090.0 132627.5 8160.0 132492.5 ;
      RECT  8090.0 133467.5 8160.0 133332.5 ;
      RECT  8090.0 133010.0 8160.0 132875.0 ;
      RECT  8090.0 133927.5 8160.0 134632.5 ;
      RECT  7710.0 134282.5 7780.0 134352.5 ;
      RECT  8090.0 134282.5 8160.0 134352.5 ;
      RECT  7710.0 134317.5 7780.0 134632.5 ;
      RECT  7745.0 134282.5 8125.0 134352.5 ;
      RECT  8090.0 133927.5 8160.0 134317.5 ;
      RECT  7710.0 134632.5 7780.0 134767.5 ;
      RECT  8090.0 134632.5 8160.0 134767.5 ;
      RECT  8090.0 133792.5 8160.0 133927.5 ;
      RECT  8090.0 134250.0 8160.0 134385.0 ;
      RECT  8090.0 136022.5 8160.0 135317.5 ;
      RECT  7710.0 135667.5 7780.0 135597.5 ;
      RECT  8090.0 135667.5 8160.0 135597.5 ;
      RECT  7710.0 135632.5 7780.0 135317.5 ;
      RECT  7745.0 135667.5 8125.0 135597.5 ;
      RECT  8090.0 136022.5 8160.0 135632.5 ;
      RECT  7710.0 135317.5 7780.0 135182.5 ;
      RECT  8090.0 135317.5 8160.0 135182.5 ;
      RECT  8090.0 136157.5 8160.0 136022.5 ;
      RECT  8090.0 135700.0 8160.0 135565.0 ;
      RECT  8090.0 136617.5 8160.0 137322.5 ;
      RECT  7710.0 136972.5 7780.0 137042.5 ;
      RECT  8090.0 136972.5 8160.0 137042.5 ;
      RECT  7710.0 137007.5 7780.0 137322.5 ;
      RECT  7745.0 136972.5 8125.0 137042.5 ;
      RECT  8090.0 136617.5 8160.0 137007.5 ;
      RECT  7710.0 137322.5 7780.0 137457.5 ;
      RECT  8090.0 137322.5 8160.0 137457.5 ;
      RECT  8090.0 136482.5 8160.0 136617.5 ;
      RECT  8090.0 136940.0 8160.0 137075.0 ;
      RECT  8090.0 138712.5 8160.0 138007.5 ;
      RECT  7710.0 138357.5 7780.0 138287.5 ;
      RECT  8090.0 138357.5 8160.0 138287.5 ;
      RECT  7710.0 138322.5 7780.0 138007.5 ;
      RECT  7745.0 138357.5 8125.0 138287.5 ;
      RECT  8090.0 138712.5 8160.0 138322.5 ;
      RECT  7710.0 138007.5 7780.0 137872.5 ;
      RECT  8090.0 138007.5 8160.0 137872.5 ;
      RECT  8090.0 138847.5 8160.0 138712.5 ;
      RECT  8090.0 138390.0 8160.0 138255.0 ;
      RECT  8090.0 139307.5 8160.0 140012.5 ;
      RECT  7710.0 139662.5 7780.0 139732.5 ;
      RECT  8090.0 139662.5 8160.0 139732.5 ;
      RECT  7710.0 139697.5 7780.0 140012.5 ;
      RECT  7745.0 139662.5 8125.0 139732.5 ;
      RECT  8090.0 139307.5 8160.0 139697.5 ;
      RECT  7710.0 140012.5 7780.0 140147.5 ;
      RECT  8090.0 140012.5 8160.0 140147.5 ;
      RECT  8090.0 139172.5 8160.0 139307.5 ;
      RECT  8090.0 139630.0 8160.0 139765.0 ;
      RECT  8090.0 141402.5 8160.0 140697.5 ;
      RECT  7710.0 141047.5 7780.0 140977.5 ;
      RECT  8090.0 141047.5 8160.0 140977.5 ;
      RECT  7710.0 141012.5 7780.0 140697.5 ;
      RECT  7745.0 141047.5 8125.0 140977.5 ;
      RECT  8090.0 141402.5 8160.0 141012.5 ;
      RECT  7710.0 140697.5 7780.0 140562.5 ;
      RECT  8090.0 140697.5 8160.0 140562.5 ;
      RECT  8090.0 141537.5 8160.0 141402.5 ;
      RECT  8090.0 141080.0 8160.0 140945.0 ;
      RECT  8090.0 141997.5 8160.0 142702.5 ;
      RECT  7710.0 142352.5 7780.0 142422.5 ;
      RECT  8090.0 142352.5 8160.0 142422.5 ;
      RECT  7710.0 142387.5 7780.0 142702.5 ;
      RECT  7745.0 142352.5 8125.0 142422.5 ;
      RECT  8090.0 141997.5 8160.0 142387.5 ;
      RECT  7710.0 142702.5 7780.0 142837.5 ;
      RECT  8090.0 142702.5 8160.0 142837.5 ;
      RECT  8090.0 141862.5 8160.0 141997.5 ;
      RECT  8090.0 142320.0 8160.0 142455.0 ;
      RECT  8090.0 144092.5 8160.0 143387.5 ;
      RECT  7710.0 143737.5 7780.0 143667.5 ;
      RECT  8090.0 143737.5 8160.0 143667.5 ;
      RECT  7710.0 143702.5 7780.0 143387.5 ;
      RECT  7745.0 143737.5 8125.0 143667.5 ;
      RECT  8090.0 144092.5 8160.0 143702.5 ;
      RECT  7710.0 143387.5 7780.0 143252.5 ;
      RECT  8090.0 143387.5 8160.0 143252.5 ;
      RECT  8090.0 144227.5 8160.0 144092.5 ;
      RECT  8090.0 143770.0 8160.0 143635.0 ;
      RECT  8090.0 144687.5 8160.0 145392.5 ;
      RECT  7710.0 145042.5 7780.0 145112.5 ;
      RECT  8090.0 145042.5 8160.0 145112.5 ;
      RECT  7710.0 145077.5 7780.0 145392.5 ;
      RECT  7745.0 145042.5 8125.0 145112.5 ;
      RECT  8090.0 144687.5 8160.0 145077.5 ;
      RECT  7710.0 145392.5 7780.0 145527.5 ;
      RECT  8090.0 145392.5 8160.0 145527.5 ;
      RECT  8090.0 144552.5 8160.0 144687.5 ;
      RECT  8090.0 145010.0 8160.0 145145.0 ;
      RECT  8090.0 146782.5 8160.0 146077.5 ;
      RECT  7710.0 146427.5 7780.0 146357.5 ;
      RECT  8090.0 146427.5 8160.0 146357.5 ;
      RECT  7710.0 146392.5 7780.0 146077.5 ;
      RECT  7745.0 146427.5 8125.0 146357.5 ;
      RECT  8090.0 146782.5 8160.0 146392.5 ;
      RECT  7710.0 146077.5 7780.0 145942.5 ;
      RECT  8090.0 146077.5 8160.0 145942.5 ;
      RECT  8090.0 146917.5 8160.0 146782.5 ;
      RECT  8090.0 146460.0 8160.0 146325.0 ;
      RECT  8090.0 147377.5 8160.0 148082.5 ;
      RECT  7710.0 147732.5 7780.0 147802.5 ;
      RECT  8090.0 147732.5 8160.0 147802.5 ;
      RECT  7710.0 147767.5 7780.0 148082.5 ;
      RECT  7745.0 147732.5 8125.0 147802.5 ;
      RECT  8090.0 147377.5 8160.0 147767.5 ;
      RECT  7710.0 148082.5 7780.0 148217.5 ;
      RECT  8090.0 148082.5 8160.0 148217.5 ;
      RECT  8090.0 147242.5 8160.0 147377.5 ;
      RECT  8090.0 147700.0 8160.0 147835.0 ;
      RECT  8090.0 149472.5 8160.0 148767.5 ;
      RECT  7710.0 149117.5 7780.0 149047.5 ;
      RECT  8090.0 149117.5 8160.0 149047.5 ;
      RECT  7710.0 149082.5 7780.0 148767.5 ;
      RECT  7745.0 149117.5 8125.0 149047.5 ;
      RECT  8090.0 149472.5 8160.0 149082.5 ;
      RECT  7710.0 148767.5 7780.0 148632.5 ;
      RECT  8090.0 148767.5 8160.0 148632.5 ;
      RECT  8090.0 149607.5 8160.0 149472.5 ;
      RECT  8090.0 149150.0 8160.0 149015.0 ;
      RECT  8090.0 150067.5 8160.0 150772.5 ;
      RECT  7710.0 150422.5 7780.0 150492.5 ;
      RECT  8090.0 150422.5 8160.0 150492.5 ;
      RECT  7710.0 150457.5 7780.0 150772.5 ;
      RECT  7745.0 150422.5 8125.0 150492.5 ;
      RECT  8090.0 150067.5 8160.0 150457.5 ;
      RECT  7710.0 150772.5 7780.0 150907.5 ;
      RECT  8090.0 150772.5 8160.0 150907.5 ;
      RECT  8090.0 149932.5 8160.0 150067.5 ;
      RECT  8090.0 150390.0 8160.0 150525.0 ;
      RECT  8090.0 152162.5 8160.0 151457.5 ;
      RECT  7710.0 151807.5 7780.0 151737.5 ;
      RECT  8090.0 151807.5 8160.0 151737.5 ;
      RECT  7710.0 151772.5 7780.0 151457.5 ;
      RECT  7745.0 151807.5 8125.0 151737.5 ;
      RECT  8090.0 152162.5 8160.0 151772.5 ;
      RECT  7710.0 151457.5 7780.0 151322.5 ;
      RECT  8090.0 151457.5 8160.0 151322.5 ;
      RECT  8090.0 152297.5 8160.0 152162.5 ;
      RECT  8090.0 151840.0 8160.0 151705.0 ;
      RECT  8090.0 152757.5 8160.0 153462.5 ;
      RECT  7710.0 153112.5 7780.0 153182.5 ;
      RECT  8090.0 153112.5 8160.0 153182.5 ;
      RECT  7710.0 153147.5 7780.0 153462.5 ;
      RECT  7745.0 153112.5 8125.0 153182.5 ;
      RECT  8090.0 152757.5 8160.0 153147.5 ;
      RECT  7710.0 153462.5 7780.0 153597.5 ;
      RECT  8090.0 153462.5 8160.0 153597.5 ;
      RECT  8090.0 152622.5 8160.0 152757.5 ;
      RECT  8090.0 153080.0 8160.0 153215.0 ;
      RECT  8090.0 154852.5 8160.0 154147.5 ;
      RECT  7710.0 154497.5 7780.0 154427.5 ;
      RECT  8090.0 154497.5 8160.0 154427.5 ;
      RECT  7710.0 154462.5 7780.0 154147.5 ;
      RECT  7745.0 154497.5 8125.0 154427.5 ;
      RECT  8090.0 154852.5 8160.0 154462.5 ;
      RECT  7710.0 154147.5 7780.0 154012.5 ;
      RECT  8090.0 154147.5 8160.0 154012.5 ;
      RECT  8090.0 154987.5 8160.0 154852.5 ;
      RECT  8090.0 154530.0 8160.0 154395.0 ;
      RECT  8090.0 155447.5 8160.0 156152.5 ;
      RECT  7710.0 155802.5 7780.0 155872.5 ;
      RECT  8090.0 155802.5 8160.0 155872.5 ;
      RECT  7710.0 155837.5 7780.0 156152.5 ;
      RECT  7745.0 155802.5 8125.0 155872.5 ;
      RECT  8090.0 155447.5 8160.0 155837.5 ;
      RECT  7710.0 156152.5 7780.0 156287.5 ;
      RECT  8090.0 156152.5 8160.0 156287.5 ;
      RECT  8090.0 155312.5 8160.0 155447.5 ;
      RECT  8090.0 155770.0 8160.0 155905.0 ;
      RECT  8090.0 157542.5 8160.0 156837.5 ;
      RECT  7710.0 157187.5 7780.0 157117.5 ;
      RECT  8090.0 157187.5 8160.0 157117.5 ;
      RECT  7710.0 157152.5 7780.0 156837.5 ;
      RECT  7745.0 157187.5 8125.0 157117.5 ;
      RECT  8090.0 157542.5 8160.0 157152.5 ;
      RECT  7710.0 156837.5 7780.0 156702.5 ;
      RECT  8090.0 156837.5 8160.0 156702.5 ;
      RECT  8090.0 157677.5 8160.0 157542.5 ;
      RECT  8090.0 157220.0 8160.0 157085.0 ;
      RECT  8090.0 158137.5 8160.0 158842.5 ;
      RECT  7710.0 158492.5 7780.0 158562.5 ;
      RECT  8090.0 158492.5 8160.0 158562.5 ;
      RECT  7710.0 158527.5 7780.0 158842.5 ;
      RECT  7745.0 158492.5 8125.0 158562.5 ;
      RECT  8090.0 158137.5 8160.0 158527.5 ;
      RECT  7710.0 158842.5 7780.0 158977.5 ;
      RECT  8090.0 158842.5 8160.0 158977.5 ;
      RECT  8090.0 158002.5 8160.0 158137.5 ;
      RECT  8090.0 158460.0 8160.0 158595.0 ;
      RECT  8090.0 160232.5 8160.0 159527.5 ;
      RECT  7710.0 159877.5 7780.0 159807.5 ;
      RECT  8090.0 159877.5 8160.0 159807.5 ;
      RECT  7710.0 159842.5 7780.0 159527.5 ;
      RECT  7745.0 159877.5 8125.0 159807.5 ;
      RECT  8090.0 160232.5 8160.0 159842.5 ;
      RECT  7710.0 159527.5 7780.0 159392.5 ;
      RECT  8090.0 159527.5 8160.0 159392.5 ;
      RECT  8090.0 160367.5 8160.0 160232.5 ;
      RECT  8090.0 159910.0 8160.0 159775.0 ;
      RECT  8090.0 160827.5 8160.0 161532.5 ;
      RECT  7710.0 161182.5 7780.0 161252.5 ;
      RECT  8090.0 161182.5 8160.0 161252.5 ;
      RECT  7710.0 161217.5 7780.0 161532.5 ;
      RECT  7745.0 161182.5 8125.0 161252.5 ;
      RECT  8090.0 160827.5 8160.0 161217.5 ;
      RECT  7710.0 161532.5 7780.0 161667.5 ;
      RECT  8090.0 161532.5 8160.0 161667.5 ;
      RECT  8090.0 160692.5 8160.0 160827.5 ;
      RECT  8090.0 161150.0 8160.0 161285.0 ;
      RECT  8090.0 162922.5 8160.0 162217.5 ;
      RECT  7710.0 162567.5 7780.0 162497.5 ;
      RECT  8090.0 162567.5 8160.0 162497.5 ;
      RECT  7710.0 162532.5 7780.0 162217.5 ;
      RECT  7745.0 162567.5 8125.0 162497.5 ;
      RECT  8090.0 162922.5 8160.0 162532.5 ;
      RECT  7710.0 162217.5 7780.0 162082.5 ;
      RECT  8090.0 162217.5 8160.0 162082.5 ;
      RECT  8090.0 163057.5 8160.0 162922.5 ;
      RECT  8090.0 162600.0 8160.0 162465.0 ;
      RECT  8090.0 163517.5 8160.0 164222.5 ;
      RECT  7710.0 163872.5 7780.0 163942.5 ;
      RECT  8090.0 163872.5 8160.0 163942.5 ;
      RECT  7710.0 163907.5 7780.0 164222.5 ;
      RECT  7745.0 163872.5 8125.0 163942.5 ;
      RECT  8090.0 163517.5 8160.0 163907.5 ;
      RECT  7710.0 164222.5 7780.0 164357.5 ;
      RECT  8090.0 164222.5 8160.0 164357.5 ;
      RECT  8090.0 163382.5 8160.0 163517.5 ;
      RECT  8090.0 163840.0 8160.0 163975.0 ;
      RECT  8090.0 165612.5 8160.0 164907.5 ;
      RECT  7710.0 165257.5 7780.0 165187.5 ;
      RECT  8090.0 165257.5 8160.0 165187.5 ;
      RECT  7710.0 165222.5 7780.0 164907.5 ;
      RECT  7745.0 165257.5 8125.0 165187.5 ;
      RECT  8090.0 165612.5 8160.0 165222.5 ;
      RECT  7710.0 164907.5 7780.0 164772.5 ;
      RECT  8090.0 164907.5 8160.0 164772.5 ;
      RECT  8090.0 165747.5 8160.0 165612.5 ;
      RECT  8090.0 165290.0 8160.0 165155.0 ;
      RECT  8090.0 166207.5 8160.0 166912.5 ;
      RECT  7710.0 166562.5 7780.0 166632.5 ;
      RECT  8090.0 166562.5 8160.0 166632.5 ;
      RECT  7710.0 166597.5 7780.0 166912.5 ;
      RECT  7745.0 166562.5 8125.0 166632.5 ;
      RECT  8090.0 166207.5 8160.0 166597.5 ;
      RECT  7710.0 166912.5 7780.0 167047.5 ;
      RECT  8090.0 166912.5 8160.0 167047.5 ;
      RECT  8090.0 166072.5 8160.0 166207.5 ;
      RECT  8090.0 166530.0 8160.0 166665.0 ;
      RECT  8090.0 168302.5 8160.0 167597.5 ;
      RECT  7710.0 167947.5 7780.0 167877.5 ;
      RECT  8090.0 167947.5 8160.0 167877.5 ;
      RECT  7710.0 167912.5 7780.0 167597.5 ;
      RECT  7745.0 167947.5 8125.0 167877.5 ;
      RECT  8090.0 168302.5 8160.0 167912.5 ;
      RECT  7710.0 167597.5 7780.0 167462.5 ;
      RECT  8090.0 167597.5 8160.0 167462.5 ;
      RECT  8090.0 168437.5 8160.0 168302.5 ;
      RECT  8090.0 167980.0 8160.0 167845.0 ;
      RECT  8090.0 168897.5 8160.0 169602.5 ;
      RECT  7710.0 169252.5 7780.0 169322.5 ;
      RECT  8090.0 169252.5 8160.0 169322.5 ;
      RECT  7710.0 169287.5 7780.0 169602.5 ;
      RECT  7745.0 169252.5 8125.0 169322.5 ;
      RECT  8090.0 168897.5 8160.0 169287.5 ;
      RECT  7710.0 169602.5 7780.0 169737.5 ;
      RECT  8090.0 169602.5 8160.0 169737.5 ;
      RECT  8090.0 168762.5 8160.0 168897.5 ;
      RECT  8090.0 169220.0 8160.0 169355.0 ;
      RECT  8090.0 170992.5 8160.0 170287.5 ;
      RECT  7710.0 170637.5 7780.0 170567.5 ;
      RECT  8090.0 170637.5 8160.0 170567.5 ;
      RECT  7710.0 170602.5 7780.0 170287.5 ;
      RECT  7745.0 170637.5 8125.0 170567.5 ;
      RECT  8090.0 170992.5 8160.0 170602.5 ;
      RECT  7710.0 170287.5 7780.0 170152.5 ;
      RECT  8090.0 170287.5 8160.0 170152.5 ;
      RECT  8090.0 171127.5 8160.0 170992.5 ;
      RECT  8090.0 170670.0 8160.0 170535.0 ;
      RECT  8090.0 171587.5 8160.0 172292.5 ;
      RECT  7710.0 171942.5 7780.0 172012.5 ;
      RECT  8090.0 171942.5 8160.0 172012.5 ;
      RECT  7710.0 171977.5 7780.0 172292.5 ;
      RECT  7745.0 171942.5 8125.0 172012.5 ;
      RECT  8090.0 171587.5 8160.0 171977.5 ;
      RECT  7710.0 172292.5 7780.0 172427.5 ;
      RECT  8090.0 172292.5 8160.0 172427.5 ;
      RECT  8090.0 171452.5 8160.0 171587.5 ;
      RECT  8090.0 171910.0 8160.0 172045.0 ;
      RECT  8090.0 173682.5 8160.0 172977.5 ;
      RECT  7710.0 173327.5 7780.0 173257.5 ;
      RECT  8090.0 173327.5 8160.0 173257.5 ;
      RECT  7710.0 173292.5 7780.0 172977.5 ;
      RECT  7745.0 173327.5 8125.0 173257.5 ;
      RECT  8090.0 173682.5 8160.0 173292.5 ;
      RECT  7710.0 172977.5 7780.0 172842.5 ;
      RECT  8090.0 172977.5 8160.0 172842.5 ;
      RECT  8090.0 173817.5 8160.0 173682.5 ;
      RECT  8090.0 173360.0 8160.0 173225.0 ;
      RECT  8090.0 174277.5 8160.0 174982.5 ;
      RECT  7710.0 174632.5 7780.0 174702.5 ;
      RECT  8090.0 174632.5 8160.0 174702.5 ;
      RECT  7710.0 174667.5 7780.0 174982.5 ;
      RECT  7745.0 174632.5 8125.0 174702.5 ;
      RECT  8090.0 174277.5 8160.0 174667.5 ;
      RECT  7710.0 174982.5 7780.0 175117.5 ;
      RECT  8090.0 174982.5 8160.0 175117.5 ;
      RECT  8090.0 174142.5 8160.0 174277.5 ;
      RECT  8090.0 174600.0 8160.0 174735.0 ;
      RECT  8090.0 176372.5 8160.0 175667.5 ;
      RECT  7710.0 176017.5 7780.0 175947.5 ;
      RECT  8090.0 176017.5 8160.0 175947.5 ;
      RECT  7710.0 175982.5 7780.0 175667.5 ;
      RECT  7745.0 176017.5 8125.0 175947.5 ;
      RECT  8090.0 176372.5 8160.0 175982.5 ;
      RECT  7710.0 175667.5 7780.0 175532.5 ;
      RECT  8090.0 175667.5 8160.0 175532.5 ;
      RECT  8090.0 176507.5 8160.0 176372.5 ;
      RECT  8090.0 176050.0 8160.0 175915.0 ;
      RECT  8090.0 176967.5 8160.0 177672.5 ;
      RECT  7710.0 177322.5 7780.0 177392.5 ;
      RECT  8090.0 177322.5 8160.0 177392.5 ;
      RECT  7710.0 177357.5 7780.0 177672.5 ;
      RECT  7745.0 177322.5 8125.0 177392.5 ;
      RECT  8090.0 176967.5 8160.0 177357.5 ;
      RECT  7710.0 177672.5 7780.0 177807.5 ;
      RECT  8090.0 177672.5 8160.0 177807.5 ;
      RECT  8090.0 176832.5 8160.0 176967.5 ;
      RECT  8090.0 177290.0 8160.0 177425.0 ;
      RECT  8090.0 179062.5 8160.0 178357.5 ;
      RECT  7710.0 178707.5 7780.0 178637.5 ;
      RECT  8090.0 178707.5 8160.0 178637.5 ;
      RECT  7710.0 178672.5 7780.0 178357.5 ;
      RECT  7745.0 178707.5 8125.0 178637.5 ;
      RECT  8090.0 179062.5 8160.0 178672.5 ;
      RECT  7710.0 178357.5 7780.0 178222.5 ;
      RECT  8090.0 178357.5 8160.0 178222.5 ;
      RECT  8090.0 179197.5 8160.0 179062.5 ;
      RECT  8090.0 178740.0 8160.0 178605.0 ;
      RECT  8090.0 179657.5 8160.0 180362.5 ;
      RECT  7710.0 180012.5 7780.0 180082.5 ;
      RECT  8090.0 180012.5 8160.0 180082.5 ;
      RECT  7710.0 180047.5 7780.0 180362.5 ;
      RECT  7745.0 180012.5 8125.0 180082.5 ;
      RECT  8090.0 179657.5 8160.0 180047.5 ;
      RECT  7710.0 180362.5 7780.0 180497.5 ;
      RECT  8090.0 180362.5 8160.0 180497.5 ;
      RECT  8090.0 179522.5 8160.0 179657.5 ;
      RECT  8090.0 179980.0 8160.0 180115.0 ;
      RECT  8090.0 181752.5 8160.0 181047.5 ;
      RECT  7710.0 181397.5 7780.0 181327.5 ;
      RECT  8090.0 181397.5 8160.0 181327.5 ;
      RECT  7710.0 181362.5 7780.0 181047.5 ;
      RECT  7745.0 181397.5 8125.0 181327.5 ;
      RECT  8090.0 181752.5 8160.0 181362.5 ;
      RECT  7710.0 181047.5 7780.0 180912.5 ;
      RECT  8090.0 181047.5 8160.0 180912.5 ;
      RECT  8090.0 181887.5 8160.0 181752.5 ;
      RECT  8090.0 181430.0 8160.0 181295.0 ;
      RECT  8090.0 182347.5 8160.0 183052.5 ;
      RECT  7710.0 182702.5 7780.0 182772.5 ;
      RECT  8090.0 182702.5 8160.0 182772.5 ;
      RECT  7710.0 182737.5 7780.0 183052.5 ;
      RECT  7745.0 182702.5 8125.0 182772.5 ;
      RECT  8090.0 182347.5 8160.0 182737.5 ;
      RECT  7710.0 183052.5 7780.0 183187.5 ;
      RECT  8090.0 183052.5 8160.0 183187.5 ;
      RECT  8090.0 182212.5 8160.0 182347.5 ;
      RECT  8090.0 182670.0 8160.0 182805.0 ;
      RECT  8090.0 184442.5 8160.0 183737.5 ;
      RECT  7710.0 184087.5 7780.0 184017.5 ;
      RECT  8090.0 184087.5 8160.0 184017.5 ;
      RECT  7710.0 184052.5 7780.0 183737.5 ;
      RECT  7745.0 184087.5 8125.0 184017.5 ;
      RECT  8090.0 184442.5 8160.0 184052.5 ;
      RECT  7710.0 183737.5 7780.0 183602.5 ;
      RECT  8090.0 183737.5 8160.0 183602.5 ;
      RECT  8090.0 184577.5 8160.0 184442.5 ;
      RECT  8090.0 184120.0 8160.0 183985.0 ;
      RECT  8090.0 185037.5 8160.0 185742.5 ;
      RECT  7710.0 185392.5 7780.0 185462.5 ;
      RECT  8090.0 185392.5 8160.0 185462.5 ;
      RECT  7710.0 185427.5 7780.0 185742.5 ;
      RECT  7745.0 185392.5 8125.0 185462.5 ;
      RECT  8090.0 185037.5 8160.0 185427.5 ;
      RECT  7710.0 185742.5 7780.0 185877.5 ;
      RECT  8090.0 185742.5 8160.0 185877.5 ;
      RECT  8090.0 184902.5 8160.0 185037.5 ;
      RECT  8090.0 185360.0 8160.0 185495.0 ;
      RECT  8090.0 187132.5 8160.0 186427.5 ;
      RECT  7710.0 186777.5 7780.0 186707.5 ;
      RECT  8090.0 186777.5 8160.0 186707.5 ;
      RECT  7710.0 186742.5 7780.0 186427.5 ;
      RECT  7745.0 186777.5 8125.0 186707.5 ;
      RECT  8090.0 187132.5 8160.0 186742.5 ;
      RECT  7710.0 186427.5 7780.0 186292.5 ;
      RECT  8090.0 186427.5 8160.0 186292.5 ;
      RECT  8090.0 187267.5 8160.0 187132.5 ;
      RECT  8090.0 186810.0 8160.0 186675.0 ;
      RECT  8090.0 187727.5 8160.0 188432.5 ;
      RECT  7710.0 188082.5 7780.0 188152.5 ;
      RECT  8090.0 188082.5 8160.0 188152.5 ;
      RECT  7710.0 188117.5 7780.0 188432.5 ;
      RECT  7745.0 188082.5 8125.0 188152.5 ;
      RECT  8090.0 187727.5 8160.0 188117.5 ;
      RECT  7710.0 188432.5 7780.0 188567.5 ;
      RECT  8090.0 188432.5 8160.0 188567.5 ;
      RECT  8090.0 187592.5 8160.0 187727.5 ;
      RECT  8090.0 188050.0 8160.0 188185.0 ;
      RECT  8090.0 189822.5 8160.0 189117.5 ;
      RECT  7710.0 189467.5 7780.0 189397.5 ;
      RECT  8090.0 189467.5 8160.0 189397.5 ;
      RECT  7710.0 189432.5 7780.0 189117.5 ;
      RECT  7745.0 189467.5 8125.0 189397.5 ;
      RECT  8090.0 189822.5 8160.0 189432.5 ;
      RECT  7710.0 189117.5 7780.0 188982.5 ;
      RECT  8090.0 189117.5 8160.0 188982.5 ;
      RECT  8090.0 189957.5 8160.0 189822.5 ;
      RECT  8090.0 189500.0 8160.0 189365.0 ;
      RECT  8090.0 190417.5 8160.0 191122.5 ;
      RECT  7710.0 190772.5 7780.0 190842.5 ;
      RECT  8090.0 190772.5 8160.0 190842.5 ;
      RECT  7710.0 190807.5 7780.0 191122.5 ;
      RECT  7745.0 190772.5 8125.0 190842.5 ;
      RECT  8090.0 190417.5 8160.0 190807.5 ;
      RECT  7710.0 191122.5 7780.0 191257.5 ;
      RECT  8090.0 191122.5 8160.0 191257.5 ;
      RECT  8090.0 190282.5 8160.0 190417.5 ;
      RECT  8090.0 190740.0 8160.0 190875.0 ;
      RECT  8090.0 192512.5 8160.0 191807.5 ;
      RECT  7710.0 192157.5 7780.0 192087.5 ;
      RECT  8090.0 192157.5 8160.0 192087.5 ;
      RECT  7710.0 192122.5 7780.0 191807.5 ;
      RECT  7745.0 192157.5 8125.0 192087.5 ;
      RECT  8090.0 192512.5 8160.0 192122.5 ;
      RECT  7710.0 191807.5 7780.0 191672.5 ;
      RECT  8090.0 191807.5 8160.0 191672.5 ;
      RECT  8090.0 192647.5 8160.0 192512.5 ;
      RECT  8090.0 192190.0 8160.0 192055.0 ;
      RECT  8090.0 193107.5 8160.0 193812.5 ;
      RECT  7710.0 193462.5 7780.0 193532.5 ;
      RECT  8090.0 193462.5 8160.0 193532.5 ;
      RECT  7710.0 193497.5 7780.0 193812.5 ;
      RECT  7745.0 193462.5 8125.0 193532.5 ;
      RECT  8090.0 193107.5 8160.0 193497.5 ;
      RECT  7710.0 193812.5 7780.0 193947.5 ;
      RECT  8090.0 193812.5 8160.0 193947.5 ;
      RECT  8090.0 192972.5 8160.0 193107.5 ;
      RECT  8090.0 193430.0 8160.0 193565.0 ;
      RECT  8090.0 195202.5 8160.0 194497.5 ;
      RECT  7710.0 194847.5 7780.0 194777.5 ;
      RECT  8090.0 194847.5 8160.0 194777.5 ;
      RECT  7710.0 194812.5 7780.0 194497.5 ;
      RECT  7745.0 194847.5 8125.0 194777.5 ;
      RECT  8090.0 195202.5 8160.0 194812.5 ;
      RECT  7710.0 194497.5 7780.0 194362.5 ;
      RECT  8090.0 194497.5 8160.0 194362.5 ;
      RECT  8090.0 195337.5 8160.0 195202.5 ;
      RECT  8090.0 194880.0 8160.0 194745.0 ;
      RECT  8090.0 195797.5 8160.0 196502.5 ;
      RECT  7710.0 196152.5 7780.0 196222.5 ;
      RECT  8090.0 196152.5 8160.0 196222.5 ;
      RECT  7710.0 196187.5 7780.0 196502.5 ;
      RECT  7745.0 196152.5 8125.0 196222.5 ;
      RECT  8090.0 195797.5 8160.0 196187.5 ;
      RECT  7710.0 196502.5 7780.0 196637.5 ;
      RECT  8090.0 196502.5 8160.0 196637.5 ;
      RECT  8090.0 195662.5 8160.0 195797.5 ;
      RECT  8090.0 196120.0 8160.0 196255.0 ;
      RECT  8090.0 197892.5 8160.0 197187.5 ;
      RECT  7710.0 197537.5 7780.0 197467.5 ;
      RECT  8090.0 197537.5 8160.0 197467.5 ;
      RECT  7710.0 197502.5 7780.0 197187.5 ;
      RECT  7745.0 197537.5 8125.0 197467.5 ;
      RECT  8090.0 197892.5 8160.0 197502.5 ;
      RECT  7710.0 197187.5 7780.0 197052.5 ;
      RECT  8090.0 197187.5 8160.0 197052.5 ;
      RECT  8090.0 198027.5 8160.0 197892.5 ;
      RECT  8090.0 197570.0 8160.0 197435.0 ;
      RECT  8090.0 198487.5 8160.0 199192.5 ;
      RECT  7710.0 198842.5 7780.0 198912.5 ;
      RECT  8090.0 198842.5 8160.0 198912.5 ;
      RECT  7710.0 198877.5 7780.0 199192.5 ;
      RECT  7745.0 198842.5 8125.0 198912.5 ;
      RECT  8090.0 198487.5 8160.0 198877.5 ;
      RECT  7710.0 199192.5 7780.0 199327.5 ;
      RECT  8090.0 199192.5 8160.0 199327.5 ;
      RECT  8090.0 198352.5 8160.0 198487.5 ;
      RECT  8090.0 198810.0 8160.0 198945.0 ;
      RECT  8090.0 200582.5 8160.0 199877.5 ;
      RECT  7710.0 200227.5 7780.0 200157.5 ;
      RECT  8090.0 200227.5 8160.0 200157.5 ;
      RECT  7710.0 200192.5 7780.0 199877.5 ;
      RECT  7745.0 200227.5 8125.0 200157.5 ;
      RECT  8090.0 200582.5 8160.0 200192.5 ;
      RECT  7710.0 199877.5 7780.0 199742.5 ;
      RECT  8090.0 199877.5 8160.0 199742.5 ;
      RECT  8090.0 200717.5 8160.0 200582.5 ;
      RECT  8090.0 200260.0 8160.0 200125.0 ;
      RECT  8090.0 201177.5 8160.0 201882.5 ;
      RECT  7710.0 201532.5 7780.0 201602.5 ;
      RECT  8090.0 201532.5 8160.0 201602.5 ;
      RECT  7710.0 201567.5 7780.0 201882.5 ;
      RECT  7745.0 201532.5 8125.0 201602.5 ;
      RECT  8090.0 201177.5 8160.0 201567.5 ;
      RECT  7710.0 201882.5 7780.0 202017.5 ;
      RECT  8090.0 201882.5 8160.0 202017.5 ;
      RECT  8090.0 201042.5 8160.0 201177.5 ;
      RECT  8090.0 201500.0 8160.0 201635.0 ;
      RECT  8090.0 203272.5 8160.0 202567.5 ;
      RECT  7710.0 202917.5 7780.0 202847.5 ;
      RECT  8090.0 202917.5 8160.0 202847.5 ;
      RECT  7710.0 202882.5 7780.0 202567.5 ;
      RECT  7745.0 202917.5 8125.0 202847.5 ;
      RECT  8090.0 203272.5 8160.0 202882.5 ;
      RECT  7710.0 202567.5 7780.0 202432.5 ;
      RECT  8090.0 202567.5 8160.0 202432.5 ;
      RECT  8090.0 203407.5 8160.0 203272.5 ;
      RECT  8090.0 202950.0 8160.0 202815.0 ;
      RECT  8090.0 203867.5 8160.0 204572.5 ;
      RECT  7710.0 204222.5 7780.0 204292.5 ;
      RECT  8090.0 204222.5 8160.0 204292.5 ;
      RECT  7710.0 204257.5 7780.0 204572.5 ;
      RECT  7745.0 204222.5 8125.0 204292.5 ;
      RECT  8090.0 203867.5 8160.0 204257.5 ;
      RECT  7710.0 204572.5 7780.0 204707.5 ;
      RECT  8090.0 204572.5 8160.0 204707.5 ;
      RECT  8090.0 203732.5 8160.0 203867.5 ;
      RECT  8090.0 204190.0 8160.0 204325.0 ;
      RECT  8090.0 205962.5 8160.0 205257.5 ;
      RECT  7710.0 205607.5 7780.0 205537.5 ;
      RECT  8090.0 205607.5 8160.0 205537.5 ;
      RECT  7710.0 205572.5 7780.0 205257.5 ;
      RECT  7745.0 205607.5 8125.0 205537.5 ;
      RECT  8090.0 205962.5 8160.0 205572.5 ;
      RECT  7710.0 205257.5 7780.0 205122.5 ;
      RECT  8090.0 205257.5 8160.0 205122.5 ;
      RECT  8090.0 206097.5 8160.0 205962.5 ;
      RECT  8090.0 205640.0 8160.0 205505.0 ;
      RECT  4757.5 13172.5 4622.5 13242.5 ;
      RECT  4932.5 14607.5 4797.5 14677.5 ;
      RECT  5107.5 15862.5 4972.5 15932.5 ;
      RECT  5282.5 17297.5 5147.5 17367.5 ;
      RECT  5457.5 18552.5 5322.5 18622.5 ;
      RECT  5632.5 19987.5 5497.5 20057.5 ;
      RECT  5807.5 21242.5 5672.5 21312.5 ;
      RECT  5982.5 22677.5 5847.5 22747.5 ;
      RECT  6157.5 23932.5 6022.5 24002.5 ;
      RECT  6332.5 25367.5 6197.5 25437.5 ;
      RECT  6507.5 26622.5 6372.5 26692.5 ;
      RECT  6682.5 28057.5 6547.5 28127.5 ;
      RECT  6857.5 29312.5 6722.5 29382.5 ;
      RECT  7032.5 30747.5 6897.5 30817.5 ;
      RECT  7207.5 32002.5 7072.5 32072.5 ;
      RECT  7382.5 33437.5 7247.5 33507.5 ;
      RECT  4757.5 34752.5 4622.5 34822.5 ;
      RECT  5457.5 34612.5 5322.5 34682.5 ;
      RECT  6157.5 34472.5 6022.5 34542.5 ;
      RECT  4757.5 36067.5 4622.5 36137.5 ;
      RECT  5457.5 36207.5 5322.5 36277.5 ;
      RECT  6332.5 36347.5 6197.5 36417.5 ;
      RECT  4757.5 37442.5 4622.5 37512.5 ;
      RECT  5457.5 37302.5 5322.5 37372.5 ;
      RECT  6507.5 37162.5 6372.5 37232.5 ;
      RECT  4757.5 38757.5 4622.5 38827.5 ;
      RECT  5457.5 38897.5 5322.5 38967.5 ;
      RECT  6682.5 39037.5 6547.5 39107.5 ;
      RECT  4757.5 40132.5 4622.5 40202.5 ;
      RECT  5457.5 39992.5 5322.5 40062.5 ;
      RECT  6857.5 39852.5 6722.5 39922.5 ;
      RECT  4757.5 41447.5 4622.5 41517.5 ;
      RECT  5457.5 41587.5 5322.5 41657.5 ;
      RECT  7032.5 41727.5 6897.5 41797.5 ;
      RECT  4757.5 42822.5 4622.5 42892.5 ;
      RECT  5457.5 42682.5 5322.5 42752.5 ;
      RECT  7207.5 42542.5 7072.5 42612.5 ;
      RECT  4757.5 44137.5 4622.5 44207.5 ;
      RECT  5457.5 44277.5 5322.5 44347.5 ;
      RECT  7382.5 44417.5 7247.5 44487.5 ;
      RECT  4757.5 45512.5 4622.5 45582.5 ;
      RECT  5632.5 45372.5 5497.5 45442.5 ;
      RECT  6157.5 45232.5 6022.5 45302.5 ;
      RECT  4757.5 46827.5 4622.5 46897.5 ;
      RECT  5632.5 46967.5 5497.5 47037.5 ;
      RECT  6332.5 47107.5 6197.5 47177.5 ;
      RECT  4757.5 48202.5 4622.5 48272.5 ;
      RECT  5632.5 48062.5 5497.5 48132.5 ;
      RECT  6507.5 47922.5 6372.5 47992.5 ;
      RECT  4757.5 49517.5 4622.5 49587.5 ;
      RECT  5632.5 49657.5 5497.5 49727.5 ;
      RECT  6682.5 49797.5 6547.5 49867.5 ;
      RECT  4757.5 50892.5 4622.5 50962.5 ;
      RECT  5632.5 50752.5 5497.5 50822.5 ;
      RECT  6857.5 50612.5 6722.5 50682.5 ;
      RECT  4757.5 52207.5 4622.5 52277.5 ;
      RECT  5632.5 52347.5 5497.5 52417.5 ;
      RECT  7032.5 52487.5 6897.5 52557.5 ;
      RECT  4757.5 53582.5 4622.5 53652.5 ;
      RECT  5632.5 53442.5 5497.5 53512.5 ;
      RECT  7207.5 53302.5 7072.5 53372.5 ;
      RECT  4757.5 54897.5 4622.5 54967.5 ;
      RECT  5632.5 55037.5 5497.5 55107.5 ;
      RECT  7382.5 55177.5 7247.5 55247.5 ;
      RECT  4757.5 56272.5 4622.5 56342.5 ;
      RECT  5807.5 56132.5 5672.5 56202.5 ;
      RECT  6157.5 55992.5 6022.5 56062.5 ;
      RECT  4757.5 57587.5 4622.5 57657.5 ;
      RECT  5807.5 57727.5 5672.5 57797.5 ;
      RECT  6332.5 57867.5 6197.5 57937.5 ;
      RECT  4757.5 58962.5 4622.5 59032.5 ;
      RECT  5807.5 58822.5 5672.5 58892.5 ;
      RECT  6507.5 58682.5 6372.5 58752.5 ;
      RECT  4757.5 60277.5 4622.5 60347.5 ;
      RECT  5807.5 60417.5 5672.5 60487.5 ;
      RECT  6682.5 60557.5 6547.5 60627.5 ;
      RECT  4757.5 61652.5 4622.5 61722.5 ;
      RECT  5807.5 61512.5 5672.5 61582.5 ;
      RECT  6857.5 61372.5 6722.5 61442.5 ;
      RECT  4757.5 62967.5 4622.5 63037.5 ;
      RECT  5807.5 63107.5 5672.5 63177.5 ;
      RECT  7032.5 63247.5 6897.5 63317.5 ;
      RECT  4757.5 64342.5 4622.5 64412.5 ;
      RECT  5807.5 64202.5 5672.5 64272.5 ;
      RECT  7207.5 64062.5 7072.5 64132.5 ;
      RECT  4757.5 65657.5 4622.5 65727.5 ;
      RECT  5807.5 65797.5 5672.5 65867.5 ;
      RECT  7382.5 65937.5 7247.5 66007.5 ;
      RECT  4757.5 67032.5 4622.5 67102.5 ;
      RECT  5982.5 66892.5 5847.5 66962.5 ;
      RECT  6157.5 66752.5 6022.5 66822.5 ;
      RECT  4757.5 68347.5 4622.5 68417.5 ;
      RECT  5982.5 68487.5 5847.5 68557.5 ;
      RECT  6332.5 68627.5 6197.5 68697.5 ;
      RECT  4757.5 69722.5 4622.5 69792.5 ;
      RECT  5982.5 69582.5 5847.5 69652.5 ;
      RECT  6507.5 69442.5 6372.5 69512.5 ;
      RECT  4757.5 71037.5 4622.5 71107.5 ;
      RECT  5982.5 71177.5 5847.5 71247.5 ;
      RECT  6682.5 71317.5 6547.5 71387.5 ;
      RECT  4757.5 72412.5 4622.5 72482.5 ;
      RECT  5982.5 72272.5 5847.5 72342.5 ;
      RECT  6857.5 72132.5 6722.5 72202.5 ;
      RECT  4757.5 73727.5 4622.5 73797.5 ;
      RECT  5982.5 73867.5 5847.5 73937.5 ;
      RECT  7032.5 74007.5 6897.5 74077.5 ;
      RECT  4757.5 75102.5 4622.5 75172.5 ;
      RECT  5982.5 74962.5 5847.5 75032.5 ;
      RECT  7207.5 74822.5 7072.5 74892.5 ;
      RECT  4757.5 76417.5 4622.5 76487.5 ;
      RECT  5982.5 76557.5 5847.5 76627.5 ;
      RECT  7382.5 76697.5 7247.5 76767.5 ;
      RECT  4932.5 77792.5 4797.5 77862.5 ;
      RECT  5457.5 77652.5 5322.5 77722.5 ;
      RECT  6157.5 77512.5 6022.5 77582.5 ;
      RECT  4932.5 79107.5 4797.5 79177.5 ;
      RECT  5457.5 79247.5 5322.5 79317.5 ;
      RECT  6332.5 79387.5 6197.5 79457.5 ;
      RECT  4932.5 80482.5 4797.5 80552.5 ;
      RECT  5457.5 80342.5 5322.5 80412.5 ;
      RECT  6507.5 80202.5 6372.5 80272.5 ;
      RECT  4932.5 81797.5 4797.5 81867.5 ;
      RECT  5457.5 81937.5 5322.5 82007.5 ;
      RECT  6682.5 82077.5 6547.5 82147.5 ;
      RECT  4932.5 83172.5 4797.5 83242.5 ;
      RECT  5457.5 83032.5 5322.5 83102.5 ;
      RECT  6857.5 82892.5 6722.5 82962.5 ;
      RECT  4932.5 84487.5 4797.5 84557.5 ;
      RECT  5457.5 84627.5 5322.5 84697.5 ;
      RECT  7032.5 84767.5 6897.5 84837.5 ;
      RECT  4932.5 85862.5 4797.5 85932.5 ;
      RECT  5457.5 85722.5 5322.5 85792.5 ;
      RECT  7207.5 85582.5 7072.5 85652.5 ;
      RECT  4932.5 87177.5 4797.5 87247.5 ;
      RECT  5457.5 87317.5 5322.5 87387.5 ;
      RECT  7382.5 87457.5 7247.5 87527.5 ;
      RECT  4932.5 88552.5 4797.5 88622.5 ;
      RECT  5632.5 88412.5 5497.5 88482.5 ;
      RECT  6157.5 88272.5 6022.5 88342.5 ;
      RECT  4932.5 89867.5 4797.5 89937.5 ;
      RECT  5632.5 90007.5 5497.5 90077.5 ;
      RECT  6332.5 90147.5 6197.5 90217.5 ;
      RECT  4932.5 91242.5 4797.5 91312.5 ;
      RECT  5632.5 91102.5 5497.5 91172.5 ;
      RECT  6507.5 90962.5 6372.5 91032.5 ;
      RECT  4932.5 92557.5 4797.5 92627.5 ;
      RECT  5632.5 92697.5 5497.5 92767.5 ;
      RECT  6682.5 92837.5 6547.5 92907.5 ;
      RECT  4932.5 93932.5 4797.5 94002.5 ;
      RECT  5632.5 93792.5 5497.5 93862.5 ;
      RECT  6857.5 93652.5 6722.5 93722.5 ;
      RECT  4932.5 95247.5 4797.5 95317.5 ;
      RECT  5632.5 95387.5 5497.5 95457.5 ;
      RECT  7032.5 95527.5 6897.5 95597.5 ;
      RECT  4932.5 96622.5 4797.5 96692.5 ;
      RECT  5632.5 96482.5 5497.5 96552.5 ;
      RECT  7207.5 96342.5 7072.5 96412.5 ;
      RECT  4932.5 97937.5 4797.5 98007.5 ;
      RECT  5632.5 98077.5 5497.5 98147.5 ;
      RECT  7382.5 98217.5 7247.5 98287.5 ;
      RECT  4932.5 99312.5 4797.5 99382.5 ;
      RECT  5807.5 99172.5 5672.5 99242.5 ;
      RECT  6157.5 99032.5 6022.5 99102.5 ;
      RECT  4932.5 100627.5 4797.5 100697.5 ;
      RECT  5807.5 100767.5 5672.5 100837.5 ;
      RECT  6332.5 100907.5 6197.5 100977.5 ;
      RECT  4932.5 102002.5 4797.5 102072.5 ;
      RECT  5807.5 101862.5 5672.5 101932.5 ;
      RECT  6507.5 101722.5 6372.5 101792.5 ;
      RECT  4932.5 103317.5 4797.5 103387.5 ;
      RECT  5807.5 103457.5 5672.5 103527.5 ;
      RECT  6682.5 103597.5 6547.5 103667.5 ;
      RECT  4932.5 104692.5 4797.5 104762.5 ;
      RECT  5807.5 104552.5 5672.5 104622.5 ;
      RECT  6857.5 104412.5 6722.5 104482.5 ;
      RECT  4932.5 106007.5 4797.5 106077.5 ;
      RECT  5807.5 106147.5 5672.5 106217.5 ;
      RECT  7032.5 106287.5 6897.5 106357.5 ;
      RECT  4932.5 107382.5 4797.5 107452.5 ;
      RECT  5807.5 107242.5 5672.5 107312.5 ;
      RECT  7207.5 107102.5 7072.5 107172.5 ;
      RECT  4932.5 108697.5 4797.5 108767.5 ;
      RECT  5807.5 108837.5 5672.5 108907.5 ;
      RECT  7382.5 108977.5 7247.5 109047.5 ;
      RECT  4932.5 110072.5 4797.5 110142.5 ;
      RECT  5982.5 109932.5 5847.5 110002.5 ;
      RECT  6157.5 109792.5 6022.5 109862.5 ;
      RECT  4932.5 111387.5 4797.5 111457.5 ;
      RECT  5982.5 111527.5 5847.5 111597.5 ;
      RECT  6332.5 111667.5 6197.5 111737.5 ;
      RECT  4932.5 112762.5 4797.5 112832.5 ;
      RECT  5982.5 112622.5 5847.5 112692.5 ;
      RECT  6507.5 112482.5 6372.5 112552.5 ;
      RECT  4932.5 114077.5 4797.5 114147.5 ;
      RECT  5982.5 114217.5 5847.5 114287.5 ;
      RECT  6682.5 114357.5 6547.5 114427.5 ;
      RECT  4932.5 115452.5 4797.5 115522.5 ;
      RECT  5982.5 115312.5 5847.5 115382.5 ;
      RECT  6857.5 115172.5 6722.5 115242.5 ;
      RECT  4932.5 116767.5 4797.5 116837.5 ;
      RECT  5982.5 116907.5 5847.5 116977.5 ;
      RECT  7032.5 117047.5 6897.5 117117.5 ;
      RECT  4932.5 118142.5 4797.5 118212.5 ;
      RECT  5982.5 118002.5 5847.5 118072.5 ;
      RECT  7207.5 117862.5 7072.5 117932.5 ;
      RECT  4932.5 119457.5 4797.5 119527.5 ;
      RECT  5982.5 119597.5 5847.5 119667.5 ;
      RECT  7382.5 119737.5 7247.5 119807.5 ;
      RECT  5107.5 120832.5 4972.5 120902.5 ;
      RECT  5457.5 120692.5 5322.5 120762.5 ;
      RECT  6157.5 120552.5 6022.5 120622.5 ;
      RECT  5107.5 122147.5 4972.5 122217.5 ;
      RECT  5457.5 122287.5 5322.5 122357.5 ;
      RECT  6332.5 122427.5 6197.5 122497.5 ;
      RECT  5107.5 123522.5 4972.5 123592.5 ;
      RECT  5457.5 123382.5 5322.5 123452.5 ;
      RECT  6507.5 123242.5 6372.5 123312.5 ;
      RECT  5107.5 124837.5 4972.5 124907.5 ;
      RECT  5457.5 124977.5 5322.5 125047.5 ;
      RECT  6682.5 125117.5 6547.5 125187.5 ;
      RECT  5107.5 126212.5 4972.5 126282.5 ;
      RECT  5457.5 126072.5 5322.5 126142.5 ;
      RECT  6857.5 125932.5 6722.5 126002.5 ;
      RECT  5107.5 127527.5 4972.5 127597.5 ;
      RECT  5457.5 127667.5 5322.5 127737.5 ;
      RECT  7032.5 127807.5 6897.5 127877.5 ;
      RECT  5107.5 128902.5 4972.5 128972.5 ;
      RECT  5457.5 128762.5 5322.5 128832.5 ;
      RECT  7207.5 128622.5 7072.5 128692.5 ;
      RECT  5107.5 130217.5 4972.5 130287.5 ;
      RECT  5457.5 130357.5 5322.5 130427.5 ;
      RECT  7382.5 130497.5 7247.5 130567.5 ;
      RECT  5107.5 131592.5 4972.5 131662.5 ;
      RECT  5632.5 131452.5 5497.5 131522.5 ;
      RECT  6157.5 131312.5 6022.5 131382.5 ;
      RECT  5107.5 132907.5 4972.5 132977.5 ;
      RECT  5632.5 133047.5 5497.5 133117.5 ;
      RECT  6332.5 133187.5 6197.5 133257.5 ;
      RECT  5107.5 134282.5 4972.5 134352.5 ;
      RECT  5632.5 134142.5 5497.5 134212.5 ;
      RECT  6507.5 134002.5 6372.5 134072.5 ;
      RECT  5107.5 135597.5 4972.5 135667.5 ;
      RECT  5632.5 135737.5 5497.5 135807.5 ;
      RECT  6682.5 135877.5 6547.5 135947.5 ;
      RECT  5107.5 136972.5 4972.5 137042.5 ;
      RECT  5632.5 136832.5 5497.5 136902.5 ;
      RECT  6857.5 136692.5 6722.5 136762.5 ;
      RECT  5107.5 138287.5 4972.5 138357.5 ;
      RECT  5632.5 138427.5 5497.5 138497.5 ;
      RECT  7032.5 138567.5 6897.5 138637.5 ;
      RECT  5107.5 139662.5 4972.5 139732.5 ;
      RECT  5632.5 139522.5 5497.5 139592.5 ;
      RECT  7207.5 139382.5 7072.5 139452.5 ;
      RECT  5107.5 140977.5 4972.5 141047.5 ;
      RECT  5632.5 141117.5 5497.5 141187.5 ;
      RECT  7382.5 141257.5 7247.5 141327.5 ;
      RECT  5107.5 142352.5 4972.5 142422.5 ;
      RECT  5807.5 142212.5 5672.5 142282.5 ;
      RECT  6157.5 142072.5 6022.5 142142.5 ;
      RECT  5107.5 143667.5 4972.5 143737.5 ;
      RECT  5807.5 143807.5 5672.5 143877.5 ;
      RECT  6332.5 143947.5 6197.5 144017.5 ;
      RECT  5107.5 145042.5 4972.5 145112.5 ;
      RECT  5807.5 144902.5 5672.5 144972.5 ;
      RECT  6507.5 144762.5 6372.5 144832.5 ;
      RECT  5107.5 146357.5 4972.5 146427.5 ;
      RECT  5807.5 146497.5 5672.5 146567.5 ;
      RECT  6682.5 146637.5 6547.5 146707.5 ;
      RECT  5107.5 147732.5 4972.5 147802.5 ;
      RECT  5807.5 147592.5 5672.5 147662.5 ;
      RECT  6857.5 147452.5 6722.5 147522.5 ;
      RECT  5107.5 149047.5 4972.5 149117.5 ;
      RECT  5807.5 149187.5 5672.5 149257.5 ;
      RECT  7032.5 149327.5 6897.5 149397.5 ;
      RECT  5107.5 150422.5 4972.5 150492.5 ;
      RECT  5807.5 150282.5 5672.5 150352.5 ;
      RECT  7207.5 150142.5 7072.5 150212.5 ;
      RECT  5107.5 151737.5 4972.5 151807.5 ;
      RECT  5807.5 151877.5 5672.5 151947.5 ;
      RECT  7382.5 152017.5 7247.5 152087.5 ;
      RECT  5107.5 153112.5 4972.5 153182.5 ;
      RECT  5982.5 152972.5 5847.5 153042.5 ;
      RECT  6157.5 152832.5 6022.5 152902.5 ;
      RECT  5107.5 154427.5 4972.5 154497.5 ;
      RECT  5982.5 154567.5 5847.5 154637.5 ;
      RECT  6332.5 154707.5 6197.5 154777.5 ;
      RECT  5107.5 155802.5 4972.5 155872.5 ;
      RECT  5982.5 155662.5 5847.5 155732.5 ;
      RECT  6507.5 155522.5 6372.5 155592.5 ;
      RECT  5107.5 157117.5 4972.5 157187.5 ;
      RECT  5982.5 157257.5 5847.5 157327.5 ;
      RECT  6682.5 157397.5 6547.5 157467.5 ;
      RECT  5107.5 158492.5 4972.5 158562.5 ;
      RECT  5982.5 158352.5 5847.5 158422.5 ;
      RECT  6857.5 158212.5 6722.5 158282.5 ;
      RECT  5107.5 159807.5 4972.5 159877.5 ;
      RECT  5982.5 159947.5 5847.5 160017.5 ;
      RECT  7032.5 160087.5 6897.5 160157.5 ;
      RECT  5107.5 161182.5 4972.5 161252.5 ;
      RECT  5982.5 161042.5 5847.5 161112.5 ;
      RECT  7207.5 160902.5 7072.5 160972.5 ;
      RECT  5107.5 162497.5 4972.5 162567.5 ;
      RECT  5982.5 162637.5 5847.5 162707.5 ;
      RECT  7382.5 162777.5 7247.5 162847.5 ;
      RECT  5282.5 163872.5 5147.5 163942.5 ;
      RECT  5457.5 163732.5 5322.5 163802.5 ;
      RECT  6157.5 163592.5 6022.5 163662.5 ;
      RECT  5282.5 165187.5 5147.5 165257.5 ;
      RECT  5457.5 165327.5 5322.5 165397.5 ;
      RECT  6332.5 165467.5 6197.5 165537.5 ;
      RECT  5282.5 166562.5 5147.5 166632.5 ;
      RECT  5457.5 166422.5 5322.5 166492.5 ;
      RECT  6507.5 166282.5 6372.5 166352.5 ;
      RECT  5282.5 167877.5 5147.5 167947.5 ;
      RECT  5457.5 168017.5 5322.5 168087.5 ;
      RECT  6682.5 168157.5 6547.5 168227.5 ;
      RECT  5282.5 169252.5 5147.5 169322.5 ;
      RECT  5457.5 169112.5 5322.5 169182.5 ;
      RECT  6857.5 168972.5 6722.5 169042.5 ;
      RECT  5282.5 170567.5 5147.5 170637.5 ;
      RECT  5457.5 170707.5 5322.5 170777.5 ;
      RECT  7032.5 170847.5 6897.5 170917.5 ;
      RECT  5282.5 171942.5 5147.5 172012.5 ;
      RECT  5457.5 171802.5 5322.5 171872.5 ;
      RECT  7207.5 171662.5 7072.5 171732.5 ;
      RECT  5282.5 173257.5 5147.5 173327.5 ;
      RECT  5457.5 173397.5 5322.5 173467.5 ;
      RECT  7382.5 173537.5 7247.5 173607.5 ;
      RECT  5282.5 174632.5 5147.5 174702.5 ;
      RECT  5632.5 174492.5 5497.5 174562.5 ;
      RECT  6157.5 174352.5 6022.5 174422.5 ;
      RECT  5282.5 175947.5 5147.5 176017.5 ;
      RECT  5632.5 176087.5 5497.5 176157.5 ;
      RECT  6332.5 176227.5 6197.5 176297.5 ;
      RECT  5282.5 177322.5 5147.5 177392.5 ;
      RECT  5632.5 177182.5 5497.5 177252.5 ;
      RECT  6507.5 177042.5 6372.5 177112.5 ;
      RECT  5282.5 178637.5 5147.5 178707.5 ;
      RECT  5632.5 178777.5 5497.5 178847.5 ;
      RECT  6682.5 178917.5 6547.5 178987.5 ;
      RECT  5282.5 180012.5 5147.5 180082.5 ;
      RECT  5632.5 179872.5 5497.5 179942.5 ;
      RECT  6857.5 179732.5 6722.5 179802.5 ;
      RECT  5282.5 181327.5 5147.5 181397.5 ;
      RECT  5632.5 181467.5 5497.5 181537.5 ;
      RECT  7032.5 181607.5 6897.5 181677.5 ;
      RECT  5282.5 182702.5 5147.5 182772.5 ;
      RECT  5632.5 182562.5 5497.5 182632.5 ;
      RECT  7207.5 182422.5 7072.5 182492.5 ;
      RECT  5282.5 184017.5 5147.5 184087.5 ;
      RECT  5632.5 184157.5 5497.5 184227.5 ;
      RECT  7382.5 184297.5 7247.5 184367.5 ;
      RECT  5282.5 185392.5 5147.5 185462.5 ;
      RECT  5807.5 185252.5 5672.5 185322.5 ;
      RECT  6157.5 185112.5 6022.5 185182.5 ;
      RECT  5282.5 186707.5 5147.5 186777.5 ;
      RECT  5807.5 186847.5 5672.5 186917.5 ;
      RECT  6332.5 186987.5 6197.5 187057.5 ;
      RECT  5282.5 188082.5 5147.5 188152.5 ;
      RECT  5807.5 187942.5 5672.5 188012.5 ;
      RECT  6507.5 187802.5 6372.5 187872.5 ;
      RECT  5282.5 189397.5 5147.5 189467.5 ;
      RECT  5807.5 189537.5 5672.5 189607.5 ;
      RECT  6682.5 189677.5 6547.5 189747.5 ;
      RECT  5282.5 190772.5 5147.5 190842.5 ;
      RECT  5807.5 190632.5 5672.5 190702.5 ;
      RECT  6857.5 190492.5 6722.5 190562.5 ;
      RECT  5282.5 192087.5 5147.5 192157.5 ;
      RECT  5807.5 192227.5 5672.5 192297.5 ;
      RECT  7032.5 192367.5 6897.5 192437.5 ;
      RECT  5282.5 193462.5 5147.5 193532.5 ;
      RECT  5807.5 193322.5 5672.5 193392.5 ;
      RECT  7207.5 193182.5 7072.5 193252.5 ;
      RECT  5282.5 194777.5 5147.5 194847.5 ;
      RECT  5807.5 194917.5 5672.5 194987.5 ;
      RECT  7382.5 195057.5 7247.5 195127.5 ;
      RECT  5282.5 196152.5 5147.5 196222.5 ;
      RECT  5982.5 196012.5 5847.5 196082.5 ;
      RECT  6157.5 195872.5 6022.5 195942.5 ;
      RECT  5282.5 197467.5 5147.5 197537.5 ;
      RECT  5982.5 197607.5 5847.5 197677.5 ;
      RECT  6332.5 197747.5 6197.5 197817.5 ;
      RECT  5282.5 198842.5 5147.5 198912.5 ;
      RECT  5982.5 198702.5 5847.5 198772.5 ;
      RECT  6507.5 198562.5 6372.5 198632.5 ;
      RECT  5282.5 200157.5 5147.5 200227.5 ;
      RECT  5982.5 200297.5 5847.5 200367.5 ;
      RECT  6682.5 200437.5 6547.5 200507.5 ;
      RECT  5282.5 201532.5 5147.5 201602.5 ;
      RECT  5982.5 201392.5 5847.5 201462.5 ;
      RECT  6857.5 201252.5 6722.5 201322.5 ;
      RECT  5282.5 202847.5 5147.5 202917.5 ;
      RECT  5982.5 202987.5 5847.5 203057.5 ;
      RECT  7032.5 203127.5 6897.5 203197.5 ;
      RECT  5282.5 204222.5 5147.5 204292.5 ;
      RECT  5982.5 204082.5 5847.5 204152.5 ;
      RECT  7207.5 203942.5 7072.5 204012.5 ;
      RECT  5282.5 205537.5 5147.5 205607.5 ;
      RECT  5982.5 205677.5 5847.5 205747.5 ;
      RECT  7382.5 205817.5 7247.5 205887.5 ;
      RECT  11350.0 12580.0 11420.0 17820.0 ;
      RECT  11075.0 12580.0 11145.0 17820.0 ;
      RECT  11350.0 17960.0 11420.0 23200.0 ;
      RECT  11075.0 17960.0 11145.0 23200.0 ;
      RECT  12265.0 23340.0 12335.0 33960.0 ;
      RECT  11990.0 23340.0 12060.0 33960.0 ;
      RECT  11715.0 23340.0 11785.0 33960.0 ;
      RECT  9360.0 34490.0 9430.0 34560.0 ;
      RECT  9360.0 34455.0 9430.0 34525.0 ;
      RECT  9395.0 34490.0 10357.5 34560.0 ;
      RECT  9360.0 36330.0 9430.0 36400.0 ;
      RECT  9360.0 36365.0 9430.0 36435.0 ;
      RECT  9395.0 36330.0 10357.5 36400.0 ;
      RECT  9360.0 37180.0 9430.0 37250.0 ;
      RECT  9360.0 37145.0 9430.0 37215.0 ;
      RECT  9395.0 37180.0 10357.5 37250.0 ;
      RECT  9360.0 39020.0 9430.0 39090.0 ;
      RECT  9360.0 39055.0 9430.0 39125.0 ;
      RECT  9395.0 39020.0 10357.5 39090.0 ;
      RECT  9360.0 39870.0 9430.0 39940.0 ;
      RECT  9360.0 39835.0 9430.0 39905.0 ;
      RECT  9395.0 39870.0 10357.5 39940.0 ;
      RECT  9360.0 41710.0 9430.0 41780.0 ;
      RECT  9360.0 41745.0 9430.0 41815.0 ;
      RECT  9395.0 41710.0 10357.5 41780.0 ;
      RECT  9360.0 42560.0 9430.0 42630.0 ;
      RECT  9360.0 42525.0 9430.0 42595.0 ;
      RECT  9395.0 42560.0 10357.5 42630.0 ;
      RECT  9360.0 44400.0 9430.0 44470.0 ;
      RECT  9360.0 44435.0 9430.0 44505.0 ;
      RECT  9395.0 44400.0 10357.5 44470.0 ;
      RECT  9360.0 45250.0 9430.0 45320.0 ;
      RECT  9360.0 45215.0 9430.0 45285.0 ;
      RECT  9395.0 45250.0 10357.5 45320.0 ;
      RECT  9360.0 47090.0 9430.0 47160.0 ;
      RECT  9360.0 47125.0 9430.0 47195.0 ;
      RECT  9395.0 47090.0 10357.5 47160.0 ;
      RECT  9360.0 47940.0 9430.0 48010.0 ;
      RECT  9360.0 47905.0 9430.0 47975.0 ;
      RECT  9395.0 47940.0 10357.5 48010.0 ;
      RECT  9360.0 49780.0 9430.0 49850.0 ;
      RECT  9360.0 49815.0 9430.0 49885.0 ;
      RECT  9395.0 49780.0 10357.5 49850.0 ;
      RECT  9360.0 50630.0 9430.0 50700.0 ;
      RECT  9360.0 50595.0 9430.0 50665.0 ;
      RECT  9395.0 50630.0 10357.5 50700.0 ;
      RECT  9360.0 52470.0 9430.0 52540.0 ;
      RECT  9360.0 52505.0 9430.0 52575.0 ;
      RECT  9395.0 52470.0 10357.5 52540.0 ;
      RECT  9360.0 53320.0 9430.0 53390.0 ;
      RECT  9360.0 53285.0 9430.0 53355.0 ;
      RECT  9395.0 53320.0 10357.5 53390.0 ;
      RECT  9360.0 55160.0 9430.0 55230.0 ;
      RECT  9360.0 55195.0 9430.0 55265.0 ;
      RECT  9395.0 55160.0 10357.5 55230.0 ;
      RECT  9360.0 56010.0 9430.0 56080.0 ;
      RECT  9360.0 55975.0 9430.0 56045.0 ;
      RECT  9395.0 56010.0 10357.5 56080.0 ;
      RECT  9360.0 57850.0 9430.0 57920.0 ;
      RECT  9360.0 57885.0 9430.0 57955.0 ;
      RECT  9395.0 57850.0 10357.5 57920.0 ;
      RECT  9360.0 58700.0 9430.0 58770.0 ;
      RECT  9360.0 58665.0 9430.0 58735.0 ;
      RECT  9395.0 58700.0 10357.5 58770.0 ;
      RECT  9360.0 60540.0 9430.0 60610.0 ;
      RECT  9360.0 60575.0 9430.0 60645.0 ;
      RECT  9395.0 60540.0 10357.5 60610.0 ;
      RECT  9360.0 61390.0 9430.0 61460.0 ;
      RECT  9360.0 61355.0 9430.0 61425.0 ;
      RECT  9395.0 61390.0 10357.5 61460.0 ;
      RECT  9360.0 63230.0 9430.0 63300.0 ;
      RECT  9360.0 63265.0 9430.0 63335.0 ;
      RECT  9395.0 63230.0 10357.5 63300.0 ;
      RECT  9360.0 64080.0 9430.0 64150.0 ;
      RECT  9360.0 64045.0 9430.0 64115.0 ;
      RECT  9395.0 64080.0 10357.5 64150.0 ;
      RECT  9360.0 65920.0 9430.0 65990.0 ;
      RECT  9360.0 65955.0 9430.0 66025.0 ;
      RECT  9395.0 65920.0 10357.5 65990.0 ;
      RECT  9360.0 66770.0 9430.0 66840.0 ;
      RECT  9360.0 66735.0 9430.0 66805.0 ;
      RECT  9395.0 66770.0 10357.5 66840.0 ;
      RECT  9360.0 68610.0 9430.0 68680.0 ;
      RECT  9360.0 68645.0 9430.0 68715.0 ;
      RECT  9395.0 68610.0 10357.5 68680.0 ;
      RECT  9360.0 69460.0 9430.0 69530.0 ;
      RECT  9360.0 69425.0 9430.0 69495.0 ;
      RECT  9395.0 69460.0 10357.5 69530.0 ;
      RECT  9360.0 71300.0 9430.0 71370.0 ;
      RECT  9360.0 71335.0 9430.0 71405.0 ;
      RECT  9395.0 71300.0 10357.5 71370.0 ;
      RECT  9360.0 72150.0 9430.0 72220.0 ;
      RECT  9360.0 72115.0 9430.0 72185.0 ;
      RECT  9395.0 72150.0 10357.5 72220.0 ;
      RECT  9360.0 73990.0 9430.0 74060.0 ;
      RECT  9360.0 74025.0 9430.0 74095.0 ;
      RECT  9395.0 73990.0 10357.5 74060.0 ;
      RECT  9360.0 74840.0 9430.0 74910.0 ;
      RECT  9360.0 74805.0 9430.0 74875.0 ;
      RECT  9395.0 74840.0 10357.5 74910.0 ;
      RECT  9360.0 76680.0 9430.0 76750.0 ;
      RECT  9360.0 76715.0 9430.0 76785.0 ;
      RECT  9395.0 76680.0 10357.5 76750.0 ;
      RECT  9360.0 77530.0 9430.0 77600.0 ;
      RECT  9360.0 77495.0 9430.0 77565.0 ;
      RECT  9395.0 77530.0 10357.5 77600.0 ;
      RECT  9360.0 79370.0 9430.0 79440.0 ;
      RECT  9360.0 79405.0 9430.0 79475.0 ;
      RECT  9395.0 79370.0 10357.5 79440.0 ;
      RECT  9360.0 80220.0 9430.0 80290.0 ;
      RECT  9360.0 80185.0 9430.0 80255.0 ;
      RECT  9395.0 80220.0 10357.5 80290.0 ;
      RECT  9360.0 82060.0 9430.0 82130.0 ;
      RECT  9360.0 82095.0 9430.0 82165.0 ;
      RECT  9395.0 82060.0 10357.5 82130.0 ;
      RECT  9360.0 82910.0 9430.0 82980.0 ;
      RECT  9360.0 82875.0 9430.0 82945.0 ;
      RECT  9395.0 82910.0 10357.5 82980.0 ;
      RECT  9360.0 84750.0 9430.0 84820.0 ;
      RECT  9360.0 84785.0 9430.0 84855.0 ;
      RECT  9395.0 84750.0 10357.5 84820.0 ;
      RECT  9360.0 85600.0 9430.0 85670.0 ;
      RECT  9360.0 85565.0 9430.0 85635.0 ;
      RECT  9395.0 85600.0 10357.5 85670.0 ;
      RECT  9360.0 87440.0 9430.0 87510.0 ;
      RECT  9360.0 87475.0 9430.0 87545.0 ;
      RECT  9395.0 87440.0 10357.5 87510.0 ;
      RECT  9360.0 88290.0 9430.0 88360.0 ;
      RECT  9360.0 88255.0 9430.0 88325.0 ;
      RECT  9395.0 88290.0 10357.5 88360.0 ;
      RECT  9360.0 90130.0 9430.0 90200.0 ;
      RECT  9360.0 90165.0 9430.0 90235.0 ;
      RECT  9395.0 90130.0 10357.5 90200.0 ;
      RECT  9360.0 90980.0 9430.0 91050.0 ;
      RECT  9360.0 90945.0 9430.0 91015.0 ;
      RECT  9395.0 90980.0 10357.5 91050.0 ;
      RECT  9360.0 92820.0 9430.0 92890.0 ;
      RECT  9360.0 92855.0 9430.0 92925.0 ;
      RECT  9395.0 92820.0 10357.5 92890.0 ;
      RECT  9360.0 93670.0 9430.0 93740.0 ;
      RECT  9360.0 93635.0 9430.0 93705.0 ;
      RECT  9395.0 93670.0 10357.5 93740.0 ;
      RECT  9360.0 95510.0 9430.0 95580.0 ;
      RECT  9360.0 95545.0 9430.0 95615.0 ;
      RECT  9395.0 95510.0 10357.5 95580.0 ;
      RECT  9360.0 96360.0 9430.0 96430.0 ;
      RECT  9360.0 96325.0 9430.0 96395.0 ;
      RECT  9395.0 96360.0 10357.5 96430.0 ;
      RECT  9360.0 98200.0 9430.0 98270.0 ;
      RECT  9360.0 98235.0 9430.0 98305.0 ;
      RECT  9395.0 98200.0 10357.5 98270.0 ;
      RECT  9360.0 99050.0 9430.0 99120.0 ;
      RECT  9360.0 99015.0 9430.0 99085.0 ;
      RECT  9395.0 99050.0 10357.5 99120.0 ;
      RECT  9360.0 100890.0 9430.0 100960.0 ;
      RECT  9360.0 100925.0 9430.0 100995.0 ;
      RECT  9395.0 100890.0 10357.5 100960.0 ;
      RECT  9360.0 101740.0 9430.0 101810.0 ;
      RECT  9360.0 101705.0 9430.0 101775.0 ;
      RECT  9395.0 101740.0 10357.5 101810.0 ;
      RECT  9360.0 103580.0 9430.0 103650.0 ;
      RECT  9360.0 103615.0 9430.0 103685.0 ;
      RECT  9395.0 103580.0 10357.5 103650.0 ;
      RECT  9360.0 104430.0 9430.0 104500.0 ;
      RECT  9360.0 104395.0 9430.0 104465.0 ;
      RECT  9395.0 104430.0 10357.5 104500.0 ;
      RECT  9360.0 106270.0 9430.0 106340.0 ;
      RECT  9360.0 106305.0 9430.0 106375.0 ;
      RECT  9395.0 106270.0 10357.5 106340.0 ;
      RECT  9360.0 107120.0 9430.0 107190.0 ;
      RECT  9360.0 107085.0 9430.0 107155.0 ;
      RECT  9395.0 107120.0 10357.5 107190.0 ;
      RECT  9360.0 108960.0 9430.0 109030.0 ;
      RECT  9360.0 108995.0 9430.0 109065.0 ;
      RECT  9395.0 108960.0 10357.5 109030.0 ;
      RECT  9360.0 109810.0 9430.0 109880.0 ;
      RECT  9360.0 109775.0 9430.0 109845.0 ;
      RECT  9395.0 109810.0 10357.5 109880.0 ;
      RECT  9360.0 111650.0 9430.0 111720.0 ;
      RECT  9360.0 111685.0 9430.0 111755.0 ;
      RECT  9395.0 111650.0 10357.5 111720.0 ;
      RECT  9360.0 112500.0 9430.0 112570.0 ;
      RECT  9360.0 112465.0 9430.0 112535.0 ;
      RECT  9395.0 112500.0 10357.5 112570.0 ;
      RECT  9360.0 114340.0 9430.0 114410.0 ;
      RECT  9360.0 114375.0 9430.0 114445.0 ;
      RECT  9395.0 114340.0 10357.5 114410.0 ;
      RECT  9360.0 115190.0 9430.0 115260.0 ;
      RECT  9360.0 115155.0 9430.0 115225.0 ;
      RECT  9395.0 115190.0 10357.5 115260.0 ;
      RECT  9360.0 117030.0 9430.0 117100.0 ;
      RECT  9360.0 117065.0 9430.0 117135.0 ;
      RECT  9395.0 117030.0 10357.5 117100.0 ;
      RECT  9360.0 117880.0 9430.0 117950.0 ;
      RECT  9360.0 117845.0 9430.0 117915.0 ;
      RECT  9395.0 117880.0 10357.5 117950.0 ;
      RECT  9360.0 119720.0 9430.0 119790.0 ;
      RECT  9360.0 119755.0 9430.0 119825.0 ;
      RECT  9395.0 119720.0 10357.5 119790.0 ;
      RECT  9360.0 120570.0 9430.0 120640.0 ;
      RECT  9360.0 120535.0 9430.0 120605.0 ;
      RECT  9395.0 120570.0 10357.5 120640.0 ;
      RECT  9360.0 122410.0 9430.0 122480.0 ;
      RECT  9360.0 122445.0 9430.0 122515.0 ;
      RECT  9395.0 122410.0 10357.5 122480.0 ;
      RECT  9360.0 123260.0 9430.0 123330.0 ;
      RECT  9360.0 123225.0 9430.0 123295.0 ;
      RECT  9395.0 123260.0 10357.5 123330.0 ;
      RECT  9360.0 125100.0 9430.0 125170.0 ;
      RECT  9360.0 125135.0 9430.0 125205.0 ;
      RECT  9395.0 125100.0 10357.5 125170.0 ;
      RECT  9360.0 125950.0 9430.0 126020.0 ;
      RECT  9360.0 125915.0 9430.0 125985.0 ;
      RECT  9395.0 125950.0 10357.5 126020.0 ;
      RECT  9360.0 127790.0 9430.0 127860.0 ;
      RECT  9360.0 127825.0 9430.0 127895.0 ;
      RECT  9395.0 127790.0 10357.5 127860.0 ;
      RECT  9360.0 128640.0 9430.0 128710.0 ;
      RECT  9360.0 128605.0 9430.0 128675.0 ;
      RECT  9395.0 128640.0 10357.5 128710.0 ;
      RECT  9360.0 130480.0 9430.0 130550.0 ;
      RECT  9360.0 130515.0 9430.0 130585.0 ;
      RECT  9395.0 130480.0 10357.5 130550.0 ;
      RECT  9360.0 131330.0 9430.0 131400.0 ;
      RECT  9360.0 131295.0 9430.0 131365.0 ;
      RECT  9395.0 131330.0 10357.5 131400.0 ;
      RECT  9360.0 133170.0 9430.0 133240.0 ;
      RECT  9360.0 133205.0 9430.0 133275.0 ;
      RECT  9395.0 133170.0 10357.5 133240.0 ;
      RECT  9360.0 134020.0 9430.0 134090.0 ;
      RECT  9360.0 133985.0 9430.0 134055.0 ;
      RECT  9395.0 134020.0 10357.5 134090.0 ;
      RECT  9360.0 135860.0 9430.0 135930.0 ;
      RECT  9360.0 135895.0 9430.0 135965.0 ;
      RECT  9395.0 135860.0 10357.5 135930.0 ;
      RECT  9360.0 136710.0 9430.0 136780.0 ;
      RECT  9360.0 136675.0 9430.0 136745.0 ;
      RECT  9395.0 136710.0 10357.5 136780.0 ;
      RECT  9360.0 138550.0 9430.0 138620.0 ;
      RECT  9360.0 138585.0 9430.0 138655.0 ;
      RECT  9395.0 138550.0 10357.5 138620.0 ;
      RECT  9360.0 139400.0 9430.0 139470.0 ;
      RECT  9360.0 139365.0 9430.0 139435.0 ;
      RECT  9395.0 139400.0 10357.5 139470.0 ;
      RECT  9360.0 141240.0 9430.0 141310.0 ;
      RECT  9360.0 141275.0 9430.0 141345.0 ;
      RECT  9395.0 141240.0 10357.5 141310.0 ;
      RECT  9360.0 142090.0 9430.0 142160.0 ;
      RECT  9360.0 142055.0 9430.0 142125.0 ;
      RECT  9395.0 142090.0 10357.5 142160.0 ;
      RECT  9360.0 143930.0 9430.0 144000.0 ;
      RECT  9360.0 143965.0 9430.0 144035.0 ;
      RECT  9395.0 143930.0 10357.5 144000.0 ;
      RECT  9360.0 144780.0 9430.0 144850.0 ;
      RECT  9360.0 144745.0 9430.0 144815.0 ;
      RECT  9395.0 144780.0 10357.5 144850.0 ;
      RECT  9360.0 146620.0 9430.0 146690.0 ;
      RECT  9360.0 146655.0 9430.0 146725.0 ;
      RECT  9395.0 146620.0 10357.5 146690.0 ;
      RECT  9360.0 147470.0 9430.0 147540.0 ;
      RECT  9360.0 147435.0 9430.0 147505.0 ;
      RECT  9395.0 147470.0 10357.5 147540.0 ;
      RECT  9360.0 149310.0 9430.0 149380.0 ;
      RECT  9360.0 149345.0 9430.0 149415.0 ;
      RECT  9395.0 149310.0 10357.5 149380.0 ;
      RECT  9360.0 150160.0 9430.0 150230.0 ;
      RECT  9360.0 150125.0 9430.0 150195.0 ;
      RECT  9395.0 150160.0 10357.5 150230.0 ;
      RECT  9360.0 152000.0 9430.0 152070.0 ;
      RECT  9360.0 152035.0 9430.0 152105.0 ;
      RECT  9395.0 152000.0 10357.5 152070.0 ;
      RECT  9360.0 152850.0 9430.0 152920.0 ;
      RECT  9360.0 152815.0 9430.0 152885.0 ;
      RECT  9395.0 152850.0 10357.5 152920.0 ;
      RECT  9360.0 154690.0 9430.0 154760.0 ;
      RECT  9360.0 154725.0 9430.0 154795.0 ;
      RECT  9395.0 154690.0 10357.5 154760.0 ;
      RECT  9360.0 155540.0 9430.0 155610.0 ;
      RECT  9360.0 155505.0 9430.0 155575.0 ;
      RECT  9395.0 155540.0 10357.5 155610.0 ;
      RECT  9360.0 157380.0 9430.0 157450.0 ;
      RECT  9360.0 157415.0 9430.0 157485.0 ;
      RECT  9395.0 157380.0 10357.5 157450.0 ;
      RECT  9360.0 158230.0 9430.0 158300.0 ;
      RECT  9360.0 158195.0 9430.0 158265.0 ;
      RECT  9395.0 158230.0 10357.5 158300.0 ;
      RECT  9360.0 160070.0 9430.0 160140.0 ;
      RECT  9360.0 160105.0 9430.0 160175.0 ;
      RECT  9395.0 160070.0 10357.5 160140.0 ;
      RECT  9360.0 160920.0 9430.0 160990.0 ;
      RECT  9360.0 160885.0 9430.0 160955.0 ;
      RECT  9395.0 160920.0 10357.5 160990.0 ;
      RECT  9360.0 162760.0 9430.0 162830.0 ;
      RECT  9360.0 162795.0 9430.0 162865.0 ;
      RECT  9395.0 162760.0 10357.5 162830.0 ;
      RECT  9360.0 163610.0 9430.0 163680.0 ;
      RECT  9360.0 163575.0 9430.0 163645.0 ;
      RECT  9395.0 163610.0 10357.5 163680.0 ;
      RECT  9360.0 165450.0 9430.0 165520.0 ;
      RECT  9360.0 165485.0 9430.0 165555.0 ;
      RECT  9395.0 165450.0 10357.5 165520.0 ;
      RECT  9360.0 166300.0 9430.0 166370.0 ;
      RECT  9360.0 166265.0 9430.0 166335.0 ;
      RECT  9395.0 166300.0 10357.5 166370.0 ;
      RECT  9360.0 168140.0 9430.0 168210.0 ;
      RECT  9360.0 168175.0 9430.0 168245.0 ;
      RECT  9395.0 168140.0 10357.5 168210.0 ;
      RECT  9360.0 168990.0 9430.0 169060.0 ;
      RECT  9360.0 168955.0 9430.0 169025.0 ;
      RECT  9395.0 168990.0 10357.5 169060.0 ;
      RECT  9360.0 170830.0 9430.0 170900.0 ;
      RECT  9360.0 170865.0 9430.0 170935.0 ;
      RECT  9395.0 170830.0 10357.5 170900.0 ;
      RECT  9360.0 171680.0 9430.0 171750.0 ;
      RECT  9360.0 171645.0 9430.0 171715.0 ;
      RECT  9395.0 171680.0 10357.5 171750.0 ;
      RECT  9360.0 173520.0 9430.0 173590.0 ;
      RECT  9360.0 173555.0 9430.0 173625.0 ;
      RECT  9395.0 173520.0 10357.5 173590.0 ;
      RECT  9360.0 174370.0 9430.0 174440.0 ;
      RECT  9360.0 174335.0 9430.0 174405.0 ;
      RECT  9395.0 174370.0 10357.5 174440.0 ;
      RECT  9360.0 176210.0 9430.0 176280.0 ;
      RECT  9360.0 176245.0 9430.0 176315.0 ;
      RECT  9395.0 176210.0 10357.5 176280.0 ;
      RECT  9360.0 177060.0 9430.0 177130.0 ;
      RECT  9360.0 177025.0 9430.0 177095.0 ;
      RECT  9395.0 177060.0 10357.5 177130.0 ;
      RECT  9360.0 178900.0 9430.0 178970.0 ;
      RECT  9360.0 178935.0 9430.0 179005.0 ;
      RECT  9395.0 178900.0 10357.5 178970.0 ;
      RECT  9360.0 179750.0 9430.0 179820.0 ;
      RECT  9360.0 179715.0 9430.0 179785.0 ;
      RECT  9395.0 179750.0 10357.5 179820.0 ;
      RECT  9360.0 181590.0 9430.0 181660.0 ;
      RECT  9360.0 181625.0 9430.0 181695.0 ;
      RECT  9395.0 181590.0 10357.5 181660.0 ;
      RECT  9360.0 182440.0 9430.0 182510.0 ;
      RECT  9360.0 182405.0 9430.0 182475.0 ;
      RECT  9395.0 182440.0 10357.5 182510.0 ;
      RECT  9360.0 184280.0 9430.0 184350.0 ;
      RECT  9360.0 184315.0 9430.0 184385.0 ;
      RECT  9395.0 184280.0 10357.5 184350.0 ;
      RECT  9360.0 185130.0 9430.0 185200.0 ;
      RECT  9360.0 185095.0 9430.0 185165.0 ;
      RECT  9395.0 185130.0 10357.5 185200.0 ;
      RECT  9360.0 186970.0 9430.0 187040.0 ;
      RECT  9360.0 187005.0 9430.0 187075.0 ;
      RECT  9395.0 186970.0 10357.5 187040.0 ;
      RECT  9360.0 187820.0 9430.0 187890.0 ;
      RECT  9360.0 187785.0 9430.0 187855.0 ;
      RECT  9395.0 187820.0 10357.5 187890.0 ;
      RECT  9360.0 189660.0 9430.0 189730.0 ;
      RECT  9360.0 189695.0 9430.0 189765.0 ;
      RECT  9395.0 189660.0 10357.5 189730.0 ;
      RECT  9360.0 190510.0 9430.0 190580.0 ;
      RECT  9360.0 190475.0 9430.0 190545.0 ;
      RECT  9395.0 190510.0 10357.5 190580.0 ;
      RECT  9360.0 192350.0 9430.0 192420.0 ;
      RECT  9360.0 192385.0 9430.0 192455.0 ;
      RECT  9395.0 192350.0 10357.5 192420.0 ;
      RECT  9360.0 193200.0 9430.0 193270.0 ;
      RECT  9360.0 193165.0 9430.0 193235.0 ;
      RECT  9395.0 193200.0 10357.5 193270.0 ;
      RECT  9360.0 195040.0 9430.0 195110.0 ;
      RECT  9360.0 195075.0 9430.0 195145.0 ;
      RECT  9395.0 195040.0 10357.5 195110.0 ;
      RECT  9360.0 195890.0 9430.0 195960.0 ;
      RECT  9360.0 195855.0 9430.0 195925.0 ;
      RECT  9395.0 195890.0 10357.5 195960.0 ;
      RECT  9360.0 197730.0 9430.0 197800.0 ;
      RECT  9360.0 197765.0 9430.0 197835.0 ;
      RECT  9395.0 197730.0 10357.5 197800.0 ;
      RECT  9360.0 198580.0 9430.0 198650.0 ;
      RECT  9360.0 198545.0 9430.0 198615.0 ;
      RECT  9395.0 198580.0 10357.5 198650.0 ;
      RECT  9360.0 200420.0 9430.0 200490.0 ;
      RECT  9360.0 200455.0 9430.0 200525.0 ;
      RECT  9395.0 200420.0 10357.5 200490.0 ;
      RECT  9360.0 201270.0 9430.0 201340.0 ;
      RECT  9360.0 201235.0 9430.0 201305.0 ;
      RECT  9395.0 201270.0 10357.5 201340.0 ;
      RECT  9360.0 203110.0 9430.0 203180.0 ;
      RECT  9360.0 203145.0 9430.0 203215.0 ;
      RECT  9395.0 203110.0 10357.5 203180.0 ;
      RECT  9360.0 203960.0 9430.0 204030.0 ;
      RECT  9360.0 203925.0 9430.0 203995.0 ;
      RECT  9395.0 203960.0 10357.5 204030.0 ;
      RECT  9360.0 205800.0 9430.0 205870.0 ;
      RECT  9360.0 205835.0 9430.0 205905.0 ;
      RECT  9395.0 205800.0 10357.5 205870.0 ;
      RECT  10295.0 34705.0 10365.0 34775.0 ;
      RECT  10485.0 34705.0 10555.0 34775.0 ;
      RECT  10295.0 34740.0 10365.0 35102.5 ;
      RECT  10330.0 34705.0 10520.0 34775.0 ;
      RECT  10485.0 34397.5 10555.0 34740.0 ;
      RECT  10295.0 35102.5 10365.0 35237.5 ;
      RECT  10485.0 34262.5 10555.0 34397.5 ;
      RECT  10587.5 34705.0 10452.5 34775.0 ;
      RECT  9220.0 34660.0 9290.0 34795.0 ;
      RECT  9360.0 34387.5 9430.0 34522.5 ;
      RECT  10357.5 34490.0 10222.5 34560.0 ;
      RECT  10295.0 36185.0 10365.0 36115.0 ;
      RECT  10485.0 36185.0 10555.0 36115.0 ;
      RECT  10295.0 36150.0 10365.0 35787.5 ;
      RECT  10330.0 36185.0 10520.0 36115.0 ;
      RECT  10485.0 36492.5 10555.0 36150.0 ;
      RECT  10295.0 35787.5 10365.0 35652.5 ;
      RECT  10485.0 36627.5 10555.0 36492.5 ;
      RECT  10587.5 36185.0 10452.5 36115.0 ;
      RECT  9220.0 36095.0 9290.0 36230.0 ;
      RECT  9360.0 36367.5 9430.0 36502.5 ;
      RECT  10357.5 36330.0 10222.5 36400.0 ;
      RECT  10295.0 37395.0 10365.0 37465.0 ;
      RECT  10485.0 37395.0 10555.0 37465.0 ;
      RECT  10295.0 37430.0 10365.0 37792.5 ;
      RECT  10330.0 37395.0 10520.0 37465.0 ;
      RECT  10485.0 37087.5 10555.0 37430.0 ;
      RECT  10295.0 37792.5 10365.0 37927.5 ;
      RECT  10485.0 36952.5 10555.0 37087.5 ;
      RECT  10587.5 37395.0 10452.5 37465.0 ;
      RECT  9220.0 37350.0 9290.0 37485.0 ;
      RECT  9360.0 37077.5 9430.0 37212.5 ;
      RECT  10357.5 37180.0 10222.5 37250.0 ;
      RECT  10295.0 38875.0 10365.0 38805.0 ;
      RECT  10485.0 38875.0 10555.0 38805.0 ;
      RECT  10295.0 38840.0 10365.0 38477.5 ;
      RECT  10330.0 38875.0 10520.0 38805.0 ;
      RECT  10485.0 39182.5 10555.0 38840.0 ;
      RECT  10295.0 38477.5 10365.0 38342.5 ;
      RECT  10485.0 39317.5 10555.0 39182.5 ;
      RECT  10587.5 38875.0 10452.5 38805.0 ;
      RECT  9220.0 38785.0 9290.0 38920.0 ;
      RECT  9360.0 39057.5 9430.0 39192.5 ;
      RECT  10357.5 39020.0 10222.5 39090.0 ;
      RECT  10295.0 40085.0 10365.0 40155.0 ;
      RECT  10485.0 40085.0 10555.0 40155.0 ;
      RECT  10295.0 40120.0 10365.0 40482.5 ;
      RECT  10330.0 40085.0 10520.0 40155.0 ;
      RECT  10485.0 39777.5 10555.0 40120.0 ;
      RECT  10295.0 40482.5 10365.0 40617.5 ;
      RECT  10485.0 39642.5 10555.0 39777.5 ;
      RECT  10587.5 40085.0 10452.5 40155.0 ;
      RECT  9220.0 40040.0 9290.0 40175.0 ;
      RECT  9360.0 39767.5 9430.0 39902.5 ;
      RECT  10357.5 39870.0 10222.5 39940.0 ;
      RECT  10295.0 41565.0 10365.0 41495.0 ;
      RECT  10485.0 41565.0 10555.0 41495.0 ;
      RECT  10295.0 41530.0 10365.0 41167.5 ;
      RECT  10330.0 41565.0 10520.0 41495.0 ;
      RECT  10485.0 41872.5 10555.0 41530.0 ;
      RECT  10295.0 41167.5 10365.0 41032.5 ;
      RECT  10485.0 42007.5 10555.0 41872.5 ;
      RECT  10587.5 41565.0 10452.5 41495.0 ;
      RECT  9220.0 41475.0 9290.0 41610.0 ;
      RECT  9360.0 41747.5 9430.0 41882.5 ;
      RECT  10357.5 41710.0 10222.5 41780.0 ;
      RECT  10295.0 42775.0 10365.0 42845.0 ;
      RECT  10485.0 42775.0 10555.0 42845.0 ;
      RECT  10295.0 42810.0 10365.0 43172.5 ;
      RECT  10330.0 42775.0 10520.0 42845.0 ;
      RECT  10485.0 42467.5 10555.0 42810.0 ;
      RECT  10295.0 43172.5 10365.0 43307.5 ;
      RECT  10485.0 42332.5 10555.0 42467.5 ;
      RECT  10587.5 42775.0 10452.5 42845.0 ;
      RECT  9220.0 42730.0 9290.0 42865.0 ;
      RECT  9360.0 42457.5 9430.0 42592.5 ;
      RECT  10357.5 42560.0 10222.5 42630.0 ;
      RECT  10295.0 44255.0 10365.0 44185.0 ;
      RECT  10485.0 44255.0 10555.0 44185.0 ;
      RECT  10295.0 44220.0 10365.0 43857.5 ;
      RECT  10330.0 44255.0 10520.0 44185.0 ;
      RECT  10485.0 44562.5 10555.0 44220.0 ;
      RECT  10295.0 43857.5 10365.0 43722.5 ;
      RECT  10485.0 44697.5 10555.0 44562.5 ;
      RECT  10587.5 44255.0 10452.5 44185.0 ;
      RECT  9220.0 44165.0 9290.0 44300.0 ;
      RECT  9360.0 44437.5 9430.0 44572.5 ;
      RECT  10357.5 44400.0 10222.5 44470.0 ;
      RECT  10295.0 45465.0 10365.0 45535.0 ;
      RECT  10485.0 45465.0 10555.0 45535.0 ;
      RECT  10295.0 45500.0 10365.0 45862.5 ;
      RECT  10330.0 45465.0 10520.0 45535.0 ;
      RECT  10485.0 45157.5 10555.0 45500.0 ;
      RECT  10295.0 45862.5 10365.0 45997.5 ;
      RECT  10485.0 45022.5 10555.0 45157.5 ;
      RECT  10587.5 45465.0 10452.5 45535.0 ;
      RECT  9220.0 45420.0 9290.0 45555.0 ;
      RECT  9360.0 45147.5 9430.0 45282.5 ;
      RECT  10357.5 45250.0 10222.5 45320.0 ;
      RECT  10295.0 46945.0 10365.0 46875.0 ;
      RECT  10485.0 46945.0 10555.0 46875.0 ;
      RECT  10295.0 46910.0 10365.0 46547.5 ;
      RECT  10330.0 46945.0 10520.0 46875.0 ;
      RECT  10485.0 47252.5 10555.0 46910.0 ;
      RECT  10295.0 46547.5 10365.0 46412.5 ;
      RECT  10485.0 47387.5 10555.0 47252.5 ;
      RECT  10587.5 46945.0 10452.5 46875.0 ;
      RECT  9220.0 46855.0 9290.0 46990.0 ;
      RECT  9360.0 47127.5 9430.0 47262.5 ;
      RECT  10357.5 47090.0 10222.5 47160.0 ;
      RECT  10295.0 48155.0 10365.0 48225.0 ;
      RECT  10485.0 48155.0 10555.0 48225.0 ;
      RECT  10295.0 48190.0 10365.0 48552.5 ;
      RECT  10330.0 48155.0 10520.0 48225.0 ;
      RECT  10485.0 47847.5 10555.0 48190.0 ;
      RECT  10295.0 48552.5 10365.0 48687.5 ;
      RECT  10485.0 47712.5 10555.0 47847.5 ;
      RECT  10587.5 48155.0 10452.5 48225.0 ;
      RECT  9220.0 48110.0 9290.0 48245.0 ;
      RECT  9360.0 47837.5 9430.0 47972.5 ;
      RECT  10357.5 47940.0 10222.5 48010.0 ;
      RECT  10295.0 49635.0 10365.0 49565.0 ;
      RECT  10485.0 49635.0 10555.0 49565.0 ;
      RECT  10295.0 49600.0 10365.0 49237.5 ;
      RECT  10330.0 49635.0 10520.0 49565.0 ;
      RECT  10485.0 49942.5 10555.0 49600.0 ;
      RECT  10295.0 49237.5 10365.0 49102.5 ;
      RECT  10485.0 50077.5 10555.0 49942.5 ;
      RECT  10587.5 49635.0 10452.5 49565.0 ;
      RECT  9220.0 49545.0 9290.0 49680.0 ;
      RECT  9360.0 49817.5 9430.0 49952.5 ;
      RECT  10357.5 49780.0 10222.5 49850.0 ;
      RECT  10295.0 50845.0 10365.0 50915.0 ;
      RECT  10485.0 50845.0 10555.0 50915.0 ;
      RECT  10295.0 50880.0 10365.0 51242.5 ;
      RECT  10330.0 50845.0 10520.0 50915.0 ;
      RECT  10485.0 50537.5 10555.0 50880.0 ;
      RECT  10295.0 51242.5 10365.0 51377.5 ;
      RECT  10485.0 50402.5 10555.0 50537.5 ;
      RECT  10587.5 50845.0 10452.5 50915.0 ;
      RECT  9220.0 50800.0 9290.0 50935.0 ;
      RECT  9360.0 50527.5 9430.0 50662.5 ;
      RECT  10357.5 50630.0 10222.5 50700.0 ;
      RECT  10295.0 52325.0 10365.0 52255.0 ;
      RECT  10485.0 52325.0 10555.0 52255.0 ;
      RECT  10295.0 52290.0 10365.0 51927.5 ;
      RECT  10330.0 52325.0 10520.0 52255.0 ;
      RECT  10485.0 52632.5 10555.0 52290.0 ;
      RECT  10295.0 51927.5 10365.0 51792.5 ;
      RECT  10485.0 52767.5 10555.0 52632.5 ;
      RECT  10587.5 52325.0 10452.5 52255.0 ;
      RECT  9220.0 52235.0 9290.0 52370.0 ;
      RECT  9360.0 52507.5 9430.0 52642.5 ;
      RECT  10357.5 52470.0 10222.5 52540.0 ;
      RECT  10295.0 53535.0 10365.0 53605.0 ;
      RECT  10485.0 53535.0 10555.0 53605.0 ;
      RECT  10295.0 53570.0 10365.0 53932.5 ;
      RECT  10330.0 53535.0 10520.0 53605.0 ;
      RECT  10485.0 53227.5 10555.0 53570.0 ;
      RECT  10295.0 53932.5 10365.0 54067.5 ;
      RECT  10485.0 53092.5 10555.0 53227.5 ;
      RECT  10587.5 53535.0 10452.5 53605.0 ;
      RECT  9220.0 53490.0 9290.0 53625.0 ;
      RECT  9360.0 53217.5 9430.0 53352.5 ;
      RECT  10357.5 53320.0 10222.5 53390.0 ;
      RECT  10295.0 55015.0 10365.0 54945.0 ;
      RECT  10485.0 55015.0 10555.0 54945.0 ;
      RECT  10295.0 54980.0 10365.0 54617.5 ;
      RECT  10330.0 55015.0 10520.0 54945.0 ;
      RECT  10485.0 55322.5 10555.0 54980.0 ;
      RECT  10295.0 54617.5 10365.0 54482.5 ;
      RECT  10485.0 55457.5 10555.0 55322.5 ;
      RECT  10587.5 55015.0 10452.5 54945.0 ;
      RECT  9220.0 54925.0 9290.0 55060.0 ;
      RECT  9360.0 55197.5 9430.0 55332.5 ;
      RECT  10357.5 55160.0 10222.5 55230.0 ;
      RECT  10295.0 56225.0 10365.0 56295.0 ;
      RECT  10485.0 56225.0 10555.0 56295.0 ;
      RECT  10295.0 56260.0 10365.0 56622.5 ;
      RECT  10330.0 56225.0 10520.0 56295.0 ;
      RECT  10485.0 55917.5 10555.0 56260.0 ;
      RECT  10295.0 56622.5 10365.0 56757.5 ;
      RECT  10485.0 55782.5 10555.0 55917.5 ;
      RECT  10587.5 56225.0 10452.5 56295.0 ;
      RECT  9220.0 56180.0 9290.0 56315.0 ;
      RECT  9360.0 55907.5 9430.0 56042.5 ;
      RECT  10357.5 56010.0 10222.5 56080.0 ;
      RECT  10295.0 57705.0 10365.0 57635.0 ;
      RECT  10485.0 57705.0 10555.0 57635.0 ;
      RECT  10295.0 57670.0 10365.0 57307.5 ;
      RECT  10330.0 57705.0 10520.0 57635.0 ;
      RECT  10485.0 58012.5 10555.0 57670.0 ;
      RECT  10295.0 57307.5 10365.0 57172.5 ;
      RECT  10485.0 58147.5 10555.0 58012.5 ;
      RECT  10587.5 57705.0 10452.5 57635.0 ;
      RECT  9220.0 57615.0 9290.0 57750.0 ;
      RECT  9360.0 57887.5 9430.0 58022.5 ;
      RECT  10357.5 57850.0 10222.5 57920.0 ;
      RECT  10295.0 58915.0 10365.0 58985.0 ;
      RECT  10485.0 58915.0 10555.0 58985.0 ;
      RECT  10295.0 58950.0 10365.0 59312.5 ;
      RECT  10330.0 58915.0 10520.0 58985.0 ;
      RECT  10485.0 58607.5 10555.0 58950.0 ;
      RECT  10295.0 59312.5 10365.0 59447.5 ;
      RECT  10485.0 58472.5 10555.0 58607.5 ;
      RECT  10587.5 58915.0 10452.5 58985.0 ;
      RECT  9220.0 58870.0 9290.0 59005.0 ;
      RECT  9360.0 58597.5 9430.0 58732.5 ;
      RECT  10357.5 58700.0 10222.5 58770.0 ;
      RECT  10295.0 60395.0 10365.0 60325.0 ;
      RECT  10485.0 60395.0 10555.0 60325.0 ;
      RECT  10295.0 60360.0 10365.0 59997.5 ;
      RECT  10330.0 60395.0 10520.0 60325.0 ;
      RECT  10485.0 60702.5 10555.0 60360.0 ;
      RECT  10295.0 59997.5 10365.0 59862.5 ;
      RECT  10485.0 60837.5 10555.0 60702.5 ;
      RECT  10587.5 60395.0 10452.5 60325.0 ;
      RECT  9220.0 60305.0 9290.0 60440.0 ;
      RECT  9360.0 60577.5 9430.0 60712.5 ;
      RECT  10357.5 60540.0 10222.5 60610.0 ;
      RECT  10295.0 61605.0 10365.0 61675.0 ;
      RECT  10485.0 61605.0 10555.0 61675.0 ;
      RECT  10295.0 61640.0 10365.0 62002.5 ;
      RECT  10330.0 61605.0 10520.0 61675.0 ;
      RECT  10485.0 61297.5 10555.0 61640.0 ;
      RECT  10295.0 62002.5 10365.0 62137.5 ;
      RECT  10485.0 61162.5 10555.0 61297.5 ;
      RECT  10587.5 61605.0 10452.5 61675.0 ;
      RECT  9220.0 61560.0 9290.0 61695.0 ;
      RECT  9360.0 61287.5 9430.0 61422.5 ;
      RECT  10357.5 61390.0 10222.5 61460.0 ;
      RECT  10295.0 63085.0 10365.0 63015.0 ;
      RECT  10485.0 63085.0 10555.0 63015.0 ;
      RECT  10295.0 63050.0 10365.0 62687.5 ;
      RECT  10330.0 63085.0 10520.0 63015.0 ;
      RECT  10485.0 63392.5 10555.0 63050.0 ;
      RECT  10295.0 62687.5 10365.0 62552.5 ;
      RECT  10485.0 63527.5 10555.0 63392.5 ;
      RECT  10587.5 63085.0 10452.5 63015.0 ;
      RECT  9220.0 62995.0 9290.0 63130.0 ;
      RECT  9360.0 63267.5 9430.0 63402.5 ;
      RECT  10357.5 63230.0 10222.5 63300.0 ;
      RECT  10295.0 64295.0 10365.0 64365.0 ;
      RECT  10485.0 64295.0 10555.0 64365.0 ;
      RECT  10295.0 64330.0 10365.0 64692.5 ;
      RECT  10330.0 64295.0 10520.0 64365.0 ;
      RECT  10485.0 63987.5 10555.0 64330.0 ;
      RECT  10295.0 64692.5 10365.0 64827.5 ;
      RECT  10485.0 63852.5 10555.0 63987.5 ;
      RECT  10587.5 64295.0 10452.5 64365.0 ;
      RECT  9220.0 64250.0 9290.0 64385.0 ;
      RECT  9360.0 63977.5 9430.0 64112.5 ;
      RECT  10357.5 64080.0 10222.5 64150.0 ;
      RECT  10295.0 65775.0 10365.0 65705.0 ;
      RECT  10485.0 65775.0 10555.0 65705.0 ;
      RECT  10295.0 65740.0 10365.0 65377.5 ;
      RECT  10330.0 65775.0 10520.0 65705.0 ;
      RECT  10485.0 66082.5 10555.0 65740.0 ;
      RECT  10295.0 65377.5 10365.0 65242.5 ;
      RECT  10485.0 66217.5 10555.0 66082.5 ;
      RECT  10587.5 65775.0 10452.5 65705.0 ;
      RECT  9220.0 65685.0 9290.0 65820.0 ;
      RECT  9360.0 65957.5 9430.0 66092.5 ;
      RECT  10357.5 65920.0 10222.5 65990.0 ;
      RECT  10295.0 66985.0 10365.0 67055.0 ;
      RECT  10485.0 66985.0 10555.0 67055.0 ;
      RECT  10295.0 67020.0 10365.0 67382.5 ;
      RECT  10330.0 66985.0 10520.0 67055.0 ;
      RECT  10485.0 66677.5 10555.0 67020.0 ;
      RECT  10295.0 67382.5 10365.0 67517.5 ;
      RECT  10485.0 66542.5 10555.0 66677.5 ;
      RECT  10587.5 66985.0 10452.5 67055.0 ;
      RECT  9220.0 66940.0 9290.0 67075.0 ;
      RECT  9360.0 66667.5 9430.0 66802.5 ;
      RECT  10357.5 66770.0 10222.5 66840.0 ;
      RECT  10295.0 68465.0 10365.0 68395.0 ;
      RECT  10485.0 68465.0 10555.0 68395.0 ;
      RECT  10295.0 68430.0 10365.0 68067.5 ;
      RECT  10330.0 68465.0 10520.0 68395.0 ;
      RECT  10485.0 68772.5 10555.0 68430.0 ;
      RECT  10295.0 68067.5 10365.0 67932.5 ;
      RECT  10485.0 68907.5 10555.0 68772.5 ;
      RECT  10587.5 68465.0 10452.5 68395.0 ;
      RECT  9220.0 68375.0 9290.0 68510.0 ;
      RECT  9360.0 68647.5 9430.0 68782.5 ;
      RECT  10357.5 68610.0 10222.5 68680.0 ;
      RECT  10295.0 69675.0 10365.0 69745.0 ;
      RECT  10485.0 69675.0 10555.0 69745.0 ;
      RECT  10295.0 69710.0 10365.0 70072.5 ;
      RECT  10330.0 69675.0 10520.0 69745.0 ;
      RECT  10485.0 69367.5 10555.0 69710.0 ;
      RECT  10295.0 70072.5 10365.0 70207.5 ;
      RECT  10485.0 69232.5 10555.0 69367.5 ;
      RECT  10587.5 69675.0 10452.5 69745.0 ;
      RECT  9220.0 69630.0 9290.0 69765.0 ;
      RECT  9360.0 69357.5 9430.0 69492.5 ;
      RECT  10357.5 69460.0 10222.5 69530.0 ;
      RECT  10295.0 71155.0 10365.0 71085.0 ;
      RECT  10485.0 71155.0 10555.0 71085.0 ;
      RECT  10295.0 71120.0 10365.0 70757.5 ;
      RECT  10330.0 71155.0 10520.0 71085.0 ;
      RECT  10485.0 71462.5 10555.0 71120.0 ;
      RECT  10295.0 70757.5 10365.0 70622.5 ;
      RECT  10485.0 71597.5 10555.0 71462.5 ;
      RECT  10587.5 71155.0 10452.5 71085.0 ;
      RECT  9220.0 71065.0 9290.0 71200.0 ;
      RECT  9360.0 71337.5 9430.0 71472.5 ;
      RECT  10357.5 71300.0 10222.5 71370.0 ;
      RECT  10295.0 72365.0 10365.0 72435.0 ;
      RECT  10485.0 72365.0 10555.0 72435.0 ;
      RECT  10295.0 72400.0 10365.0 72762.5 ;
      RECT  10330.0 72365.0 10520.0 72435.0 ;
      RECT  10485.0 72057.5 10555.0 72400.0 ;
      RECT  10295.0 72762.5 10365.0 72897.5 ;
      RECT  10485.0 71922.5 10555.0 72057.5 ;
      RECT  10587.5 72365.0 10452.5 72435.0 ;
      RECT  9220.0 72320.0 9290.0 72455.0 ;
      RECT  9360.0 72047.5 9430.0 72182.5 ;
      RECT  10357.5 72150.0 10222.5 72220.0 ;
      RECT  10295.0 73845.0 10365.0 73775.0 ;
      RECT  10485.0 73845.0 10555.0 73775.0 ;
      RECT  10295.0 73810.0 10365.0 73447.5 ;
      RECT  10330.0 73845.0 10520.0 73775.0 ;
      RECT  10485.0 74152.5 10555.0 73810.0 ;
      RECT  10295.0 73447.5 10365.0 73312.5 ;
      RECT  10485.0 74287.5 10555.0 74152.5 ;
      RECT  10587.5 73845.0 10452.5 73775.0 ;
      RECT  9220.0 73755.0 9290.0 73890.0 ;
      RECT  9360.0 74027.5 9430.0 74162.5 ;
      RECT  10357.5 73990.0 10222.5 74060.0 ;
      RECT  10295.0 75055.0 10365.0 75125.0 ;
      RECT  10485.0 75055.0 10555.0 75125.0 ;
      RECT  10295.0 75090.0 10365.0 75452.5 ;
      RECT  10330.0 75055.0 10520.0 75125.0 ;
      RECT  10485.0 74747.5 10555.0 75090.0 ;
      RECT  10295.0 75452.5 10365.0 75587.5 ;
      RECT  10485.0 74612.5 10555.0 74747.5 ;
      RECT  10587.5 75055.0 10452.5 75125.0 ;
      RECT  9220.0 75010.0 9290.0 75145.0 ;
      RECT  9360.0 74737.5 9430.0 74872.5 ;
      RECT  10357.5 74840.0 10222.5 74910.0 ;
      RECT  10295.0 76535.0 10365.0 76465.0 ;
      RECT  10485.0 76535.0 10555.0 76465.0 ;
      RECT  10295.0 76500.0 10365.0 76137.5 ;
      RECT  10330.0 76535.0 10520.0 76465.0 ;
      RECT  10485.0 76842.5 10555.0 76500.0 ;
      RECT  10295.0 76137.5 10365.0 76002.5 ;
      RECT  10485.0 76977.5 10555.0 76842.5 ;
      RECT  10587.5 76535.0 10452.5 76465.0 ;
      RECT  9220.0 76445.0 9290.0 76580.0 ;
      RECT  9360.0 76717.5 9430.0 76852.5 ;
      RECT  10357.5 76680.0 10222.5 76750.0 ;
      RECT  10295.0 77745.0 10365.0 77815.0 ;
      RECT  10485.0 77745.0 10555.0 77815.0 ;
      RECT  10295.0 77780.0 10365.0 78142.5 ;
      RECT  10330.0 77745.0 10520.0 77815.0 ;
      RECT  10485.0 77437.5 10555.0 77780.0 ;
      RECT  10295.0 78142.5 10365.0 78277.5 ;
      RECT  10485.0 77302.5 10555.0 77437.5 ;
      RECT  10587.5 77745.0 10452.5 77815.0 ;
      RECT  9220.0 77700.0 9290.0 77835.0 ;
      RECT  9360.0 77427.5 9430.0 77562.5 ;
      RECT  10357.5 77530.0 10222.5 77600.0 ;
      RECT  10295.0 79225.0 10365.0 79155.0 ;
      RECT  10485.0 79225.0 10555.0 79155.0 ;
      RECT  10295.0 79190.0 10365.0 78827.5 ;
      RECT  10330.0 79225.0 10520.0 79155.0 ;
      RECT  10485.0 79532.5 10555.0 79190.0 ;
      RECT  10295.0 78827.5 10365.0 78692.5 ;
      RECT  10485.0 79667.5 10555.0 79532.5 ;
      RECT  10587.5 79225.0 10452.5 79155.0 ;
      RECT  9220.0 79135.0 9290.0 79270.0 ;
      RECT  9360.0 79407.5 9430.0 79542.5 ;
      RECT  10357.5 79370.0 10222.5 79440.0 ;
      RECT  10295.0 80435.0 10365.0 80505.0 ;
      RECT  10485.0 80435.0 10555.0 80505.0 ;
      RECT  10295.0 80470.0 10365.0 80832.5 ;
      RECT  10330.0 80435.0 10520.0 80505.0 ;
      RECT  10485.0 80127.5 10555.0 80470.0 ;
      RECT  10295.0 80832.5 10365.0 80967.5 ;
      RECT  10485.0 79992.5 10555.0 80127.5 ;
      RECT  10587.5 80435.0 10452.5 80505.0 ;
      RECT  9220.0 80390.0 9290.0 80525.0 ;
      RECT  9360.0 80117.5 9430.0 80252.5 ;
      RECT  10357.5 80220.0 10222.5 80290.0 ;
      RECT  10295.0 81915.0 10365.0 81845.0 ;
      RECT  10485.0 81915.0 10555.0 81845.0 ;
      RECT  10295.0 81880.0 10365.0 81517.5 ;
      RECT  10330.0 81915.0 10520.0 81845.0 ;
      RECT  10485.0 82222.5 10555.0 81880.0 ;
      RECT  10295.0 81517.5 10365.0 81382.5 ;
      RECT  10485.0 82357.5 10555.0 82222.5 ;
      RECT  10587.5 81915.0 10452.5 81845.0 ;
      RECT  9220.0 81825.0 9290.0 81960.0 ;
      RECT  9360.0 82097.5 9430.0 82232.5 ;
      RECT  10357.5 82060.0 10222.5 82130.0 ;
      RECT  10295.0 83125.0 10365.0 83195.0 ;
      RECT  10485.0 83125.0 10555.0 83195.0 ;
      RECT  10295.0 83160.0 10365.0 83522.5 ;
      RECT  10330.0 83125.0 10520.0 83195.0 ;
      RECT  10485.0 82817.5 10555.0 83160.0 ;
      RECT  10295.0 83522.5 10365.0 83657.5 ;
      RECT  10485.0 82682.5 10555.0 82817.5 ;
      RECT  10587.5 83125.0 10452.5 83195.0 ;
      RECT  9220.0 83080.0 9290.0 83215.0 ;
      RECT  9360.0 82807.5 9430.0 82942.5 ;
      RECT  10357.5 82910.0 10222.5 82980.0 ;
      RECT  10295.0 84605.0 10365.0 84535.0 ;
      RECT  10485.0 84605.0 10555.0 84535.0 ;
      RECT  10295.0 84570.0 10365.0 84207.5 ;
      RECT  10330.0 84605.0 10520.0 84535.0 ;
      RECT  10485.0 84912.5 10555.0 84570.0 ;
      RECT  10295.0 84207.5 10365.0 84072.5 ;
      RECT  10485.0 85047.5 10555.0 84912.5 ;
      RECT  10587.5 84605.0 10452.5 84535.0 ;
      RECT  9220.0 84515.0 9290.0 84650.0 ;
      RECT  9360.0 84787.5 9430.0 84922.5 ;
      RECT  10357.5 84750.0 10222.5 84820.0 ;
      RECT  10295.0 85815.0 10365.0 85885.0 ;
      RECT  10485.0 85815.0 10555.0 85885.0 ;
      RECT  10295.0 85850.0 10365.0 86212.5 ;
      RECT  10330.0 85815.0 10520.0 85885.0 ;
      RECT  10485.0 85507.5 10555.0 85850.0 ;
      RECT  10295.0 86212.5 10365.0 86347.5 ;
      RECT  10485.0 85372.5 10555.0 85507.5 ;
      RECT  10587.5 85815.0 10452.5 85885.0 ;
      RECT  9220.0 85770.0 9290.0 85905.0 ;
      RECT  9360.0 85497.5 9430.0 85632.5 ;
      RECT  10357.5 85600.0 10222.5 85670.0 ;
      RECT  10295.0 87295.0 10365.0 87225.0 ;
      RECT  10485.0 87295.0 10555.0 87225.0 ;
      RECT  10295.0 87260.0 10365.0 86897.5 ;
      RECT  10330.0 87295.0 10520.0 87225.0 ;
      RECT  10485.0 87602.5 10555.0 87260.0 ;
      RECT  10295.0 86897.5 10365.0 86762.5 ;
      RECT  10485.0 87737.5 10555.0 87602.5 ;
      RECT  10587.5 87295.0 10452.5 87225.0 ;
      RECT  9220.0 87205.0 9290.0 87340.0 ;
      RECT  9360.0 87477.5 9430.0 87612.5 ;
      RECT  10357.5 87440.0 10222.5 87510.0 ;
      RECT  10295.0 88505.0 10365.0 88575.0 ;
      RECT  10485.0 88505.0 10555.0 88575.0 ;
      RECT  10295.0 88540.0 10365.0 88902.5 ;
      RECT  10330.0 88505.0 10520.0 88575.0 ;
      RECT  10485.0 88197.5 10555.0 88540.0 ;
      RECT  10295.0 88902.5 10365.0 89037.5 ;
      RECT  10485.0 88062.5 10555.0 88197.5 ;
      RECT  10587.5 88505.0 10452.5 88575.0 ;
      RECT  9220.0 88460.0 9290.0 88595.0 ;
      RECT  9360.0 88187.5 9430.0 88322.5 ;
      RECT  10357.5 88290.0 10222.5 88360.0 ;
      RECT  10295.0 89985.0 10365.0 89915.0 ;
      RECT  10485.0 89985.0 10555.0 89915.0 ;
      RECT  10295.0 89950.0 10365.0 89587.5 ;
      RECT  10330.0 89985.0 10520.0 89915.0 ;
      RECT  10485.0 90292.5 10555.0 89950.0 ;
      RECT  10295.0 89587.5 10365.0 89452.5 ;
      RECT  10485.0 90427.5 10555.0 90292.5 ;
      RECT  10587.5 89985.0 10452.5 89915.0 ;
      RECT  9220.0 89895.0 9290.0 90030.0 ;
      RECT  9360.0 90167.5 9430.0 90302.5 ;
      RECT  10357.5 90130.0 10222.5 90200.0 ;
      RECT  10295.0 91195.0 10365.0 91265.0 ;
      RECT  10485.0 91195.0 10555.0 91265.0 ;
      RECT  10295.0 91230.0 10365.0 91592.5 ;
      RECT  10330.0 91195.0 10520.0 91265.0 ;
      RECT  10485.0 90887.5 10555.0 91230.0 ;
      RECT  10295.0 91592.5 10365.0 91727.5 ;
      RECT  10485.0 90752.5 10555.0 90887.5 ;
      RECT  10587.5 91195.0 10452.5 91265.0 ;
      RECT  9220.0 91150.0 9290.0 91285.0 ;
      RECT  9360.0 90877.5 9430.0 91012.5 ;
      RECT  10357.5 90980.0 10222.5 91050.0 ;
      RECT  10295.0 92675.0 10365.0 92605.0 ;
      RECT  10485.0 92675.0 10555.0 92605.0 ;
      RECT  10295.0 92640.0 10365.0 92277.5 ;
      RECT  10330.0 92675.0 10520.0 92605.0 ;
      RECT  10485.0 92982.5 10555.0 92640.0 ;
      RECT  10295.0 92277.5 10365.0 92142.5 ;
      RECT  10485.0 93117.5 10555.0 92982.5 ;
      RECT  10587.5 92675.0 10452.5 92605.0 ;
      RECT  9220.0 92585.0 9290.0 92720.0 ;
      RECT  9360.0 92857.5 9430.0 92992.5 ;
      RECT  10357.5 92820.0 10222.5 92890.0 ;
      RECT  10295.0 93885.0 10365.0 93955.0 ;
      RECT  10485.0 93885.0 10555.0 93955.0 ;
      RECT  10295.0 93920.0 10365.0 94282.5 ;
      RECT  10330.0 93885.0 10520.0 93955.0 ;
      RECT  10485.0 93577.5 10555.0 93920.0 ;
      RECT  10295.0 94282.5 10365.0 94417.5 ;
      RECT  10485.0 93442.5 10555.0 93577.5 ;
      RECT  10587.5 93885.0 10452.5 93955.0 ;
      RECT  9220.0 93840.0 9290.0 93975.0 ;
      RECT  9360.0 93567.5 9430.0 93702.5 ;
      RECT  10357.5 93670.0 10222.5 93740.0 ;
      RECT  10295.0 95365.0 10365.0 95295.0 ;
      RECT  10485.0 95365.0 10555.0 95295.0 ;
      RECT  10295.0 95330.0 10365.0 94967.5 ;
      RECT  10330.0 95365.0 10520.0 95295.0 ;
      RECT  10485.0 95672.5 10555.0 95330.0 ;
      RECT  10295.0 94967.5 10365.0 94832.5 ;
      RECT  10485.0 95807.5 10555.0 95672.5 ;
      RECT  10587.5 95365.0 10452.5 95295.0 ;
      RECT  9220.0 95275.0 9290.0 95410.0 ;
      RECT  9360.0 95547.5 9430.0 95682.5 ;
      RECT  10357.5 95510.0 10222.5 95580.0 ;
      RECT  10295.0 96575.0 10365.0 96645.0 ;
      RECT  10485.0 96575.0 10555.0 96645.0 ;
      RECT  10295.0 96610.0 10365.0 96972.5 ;
      RECT  10330.0 96575.0 10520.0 96645.0 ;
      RECT  10485.0 96267.5 10555.0 96610.0 ;
      RECT  10295.0 96972.5 10365.0 97107.5 ;
      RECT  10485.0 96132.5 10555.0 96267.5 ;
      RECT  10587.5 96575.0 10452.5 96645.0 ;
      RECT  9220.0 96530.0 9290.0 96665.0 ;
      RECT  9360.0 96257.5 9430.0 96392.5 ;
      RECT  10357.5 96360.0 10222.5 96430.0 ;
      RECT  10295.0 98055.0 10365.0 97985.0 ;
      RECT  10485.0 98055.0 10555.0 97985.0 ;
      RECT  10295.0 98020.0 10365.0 97657.5 ;
      RECT  10330.0 98055.0 10520.0 97985.0 ;
      RECT  10485.0 98362.5 10555.0 98020.0 ;
      RECT  10295.0 97657.5 10365.0 97522.5 ;
      RECT  10485.0 98497.5 10555.0 98362.5 ;
      RECT  10587.5 98055.0 10452.5 97985.0 ;
      RECT  9220.0 97965.0 9290.0 98100.0 ;
      RECT  9360.0 98237.5 9430.0 98372.5 ;
      RECT  10357.5 98200.0 10222.5 98270.0 ;
      RECT  10295.0 99265.0 10365.0 99335.0 ;
      RECT  10485.0 99265.0 10555.0 99335.0 ;
      RECT  10295.0 99300.0 10365.0 99662.5 ;
      RECT  10330.0 99265.0 10520.0 99335.0 ;
      RECT  10485.0 98957.5 10555.0 99300.0 ;
      RECT  10295.0 99662.5 10365.0 99797.5 ;
      RECT  10485.0 98822.5 10555.0 98957.5 ;
      RECT  10587.5 99265.0 10452.5 99335.0 ;
      RECT  9220.0 99220.0 9290.0 99355.0 ;
      RECT  9360.0 98947.5 9430.0 99082.5 ;
      RECT  10357.5 99050.0 10222.5 99120.0 ;
      RECT  10295.0 100745.0 10365.0 100675.0 ;
      RECT  10485.0 100745.0 10555.0 100675.0 ;
      RECT  10295.0 100710.0 10365.0 100347.5 ;
      RECT  10330.0 100745.0 10520.0 100675.0 ;
      RECT  10485.0 101052.5 10555.0 100710.0 ;
      RECT  10295.0 100347.5 10365.0 100212.5 ;
      RECT  10485.0 101187.5 10555.0 101052.5 ;
      RECT  10587.5 100745.0 10452.5 100675.0 ;
      RECT  9220.0 100655.0 9290.0 100790.0 ;
      RECT  9360.0 100927.5 9430.0 101062.5 ;
      RECT  10357.5 100890.0 10222.5 100960.0 ;
      RECT  10295.0 101955.0 10365.0 102025.0 ;
      RECT  10485.0 101955.0 10555.0 102025.0 ;
      RECT  10295.0 101990.0 10365.0 102352.5 ;
      RECT  10330.0 101955.0 10520.0 102025.0 ;
      RECT  10485.0 101647.5 10555.0 101990.0 ;
      RECT  10295.0 102352.5 10365.0 102487.5 ;
      RECT  10485.0 101512.5 10555.0 101647.5 ;
      RECT  10587.5 101955.0 10452.5 102025.0 ;
      RECT  9220.0 101910.0 9290.0 102045.0 ;
      RECT  9360.0 101637.5 9430.0 101772.5 ;
      RECT  10357.5 101740.0 10222.5 101810.0 ;
      RECT  10295.0 103435.0 10365.0 103365.0 ;
      RECT  10485.0 103435.0 10555.0 103365.0 ;
      RECT  10295.0 103400.0 10365.0 103037.5 ;
      RECT  10330.0 103435.0 10520.0 103365.0 ;
      RECT  10485.0 103742.5 10555.0 103400.0 ;
      RECT  10295.0 103037.5 10365.0 102902.5 ;
      RECT  10485.0 103877.5 10555.0 103742.5 ;
      RECT  10587.5 103435.0 10452.5 103365.0 ;
      RECT  9220.0 103345.0 9290.0 103480.0 ;
      RECT  9360.0 103617.5 9430.0 103752.5 ;
      RECT  10357.5 103580.0 10222.5 103650.0 ;
      RECT  10295.0 104645.0 10365.0 104715.0 ;
      RECT  10485.0 104645.0 10555.0 104715.0 ;
      RECT  10295.0 104680.0 10365.0 105042.5 ;
      RECT  10330.0 104645.0 10520.0 104715.0 ;
      RECT  10485.0 104337.5 10555.0 104680.0 ;
      RECT  10295.0 105042.5 10365.0 105177.5 ;
      RECT  10485.0 104202.5 10555.0 104337.5 ;
      RECT  10587.5 104645.0 10452.5 104715.0 ;
      RECT  9220.0 104600.0 9290.0 104735.0 ;
      RECT  9360.0 104327.5 9430.0 104462.5 ;
      RECT  10357.5 104430.0 10222.5 104500.0 ;
      RECT  10295.0 106125.0 10365.0 106055.0 ;
      RECT  10485.0 106125.0 10555.0 106055.0 ;
      RECT  10295.0 106090.0 10365.0 105727.5 ;
      RECT  10330.0 106125.0 10520.0 106055.0 ;
      RECT  10485.0 106432.5 10555.0 106090.0 ;
      RECT  10295.0 105727.5 10365.0 105592.5 ;
      RECT  10485.0 106567.5 10555.0 106432.5 ;
      RECT  10587.5 106125.0 10452.5 106055.0 ;
      RECT  9220.0 106035.0 9290.0 106170.0 ;
      RECT  9360.0 106307.5 9430.0 106442.5 ;
      RECT  10357.5 106270.0 10222.5 106340.0 ;
      RECT  10295.0 107335.0 10365.0 107405.0 ;
      RECT  10485.0 107335.0 10555.0 107405.0 ;
      RECT  10295.0 107370.0 10365.0 107732.5 ;
      RECT  10330.0 107335.0 10520.0 107405.0 ;
      RECT  10485.0 107027.5 10555.0 107370.0 ;
      RECT  10295.0 107732.5 10365.0 107867.5 ;
      RECT  10485.0 106892.5 10555.0 107027.5 ;
      RECT  10587.5 107335.0 10452.5 107405.0 ;
      RECT  9220.0 107290.0 9290.0 107425.0 ;
      RECT  9360.0 107017.5 9430.0 107152.5 ;
      RECT  10357.5 107120.0 10222.5 107190.0 ;
      RECT  10295.0 108815.0 10365.0 108745.0 ;
      RECT  10485.0 108815.0 10555.0 108745.0 ;
      RECT  10295.0 108780.0 10365.0 108417.5 ;
      RECT  10330.0 108815.0 10520.0 108745.0 ;
      RECT  10485.0 109122.5 10555.0 108780.0 ;
      RECT  10295.0 108417.5 10365.0 108282.5 ;
      RECT  10485.0 109257.5 10555.0 109122.5 ;
      RECT  10587.5 108815.0 10452.5 108745.0 ;
      RECT  9220.0 108725.0 9290.0 108860.0 ;
      RECT  9360.0 108997.5 9430.0 109132.5 ;
      RECT  10357.5 108960.0 10222.5 109030.0 ;
      RECT  10295.0 110025.0 10365.0 110095.0 ;
      RECT  10485.0 110025.0 10555.0 110095.0 ;
      RECT  10295.0 110060.0 10365.0 110422.5 ;
      RECT  10330.0 110025.0 10520.0 110095.0 ;
      RECT  10485.0 109717.5 10555.0 110060.0 ;
      RECT  10295.0 110422.5 10365.0 110557.5 ;
      RECT  10485.0 109582.5 10555.0 109717.5 ;
      RECT  10587.5 110025.0 10452.5 110095.0 ;
      RECT  9220.0 109980.0 9290.0 110115.0 ;
      RECT  9360.0 109707.5 9430.0 109842.5 ;
      RECT  10357.5 109810.0 10222.5 109880.0 ;
      RECT  10295.0 111505.0 10365.0 111435.0 ;
      RECT  10485.0 111505.0 10555.0 111435.0 ;
      RECT  10295.0 111470.0 10365.0 111107.5 ;
      RECT  10330.0 111505.0 10520.0 111435.0 ;
      RECT  10485.0 111812.5 10555.0 111470.0 ;
      RECT  10295.0 111107.5 10365.0 110972.5 ;
      RECT  10485.0 111947.5 10555.0 111812.5 ;
      RECT  10587.5 111505.0 10452.5 111435.0 ;
      RECT  9220.0 111415.0 9290.0 111550.0 ;
      RECT  9360.0 111687.5 9430.0 111822.5 ;
      RECT  10357.5 111650.0 10222.5 111720.0 ;
      RECT  10295.0 112715.0 10365.0 112785.0 ;
      RECT  10485.0 112715.0 10555.0 112785.0 ;
      RECT  10295.0 112750.0 10365.0 113112.5 ;
      RECT  10330.0 112715.0 10520.0 112785.0 ;
      RECT  10485.0 112407.5 10555.0 112750.0 ;
      RECT  10295.0 113112.5 10365.0 113247.5 ;
      RECT  10485.0 112272.5 10555.0 112407.5 ;
      RECT  10587.5 112715.0 10452.5 112785.0 ;
      RECT  9220.0 112670.0 9290.0 112805.0 ;
      RECT  9360.0 112397.5 9430.0 112532.5 ;
      RECT  10357.5 112500.0 10222.5 112570.0 ;
      RECT  10295.0 114195.0 10365.0 114125.0 ;
      RECT  10485.0 114195.0 10555.0 114125.0 ;
      RECT  10295.0 114160.0 10365.0 113797.5 ;
      RECT  10330.0 114195.0 10520.0 114125.0 ;
      RECT  10485.0 114502.5 10555.0 114160.0 ;
      RECT  10295.0 113797.5 10365.0 113662.5 ;
      RECT  10485.0 114637.5 10555.0 114502.5 ;
      RECT  10587.5 114195.0 10452.5 114125.0 ;
      RECT  9220.0 114105.0 9290.0 114240.0 ;
      RECT  9360.0 114377.5 9430.0 114512.5 ;
      RECT  10357.5 114340.0 10222.5 114410.0 ;
      RECT  10295.0 115405.0 10365.0 115475.0 ;
      RECT  10485.0 115405.0 10555.0 115475.0 ;
      RECT  10295.0 115440.0 10365.0 115802.5 ;
      RECT  10330.0 115405.0 10520.0 115475.0 ;
      RECT  10485.0 115097.5 10555.0 115440.0 ;
      RECT  10295.0 115802.5 10365.0 115937.5 ;
      RECT  10485.0 114962.5 10555.0 115097.5 ;
      RECT  10587.5 115405.0 10452.5 115475.0 ;
      RECT  9220.0 115360.0 9290.0 115495.0 ;
      RECT  9360.0 115087.5 9430.0 115222.5 ;
      RECT  10357.5 115190.0 10222.5 115260.0 ;
      RECT  10295.0 116885.0 10365.0 116815.0 ;
      RECT  10485.0 116885.0 10555.0 116815.0 ;
      RECT  10295.0 116850.0 10365.0 116487.5 ;
      RECT  10330.0 116885.0 10520.0 116815.0 ;
      RECT  10485.0 117192.5 10555.0 116850.0 ;
      RECT  10295.0 116487.5 10365.0 116352.5 ;
      RECT  10485.0 117327.5 10555.0 117192.5 ;
      RECT  10587.5 116885.0 10452.5 116815.0 ;
      RECT  9220.0 116795.0 9290.0 116930.0 ;
      RECT  9360.0 117067.5 9430.0 117202.5 ;
      RECT  10357.5 117030.0 10222.5 117100.0 ;
      RECT  10295.0 118095.0 10365.0 118165.0 ;
      RECT  10485.0 118095.0 10555.0 118165.0 ;
      RECT  10295.0 118130.0 10365.0 118492.5 ;
      RECT  10330.0 118095.0 10520.0 118165.0 ;
      RECT  10485.0 117787.5 10555.0 118130.0 ;
      RECT  10295.0 118492.5 10365.0 118627.5 ;
      RECT  10485.0 117652.5 10555.0 117787.5 ;
      RECT  10587.5 118095.0 10452.5 118165.0 ;
      RECT  9220.0 118050.0 9290.0 118185.0 ;
      RECT  9360.0 117777.5 9430.0 117912.5 ;
      RECT  10357.5 117880.0 10222.5 117950.0 ;
      RECT  10295.0 119575.0 10365.0 119505.0 ;
      RECT  10485.0 119575.0 10555.0 119505.0 ;
      RECT  10295.0 119540.0 10365.0 119177.5 ;
      RECT  10330.0 119575.0 10520.0 119505.0 ;
      RECT  10485.0 119882.5 10555.0 119540.0 ;
      RECT  10295.0 119177.5 10365.0 119042.5 ;
      RECT  10485.0 120017.5 10555.0 119882.5 ;
      RECT  10587.5 119575.0 10452.5 119505.0 ;
      RECT  9220.0 119485.0 9290.0 119620.0 ;
      RECT  9360.0 119757.5 9430.0 119892.5 ;
      RECT  10357.5 119720.0 10222.5 119790.0 ;
      RECT  10295.0 120785.0 10365.0 120855.0 ;
      RECT  10485.0 120785.0 10555.0 120855.0 ;
      RECT  10295.0 120820.0 10365.0 121182.5 ;
      RECT  10330.0 120785.0 10520.0 120855.0 ;
      RECT  10485.0 120477.5 10555.0 120820.0 ;
      RECT  10295.0 121182.5 10365.0 121317.5 ;
      RECT  10485.0 120342.5 10555.0 120477.5 ;
      RECT  10587.5 120785.0 10452.5 120855.0 ;
      RECT  9220.0 120740.0 9290.0 120875.0 ;
      RECT  9360.0 120467.5 9430.0 120602.5 ;
      RECT  10357.5 120570.0 10222.5 120640.0 ;
      RECT  10295.0 122265.0 10365.0 122195.0 ;
      RECT  10485.0 122265.0 10555.0 122195.0 ;
      RECT  10295.0 122230.0 10365.0 121867.5 ;
      RECT  10330.0 122265.0 10520.0 122195.0 ;
      RECT  10485.0 122572.5 10555.0 122230.0 ;
      RECT  10295.0 121867.5 10365.0 121732.5 ;
      RECT  10485.0 122707.5 10555.0 122572.5 ;
      RECT  10587.5 122265.0 10452.5 122195.0 ;
      RECT  9220.0 122175.0 9290.0 122310.0 ;
      RECT  9360.0 122447.5 9430.0 122582.5 ;
      RECT  10357.5 122410.0 10222.5 122480.0 ;
      RECT  10295.0 123475.0 10365.0 123545.0 ;
      RECT  10485.0 123475.0 10555.0 123545.0 ;
      RECT  10295.0 123510.0 10365.0 123872.5 ;
      RECT  10330.0 123475.0 10520.0 123545.0 ;
      RECT  10485.0 123167.5 10555.0 123510.0 ;
      RECT  10295.0 123872.5 10365.0 124007.5 ;
      RECT  10485.0 123032.5 10555.0 123167.5 ;
      RECT  10587.5 123475.0 10452.5 123545.0 ;
      RECT  9220.0 123430.0 9290.0 123565.0 ;
      RECT  9360.0 123157.5 9430.0 123292.5 ;
      RECT  10357.5 123260.0 10222.5 123330.0 ;
      RECT  10295.0 124955.0 10365.0 124885.0 ;
      RECT  10485.0 124955.0 10555.0 124885.0 ;
      RECT  10295.0 124920.0 10365.0 124557.5 ;
      RECT  10330.0 124955.0 10520.0 124885.0 ;
      RECT  10485.0 125262.5 10555.0 124920.0 ;
      RECT  10295.0 124557.5 10365.0 124422.5 ;
      RECT  10485.0 125397.5 10555.0 125262.5 ;
      RECT  10587.5 124955.0 10452.5 124885.0 ;
      RECT  9220.0 124865.0 9290.0 125000.0 ;
      RECT  9360.0 125137.5 9430.0 125272.5 ;
      RECT  10357.5 125100.0 10222.5 125170.0 ;
      RECT  10295.0 126165.0 10365.0 126235.0 ;
      RECT  10485.0 126165.0 10555.0 126235.0 ;
      RECT  10295.0 126200.0 10365.0 126562.5 ;
      RECT  10330.0 126165.0 10520.0 126235.0 ;
      RECT  10485.0 125857.5 10555.0 126200.0 ;
      RECT  10295.0 126562.5 10365.0 126697.5 ;
      RECT  10485.0 125722.5 10555.0 125857.5 ;
      RECT  10587.5 126165.0 10452.5 126235.0 ;
      RECT  9220.0 126120.0 9290.0 126255.0 ;
      RECT  9360.0 125847.5 9430.0 125982.5 ;
      RECT  10357.5 125950.0 10222.5 126020.0 ;
      RECT  10295.0 127645.0 10365.0 127575.0 ;
      RECT  10485.0 127645.0 10555.0 127575.0 ;
      RECT  10295.0 127610.0 10365.0 127247.5 ;
      RECT  10330.0 127645.0 10520.0 127575.0 ;
      RECT  10485.0 127952.5 10555.0 127610.0 ;
      RECT  10295.0 127247.5 10365.0 127112.5 ;
      RECT  10485.0 128087.5 10555.0 127952.5 ;
      RECT  10587.5 127645.0 10452.5 127575.0 ;
      RECT  9220.0 127555.0 9290.0 127690.0 ;
      RECT  9360.0 127827.5 9430.0 127962.5 ;
      RECT  10357.5 127790.0 10222.5 127860.0 ;
      RECT  10295.0 128855.0 10365.0 128925.0 ;
      RECT  10485.0 128855.0 10555.0 128925.0 ;
      RECT  10295.0 128890.0 10365.0 129252.5 ;
      RECT  10330.0 128855.0 10520.0 128925.0 ;
      RECT  10485.0 128547.5 10555.0 128890.0 ;
      RECT  10295.0 129252.5 10365.0 129387.5 ;
      RECT  10485.0 128412.5 10555.0 128547.5 ;
      RECT  10587.5 128855.0 10452.5 128925.0 ;
      RECT  9220.0 128810.0 9290.0 128945.0 ;
      RECT  9360.0 128537.5 9430.0 128672.5 ;
      RECT  10357.5 128640.0 10222.5 128710.0 ;
      RECT  10295.0 130335.0 10365.0 130265.0 ;
      RECT  10485.0 130335.0 10555.0 130265.0 ;
      RECT  10295.0 130300.0 10365.0 129937.5 ;
      RECT  10330.0 130335.0 10520.0 130265.0 ;
      RECT  10485.0 130642.5 10555.0 130300.0 ;
      RECT  10295.0 129937.5 10365.0 129802.5 ;
      RECT  10485.0 130777.5 10555.0 130642.5 ;
      RECT  10587.5 130335.0 10452.5 130265.0 ;
      RECT  9220.0 130245.0 9290.0 130380.0 ;
      RECT  9360.0 130517.5 9430.0 130652.5 ;
      RECT  10357.5 130480.0 10222.5 130550.0 ;
      RECT  10295.0 131545.0 10365.0 131615.0 ;
      RECT  10485.0 131545.0 10555.0 131615.0 ;
      RECT  10295.0 131580.0 10365.0 131942.5 ;
      RECT  10330.0 131545.0 10520.0 131615.0 ;
      RECT  10485.0 131237.5 10555.0 131580.0 ;
      RECT  10295.0 131942.5 10365.0 132077.5 ;
      RECT  10485.0 131102.5 10555.0 131237.5 ;
      RECT  10587.5 131545.0 10452.5 131615.0 ;
      RECT  9220.0 131500.0 9290.0 131635.0 ;
      RECT  9360.0 131227.5 9430.0 131362.5 ;
      RECT  10357.5 131330.0 10222.5 131400.0 ;
      RECT  10295.0 133025.0 10365.0 132955.0 ;
      RECT  10485.0 133025.0 10555.0 132955.0 ;
      RECT  10295.0 132990.0 10365.0 132627.5 ;
      RECT  10330.0 133025.0 10520.0 132955.0 ;
      RECT  10485.0 133332.5 10555.0 132990.0 ;
      RECT  10295.0 132627.5 10365.0 132492.5 ;
      RECT  10485.0 133467.5 10555.0 133332.5 ;
      RECT  10587.5 133025.0 10452.5 132955.0 ;
      RECT  9220.0 132935.0 9290.0 133070.0 ;
      RECT  9360.0 133207.5 9430.0 133342.5 ;
      RECT  10357.5 133170.0 10222.5 133240.0 ;
      RECT  10295.0 134235.0 10365.0 134305.0 ;
      RECT  10485.0 134235.0 10555.0 134305.0 ;
      RECT  10295.0 134270.0 10365.0 134632.5 ;
      RECT  10330.0 134235.0 10520.0 134305.0 ;
      RECT  10485.0 133927.5 10555.0 134270.0 ;
      RECT  10295.0 134632.5 10365.0 134767.5 ;
      RECT  10485.0 133792.5 10555.0 133927.5 ;
      RECT  10587.5 134235.0 10452.5 134305.0 ;
      RECT  9220.0 134190.0 9290.0 134325.0 ;
      RECT  9360.0 133917.5 9430.0 134052.5 ;
      RECT  10357.5 134020.0 10222.5 134090.0 ;
      RECT  10295.0 135715.0 10365.0 135645.0 ;
      RECT  10485.0 135715.0 10555.0 135645.0 ;
      RECT  10295.0 135680.0 10365.0 135317.5 ;
      RECT  10330.0 135715.0 10520.0 135645.0 ;
      RECT  10485.0 136022.5 10555.0 135680.0 ;
      RECT  10295.0 135317.5 10365.0 135182.5 ;
      RECT  10485.0 136157.5 10555.0 136022.5 ;
      RECT  10587.5 135715.0 10452.5 135645.0 ;
      RECT  9220.0 135625.0 9290.0 135760.0 ;
      RECT  9360.0 135897.5 9430.0 136032.5 ;
      RECT  10357.5 135860.0 10222.5 135930.0 ;
      RECT  10295.0 136925.0 10365.0 136995.0 ;
      RECT  10485.0 136925.0 10555.0 136995.0 ;
      RECT  10295.0 136960.0 10365.0 137322.5 ;
      RECT  10330.0 136925.0 10520.0 136995.0 ;
      RECT  10485.0 136617.5 10555.0 136960.0 ;
      RECT  10295.0 137322.5 10365.0 137457.5 ;
      RECT  10485.0 136482.5 10555.0 136617.5 ;
      RECT  10587.5 136925.0 10452.5 136995.0 ;
      RECT  9220.0 136880.0 9290.0 137015.0 ;
      RECT  9360.0 136607.5 9430.0 136742.5 ;
      RECT  10357.5 136710.0 10222.5 136780.0 ;
      RECT  10295.0 138405.0 10365.0 138335.0 ;
      RECT  10485.0 138405.0 10555.0 138335.0 ;
      RECT  10295.0 138370.0 10365.0 138007.5 ;
      RECT  10330.0 138405.0 10520.0 138335.0 ;
      RECT  10485.0 138712.5 10555.0 138370.0 ;
      RECT  10295.0 138007.5 10365.0 137872.5 ;
      RECT  10485.0 138847.5 10555.0 138712.5 ;
      RECT  10587.5 138405.0 10452.5 138335.0 ;
      RECT  9220.0 138315.0 9290.0 138450.0 ;
      RECT  9360.0 138587.5 9430.0 138722.5 ;
      RECT  10357.5 138550.0 10222.5 138620.0 ;
      RECT  10295.0 139615.0 10365.0 139685.0 ;
      RECT  10485.0 139615.0 10555.0 139685.0 ;
      RECT  10295.0 139650.0 10365.0 140012.5 ;
      RECT  10330.0 139615.0 10520.0 139685.0 ;
      RECT  10485.0 139307.5 10555.0 139650.0 ;
      RECT  10295.0 140012.5 10365.0 140147.5 ;
      RECT  10485.0 139172.5 10555.0 139307.5 ;
      RECT  10587.5 139615.0 10452.5 139685.0 ;
      RECT  9220.0 139570.0 9290.0 139705.0 ;
      RECT  9360.0 139297.5 9430.0 139432.5 ;
      RECT  10357.5 139400.0 10222.5 139470.0 ;
      RECT  10295.0 141095.0 10365.0 141025.0 ;
      RECT  10485.0 141095.0 10555.0 141025.0 ;
      RECT  10295.0 141060.0 10365.0 140697.5 ;
      RECT  10330.0 141095.0 10520.0 141025.0 ;
      RECT  10485.0 141402.5 10555.0 141060.0 ;
      RECT  10295.0 140697.5 10365.0 140562.5 ;
      RECT  10485.0 141537.5 10555.0 141402.5 ;
      RECT  10587.5 141095.0 10452.5 141025.0 ;
      RECT  9220.0 141005.0 9290.0 141140.0 ;
      RECT  9360.0 141277.5 9430.0 141412.5 ;
      RECT  10357.5 141240.0 10222.5 141310.0 ;
      RECT  10295.0 142305.0 10365.0 142375.0 ;
      RECT  10485.0 142305.0 10555.0 142375.0 ;
      RECT  10295.0 142340.0 10365.0 142702.5 ;
      RECT  10330.0 142305.0 10520.0 142375.0 ;
      RECT  10485.0 141997.5 10555.0 142340.0 ;
      RECT  10295.0 142702.5 10365.0 142837.5 ;
      RECT  10485.0 141862.5 10555.0 141997.5 ;
      RECT  10587.5 142305.0 10452.5 142375.0 ;
      RECT  9220.0 142260.0 9290.0 142395.0 ;
      RECT  9360.0 141987.5 9430.0 142122.5 ;
      RECT  10357.5 142090.0 10222.5 142160.0 ;
      RECT  10295.0 143785.0 10365.0 143715.0 ;
      RECT  10485.0 143785.0 10555.0 143715.0 ;
      RECT  10295.0 143750.0 10365.0 143387.5 ;
      RECT  10330.0 143785.0 10520.0 143715.0 ;
      RECT  10485.0 144092.5 10555.0 143750.0 ;
      RECT  10295.0 143387.5 10365.0 143252.5 ;
      RECT  10485.0 144227.5 10555.0 144092.5 ;
      RECT  10587.5 143785.0 10452.5 143715.0 ;
      RECT  9220.0 143695.0 9290.0 143830.0 ;
      RECT  9360.0 143967.5 9430.0 144102.5 ;
      RECT  10357.5 143930.0 10222.5 144000.0 ;
      RECT  10295.0 144995.0 10365.0 145065.0 ;
      RECT  10485.0 144995.0 10555.0 145065.0 ;
      RECT  10295.0 145030.0 10365.0 145392.5 ;
      RECT  10330.0 144995.0 10520.0 145065.0 ;
      RECT  10485.0 144687.5 10555.0 145030.0 ;
      RECT  10295.0 145392.5 10365.0 145527.5 ;
      RECT  10485.0 144552.5 10555.0 144687.5 ;
      RECT  10587.5 144995.0 10452.5 145065.0 ;
      RECT  9220.0 144950.0 9290.0 145085.0 ;
      RECT  9360.0 144677.5 9430.0 144812.5 ;
      RECT  10357.5 144780.0 10222.5 144850.0 ;
      RECT  10295.0 146475.0 10365.0 146405.0 ;
      RECT  10485.0 146475.0 10555.0 146405.0 ;
      RECT  10295.0 146440.0 10365.0 146077.5 ;
      RECT  10330.0 146475.0 10520.0 146405.0 ;
      RECT  10485.0 146782.5 10555.0 146440.0 ;
      RECT  10295.0 146077.5 10365.0 145942.5 ;
      RECT  10485.0 146917.5 10555.0 146782.5 ;
      RECT  10587.5 146475.0 10452.5 146405.0 ;
      RECT  9220.0 146385.0 9290.0 146520.0 ;
      RECT  9360.0 146657.5 9430.0 146792.5 ;
      RECT  10357.5 146620.0 10222.5 146690.0 ;
      RECT  10295.0 147685.0 10365.0 147755.0 ;
      RECT  10485.0 147685.0 10555.0 147755.0 ;
      RECT  10295.0 147720.0 10365.0 148082.5 ;
      RECT  10330.0 147685.0 10520.0 147755.0 ;
      RECT  10485.0 147377.5 10555.0 147720.0 ;
      RECT  10295.0 148082.5 10365.0 148217.5 ;
      RECT  10485.0 147242.5 10555.0 147377.5 ;
      RECT  10587.5 147685.0 10452.5 147755.0 ;
      RECT  9220.0 147640.0 9290.0 147775.0 ;
      RECT  9360.0 147367.5 9430.0 147502.5 ;
      RECT  10357.5 147470.0 10222.5 147540.0 ;
      RECT  10295.0 149165.0 10365.0 149095.0 ;
      RECT  10485.0 149165.0 10555.0 149095.0 ;
      RECT  10295.0 149130.0 10365.0 148767.5 ;
      RECT  10330.0 149165.0 10520.0 149095.0 ;
      RECT  10485.0 149472.5 10555.0 149130.0 ;
      RECT  10295.0 148767.5 10365.0 148632.5 ;
      RECT  10485.0 149607.5 10555.0 149472.5 ;
      RECT  10587.5 149165.0 10452.5 149095.0 ;
      RECT  9220.0 149075.0 9290.0 149210.0 ;
      RECT  9360.0 149347.5 9430.0 149482.5 ;
      RECT  10357.5 149310.0 10222.5 149380.0 ;
      RECT  10295.0 150375.0 10365.0 150445.0 ;
      RECT  10485.0 150375.0 10555.0 150445.0 ;
      RECT  10295.0 150410.0 10365.0 150772.5 ;
      RECT  10330.0 150375.0 10520.0 150445.0 ;
      RECT  10485.0 150067.5 10555.0 150410.0 ;
      RECT  10295.0 150772.5 10365.0 150907.5 ;
      RECT  10485.0 149932.5 10555.0 150067.5 ;
      RECT  10587.5 150375.0 10452.5 150445.0 ;
      RECT  9220.0 150330.0 9290.0 150465.0 ;
      RECT  9360.0 150057.5 9430.0 150192.5 ;
      RECT  10357.5 150160.0 10222.5 150230.0 ;
      RECT  10295.0 151855.0 10365.0 151785.0 ;
      RECT  10485.0 151855.0 10555.0 151785.0 ;
      RECT  10295.0 151820.0 10365.0 151457.5 ;
      RECT  10330.0 151855.0 10520.0 151785.0 ;
      RECT  10485.0 152162.5 10555.0 151820.0 ;
      RECT  10295.0 151457.5 10365.0 151322.5 ;
      RECT  10485.0 152297.5 10555.0 152162.5 ;
      RECT  10587.5 151855.0 10452.5 151785.0 ;
      RECT  9220.0 151765.0 9290.0 151900.0 ;
      RECT  9360.0 152037.5 9430.0 152172.5 ;
      RECT  10357.5 152000.0 10222.5 152070.0 ;
      RECT  10295.0 153065.0 10365.0 153135.0 ;
      RECT  10485.0 153065.0 10555.0 153135.0 ;
      RECT  10295.0 153100.0 10365.0 153462.5 ;
      RECT  10330.0 153065.0 10520.0 153135.0 ;
      RECT  10485.0 152757.5 10555.0 153100.0 ;
      RECT  10295.0 153462.5 10365.0 153597.5 ;
      RECT  10485.0 152622.5 10555.0 152757.5 ;
      RECT  10587.5 153065.0 10452.5 153135.0 ;
      RECT  9220.0 153020.0 9290.0 153155.0 ;
      RECT  9360.0 152747.5 9430.0 152882.5 ;
      RECT  10357.5 152850.0 10222.5 152920.0 ;
      RECT  10295.0 154545.0 10365.0 154475.0 ;
      RECT  10485.0 154545.0 10555.0 154475.0 ;
      RECT  10295.0 154510.0 10365.0 154147.5 ;
      RECT  10330.0 154545.0 10520.0 154475.0 ;
      RECT  10485.0 154852.5 10555.0 154510.0 ;
      RECT  10295.0 154147.5 10365.0 154012.5 ;
      RECT  10485.0 154987.5 10555.0 154852.5 ;
      RECT  10587.5 154545.0 10452.5 154475.0 ;
      RECT  9220.0 154455.0 9290.0 154590.0 ;
      RECT  9360.0 154727.5 9430.0 154862.5 ;
      RECT  10357.5 154690.0 10222.5 154760.0 ;
      RECT  10295.0 155755.0 10365.0 155825.0 ;
      RECT  10485.0 155755.0 10555.0 155825.0 ;
      RECT  10295.0 155790.0 10365.0 156152.5 ;
      RECT  10330.0 155755.0 10520.0 155825.0 ;
      RECT  10485.0 155447.5 10555.0 155790.0 ;
      RECT  10295.0 156152.5 10365.0 156287.5 ;
      RECT  10485.0 155312.5 10555.0 155447.5 ;
      RECT  10587.5 155755.0 10452.5 155825.0 ;
      RECT  9220.0 155710.0 9290.0 155845.0 ;
      RECT  9360.0 155437.5 9430.0 155572.5 ;
      RECT  10357.5 155540.0 10222.5 155610.0 ;
      RECT  10295.0 157235.0 10365.0 157165.0 ;
      RECT  10485.0 157235.0 10555.0 157165.0 ;
      RECT  10295.0 157200.0 10365.0 156837.5 ;
      RECT  10330.0 157235.0 10520.0 157165.0 ;
      RECT  10485.0 157542.5 10555.0 157200.0 ;
      RECT  10295.0 156837.5 10365.0 156702.5 ;
      RECT  10485.0 157677.5 10555.0 157542.5 ;
      RECT  10587.5 157235.0 10452.5 157165.0 ;
      RECT  9220.0 157145.0 9290.0 157280.0 ;
      RECT  9360.0 157417.5 9430.0 157552.5 ;
      RECT  10357.5 157380.0 10222.5 157450.0 ;
      RECT  10295.0 158445.0 10365.0 158515.0 ;
      RECT  10485.0 158445.0 10555.0 158515.0 ;
      RECT  10295.0 158480.0 10365.0 158842.5 ;
      RECT  10330.0 158445.0 10520.0 158515.0 ;
      RECT  10485.0 158137.5 10555.0 158480.0 ;
      RECT  10295.0 158842.5 10365.0 158977.5 ;
      RECT  10485.0 158002.5 10555.0 158137.5 ;
      RECT  10587.5 158445.0 10452.5 158515.0 ;
      RECT  9220.0 158400.0 9290.0 158535.0 ;
      RECT  9360.0 158127.5 9430.0 158262.5 ;
      RECT  10357.5 158230.0 10222.5 158300.0 ;
      RECT  10295.0 159925.0 10365.0 159855.0 ;
      RECT  10485.0 159925.0 10555.0 159855.0 ;
      RECT  10295.0 159890.0 10365.0 159527.5 ;
      RECT  10330.0 159925.0 10520.0 159855.0 ;
      RECT  10485.0 160232.5 10555.0 159890.0 ;
      RECT  10295.0 159527.5 10365.0 159392.5 ;
      RECT  10485.0 160367.5 10555.0 160232.5 ;
      RECT  10587.5 159925.0 10452.5 159855.0 ;
      RECT  9220.0 159835.0 9290.0 159970.0 ;
      RECT  9360.0 160107.5 9430.0 160242.5 ;
      RECT  10357.5 160070.0 10222.5 160140.0 ;
      RECT  10295.0 161135.0 10365.0 161205.0 ;
      RECT  10485.0 161135.0 10555.0 161205.0 ;
      RECT  10295.0 161170.0 10365.0 161532.5 ;
      RECT  10330.0 161135.0 10520.0 161205.0 ;
      RECT  10485.0 160827.5 10555.0 161170.0 ;
      RECT  10295.0 161532.5 10365.0 161667.5 ;
      RECT  10485.0 160692.5 10555.0 160827.5 ;
      RECT  10587.5 161135.0 10452.5 161205.0 ;
      RECT  9220.0 161090.0 9290.0 161225.0 ;
      RECT  9360.0 160817.5 9430.0 160952.5 ;
      RECT  10357.5 160920.0 10222.5 160990.0 ;
      RECT  10295.0 162615.0 10365.0 162545.0 ;
      RECT  10485.0 162615.0 10555.0 162545.0 ;
      RECT  10295.0 162580.0 10365.0 162217.5 ;
      RECT  10330.0 162615.0 10520.0 162545.0 ;
      RECT  10485.0 162922.5 10555.0 162580.0 ;
      RECT  10295.0 162217.5 10365.0 162082.5 ;
      RECT  10485.0 163057.5 10555.0 162922.5 ;
      RECT  10587.5 162615.0 10452.5 162545.0 ;
      RECT  9220.0 162525.0 9290.0 162660.0 ;
      RECT  9360.0 162797.5 9430.0 162932.5 ;
      RECT  10357.5 162760.0 10222.5 162830.0 ;
      RECT  10295.0 163825.0 10365.0 163895.0 ;
      RECT  10485.0 163825.0 10555.0 163895.0 ;
      RECT  10295.0 163860.0 10365.0 164222.5 ;
      RECT  10330.0 163825.0 10520.0 163895.0 ;
      RECT  10485.0 163517.5 10555.0 163860.0 ;
      RECT  10295.0 164222.5 10365.0 164357.5 ;
      RECT  10485.0 163382.5 10555.0 163517.5 ;
      RECT  10587.5 163825.0 10452.5 163895.0 ;
      RECT  9220.0 163780.0 9290.0 163915.0 ;
      RECT  9360.0 163507.5 9430.0 163642.5 ;
      RECT  10357.5 163610.0 10222.5 163680.0 ;
      RECT  10295.0 165305.0 10365.0 165235.0 ;
      RECT  10485.0 165305.0 10555.0 165235.0 ;
      RECT  10295.0 165270.0 10365.0 164907.5 ;
      RECT  10330.0 165305.0 10520.0 165235.0 ;
      RECT  10485.0 165612.5 10555.0 165270.0 ;
      RECT  10295.0 164907.5 10365.0 164772.5 ;
      RECT  10485.0 165747.5 10555.0 165612.5 ;
      RECT  10587.5 165305.0 10452.5 165235.0 ;
      RECT  9220.0 165215.0 9290.0 165350.0 ;
      RECT  9360.0 165487.5 9430.0 165622.5 ;
      RECT  10357.5 165450.0 10222.5 165520.0 ;
      RECT  10295.0 166515.0 10365.0 166585.0 ;
      RECT  10485.0 166515.0 10555.0 166585.0 ;
      RECT  10295.0 166550.0 10365.0 166912.5 ;
      RECT  10330.0 166515.0 10520.0 166585.0 ;
      RECT  10485.0 166207.5 10555.0 166550.0 ;
      RECT  10295.0 166912.5 10365.0 167047.5 ;
      RECT  10485.0 166072.5 10555.0 166207.5 ;
      RECT  10587.5 166515.0 10452.5 166585.0 ;
      RECT  9220.0 166470.0 9290.0 166605.0 ;
      RECT  9360.0 166197.5 9430.0 166332.5 ;
      RECT  10357.5 166300.0 10222.5 166370.0 ;
      RECT  10295.0 167995.0 10365.0 167925.0 ;
      RECT  10485.0 167995.0 10555.0 167925.0 ;
      RECT  10295.0 167960.0 10365.0 167597.5 ;
      RECT  10330.0 167995.0 10520.0 167925.0 ;
      RECT  10485.0 168302.5 10555.0 167960.0 ;
      RECT  10295.0 167597.5 10365.0 167462.5 ;
      RECT  10485.0 168437.5 10555.0 168302.5 ;
      RECT  10587.5 167995.0 10452.5 167925.0 ;
      RECT  9220.0 167905.0 9290.0 168040.0 ;
      RECT  9360.0 168177.5 9430.0 168312.5 ;
      RECT  10357.5 168140.0 10222.5 168210.0 ;
      RECT  10295.0 169205.0 10365.0 169275.0 ;
      RECT  10485.0 169205.0 10555.0 169275.0 ;
      RECT  10295.0 169240.0 10365.0 169602.5 ;
      RECT  10330.0 169205.0 10520.0 169275.0 ;
      RECT  10485.0 168897.5 10555.0 169240.0 ;
      RECT  10295.0 169602.5 10365.0 169737.5 ;
      RECT  10485.0 168762.5 10555.0 168897.5 ;
      RECT  10587.5 169205.0 10452.5 169275.0 ;
      RECT  9220.0 169160.0 9290.0 169295.0 ;
      RECT  9360.0 168887.5 9430.0 169022.5 ;
      RECT  10357.5 168990.0 10222.5 169060.0 ;
      RECT  10295.0 170685.0 10365.0 170615.0 ;
      RECT  10485.0 170685.0 10555.0 170615.0 ;
      RECT  10295.0 170650.0 10365.0 170287.5 ;
      RECT  10330.0 170685.0 10520.0 170615.0 ;
      RECT  10485.0 170992.5 10555.0 170650.0 ;
      RECT  10295.0 170287.5 10365.0 170152.5 ;
      RECT  10485.0 171127.5 10555.0 170992.5 ;
      RECT  10587.5 170685.0 10452.5 170615.0 ;
      RECT  9220.0 170595.0 9290.0 170730.0 ;
      RECT  9360.0 170867.5 9430.0 171002.5 ;
      RECT  10357.5 170830.0 10222.5 170900.0 ;
      RECT  10295.0 171895.0 10365.0 171965.0 ;
      RECT  10485.0 171895.0 10555.0 171965.0 ;
      RECT  10295.0 171930.0 10365.0 172292.5 ;
      RECT  10330.0 171895.0 10520.0 171965.0 ;
      RECT  10485.0 171587.5 10555.0 171930.0 ;
      RECT  10295.0 172292.5 10365.0 172427.5 ;
      RECT  10485.0 171452.5 10555.0 171587.5 ;
      RECT  10587.5 171895.0 10452.5 171965.0 ;
      RECT  9220.0 171850.0 9290.0 171985.0 ;
      RECT  9360.0 171577.5 9430.0 171712.5 ;
      RECT  10357.5 171680.0 10222.5 171750.0 ;
      RECT  10295.0 173375.0 10365.0 173305.0 ;
      RECT  10485.0 173375.0 10555.0 173305.0 ;
      RECT  10295.0 173340.0 10365.0 172977.5 ;
      RECT  10330.0 173375.0 10520.0 173305.0 ;
      RECT  10485.0 173682.5 10555.0 173340.0 ;
      RECT  10295.0 172977.5 10365.0 172842.5 ;
      RECT  10485.0 173817.5 10555.0 173682.5 ;
      RECT  10587.5 173375.0 10452.5 173305.0 ;
      RECT  9220.0 173285.0 9290.0 173420.0 ;
      RECT  9360.0 173557.5 9430.0 173692.5 ;
      RECT  10357.5 173520.0 10222.5 173590.0 ;
      RECT  10295.0 174585.0 10365.0 174655.0 ;
      RECT  10485.0 174585.0 10555.0 174655.0 ;
      RECT  10295.0 174620.0 10365.0 174982.5 ;
      RECT  10330.0 174585.0 10520.0 174655.0 ;
      RECT  10485.0 174277.5 10555.0 174620.0 ;
      RECT  10295.0 174982.5 10365.0 175117.5 ;
      RECT  10485.0 174142.5 10555.0 174277.5 ;
      RECT  10587.5 174585.0 10452.5 174655.0 ;
      RECT  9220.0 174540.0 9290.0 174675.0 ;
      RECT  9360.0 174267.5 9430.0 174402.5 ;
      RECT  10357.5 174370.0 10222.5 174440.0 ;
      RECT  10295.0 176065.0 10365.0 175995.0 ;
      RECT  10485.0 176065.0 10555.0 175995.0 ;
      RECT  10295.0 176030.0 10365.0 175667.5 ;
      RECT  10330.0 176065.0 10520.0 175995.0 ;
      RECT  10485.0 176372.5 10555.0 176030.0 ;
      RECT  10295.0 175667.5 10365.0 175532.5 ;
      RECT  10485.0 176507.5 10555.0 176372.5 ;
      RECT  10587.5 176065.0 10452.5 175995.0 ;
      RECT  9220.0 175975.0 9290.0 176110.0 ;
      RECT  9360.0 176247.5 9430.0 176382.5 ;
      RECT  10357.5 176210.0 10222.5 176280.0 ;
      RECT  10295.0 177275.0 10365.0 177345.0 ;
      RECT  10485.0 177275.0 10555.0 177345.0 ;
      RECT  10295.0 177310.0 10365.0 177672.5 ;
      RECT  10330.0 177275.0 10520.0 177345.0 ;
      RECT  10485.0 176967.5 10555.0 177310.0 ;
      RECT  10295.0 177672.5 10365.0 177807.5 ;
      RECT  10485.0 176832.5 10555.0 176967.5 ;
      RECT  10587.5 177275.0 10452.5 177345.0 ;
      RECT  9220.0 177230.0 9290.0 177365.0 ;
      RECT  9360.0 176957.5 9430.0 177092.5 ;
      RECT  10357.5 177060.0 10222.5 177130.0 ;
      RECT  10295.0 178755.0 10365.0 178685.0 ;
      RECT  10485.0 178755.0 10555.0 178685.0 ;
      RECT  10295.0 178720.0 10365.0 178357.5 ;
      RECT  10330.0 178755.0 10520.0 178685.0 ;
      RECT  10485.0 179062.5 10555.0 178720.0 ;
      RECT  10295.0 178357.5 10365.0 178222.5 ;
      RECT  10485.0 179197.5 10555.0 179062.5 ;
      RECT  10587.5 178755.0 10452.5 178685.0 ;
      RECT  9220.0 178665.0 9290.0 178800.0 ;
      RECT  9360.0 178937.5 9430.0 179072.5 ;
      RECT  10357.5 178900.0 10222.5 178970.0 ;
      RECT  10295.0 179965.0 10365.0 180035.0 ;
      RECT  10485.0 179965.0 10555.0 180035.0 ;
      RECT  10295.0 180000.0 10365.0 180362.5 ;
      RECT  10330.0 179965.0 10520.0 180035.0 ;
      RECT  10485.0 179657.5 10555.0 180000.0 ;
      RECT  10295.0 180362.5 10365.0 180497.5 ;
      RECT  10485.0 179522.5 10555.0 179657.5 ;
      RECT  10587.5 179965.0 10452.5 180035.0 ;
      RECT  9220.0 179920.0 9290.0 180055.0 ;
      RECT  9360.0 179647.5 9430.0 179782.5 ;
      RECT  10357.5 179750.0 10222.5 179820.0 ;
      RECT  10295.0 181445.0 10365.0 181375.0 ;
      RECT  10485.0 181445.0 10555.0 181375.0 ;
      RECT  10295.0 181410.0 10365.0 181047.5 ;
      RECT  10330.0 181445.0 10520.0 181375.0 ;
      RECT  10485.0 181752.5 10555.0 181410.0 ;
      RECT  10295.0 181047.5 10365.0 180912.5 ;
      RECT  10485.0 181887.5 10555.0 181752.5 ;
      RECT  10587.5 181445.0 10452.5 181375.0 ;
      RECT  9220.0 181355.0 9290.0 181490.0 ;
      RECT  9360.0 181627.5 9430.0 181762.5 ;
      RECT  10357.5 181590.0 10222.5 181660.0 ;
      RECT  10295.0 182655.0 10365.0 182725.0 ;
      RECT  10485.0 182655.0 10555.0 182725.0 ;
      RECT  10295.0 182690.0 10365.0 183052.5 ;
      RECT  10330.0 182655.0 10520.0 182725.0 ;
      RECT  10485.0 182347.5 10555.0 182690.0 ;
      RECT  10295.0 183052.5 10365.0 183187.5 ;
      RECT  10485.0 182212.5 10555.0 182347.5 ;
      RECT  10587.5 182655.0 10452.5 182725.0 ;
      RECT  9220.0 182610.0 9290.0 182745.0 ;
      RECT  9360.0 182337.5 9430.0 182472.5 ;
      RECT  10357.5 182440.0 10222.5 182510.0 ;
      RECT  10295.0 184135.0 10365.0 184065.0 ;
      RECT  10485.0 184135.0 10555.0 184065.0 ;
      RECT  10295.0 184100.0 10365.0 183737.5 ;
      RECT  10330.0 184135.0 10520.0 184065.0 ;
      RECT  10485.0 184442.5 10555.0 184100.0 ;
      RECT  10295.0 183737.5 10365.0 183602.5 ;
      RECT  10485.0 184577.5 10555.0 184442.5 ;
      RECT  10587.5 184135.0 10452.5 184065.0 ;
      RECT  9220.0 184045.0 9290.0 184180.0 ;
      RECT  9360.0 184317.5 9430.0 184452.5 ;
      RECT  10357.5 184280.0 10222.5 184350.0 ;
      RECT  10295.0 185345.0 10365.0 185415.0 ;
      RECT  10485.0 185345.0 10555.0 185415.0 ;
      RECT  10295.0 185380.0 10365.0 185742.5 ;
      RECT  10330.0 185345.0 10520.0 185415.0 ;
      RECT  10485.0 185037.5 10555.0 185380.0 ;
      RECT  10295.0 185742.5 10365.0 185877.5 ;
      RECT  10485.0 184902.5 10555.0 185037.5 ;
      RECT  10587.5 185345.0 10452.5 185415.0 ;
      RECT  9220.0 185300.0 9290.0 185435.0 ;
      RECT  9360.0 185027.5 9430.0 185162.5 ;
      RECT  10357.5 185130.0 10222.5 185200.0 ;
      RECT  10295.0 186825.0 10365.0 186755.0 ;
      RECT  10485.0 186825.0 10555.0 186755.0 ;
      RECT  10295.0 186790.0 10365.0 186427.5 ;
      RECT  10330.0 186825.0 10520.0 186755.0 ;
      RECT  10485.0 187132.5 10555.0 186790.0 ;
      RECT  10295.0 186427.5 10365.0 186292.5 ;
      RECT  10485.0 187267.5 10555.0 187132.5 ;
      RECT  10587.5 186825.0 10452.5 186755.0 ;
      RECT  9220.0 186735.0 9290.0 186870.0 ;
      RECT  9360.0 187007.5 9430.0 187142.5 ;
      RECT  10357.5 186970.0 10222.5 187040.0 ;
      RECT  10295.0 188035.0 10365.0 188105.0 ;
      RECT  10485.0 188035.0 10555.0 188105.0 ;
      RECT  10295.0 188070.0 10365.0 188432.5 ;
      RECT  10330.0 188035.0 10520.0 188105.0 ;
      RECT  10485.0 187727.5 10555.0 188070.0 ;
      RECT  10295.0 188432.5 10365.0 188567.5 ;
      RECT  10485.0 187592.5 10555.0 187727.5 ;
      RECT  10587.5 188035.0 10452.5 188105.0 ;
      RECT  9220.0 187990.0 9290.0 188125.0 ;
      RECT  9360.0 187717.5 9430.0 187852.5 ;
      RECT  10357.5 187820.0 10222.5 187890.0 ;
      RECT  10295.0 189515.0 10365.0 189445.0 ;
      RECT  10485.0 189515.0 10555.0 189445.0 ;
      RECT  10295.0 189480.0 10365.0 189117.5 ;
      RECT  10330.0 189515.0 10520.0 189445.0 ;
      RECT  10485.0 189822.5 10555.0 189480.0 ;
      RECT  10295.0 189117.5 10365.0 188982.5 ;
      RECT  10485.0 189957.5 10555.0 189822.5 ;
      RECT  10587.5 189515.0 10452.5 189445.0 ;
      RECT  9220.0 189425.0 9290.0 189560.0 ;
      RECT  9360.0 189697.5 9430.0 189832.5 ;
      RECT  10357.5 189660.0 10222.5 189730.0 ;
      RECT  10295.0 190725.0 10365.0 190795.0 ;
      RECT  10485.0 190725.0 10555.0 190795.0 ;
      RECT  10295.0 190760.0 10365.0 191122.5 ;
      RECT  10330.0 190725.0 10520.0 190795.0 ;
      RECT  10485.0 190417.5 10555.0 190760.0 ;
      RECT  10295.0 191122.5 10365.0 191257.5 ;
      RECT  10485.0 190282.5 10555.0 190417.5 ;
      RECT  10587.5 190725.0 10452.5 190795.0 ;
      RECT  9220.0 190680.0 9290.0 190815.0 ;
      RECT  9360.0 190407.5 9430.0 190542.5 ;
      RECT  10357.5 190510.0 10222.5 190580.0 ;
      RECT  10295.0 192205.0 10365.0 192135.0 ;
      RECT  10485.0 192205.0 10555.0 192135.0 ;
      RECT  10295.0 192170.0 10365.0 191807.5 ;
      RECT  10330.0 192205.0 10520.0 192135.0 ;
      RECT  10485.0 192512.5 10555.0 192170.0 ;
      RECT  10295.0 191807.5 10365.0 191672.5 ;
      RECT  10485.0 192647.5 10555.0 192512.5 ;
      RECT  10587.5 192205.0 10452.5 192135.0 ;
      RECT  9220.0 192115.0 9290.0 192250.0 ;
      RECT  9360.0 192387.5 9430.0 192522.5 ;
      RECT  10357.5 192350.0 10222.5 192420.0 ;
      RECT  10295.0 193415.0 10365.0 193485.0 ;
      RECT  10485.0 193415.0 10555.0 193485.0 ;
      RECT  10295.0 193450.0 10365.0 193812.5 ;
      RECT  10330.0 193415.0 10520.0 193485.0 ;
      RECT  10485.0 193107.5 10555.0 193450.0 ;
      RECT  10295.0 193812.5 10365.0 193947.5 ;
      RECT  10485.0 192972.5 10555.0 193107.5 ;
      RECT  10587.5 193415.0 10452.5 193485.0 ;
      RECT  9220.0 193370.0 9290.0 193505.0 ;
      RECT  9360.0 193097.5 9430.0 193232.5 ;
      RECT  10357.5 193200.0 10222.5 193270.0 ;
      RECT  10295.0 194895.0 10365.0 194825.0 ;
      RECT  10485.0 194895.0 10555.0 194825.0 ;
      RECT  10295.0 194860.0 10365.0 194497.5 ;
      RECT  10330.0 194895.0 10520.0 194825.0 ;
      RECT  10485.0 195202.5 10555.0 194860.0 ;
      RECT  10295.0 194497.5 10365.0 194362.5 ;
      RECT  10485.0 195337.5 10555.0 195202.5 ;
      RECT  10587.5 194895.0 10452.5 194825.0 ;
      RECT  9220.0 194805.0 9290.0 194940.0 ;
      RECT  9360.0 195077.5 9430.0 195212.5 ;
      RECT  10357.5 195040.0 10222.5 195110.0 ;
      RECT  10295.0 196105.0 10365.0 196175.0 ;
      RECT  10485.0 196105.0 10555.0 196175.0 ;
      RECT  10295.0 196140.0 10365.0 196502.5 ;
      RECT  10330.0 196105.0 10520.0 196175.0 ;
      RECT  10485.0 195797.5 10555.0 196140.0 ;
      RECT  10295.0 196502.5 10365.0 196637.5 ;
      RECT  10485.0 195662.5 10555.0 195797.5 ;
      RECT  10587.5 196105.0 10452.5 196175.0 ;
      RECT  9220.0 196060.0 9290.0 196195.0 ;
      RECT  9360.0 195787.5 9430.0 195922.5 ;
      RECT  10357.5 195890.0 10222.5 195960.0 ;
      RECT  10295.0 197585.0 10365.0 197515.0 ;
      RECT  10485.0 197585.0 10555.0 197515.0 ;
      RECT  10295.0 197550.0 10365.0 197187.5 ;
      RECT  10330.0 197585.0 10520.0 197515.0 ;
      RECT  10485.0 197892.5 10555.0 197550.0 ;
      RECT  10295.0 197187.5 10365.0 197052.5 ;
      RECT  10485.0 198027.5 10555.0 197892.5 ;
      RECT  10587.5 197585.0 10452.5 197515.0 ;
      RECT  9220.0 197495.0 9290.0 197630.0 ;
      RECT  9360.0 197767.5 9430.0 197902.5 ;
      RECT  10357.5 197730.0 10222.5 197800.0 ;
      RECT  10295.0 198795.0 10365.0 198865.0 ;
      RECT  10485.0 198795.0 10555.0 198865.0 ;
      RECT  10295.0 198830.0 10365.0 199192.5 ;
      RECT  10330.0 198795.0 10520.0 198865.0 ;
      RECT  10485.0 198487.5 10555.0 198830.0 ;
      RECT  10295.0 199192.5 10365.0 199327.5 ;
      RECT  10485.0 198352.5 10555.0 198487.5 ;
      RECT  10587.5 198795.0 10452.5 198865.0 ;
      RECT  9220.0 198750.0 9290.0 198885.0 ;
      RECT  9360.0 198477.5 9430.0 198612.5 ;
      RECT  10357.5 198580.0 10222.5 198650.0 ;
      RECT  10295.0 200275.0 10365.0 200205.0 ;
      RECT  10485.0 200275.0 10555.0 200205.0 ;
      RECT  10295.0 200240.0 10365.0 199877.5 ;
      RECT  10330.0 200275.0 10520.0 200205.0 ;
      RECT  10485.0 200582.5 10555.0 200240.0 ;
      RECT  10295.0 199877.5 10365.0 199742.5 ;
      RECT  10485.0 200717.5 10555.0 200582.5 ;
      RECT  10587.5 200275.0 10452.5 200205.0 ;
      RECT  9220.0 200185.0 9290.0 200320.0 ;
      RECT  9360.0 200457.5 9430.0 200592.5 ;
      RECT  10357.5 200420.0 10222.5 200490.0 ;
      RECT  10295.0 201485.0 10365.0 201555.0 ;
      RECT  10485.0 201485.0 10555.0 201555.0 ;
      RECT  10295.0 201520.0 10365.0 201882.5 ;
      RECT  10330.0 201485.0 10520.0 201555.0 ;
      RECT  10485.0 201177.5 10555.0 201520.0 ;
      RECT  10295.0 201882.5 10365.0 202017.5 ;
      RECT  10485.0 201042.5 10555.0 201177.5 ;
      RECT  10587.5 201485.0 10452.5 201555.0 ;
      RECT  9220.0 201440.0 9290.0 201575.0 ;
      RECT  9360.0 201167.5 9430.0 201302.5 ;
      RECT  10357.5 201270.0 10222.5 201340.0 ;
      RECT  10295.0 202965.0 10365.0 202895.0 ;
      RECT  10485.0 202965.0 10555.0 202895.0 ;
      RECT  10295.0 202930.0 10365.0 202567.5 ;
      RECT  10330.0 202965.0 10520.0 202895.0 ;
      RECT  10485.0 203272.5 10555.0 202930.0 ;
      RECT  10295.0 202567.5 10365.0 202432.5 ;
      RECT  10485.0 203407.5 10555.0 203272.5 ;
      RECT  10587.5 202965.0 10452.5 202895.0 ;
      RECT  9220.0 202875.0 9290.0 203010.0 ;
      RECT  9360.0 203147.5 9430.0 203282.5 ;
      RECT  10357.5 203110.0 10222.5 203180.0 ;
      RECT  10295.0 204175.0 10365.0 204245.0 ;
      RECT  10485.0 204175.0 10555.0 204245.0 ;
      RECT  10295.0 204210.0 10365.0 204572.5 ;
      RECT  10330.0 204175.0 10520.0 204245.0 ;
      RECT  10485.0 203867.5 10555.0 204210.0 ;
      RECT  10295.0 204572.5 10365.0 204707.5 ;
      RECT  10485.0 203732.5 10555.0 203867.5 ;
      RECT  10587.5 204175.0 10452.5 204245.0 ;
      RECT  9220.0 204130.0 9290.0 204265.0 ;
      RECT  9360.0 203857.5 9430.0 203992.5 ;
      RECT  10357.5 203960.0 10222.5 204030.0 ;
      RECT  10295.0 205655.0 10365.0 205585.0 ;
      RECT  10485.0 205655.0 10555.0 205585.0 ;
      RECT  10295.0 205620.0 10365.0 205257.5 ;
      RECT  10330.0 205655.0 10520.0 205585.0 ;
      RECT  10485.0 205962.5 10555.0 205620.0 ;
      RECT  10295.0 205257.5 10365.0 205122.5 ;
      RECT  10485.0 206097.5 10555.0 205962.5 ;
      RECT  10587.5 205655.0 10452.5 205585.0 ;
      RECT  9220.0 205565.0 9290.0 205700.0 ;
      RECT  9360.0 205837.5 9430.0 205972.5 ;
      RECT  10357.5 205800.0 10222.5 205870.0 ;
      RECT  9220.0 34100.0 9290.0 206260.0 ;
      RECT  4655.0 12170.0 11095.0 11465.0 ;
      RECT  4655.0 10760.0 11095.0 11465.0 ;
      RECT  4655.0 10760.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 5825.0 ;
      RECT  4655.0 11852.5 4800.0 11782.5 ;
      RECT  4655.0 11147.5 4800.0 11077.5 ;
      RECT  4655.0 10442.5 4800.0 10372.5 ;
      RECT  4655.0 9737.5 4800.0 9667.5 ;
      RECT  4655.0 9032.5 4800.0 8962.5 ;
      RECT  4655.0 8327.5 4800.0 8257.5 ;
      RECT  4655.0 7622.5 4800.0 7552.5 ;
      RECT  4655.0 6917.5 4800.0 6847.5 ;
      RECT  4655.0 6212.5 4800.0 6142.5 ;
      RECT  10825.0 11852.5 11095.0 11782.5 ;
      RECT  10407.5 12007.5 11095.0 11937.5 ;
      RECT  10825.0 11147.5 11095.0 11077.5 ;
      RECT  10407.5 10992.5 11095.0 10922.5 ;
      RECT  10825.0 10442.5 11095.0 10372.5 ;
      RECT  10407.5 10597.5 11095.0 10527.5 ;
      RECT  10825.0 9737.5 11095.0 9667.5 ;
      RECT  10407.5 9582.5 11095.0 9512.5 ;
      RECT  10825.0 9032.5 11095.0 8962.5 ;
      RECT  10407.5 9187.5 11095.0 9117.5 ;
      RECT  10825.0 8327.5 11095.0 8257.5 ;
      RECT  10407.5 8172.5 11095.0 8102.5 ;
      RECT  10825.0 7622.5 11095.0 7552.5 ;
      RECT  10407.5 7777.5 11095.0 7707.5 ;
      RECT  10825.0 6917.5 11095.0 6847.5 ;
      RECT  10407.5 6762.5 11095.0 6692.5 ;
      RECT  10825.0 6212.5 11095.0 6142.5 ;
      RECT  10407.5 6367.5 11095.0 6297.5 ;
      RECT  4655.0 12205.0 11095.0 12135.0 ;
      RECT  4655.0 11500.0 11095.0 11430.0 ;
      RECT  4655.0 10795.0 11095.0 10725.0 ;
      RECT  4655.0 10090.0 11095.0 10020.0 ;
      RECT  4655.0 9385.0 11095.0 9315.0 ;
      RECT  4655.0 8680.0 11095.0 8610.0 ;
      RECT  4655.0 7975.0 11095.0 7905.0 ;
      RECT  4655.0 7270.0 11095.0 7200.0 ;
      RECT  4655.0 6565.0 11095.0 6495.0 ;
      RECT  4655.0 5860.0 11095.0 5790.0 ;
      RECT  17302.5 12605.0 17372.5 12740.0 ;
      RECT  20122.5 12605.0 20192.5 12740.0 ;
      RECT  22942.5 12605.0 23012.5 12740.0 ;
      RECT  25762.5 12605.0 25832.5 12740.0 ;
      RECT  28582.5 12605.0 28652.5 12740.0 ;
      RECT  31402.5 12605.0 31472.5 12740.0 ;
      RECT  34222.5 12605.0 34292.5 12740.0 ;
      RECT  37042.5 12605.0 37112.5 12740.0 ;
      RECT  39862.5 12605.0 39932.5 12740.0 ;
      RECT  42682.5 12605.0 42752.5 12740.0 ;
      RECT  45502.5 12605.0 45572.5 12740.0 ;
      RECT  48322.5 12605.0 48392.5 12740.0 ;
      RECT  51142.5 12605.0 51212.5 12740.0 ;
      RECT  53962.5 12605.0 54032.5 12740.0 ;
      RECT  56782.5 12605.0 56852.5 12740.0 ;
      RECT  59602.5 12605.0 59672.5 12740.0 ;
      RECT  62422.5 12605.0 62492.5 12740.0 ;
      RECT  65242.5 12605.0 65312.5 12740.0 ;
      RECT  68062.5 12605.0 68132.5 12740.0 ;
      RECT  70882.5 12605.0 70952.5 12740.0 ;
      RECT  73702.5 12605.0 73772.5 12740.0 ;
      RECT  76522.5 12605.0 76592.5 12740.0 ;
      RECT  79342.5 12605.0 79412.5 12740.0 ;
      RECT  82162.5 12605.0 82232.5 12740.0 ;
      RECT  84982.5 12605.0 85052.5 12740.0 ;
      RECT  87802.5 12605.0 87872.5 12740.0 ;
      RECT  90622.5 12605.0 90692.5 12740.0 ;
      RECT  93442.5 12605.0 93512.5 12740.0 ;
      RECT  96262.5 12605.0 96332.5 12740.0 ;
      RECT  99082.5 12605.0 99152.5 12740.0 ;
      RECT  101902.5 12605.0 101972.5 12740.0 ;
      RECT  104722.5 12605.0 104792.5 12740.0 ;
      RECT  17512.5 35.0 17582.5 170.0 ;
      RECT  20332.5 35.0 20402.5 170.0 ;
      RECT  23152.5 35.0 23222.5 170.0 ;
      RECT  25972.5 35.0 26042.5 170.0 ;
      RECT  28792.5 35.0 28862.5 170.0 ;
      RECT  31612.5 35.0 31682.5 170.0 ;
      RECT  34432.5 35.0 34502.5 170.0 ;
      RECT  37252.5 35.0 37322.5 170.0 ;
      RECT  40072.5 35.0 40142.5 170.0 ;
      RECT  42892.5 35.0 42962.5 170.0 ;
      RECT  45712.5 35.0 45782.5 170.0 ;
      RECT  48532.5 35.0 48602.5 170.0 ;
      RECT  51352.5 35.0 51422.5 170.0 ;
      RECT  54172.5 35.0 54242.5 170.0 ;
      RECT  56992.5 35.0 57062.5 170.0 ;
      RECT  59812.5 35.0 59882.5 170.0 ;
      RECT  62632.5 35.0 62702.5 170.0 ;
      RECT  65452.5 35.0 65522.5 170.0 ;
      RECT  68272.5 35.0 68342.5 170.0 ;
      RECT  71092.5 35.0 71162.5 170.0 ;
      RECT  73912.5 35.0 73982.5 170.0 ;
      RECT  76732.5 35.0 76802.5 170.0 ;
      RECT  79552.5 35.0 79622.5 170.0 ;
      RECT  82372.5 35.0 82442.5 170.0 ;
      RECT  85192.5 35.0 85262.5 170.0 ;
      RECT  88012.5 35.0 88082.5 170.0 ;
      RECT  90832.5 35.0 90902.5 170.0 ;
      RECT  93652.5 35.0 93722.5 170.0 ;
      RECT  96472.5 35.0 96542.5 170.0 ;
      RECT  99292.5 35.0 99362.5 170.0 ;
      RECT  102112.5 35.0 102182.5 170.0 ;
      RECT  104932.5 35.0 105002.5 170.0 ;
      RECT  15102.5 34135.0 15237.5 34065.0 ;
      RECT  15102.5 36825.0 15237.5 36755.0 ;
      RECT  15102.5 39515.0 15237.5 39445.0 ;
      RECT  15102.5 42205.0 15237.5 42135.0 ;
      RECT  15102.5 44895.0 15237.5 44825.0 ;
      RECT  15102.5 47585.0 15237.5 47515.0 ;
      RECT  15102.5 50275.0 15237.5 50205.0 ;
      RECT  15102.5 52965.0 15237.5 52895.0 ;
      RECT  15102.5 55655.0 15237.5 55585.0 ;
      RECT  15102.5 58345.0 15237.5 58275.0 ;
      RECT  15102.5 61035.0 15237.5 60965.0 ;
      RECT  15102.5 63725.0 15237.5 63655.0 ;
      RECT  15102.5 66415.0 15237.5 66345.0 ;
      RECT  15102.5 69105.0 15237.5 69035.0 ;
      RECT  15102.5 71795.0 15237.5 71725.0 ;
      RECT  15102.5 74485.0 15237.5 74415.0 ;
      RECT  15102.5 77175.0 15237.5 77105.0 ;
      RECT  15102.5 79865.0 15237.5 79795.0 ;
      RECT  15102.5 82555.0 15237.5 82485.0 ;
      RECT  15102.5 85245.0 15237.5 85175.0 ;
      RECT  15102.5 87935.0 15237.5 87865.0 ;
      RECT  15102.5 90625.0 15237.5 90555.0 ;
      RECT  15102.5 93315.0 15237.5 93245.0 ;
      RECT  15102.5 96005.0 15237.5 95935.0 ;
      RECT  15102.5 98695.0 15237.5 98625.0 ;
      RECT  15102.5 101385.0 15237.5 101315.0 ;
      RECT  15102.5 104075.0 15237.5 104005.0 ;
      RECT  15102.5 106765.0 15237.5 106695.0 ;
      RECT  15102.5 109455.0 15237.5 109385.0 ;
      RECT  15102.5 112145.0 15237.5 112075.0 ;
      RECT  15102.5 114835.0 15237.5 114765.0 ;
      RECT  15102.5 117525.0 15237.5 117455.0 ;
      RECT  15102.5 120215.0 15237.5 120145.0 ;
      RECT  15102.5 122905.0 15237.5 122835.0 ;
      RECT  15102.5 125595.0 15237.5 125525.0 ;
      RECT  15102.5 128285.0 15237.5 128215.0 ;
      RECT  15102.5 130975.0 15237.5 130905.0 ;
      RECT  15102.5 133665.0 15237.5 133595.0 ;
      RECT  15102.5 136355.0 15237.5 136285.0 ;
      RECT  15102.5 139045.0 15237.5 138975.0 ;
      RECT  15102.5 141735.0 15237.5 141665.0 ;
      RECT  15102.5 144425.0 15237.5 144355.0 ;
      RECT  15102.5 147115.0 15237.5 147045.0 ;
      RECT  15102.5 149805.0 15237.5 149735.0 ;
      RECT  15102.5 152495.0 15237.5 152425.0 ;
      RECT  15102.5 155185.0 15237.5 155115.0 ;
      RECT  15102.5 157875.0 15237.5 157805.0 ;
      RECT  15102.5 160565.0 15237.5 160495.0 ;
      RECT  15102.5 163255.0 15237.5 163185.0 ;
      RECT  15102.5 165945.0 15237.5 165875.0 ;
      RECT  15102.5 168635.0 15237.5 168565.0 ;
      RECT  15102.5 171325.0 15237.5 171255.0 ;
      RECT  15102.5 174015.0 15237.5 173945.0 ;
      RECT  15102.5 176705.0 15237.5 176635.0 ;
      RECT  15102.5 179395.0 15237.5 179325.0 ;
      RECT  15102.5 182085.0 15237.5 182015.0 ;
      RECT  15102.5 184775.0 15237.5 184705.0 ;
      RECT  15102.5 187465.0 15237.5 187395.0 ;
      RECT  15102.5 190155.0 15237.5 190085.0 ;
      RECT  15102.5 192845.0 15237.5 192775.0 ;
      RECT  15102.5 195535.0 15237.5 195465.0 ;
      RECT  15102.5 198225.0 15237.5 198155.0 ;
      RECT  15102.5 200915.0 15237.5 200845.0 ;
      RECT  15102.5 203605.0 15237.5 203535.0 ;
      RECT  15102.5 206295.0 15237.5 206225.0 ;
      RECT  11420.0 12750.0 11285.0 12820.0 ;
      RECT  12745.0 12750.0 12610.0 12820.0 ;
      RECT  11145.0 14095.0 11010.0 14165.0 ;
      RECT  12950.0 14095.0 12815.0 14165.0 ;
      RECT  11420.0 18130.0 11285.0 18200.0 ;
      RECT  13155.0 18130.0 13020.0 18200.0 ;
      RECT  11145.0 19475.0 11010.0 19545.0 ;
      RECT  13360.0 19475.0 13225.0 19545.0 ;
      RECT  12335.0 23510.0 12200.0 23580.0 ;
      RECT  13565.0 23510.0 13430.0 23580.0 ;
      RECT  12060.0 24855.0 11925.0 24925.0 ;
      RECT  13770.0 24855.0 13635.0 24925.0 ;
      RECT  11785.0 26200.0 11650.0 26270.0 ;
      RECT  13975.0 26200.0 13840.0 26270.0 ;
      RECT  12540.0 12545.0 12405.0 12615.0 ;
      RECT  12540.0 12545.0 12405.0 12615.0 ;
      RECT  15035.0 12615.0 15170.0 12545.0 ;
      RECT  12540.0 15235.0 12405.0 15305.0 ;
      RECT  12540.0 15235.0 12405.0 15305.0 ;
      RECT  15035.0 15305.0 15170.0 15235.0 ;
      RECT  12540.0 17925.0 12405.0 17995.0 ;
      RECT  12540.0 17925.0 12405.0 17995.0 ;
      RECT  15035.0 17995.0 15170.0 17925.0 ;
      RECT  12540.0 20615.0 12405.0 20685.0 ;
      RECT  12540.0 20615.0 12405.0 20685.0 ;
      RECT  15035.0 20685.0 15170.0 20615.0 ;
      RECT  12540.0 23305.0 12405.0 23375.0 ;
      RECT  12540.0 23305.0 12405.0 23375.0 ;
      RECT  15035.0 23375.0 15170.0 23305.0 ;
      RECT  12540.0 25995.0 12405.0 26065.0 ;
      RECT  12540.0 25995.0 12405.0 26065.0 ;
      RECT  15035.0 26065.0 15170.0 25995.0 ;
      RECT  12540.0 28685.0 12405.0 28755.0 ;
      RECT  12540.0 28685.0 12405.0 28755.0 ;
      RECT  15035.0 28755.0 15170.0 28685.0 ;
      RECT  12540.0 31375.0 12405.0 31445.0 ;
      RECT  12540.0 31375.0 12405.0 31445.0 ;
      RECT  15035.0 31445.0 15170.0 31375.0 ;
      RECT  14180.0 32095.0 14045.0 32165.0 ;
      RECT  14385.0 31955.0 14250.0 32025.0 ;
      RECT  14590.0 31815.0 14455.0 31885.0 ;
      RECT  14795.0 31675.0 14660.0 31745.0 ;
      RECT  14180.0 627.5 14045.0 697.5 ;
      RECT  14385.0 2062.5 14250.0 2132.5 ;
      RECT  14590.0 3317.5 14455.0 3387.5 ;
      RECT  14795.0 4752.5 14660.0 4822.5 ;
      RECT  15102.5 70.0 15237.5 2.49800180541e-13 ;
      RECT  15102.5 2760.0 15237.5 2690.0 ;
      RECT  15102.5 5450.0 15237.5 5380.0 ;
      RECT  11162.5 6847.5 11027.5 6917.5 ;
      RECT  7960.0 5207.5 8030.0 5342.5 ;
      RECT  11162.5 6142.5 11027.5 6212.5 ;
      RECT  8235.0 5207.5 8305.0 5342.5 ;
      RECT  11162.5 11782.5 11027.5 11852.5 ;
      RECT  12745.0 11782.5 12610.0 11852.5 ;
      RECT  11162.5 11077.5 11027.5 11147.5 ;
      RECT  12950.0 11077.5 12815.0 11147.5 ;
      RECT  11162.5 10372.5 11027.5 10442.5 ;
      RECT  13155.0 10372.5 13020.0 10442.5 ;
      RECT  11162.5 9667.5 11027.5 9737.5 ;
      RECT  13360.0 9667.5 13225.0 9737.5 ;
      RECT  11162.5 8962.5 11027.5 9032.5 ;
      RECT  13565.0 8962.5 13430.0 9032.5 ;
      RECT  11162.5 8257.5 11027.5 8327.5 ;
      RECT  13770.0 8257.5 13635.0 8327.5 ;
      RECT  11162.5 7552.5 11027.5 7622.5 ;
      RECT  13975.0 7552.5 13840.0 7622.5 ;
      RECT  11230.0 12135.0 11095.0 12205.0 ;
      RECT  15237.5 12135.0 15102.5 12205.0 ;
      RECT  11230.0 11430.0 11095.0 11500.0 ;
      RECT  15237.5 11430.0 15102.5 11500.0 ;
      RECT  11230.0 10725.0 11095.0 10795.0 ;
      RECT  15237.5 10725.0 15102.5 10795.0 ;
      RECT  11230.0 10020.0 11095.0 10090.0 ;
      RECT  15237.5 10020.0 15102.5 10090.0 ;
      RECT  11230.0 9315.0 11095.0 9385.0 ;
      RECT  15237.5 9315.0 15102.5 9385.0 ;
      RECT  11230.0 8610.0 11095.0 8680.0 ;
      RECT  15237.5 8610.0 15102.5 8680.0 ;
      RECT  11230.0 7905.0 11095.0 7975.0 ;
      RECT  15237.5 7905.0 15102.5 7975.0 ;
      RECT  11230.0 7200.0 11095.0 7270.0 ;
      RECT  15237.5 7200.0 15102.5 7270.0 ;
      RECT  11230.0 6495.0 11095.0 6565.0 ;
      RECT  15237.5 6495.0 15102.5 6565.0 ;
      RECT  11230.0 5790.0 11095.0 5860.0 ;
      RECT  15237.5 5790.0 15102.5 5860.0 ;
      RECT  16375.0 15957.5 16240.0 16027.5 ;
      RECT  15965.0 13772.5 15830.0 13842.5 ;
      RECT  16170.0 15320.0 16035.0 15390.0 ;
      RECT  16375.0 207235.0 16240.0 207305.0 ;
      RECT  16580.0 22460.0 16445.0 22530.0 ;
      RECT  16785.0 26485.0 16650.0 26555.0 ;
      RECT  15760.0 12340.0 15625.0 12410.0 ;
      RECT  9322.5 206430.0 9187.5 206500.0 ;
      RECT  15760.0 206430.0 15625.0 206500.0 ;
      RECT  15452.5 15190.0 15317.5 15260.0 ;
      RECT  15452.5 26615.0 15317.5 26685.0 ;
      RECT  15452.5 16117.5 15317.5 16187.5 ;
      RECT  15452.5 23392.5 15317.5 23462.5 ;
      RECT  17512.5 35.0 17582.5 175.0 ;
      RECT  20332.5 35.0 20402.5 175.0 ;
      RECT  23152.5 35.0 23222.5 175.0 ;
      RECT  25972.5 35.0 26042.5 175.0 ;
      RECT  28792.5 35.0 28862.5 175.0 ;
      RECT  31612.5 35.0 31682.5 175.0 ;
      RECT  34432.5 35.0 34502.5 175.0 ;
      RECT  37252.5 35.0 37322.5 175.0 ;
      RECT  40072.5 35.0 40142.5 175.0 ;
      RECT  42892.5 35.0 42962.5 175.0 ;
      RECT  45712.5 35.0 45782.5 175.0 ;
      RECT  48532.5 35.0 48602.5 175.0 ;
      RECT  51352.5 35.0 51422.5 175.0 ;
      RECT  54172.5 35.0 54242.5 175.0 ;
      RECT  56992.5 35.0 57062.5 175.0 ;
      RECT  59812.5 35.0 59882.5 175.0 ;
      RECT  62632.5 35.0 62702.5 175.0 ;
      RECT  65452.5 35.0 65522.5 175.0 ;
      RECT  68272.5 35.0 68342.5 175.0 ;
      RECT  71092.5 35.0 71162.5 175.0 ;
      RECT  73912.5 35.0 73982.5 175.0 ;
      RECT  76732.5 35.0 76802.5 175.0 ;
      RECT  79552.5 35.0 79622.5 175.0 ;
      RECT  82372.5 35.0 82442.5 175.0 ;
      RECT  85192.5 35.0 85262.5 175.0 ;
      RECT  88012.5 35.0 88082.5 175.0 ;
      RECT  90832.5 35.0 90902.5 175.0 ;
      RECT  93652.5 35.0 93722.5 175.0 ;
      RECT  96472.5 35.0 96542.5 175.0 ;
      RECT  99292.5 35.0 99362.5 175.0 ;
      RECT  102112.5 35.0 102182.5 175.0 ;
      RECT  104932.5 35.0 105002.5 175.0 ;
      RECT  16682.5 35.0 16752.5 207987.5 ;
      RECT  16477.5 35.0 16547.5 207987.5 ;
      RECT  15862.5 35.0 15932.5 207987.5 ;
      RECT  16067.5 35.0 16137.5 207987.5 ;
      RECT  16272.5 35.0 16342.5 207987.5 ;
      RECT  15657.5 35.0 15727.5 207987.5 ;
      RECT  15102.5 35.0 15452.5 207987.5 ;
      RECT  4035.0 41500.0 8.881784197e-13 41570.0 ;
      RECT  4035.0 41705.0 8.881784197e-13 41775.0 ;
      RECT  4035.0 41910.0 8.881784197e-13 41980.0 ;
      RECT  4035.0 42320.0 8.881784197e-13 42390.0 ;
      RECT  3422.5 37010.0 2690.0 37080.0 ;
      RECT  2520.0 34477.5 2450.0 41125.0 ;
      RECT  4035.0 41295.0 3830.0 41365.0 ;
      RECT  2895.0 42115.0 2690.0 42185.0 ;
      RECT  1550.0 41295.0 1345.0 41365.0 ;
      RECT  205.0 42115.0 8.881784197e-13 42185.0 ;
      RECT  165.0 34240.0 870.0 40680.0 ;
      RECT  1575.0 34240.0 870.0 40680.0 ;
      RECT  1575.0 34240.0 2280.0 40680.0 ;
      RECT  482.5 34240.0 552.5 34385.0 ;
      RECT  1187.5 34240.0 1257.5 34385.0 ;
      RECT  1892.5 34240.0 1962.5 34385.0 ;
      RECT  482.5 40410.0 552.5 40680.0 ;
      RECT  327.5 39992.5 397.5 40680.0 ;
      RECT  1187.5 40410.0 1257.5 40680.0 ;
      RECT  1342.5 39992.5 1412.5 40680.0 ;
      RECT  1892.5 40410.0 1962.5 40680.0 ;
      RECT  1737.5 39992.5 1807.5 40680.0 ;
      RECT  130.0 34240.0 200.0 40680.0 ;
      RECT  835.0 34240.0 905.0 40680.0 ;
      RECT  1540.0 34240.0 1610.0 40680.0 ;
      RECT  2245.0 34240.0 2315.0 40680.0 ;
      RECT  3737.5 43570.0 3032.5 43640.0 ;
      RECT  3382.5 43190.0 3312.5 43260.0 ;
      RECT  3382.5 43570.0 3312.5 43640.0 ;
      RECT  3347.5 43190.0 3032.5 43260.0 ;
      RECT  3382.5 43225.0 3312.5 43605.0 ;
      RECT  3737.5 43570.0 3347.5 43640.0 ;
      RECT  3032.5 43190.0 2897.5 43260.0 ;
      RECT  3032.5 43570.0 2897.5 43640.0 ;
      RECT  3872.5 43570.0 3737.5 43640.0 ;
      RECT  3415.0 43570.0 3280.0 43640.0 ;
      RECT  1895.0 43380.0 1965.0 43450.0 ;
      RECT  1930.0 43380.0 2280.0 43450.0 ;
      RECT  1895.0 43415.0 1965.0 43485.0 ;
      RECT  1495.0 43380.0 1565.0 43450.0 ;
      RECT  1495.0 43257.5 1565.0 43415.0 ;
      RECT  1530.0 43380.0 1930.0 43450.0 ;
      RECT  2280.0 43380.0 2415.0 43450.0 ;
      RECT  1495.0 43292.5 1565.0 43157.5 ;
      RECT  1895.0 43552.5 1965.0 43417.5 ;
      RECT  1950.0 44335.0 2020.0 44405.0 ;
      RECT  1950.0 44525.0 2020.0 44595.0 ;
      RECT  1985.0 44335.0 2347.5 44405.0 ;
      RECT  1950.0 44370.0 2020.0 44560.0 ;
      RECT  1642.5 44525.0 1985.0 44595.0 ;
      RECT  2347.5 44335.0 2482.5 44405.0 ;
      RECT  1507.5 44525.0 1642.5 44595.0 ;
      RECT  1950.0 44627.5 2020.0 44492.5 ;
      RECT  1047.5 44130.0 342.5 44200.0 ;
      RECT  692.5 43750.0 622.5 43820.0 ;
      RECT  692.5 44130.0 622.5 44200.0 ;
      RECT  657.5 43750.0 342.5 43820.0 ;
      RECT  692.5 43785.0 622.5 44165.0 ;
      RECT  1047.5 44130.0 657.5 44200.0 ;
      RECT  342.5 43750.0 207.5 43820.0 ;
      RECT  342.5 44130.0 207.5 44200.0 ;
      RECT  1182.5 44130.0 1047.5 44200.0 ;
      RECT  725.0 44130.0 590.0 44200.0 ;
      RECT  397.5 40747.5 327.5 40612.5 ;
      RECT  397.5 42422.5 327.5 42287.5 ;
      RECT  552.5 40747.5 482.5 40612.5 ;
      RECT  552.5 41602.5 482.5 41467.5 ;
      RECT  1412.5 40747.5 1342.5 40612.5 ;
      RECT  1412.5 41807.5 1342.5 41672.5 ;
      RECT  1807.5 40747.5 1737.5 40612.5 ;
      RECT  1807.5 42012.5 1737.5 41877.5 ;
      RECT  200.0 40747.5 130.0 40612.5 ;
      RECT  200.0 41397.5 130.0 41262.5 ;
      RECT  905.0 40747.5 835.0 40612.5 ;
      RECT  905.0 41397.5 835.0 41262.5 ;
      RECT  1610.0 40747.5 1540.0 40612.5 ;
      RECT  1610.0 41397.5 1540.0 41262.5 ;
      RECT  2315.0 40747.5 2245.0 40612.5 ;
      RECT  2315.0 41397.5 2245.0 41262.5 ;
      RECT  1380.0 46905.0 1310.0 84245.0 ;
      RECT  970.0 46905.0 900.0 83935.0 ;
      RECT  265.0 46905.0 195.0 83935.0 ;
      RECT  1207.5 47072.5 1137.5 47670.0 ;
      RECT  785.0 47072.5 715.0 47352.5 ;
      RECT  3372.5 49467.5 3442.5 49862.5 ;
      RECT  3372.5 49862.5 3442.5 50422.5 ;
      RECT  3372.5 50422.5 3442.5 50982.5 ;
      RECT  3372.5 51147.5 3442.5 51542.5 ;
      RECT  3372.5 51542.5 3442.5 52102.5 ;
      RECT  3372.5 52102.5 3442.5 52662.5 ;
      RECT  2655.0 52792.5 2725.0 52862.5 ;
      RECT  2655.0 52312.5 2725.0 52382.5 ;
      RECT  2690.0 52792.5 3407.5 52862.5 ;
      RECT  2655.0 52347.5 2725.0 52827.5 ;
      RECT  1972.5 52312.5 2690.0 52382.5 ;
      RECT  1937.5 51787.5 2007.5 52347.5 ;
      RECT  1937.5 51227.5 2007.5 51787.5 ;
      RECT  1937.5 50667.5 2007.5 51062.5 ;
      RECT  1937.5 50107.5 2007.5 50667.5 ;
      RECT  1937.5 49547.5 2007.5 50107.5 ;
      RECT  3340.0 49827.5 3475.0 49897.5 ;
      RECT  3340.0 50387.5 3475.0 50457.5 ;
      RECT  3340.0 50947.5 3475.0 51017.5 ;
      RECT  3340.0 51507.5 3475.0 51577.5 ;
      RECT  3340.0 52067.5 3475.0 52137.5 ;
      RECT  3340.0 52627.5 3475.0 52697.5 ;
      RECT  1905.0 52312.5 2040.0 52382.5 ;
      RECT  1905.0 51752.5 2040.0 51822.5 ;
      RECT  1905.0 51192.5 2040.0 51262.5 ;
      RECT  1905.0 50632.5 2040.0 50702.5 ;
      RECT  1905.0 50072.5 2040.0 50142.5 ;
      RECT  1905.0 49512.5 2040.0 49582.5 ;
      RECT  3340.0 49432.5 3475.0 49502.5 ;
      RECT  3340.0 51112.5 3475.0 51182.5 ;
      RECT  3340.0 52792.5 3475.0 52862.5 ;
      RECT  1905.0 51027.5 2040.0 51097.5 ;
      RECT  935.0 48810.0 225.0 47465.0 ;
      RECT  935.0 48810.0 230.0 50155.0 ;
      RECT  935.0 51500.0 230.0 50155.0 ;
      RECT  935.0 51500.0 230.0 52845.0 ;
      RECT  935.0 54190.0 230.0 52845.0 ;
      RECT  935.0 54190.0 230.0 55535.0 ;
      RECT  935.0 56880.0 230.0 55535.0 ;
      RECT  935.0 56880.0 230.0 58225.0 ;
      RECT  935.0 59570.0 230.0 58225.0 ;
      RECT  935.0 59570.0 230.0 60915.0 ;
      RECT  935.0 62260.0 230.0 60915.0 ;
      RECT  935.0 62260.0 230.0 63605.0 ;
      RECT  935.0 64950.0 230.0 63605.0 ;
      RECT  935.0 64950.0 230.0 66295.0 ;
      RECT  935.0 67640.0 230.0 66295.0 ;
      RECT  935.0 67640.0 230.0 68985.0 ;
      RECT  935.0 70330.0 230.0 68985.0 ;
      RECT  935.0 70330.0 230.0 71675.0 ;
      RECT  935.0 73020.0 230.0 71675.0 ;
      RECT  935.0 73020.0 230.0 74365.0 ;
      RECT  935.0 75710.0 230.0 74365.0 ;
      RECT  935.0 75710.0 230.0 77055.0 ;
      RECT  935.0 78400.0 230.0 77055.0 ;
      RECT  935.0 78400.0 230.0 79745.0 ;
      RECT  935.0 81090.0 230.0 79745.0 ;
      RECT  935.0 81090.0 230.0 82435.0 ;
      RECT  935.0 83780.0 230.0 82435.0 ;
      RECT  785.0 48710.0 715.0 83935.0 ;
      RECT  450.0 48710.0 380.0 83935.0 ;
      RECT  970.0 48710.0 900.0 83935.0 ;
      RECT  265.0 48710.0 195.0 83935.0 ;
      RECT  1347.5 48882.5 1277.5 49017.5 ;
      RECT  1347.5 51292.5 1277.5 51427.5 ;
      RECT  1347.5 51572.5 1277.5 51707.5 ;
      RECT  1347.5 53982.5 1277.5 54117.5 ;
      RECT  1347.5 54262.5 1277.5 54397.5 ;
      RECT  1347.5 56672.5 1277.5 56807.5 ;
      RECT  1347.5 56952.5 1277.5 57087.5 ;
      RECT  1347.5 59362.5 1277.5 59497.5 ;
      RECT  1347.5 59642.5 1277.5 59777.5 ;
      RECT  1347.5 62052.5 1277.5 62187.5 ;
      RECT  1347.5 62332.5 1277.5 62467.5 ;
      RECT  1347.5 64742.5 1277.5 64877.5 ;
      RECT  1347.5 65022.5 1277.5 65157.5 ;
      RECT  1347.5 67432.5 1277.5 67567.5 ;
      RECT  1347.5 67712.5 1277.5 67847.5 ;
      RECT  1347.5 70122.5 1277.5 70257.5 ;
      RECT  1347.5 70402.5 1277.5 70537.5 ;
      RECT  1347.5 72812.5 1277.5 72947.5 ;
      RECT  1347.5 73092.5 1277.5 73227.5 ;
      RECT  1347.5 75502.5 1277.5 75637.5 ;
      RECT  1347.5 75782.5 1277.5 75917.5 ;
      RECT  1347.5 78192.5 1277.5 78327.5 ;
      RECT  1347.5 78472.5 1277.5 78607.5 ;
      RECT  1347.5 80882.5 1277.5 81017.5 ;
      RECT  1347.5 81162.5 1277.5 81297.5 ;
      RECT  1347.5 83572.5 1277.5 83707.5 ;
      RECT  1345.0 49145.0 1275.0 49280.0 ;
      RECT  1380.0 46770.0 1310.0 46905.0 ;
      RECT  867.5 46870.0 1002.5 46940.0 ;
      RECT  162.5 46870.0 297.5 46940.0 ;
      RECT  1105.0 47635.0 1240.0 47705.0 ;
      RECT  1105.0 47037.5 1240.0 47107.5 ;
      RECT  682.5 47037.5 817.5 47107.5 ;
      RECT  3457.5 41192.5 3387.5 41057.5 ;
      RECT  3457.5 37112.5 3387.5 36977.5 ;
      RECT  2725.0 37112.5 2655.0 36977.5 ;
      RECT  2725.0 42627.5 2655.0 42492.5 ;
      RECT  2520.0 34545.0 2450.0 34410.0 ;
      RECT  1965.0 41192.5 1895.0 41057.5 ;
      RECT  1750.0 41602.5 1680.0 41467.5 ;
      RECT  2020.0 44140.0 1950.0 44005.0 ;
      RECT  2020.0 44140.0 1950.0 44005.0 ;
      RECT  2020.0 42627.5 1950.0 42492.5 ;
      RECT  1805.0 44397.5 1735.0 44262.5 ;
      RECT  1805.0 44397.5 1735.0 44262.5 ;
      RECT  1805.0 42422.5 1735.0 42287.5 ;
      RECT  3382.5 42627.5 3312.5 42492.5 ;
      RECT  3522.5 42422.5 3452.5 42287.5 ;
      RECT  3662.5 41807.5 3592.5 41672.5 ;
      RECT  692.5 42627.5 622.5 42492.5 ;
      RECT  832.5 41807.5 762.5 41672.5 ;
      RECT  972.5 42012.5 902.5 41877.5 ;
      RECT  1997.5 43820.0 1862.5 43890.0 ;
      RECT  2052.5 44965.0 1917.5 45035.0 ;
      RECT  785.0 46150.0 650.0 46220.0 ;
      RECT  2040.0 45190.0 1905.0 45260.0 ;
      RECT  4070.0 41397.5 4000.0 41262.5 ;
      RECT  2725.0 42217.5 2655.0 42082.5 ;
      RECT  1380.0 41397.5 1310.0 41262.5 ;
      RECT  35.0 42217.5 -35.0 42082.5 ;
      RECT  4035.0 45190.0 1972.5 45260.0 ;
      RECT  4035.0 46150.0 717.5 46220.0 ;
      RECT  4035.0 43820.0 1930.0 43890.0 ;
      RECT  4035.0 44965.0 1985.0 45035.0 ;
      RECT  4035.0 42525.0 8.881784197e-13 42595.0 ;
      RECT  4035.0 41090.0 0.0 41160.0 ;
      RECT  4035.0 42115.0 8.881784197e-13 42185.0 ;
      RECT  4035.0 41295.0 0.0 41365.0 ;
      RECT  16785.0 45190.0 16650.0 45260.0 ;
      RECT  4035.0 45190.0 3900.0 45260.0 ;
      RECT  16580.0 46150.0 16445.0 46220.0 ;
      RECT  4035.0 46150.0 3900.0 46220.0 ;
      RECT  16170.0 43820.0 16035.0 43890.0 ;
      RECT  4035.0 43820.0 3900.0 43890.0 ;
      RECT  15965.0 44965.0 15830.0 45035.0 ;
      RECT  4035.0 44965.0 3900.0 45035.0 ;
      RECT  16375.0 42525.0 16240.0 42595.0 ;
      RECT  4035.0 42525.0 3900.0 42595.0 ;
      RECT  15760.0 41090.0 15625.0 41160.0 ;
      RECT  4035.0 41090.0 3900.0 41160.0 ;
      RECT  4417.5 42115.0 4282.5 42185.0 ;
      RECT  15345.0 41295.0 15210.0 41365.0 ;
      RECT  4035.0 41295.0 3900.0 41365.0 ;
   LAYER  metal3 ;
      RECT  4035.0 45190.0 16717.5 45260.0 ;
      RECT  4035.0 46150.0 16512.5 46220.0 ;
      RECT  4035.0 43820.0 16102.5 43890.0 ;
      RECT  4035.0 44965.0 15897.5 45035.0 ;
      RECT  4035.0 42525.0 16307.5 42595.0 ;
      RECT  4035.0 41090.0 15692.5 41160.0 ;
      RECT  4035.0 41295.0 15277.5 41365.0 ;
      RECT  17302.5 31150.0 17372.5 31220.0 ;
      RECT  17302.5 12640.0 17372.5 31185.0 ;
      RECT  17337.5 31150.0 17507.5 31220.0 ;
      RECT  20122.5 31150.0 20192.5 31220.0 ;
      RECT  20122.5 12640.0 20192.5 31185.0 ;
      RECT  20157.5 31150.0 20327.5 31220.0 ;
      RECT  22942.5 31150.0 23012.5 31220.0 ;
      RECT  22942.5 12640.0 23012.5 31185.0 ;
      RECT  22977.5 31150.0 23147.5 31220.0 ;
      RECT  25762.5 31150.0 25832.5 31220.0 ;
      RECT  25762.5 12640.0 25832.5 31185.0 ;
      RECT  25797.5 31150.0 25967.5 31220.0 ;
      RECT  28582.5 31150.0 28652.5 31220.0 ;
      RECT  28582.5 12640.0 28652.5 31185.0 ;
      RECT  28617.5 31150.0 28787.5 31220.0 ;
      RECT  31402.5 31150.0 31472.5 31220.0 ;
      RECT  31402.5 12640.0 31472.5 31185.0 ;
      RECT  31437.5 31150.0 31607.5 31220.0 ;
      RECT  34222.5 31150.0 34292.5 31220.0 ;
      RECT  34222.5 12640.0 34292.5 31185.0 ;
      RECT  34257.5 31150.0 34427.5 31220.0 ;
      RECT  37042.5 31150.0 37112.5 31220.0 ;
      RECT  37042.5 12640.0 37112.5 31185.0 ;
      RECT  37077.5 31150.0 37247.5 31220.0 ;
      RECT  39862.5 31150.0 39932.5 31220.0 ;
      RECT  39862.5 12640.0 39932.5 31185.0 ;
      RECT  39897.5 31150.0 40067.5 31220.0 ;
      RECT  42682.5 31150.0 42752.5 31220.0 ;
      RECT  42682.5 12640.0 42752.5 31185.0 ;
      RECT  42717.5 31150.0 42887.5 31220.0 ;
      RECT  45502.5 31150.0 45572.5 31220.0 ;
      RECT  45502.5 12640.0 45572.5 31185.0 ;
      RECT  45537.5 31150.0 45707.5 31220.0 ;
      RECT  48322.5 31150.0 48392.5 31220.0 ;
      RECT  48322.5 12640.0 48392.5 31185.0 ;
      RECT  48357.5 31150.0 48527.5 31220.0 ;
      RECT  51142.5 31150.0 51212.5 31220.0 ;
      RECT  51142.5 12640.0 51212.5 31185.0 ;
      RECT  51177.5 31150.0 51347.5 31220.0 ;
      RECT  53962.5 31150.0 54032.5 31220.0 ;
      RECT  53962.5 12640.0 54032.5 31185.0 ;
      RECT  53997.5 31150.0 54167.5 31220.0 ;
      RECT  56782.5 31150.0 56852.5 31220.0 ;
      RECT  56782.5 12640.0 56852.5 31185.0 ;
      RECT  56817.5 31150.0 56987.5 31220.0 ;
      RECT  59602.5 31150.0 59672.5 31220.0 ;
      RECT  59602.5 12640.0 59672.5 31185.0 ;
      RECT  59637.5 31150.0 59807.5 31220.0 ;
      RECT  62422.5 31150.0 62492.5 31220.0 ;
      RECT  62422.5 12640.0 62492.5 31185.0 ;
      RECT  62457.5 31150.0 62627.5 31220.0 ;
      RECT  65242.5 31150.0 65312.5 31220.0 ;
      RECT  65242.5 12640.0 65312.5 31185.0 ;
      RECT  65277.5 31150.0 65447.5 31220.0 ;
      RECT  68062.5 31150.0 68132.5 31220.0 ;
      RECT  68062.5 12640.0 68132.5 31185.0 ;
      RECT  68097.5 31150.0 68267.5 31220.0 ;
      RECT  70882.5 31150.0 70952.5 31220.0 ;
      RECT  70882.5 12640.0 70952.5 31185.0 ;
      RECT  70917.5 31150.0 71087.5 31220.0 ;
      RECT  73702.5 31150.0 73772.5 31220.0 ;
      RECT  73702.5 12640.0 73772.5 31185.0 ;
      RECT  73737.5 31150.0 73907.5 31220.0 ;
      RECT  76522.5 31150.0 76592.5 31220.0 ;
      RECT  76522.5 12640.0 76592.5 31185.0 ;
      RECT  76557.5 31150.0 76727.5 31220.0 ;
      RECT  79342.5 31150.0 79412.5 31220.0 ;
      RECT  79342.5 12640.0 79412.5 31185.0 ;
      RECT  79377.5 31150.0 79547.5 31220.0 ;
      RECT  82162.5 31150.0 82232.5 31220.0 ;
      RECT  82162.5 12640.0 82232.5 31185.0 ;
      RECT  82197.5 31150.0 82367.5 31220.0 ;
      RECT  84982.5 31150.0 85052.5 31220.0 ;
      RECT  84982.5 12640.0 85052.5 31185.0 ;
      RECT  85017.5 31150.0 85187.5 31220.0 ;
      RECT  87802.5 31150.0 87872.5 31220.0 ;
      RECT  87802.5 12640.0 87872.5 31185.0 ;
      RECT  87837.5 31150.0 88007.5 31220.0 ;
      RECT  90622.5 31150.0 90692.5 31220.0 ;
      RECT  90622.5 12640.0 90692.5 31185.0 ;
      RECT  90657.5 31150.0 90827.5 31220.0 ;
      RECT  93442.5 31150.0 93512.5 31220.0 ;
      RECT  93442.5 12640.0 93512.5 31185.0 ;
      RECT  93477.5 31150.0 93647.5 31220.0 ;
      RECT  96262.5 31150.0 96332.5 31220.0 ;
      RECT  96262.5 12640.0 96332.5 31185.0 ;
      RECT  96297.5 31150.0 96467.5 31220.0 ;
      RECT  99082.5 31150.0 99152.5 31220.0 ;
      RECT  99082.5 12640.0 99152.5 31185.0 ;
      RECT  99117.5 31150.0 99287.5 31220.0 ;
      RECT  101902.5 31150.0 101972.5 31220.0 ;
      RECT  101902.5 12640.0 101972.5 31185.0 ;
      RECT  101937.5 31150.0 102107.5 31220.0 ;
      RECT  104722.5 31150.0 104792.5 31220.0 ;
      RECT  104722.5 12640.0 104792.5 31185.0 ;
      RECT  104757.5 31150.0 104927.5 31220.0 ;
      RECT  17512.5 35.0 17582.5 15755.0 ;
      RECT  20332.5 35.0 20402.5 15755.0 ;
      RECT  23152.5 35.0 23222.5 15755.0 ;
      RECT  25972.5 35.0 26042.5 15755.0 ;
      RECT  28792.5 35.0 28862.5 15755.0 ;
      RECT  31612.5 35.0 31682.5 15755.0 ;
      RECT  34432.5 35.0 34502.5 15755.0 ;
      RECT  37252.5 35.0 37322.5 15755.0 ;
      RECT  40072.5 35.0 40142.5 15755.0 ;
      RECT  42892.5 35.0 42962.5 15755.0 ;
      RECT  45712.5 35.0 45782.5 15755.0 ;
      RECT  48532.5 35.0 48602.5 15755.0 ;
      RECT  51352.5 35.0 51422.5 15755.0 ;
      RECT  54172.5 35.0 54242.5 15755.0 ;
      RECT  56992.5 35.0 57062.5 15755.0 ;
      RECT  59812.5 35.0 59882.5 15755.0 ;
      RECT  62632.5 35.0 62702.5 15755.0 ;
      RECT  65452.5 35.0 65522.5 15755.0 ;
      RECT  68272.5 35.0 68342.5 15755.0 ;
      RECT  71092.5 35.0 71162.5 15755.0 ;
      RECT  73912.5 35.0 73982.5 15755.0 ;
      RECT  76732.5 35.0 76802.5 15755.0 ;
      RECT  79552.5 35.0 79622.5 15755.0 ;
      RECT  82372.5 35.0 82442.5 15755.0 ;
      RECT  85192.5 35.0 85262.5 15755.0 ;
      RECT  88012.5 35.0 88082.5 15755.0 ;
      RECT  90832.5 35.0 90902.5 15755.0 ;
      RECT  93652.5 35.0 93722.5 15755.0 ;
      RECT  96472.5 35.0 96542.5 15755.0 ;
      RECT  99292.5 35.0 99362.5 15755.0 ;
      RECT  102112.5 35.0 102182.5 15755.0 ;
      RECT  104932.5 35.0 105002.5 15755.0 ;
      RECT  12472.5 12545.0 15102.5 12615.0 ;
      RECT  12472.5 15235.0 15102.5 15305.0 ;
      RECT  12472.5 17925.0 15102.5 17995.0 ;
      RECT  12472.5 20615.0 15102.5 20685.0 ;
      RECT  12472.5 23305.0 15102.5 23375.0 ;
      RECT  12472.5 25995.0 15102.5 26065.0 ;
      RECT  12472.5 28685.0 15102.5 28755.0 ;
      RECT  12472.5 31375.0 15102.5 31445.0 ;
      RECT  7960.0 6847.5 8030.0 6917.5 ;
      RECT  7995.0 6847.5 11095.0 6917.5 ;
      RECT  7960.0 5275.0 8030.0 6882.5 ;
      RECT  8235.0 6142.5 8305.0 6212.5 ;
      RECT  8270.0 6142.5 11095.0 6212.5 ;
      RECT  8235.0 5275.0 8305.0 6177.5 ;
      RECT  17507.5 31115.0 17577.5 31255.0 ;
      RECT  20327.5 31115.0 20397.5 31255.0 ;
      RECT  23147.5 31115.0 23217.5 31255.0 ;
      RECT  25967.5 31115.0 26037.5 31255.0 ;
      RECT  28787.5 31115.0 28857.5 31255.0 ;
      RECT  31607.5 31115.0 31677.5 31255.0 ;
      RECT  34427.5 31115.0 34497.5 31255.0 ;
      RECT  37247.5 31115.0 37317.5 31255.0 ;
      RECT  40067.5 31115.0 40137.5 31255.0 ;
      RECT  42887.5 31115.0 42957.5 31255.0 ;
      RECT  45707.5 31115.0 45777.5 31255.0 ;
      RECT  48527.5 31115.0 48597.5 31255.0 ;
      RECT  51347.5 31115.0 51417.5 31255.0 ;
      RECT  54167.5 31115.0 54237.5 31255.0 ;
      RECT  56987.5 31115.0 57057.5 31255.0 ;
      RECT  59807.5 31115.0 59877.5 31255.0 ;
      RECT  62627.5 31115.0 62697.5 31255.0 ;
      RECT  65447.5 31115.0 65517.5 31255.0 ;
      RECT  68267.5 31115.0 68337.5 31255.0 ;
      RECT  71087.5 31115.0 71157.5 31255.0 ;
      RECT  73907.5 31115.0 73977.5 31255.0 ;
      RECT  76727.5 31115.0 76797.5 31255.0 ;
      RECT  79547.5 31115.0 79617.5 31255.0 ;
      RECT  82367.5 31115.0 82437.5 31255.0 ;
      RECT  85187.5 31115.0 85257.5 31255.0 ;
      RECT  88007.5 31115.0 88077.5 31255.0 ;
      RECT  90827.5 31115.0 90897.5 31255.0 ;
      RECT  93647.5 31115.0 93717.5 31255.0 ;
      RECT  96467.5 31115.0 96537.5 31255.0 ;
      RECT  99287.5 31115.0 99357.5 31255.0 ;
      RECT  102107.5 31115.0 102177.5 31255.0 ;
      RECT  104927.5 31115.0 104997.5 31255.0 ;
      RECT  17512.5 15755.0 17582.5 15895.0 ;
      RECT  20332.5 15755.0 20402.5 15895.0 ;
      RECT  23152.5 15755.0 23222.5 15895.0 ;
      RECT  25972.5 15755.0 26042.5 15895.0 ;
      RECT  28792.5 15755.0 28862.5 15895.0 ;
      RECT  31612.5 15755.0 31682.5 15895.0 ;
      RECT  34432.5 15755.0 34502.5 15895.0 ;
      RECT  37252.5 15755.0 37322.5 15895.0 ;
      RECT  40072.5 15755.0 40142.5 15895.0 ;
      RECT  42892.5 15755.0 42962.5 15895.0 ;
      RECT  45712.5 15755.0 45782.5 15895.0 ;
      RECT  48532.5 15755.0 48602.5 15895.0 ;
      RECT  51352.5 15755.0 51422.5 15895.0 ;
      RECT  54172.5 15755.0 54242.5 15895.0 ;
      RECT  56992.5 15755.0 57062.5 15895.0 ;
      RECT  59812.5 15755.0 59882.5 15895.0 ;
      RECT  62632.5 15755.0 62702.5 15895.0 ;
      RECT  65452.5 15755.0 65522.5 15895.0 ;
      RECT  68272.5 15755.0 68342.5 15895.0 ;
      RECT  71092.5 15755.0 71162.5 15895.0 ;
      RECT  73912.5 15755.0 73982.5 15895.0 ;
      RECT  76732.5 15755.0 76802.5 15895.0 ;
      RECT  79552.5 15755.0 79622.5 15895.0 ;
      RECT  82372.5 15755.0 82442.5 15895.0 ;
      RECT  85192.5 15755.0 85262.5 15895.0 ;
      RECT  88012.5 15755.0 88082.5 15895.0 ;
      RECT  90832.5 15755.0 90902.5 15895.0 ;
      RECT  93652.5 15755.0 93722.5 15895.0 ;
      RECT  96472.5 15755.0 96542.5 15895.0 ;
      RECT  99292.5 15755.0 99362.5 15895.0 ;
      RECT  102112.5 15755.0 102182.5 15895.0 ;
      RECT  104932.5 15755.0 105002.5 15895.0 ;
      RECT  4655.0 11852.5 4795.0 11782.5 ;
      RECT  4655.0 11147.5 4795.0 11077.5 ;
      RECT  4655.0 10442.5 4795.0 10372.5 ;
      RECT  4655.0 9737.5 4795.0 9667.5 ;
      RECT  4655.0 9032.5 4795.0 8962.5 ;
      RECT  4655.0 8327.5 4795.0 8257.5 ;
      RECT  4655.0 7622.5 4795.0 7552.5 ;
      RECT  4655.0 6917.5 4795.0 6847.5 ;
      RECT  4655.0 6212.5 4795.0 6142.5 ;
      RECT  17302.5 12605.0 17372.5 12740.0 ;
      RECT  20122.5 12605.0 20192.5 12740.0 ;
      RECT  22942.5 12605.0 23012.5 12740.0 ;
      RECT  25762.5 12605.0 25832.5 12740.0 ;
      RECT  28582.5 12605.0 28652.5 12740.0 ;
      RECT  31402.5 12605.0 31472.5 12740.0 ;
      RECT  34222.5 12605.0 34292.5 12740.0 ;
      RECT  37042.5 12605.0 37112.5 12740.0 ;
      RECT  39862.5 12605.0 39932.5 12740.0 ;
      RECT  42682.5 12605.0 42752.5 12740.0 ;
      RECT  45502.5 12605.0 45572.5 12740.0 ;
      RECT  48322.5 12605.0 48392.5 12740.0 ;
      RECT  51142.5 12605.0 51212.5 12740.0 ;
      RECT  53962.5 12605.0 54032.5 12740.0 ;
      RECT  56782.5 12605.0 56852.5 12740.0 ;
      RECT  59602.5 12605.0 59672.5 12740.0 ;
      RECT  62422.5 12605.0 62492.5 12740.0 ;
      RECT  65242.5 12605.0 65312.5 12740.0 ;
      RECT  68062.5 12605.0 68132.5 12740.0 ;
      RECT  70882.5 12605.0 70952.5 12740.0 ;
      RECT  73702.5 12605.0 73772.5 12740.0 ;
      RECT  76522.5 12605.0 76592.5 12740.0 ;
      RECT  79342.5 12605.0 79412.5 12740.0 ;
      RECT  82162.5 12605.0 82232.5 12740.0 ;
      RECT  84982.5 12605.0 85052.5 12740.0 ;
      RECT  87802.5 12605.0 87872.5 12740.0 ;
      RECT  90622.5 12605.0 90692.5 12740.0 ;
      RECT  93442.5 12605.0 93512.5 12740.0 ;
      RECT  96262.5 12605.0 96332.5 12740.0 ;
      RECT  99082.5 12605.0 99152.5 12740.0 ;
      RECT  101902.5 12605.0 101972.5 12740.0 ;
      RECT  104722.5 12605.0 104792.5 12740.0 ;
      RECT  17512.5 35.0 17582.5 170.0 ;
      RECT  20332.5 35.0 20402.5 170.0 ;
      RECT  23152.5 35.0 23222.5 170.0 ;
      RECT  25972.5 35.0 26042.5 170.0 ;
      RECT  28792.5 35.0 28862.5 170.0 ;
      RECT  31612.5 35.0 31682.5 170.0 ;
      RECT  34432.5 35.0 34502.5 170.0 ;
      RECT  37252.5 35.0 37322.5 170.0 ;
      RECT  40072.5 35.0 40142.5 170.0 ;
      RECT  42892.5 35.0 42962.5 170.0 ;
      RECT  45712.5 35.0 45782.5 170.0 ;
      RECT  48532.5 35.0 48602.5 170.0 ;
      RECT  51352.5 35.0 51422.5 170.0 ;
      RECT  54172.5 35.0 54242.5 170.0 ;
      RECT  56992.5 35.0 57062.5 170.0 ;
      RECT  59812.5 35.0 59882.5 170.0 ;
      RECT  62632.5 35.0 62702.5 170.0 ;
      RECT  65452.5 35.0 65522.5 170.0 ;
      RECT  68272.5 35.0 68342.5 170.0 ;
      RECT  71092.5 35.0 71162.5 170.0 ;
      RECT  73912.5 35.0 73982.5 170.0 ;
      RECT  76732.5 35.0 76802.5 170.0 ;
      RECT  79552.5 35.0 79622.5 170.0 ;
      RECT  82372.5 35.0 82442.5 170.0 ;
      RECT  85192.5 35.0 85262.5 170.0 ;
      RECT  88012.5 35.0 88082.5 170.0 ;
      RECT  90832.5 35.0 90902.5 170.0 ;
      RECT  93652.5 35.0 93722.5 170.0 ;
      RECT  96472.5 35.0 96542.5 170.0 ;
      RECT  99292.5 35.0 99362.5 170.0 ;
      RECT  102112.5 35.0 102182.5 170.0 ;
      RECT  104932.5 35.0 105002.5 170.0 ;
      RECT  12540.0 12545.0 12405.0 12615.0 ;
      RECT  15035.0 12615.0 15170.0 12545.0 ;
      RECT  12540.0 15235.0 12405.0 15305.0 ;
      RECT  15035.0 15305.0 15170.0 15235.0 ;
      RECT  12540.0 17925.0 12405.0 17995.0 ;
      RECT  15035.0 17995.0 15170.0 17925.0 ;
      RECT  12540.0 20615.0 12405.0 20685.0 ;
      RECT  15035.0 20685.0 15170.0 20615.0 ;
      RECT  12540.0 23305.0 12405.0 23375.0 ;
      RECT  15035.0 23375.0 15170.0 23305.0 ;
      RECT  12540.0 25995.0 12405.0 26065.0 ;
      RECT  15035.0 26065.0 15170.0 25995.0 ;
      RECT  12540.0 28685.0 12405.0 28755.0 ;
      RECT  15035.0 28755.0 15170.0 28685.0 ;
      RECT  12540.0 31375.0 12405.0 31445.0 ;
      RECT  15035.0 31445.0 15170.0 31375.0 ;
      RECT  11162.5 6847.5 11027.5 6917.5 ;
      RECT  7960.0 5207.5 8030.0 5342.5 ;
      RECT  11162.5 6142.5 11027.5 6212.5 ;
      RECT  8235.0 5207.5 8305.0 5342.5 ;
      RECT  4175.0 11782.5 4655.0 11852.5 ;
      RECT  4175.0 11077.5 4655.0 11147.5 ;
      RECT  4175.0 10372.5 4655.0 10442.5 ;
      RECT  4175.0 9667.5 4655.0 9737.5 ;
      RECT  4175.0 8962.5 4655.0 9032.5 ;
      RECT  4175.0 8257.5 4655.0 8327.5 ;
      RECT  4175.0 7552.5 4655.0 7622.5 ;
      RECT  4175.0 6847.5 4655.0 6917.5 ;
      RECT  4175.0 6142.5 4655.0 6212.5 ;
      RECT  397.5 40680.0 327.5 42355.0 ;
      RECT  552.5 40680.0 482.5 41535.0 ;
      RECT  1412.5 40680.0 1342.5 41740.0 ;
      RECT  1807.5 40680.0 1737.5 41945.0 ;
      RECT  200.0 40680.0 130.0 41330.0 ;
      RECT  905.0 40680.0 835.0 41330.0 ;
      RECT  1610.0 40680.0 1540.0 41330.0 ;
      RECT  2315.0 40680.0 2245.0 41330.0 ;
      RECT  2725.0 37045.0 2655.0 42560.0 ;
      RECT  2020.0 42560.0 1950.0 44072.5 ;
      RECT  1805.0 42355.0 1735.0 44330.0 ;
      RECT  482.5 34240.0 552.5 34380.0 ;
      RECT  1187.5 34240.0 1257.5 34380.0 ;
      RECT  1892.5 34240.0 1962.5 34380.0 ;
      RECT  397.5 40747.5 327.5 40612.5 ;
      RECT  397.5 42422.5 327.5 42287.5 ;
      RECT  552.5 40747.5 482.5 40612.5 ;
      RECT  552.5 41602.5 482.5 41467.5 ;
      RECT  1412.5 40747.5 1342.5 40612.5 ;
      RECT  1412.5 41807.5 1342.5 41672.5 ;
      RECT  1807.5 40747.5 1737.5 40612.5 ;
      RECT  1807.5 42012.5 1737.5 41877.5 ;
      RECT  200.0 40747.5 130.0 40612.5 ;
      RECT  200.0 41397.5 130.0 41262.5 ;
      RECT  905.0 40747.5 835.0 40612.5 ;
      RECT  905.0 41397.5 835.0 41262.5 ;
      RECT  1610.0 40747.5 1540.0 40612.5 ;
      RECT  1610.0 41397.5 1540.0 41262.5 ;
      RECT  2315.0 40747.5 2245.0 40612.5 ;
      RECT  2315.0 41397.5 2245.0 41262.5 ;
      RECT  2725.0 37112.5 2655.0 36977.5 ;
      RECT  2725.0 42627.5 2655.0 42492.5 ;
      RECT  2020.0 44140.0 1950.0 44005.0 ;
      RECT  2020.0 42627.5 1950.0 42492.5 ;
      RECT  1805.0 44397.5 1735.0 44262.5 ;
      RECT  1805.0 42422.5 1735.0 42287.5 ;
      RECT  1257.5 34240.0 1187.5 34380.0 ;
      RECT  1962.5 34240.0 1892.5 34380.0 ;
      RECT  552.5 34240.0 482.5 34380.0 ;
      RECT  16785.0 45190.0 16650.0 45260.0 ;
      RECT  4035.0 45190.0 3900.0 45260.0 ;
      RECT  16580.0 46150.0 16445.0 46220.0 ;
      RECT  4035.0 46150.0 3900.0 46220.0 ;
      RECT  16170.0 43820.0 16035.0 43890.0 ;
      RECT  4035.0 43820.0 3900.0 43890.0 ;
      RECT  15965.0 44965.0 15830.0 45035.0 ;
      RECT  4035.0 44965.0 3900.0 45035.0 ;
      RECT  16375.0 42525.0 16240.0 42595.0 ;
      RECT  4035.0 42525.0 3900.0 42595.0 ;
      RECT  15760.0 41090.0 15625.0 41160.0 ;
      RECT  4035.0 41090.0 3900.0 41160.0 ;
      RECT  15345.0 41295.0 15210.0 41365.0 ;
      RECT  4035.0 41295.0 3900.0 41365.0 ;
   END
   END    sram_1rw_32b_512w_1bank_freepdk45
END    LIBRARY
