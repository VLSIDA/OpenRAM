VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 1534200.0 by 2165400.0 ;
END  MacroSite
MACRO sram_1rw_32b_512w_1bank_scn3me_subm
   CLASS BLOCK ;
   SIZE 1534200.0 BY 2165400.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  225900.0 600.0 226800.0 2400.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  266700.0 600.0 267600.0 2400.0 ;
      END
   END DATA[1]
   PIN DATA[2]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  307500.0 600.0 308400.0 2400.0 ;
      END
   END DATA[2]
   PIN DATA[3]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  348300.0 600.0 349200.0 2400.0 ;
      END
   END DATA[3]
   PIN DATA[4]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  389100.0 600.0 390000.0 2400.0 ;
      END
   END DATA[4]
   PIN DATA[5]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  429900.0 600.0 430800.0 2400.0 ;
      END
   END DATA[5]
   PIN DATA[6]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  470700.0 600.0 471600.0 2400.0 ;
      END
   END DATA[6]
   PIN DATA[7]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  511500.0 600.0 512400.0 2400.0 ;
      END
   END DATA[7]
   PIN DATA[8]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  552300.0 600.0 553200.0 2400.0 ;
      END
   END DATA[8]
   PIN DATA[9]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  593100.0 600.0 594000.0 2400.0 ;
      END
   END DATA[9]
   PIN DATA[10]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  633900.0 600.0 634800.0 2400.0 ;
      END
   END DATA[10]
   PIN DATA[11]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  674700.0 600.0 675600.0 2400.0 ;
      END
   END DATA[11]
   PIN DATA[12]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  715500.0 600.0 716400.0 2400.0 ;
      END
   END DATA[12]
   PIN DATA[13]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  756300.0 600.0 757200.0 2400.0 ;
      END
   END DATA[13]
   PIN DATA[14]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  797100.0 600.0 798000.0 2400.0 ;
      END
   END DATA[14]
   PIN DATA[15]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  837900.0 600.0 838800.0 2400.0 ;
      END
   END DATA[15]
   PIN DATA[16]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  878700.0 600.0 879600.0 2400.0 ;
      END
   END DATA[16]
   PIN DATA[17]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  919500.0 600.0 920400.0 2400.0 ;
      END
   END DATA[17]
   PIN DATA[18]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  960300.0 600.0 961200.0 2400.0 ;
      END
   END DATA[18]
   PIN DATA[19]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1001100.0 600.0 1002000.0 2400.0 ;
      END
   END DATA[19]
   PIN DATA[20]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1041900.0 600.0 1042800.0 2400.0 ;
      END
   END DATA[20]
   PIN DATA[21]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1082700.0 600.0 1083600.0 2400.0 ;
      END
   END DATA[21]
   PIN DATA[22]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1123500.0 600.0 1124400.0 2400.0 ;
      END
   END DATA[22]
   PIN DATA[23]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1164300.0 600.0 1165200.0 2400.0 ;
      END
   END DATA[23]
   PIN DATA[24]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1205100.0 600.0 1206000.0 2400.0 ;
      END
   END DATA[24]
   PIN DATA[25]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1245900.0 600.0 1246800.0 2400.0 ;
      END
   END DATA[25]
   PIN DATA[26]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1286700.0 600.0 1287600.0 2400.0 ;
      END
   END DATA[26]
   PIN DATA[27]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1327500.0 600.0 1328400.0 2400.0 ;
      END
   END DATA[27]
   PIN DATA[28]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1368300.0 600.0 1369200.0 2400.0 ;
      END
   END DATA[28]
   PIN DATA[29]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1409100.0 600.0 1410000.0 2400.0 ;
      END
   END DATA[29]
   PIN DATA[30]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1449900.0 600.0 1450800.0 2400.0 ;
      END
   END DATA[30]
   PIN DATA[31]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  1490700.0 600.0 1491600.0 2400.0 ;
      END
   END DATA[31]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 147000.0 60000.0 148500.0 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 136800.0 60000.0 138300.0 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 126600.0 60000.0 128100.0 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 116400.0 60000.0 117900.0 ;
      END
   END ADDR[3]
   PIN ADDR[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 106200.0 60000.0 107700.0 ;
      END
   END ADDR[4]
   PIN ADDR[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 96000.0 60000.0 97500.0 ;
      END
   END ADDR[5]
   PIN ADDR[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 85800.0 60000.0 87300.0 ;
      END
   END ADDR[6]
   PIN ADDR[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 75600.0 60000.0 77100.0 ;
      END
   END ADDR[7]
   PIN ADDR[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 65400.0 60000.0 66900.0 ;
      END
   END ADDR[8]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14400.0 383100.0 16200.0 384900.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24600.0 383100.0 26400.0 384900.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4200.0 383100.0 6000.0 384900.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  42600.0 382200.0 43800.0 385800.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  1529700.0 600.0 1534200.0 2166000.0 ;
         LAYER metal1 ;
         RECT  52800.0 600.0 57300.0 2166000.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  193950.0 600.0 198450.0 2166000.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  54600.0 475650.0 55500.0 478350.0 ;
      RECT  115500.0 385350.0 116400.0 386250.0 ;
      RECT  115500.0 382950.0 116400.0 383850.0 ;
      RECT  114150.0 385350.0 115950.0 386250.0 ;
      RECT  115500.0 383400.0 116400.0 385800.0 ;
      RECT  115950.0 382950.0 117900.0 383850.0 ;
      RECT  186900.0 385350.0 187800.0 386250.0 ;
      RECT  186900.0 380850.0 187800.0 381750.0 ;
      RECT  154050.0 385350.0 187350.0 386250.0 ;
      RECT  186900.0 381300.0 187800.0 385800.0 ;
      RECT  187350.0 380850.0 220800.0 381750.0 ;
      RECT  115500.0 399750.0 116400.0 400650.0 ;
      RECT  115500.0 402150.0 116400.0 403050.0 ;
      RECT  114150.0 399750.0 115950.0 400650.0 ;
      RECT  115500.0 400200.0 116400.0 402600.0 ;
      RECT  115950.0 402150.0 117900.0 403050.0 ;
      RECT  186900.0 399750.0 187800.0 400650.0 ;
      RECT  186900.0 404250.0 187800.0 405150.0 ;
      RECT  154050.0 399750.0 187350.0 400650.0 ;
      RECT  186900.0 400200.0 187800.0 404700.0 ;
      RECT  187350.0 404250.0 220800.0 405150.0 ;
      RECT  115500.0 412950.0 116400.0 413850.0 ;
      RECT  115500.0 410550.0 116400.0 411450.0 ;
      RECT  114150.0 412950.0 115950.0 413850.0 ;
      RECT  115500.0 411000.0 116400.0 413400.0 ;
      RECT  115950.0 410550.0 117900.0 411450.0 ;
      RECT  186900.0 412950.0 187800.0 413850.0 ;
      RECT  186900.0 408450.0 187800.0 409350.0 ;
      RECT  154050.0 412950.0 187350.0 413850.0 ;
      RECT  186900.0 408900.0 187800.0 413400.0 ;
      RECT  187350.0 408450.0 220800.0 409350.0 ;
      RECT  115500.0 427350.0 116400.0 428250.0 ;
      RECT  115500.0 429750.0 116400.0 430650.0 ;
      RECT  114150.0 427350.0 115950.0 428250.0 ;
      RECT  115500.0 427800.0 116400.0 430200.0 ;
      RECT  115950.0 429750.0 117900.0 430650.0 ;
      RECT  186900.0 427350.0 187800.0 428250.0 ;
      RECT  186900.0 431850.0 187800.0 432750.0 ;
      RECT  154050.0 427350.0 187350.0 428250.0 ;
      RECT  186900.0 427800.0 187800.0 432300.0 ;
      RECT  187350.0 431850.0 220800.0 432750.0 ;
      RECT  115500.0 440550.0 116400.0 441450.0 ;
      RECT  115500.0 438150.0 116400.0 439050.0 ;
      RECT  114150.0 440550.0 115950.0 441450.0 ;
      RECT  115500.0 438600.0 116400.0 441000.0 ;
      RECT  115950.0 438150.0 117900.0 439050.0 ;
      RECT  186900.0 440550.0 187800.0 441450.0 ;
      RECT  186900.0 436050.0 187800.0 436950.0 ;
      RECT  154050.0 440550.0 187350.0 441450.0 ;
      RECT  186900.0 436500.0 187800.0 441000.0 ;
      RECT  187350.0 436050.0 220800.0 436950.0 ;
      RECT  115500.0 454950.0 116400.0 455850.0 ;
      RECT  115500.0 457350.0 116400.0 458250.0 ;
      RECT  114150.0 454950.0 115950.0 455850.0 ;
      RECT  115500.0 455400.0 116400.0 457800.0 ;
      RECT  115950.0 457350.0 117900.0 458250.0 ;
      RECT  186900.0 454950.0 187800.0 455850.0 ;
      RECT  186900.0 459450.0 187800.0 460350.0 ;
      RECT  154050.0 454950.0 187350.0 455850.0 ;
      RECT  186900.0 455400.0 187800.0 459900.0 ;
      RECT  187350.0 459450.0 220800.0 460350.0 ;
      RECT  115500.0 468150.0 116400.0 469050.0 ;
      RECT  115500.0 465750.0 116400.0 466650.0 ;
      RECT  114150.0 468150.0 115950.0 469050.0 ;
      RECT  115500.0 466200.0 116400.0 468600.0 ;
      RECT  115950.0 465750.0 117900.0 466650.0 ;
      RECT  186900.0 468150.0 187800.0 469050.0 ;
      RECT  186900.0 463650.0 187800.0 464550.0 ;
      RECT  154050.0 468150.0 187350.0 469050.0 ;
      RECT  186900.0 464100.0 187800.0 468600.0 ;
      RECT  187350.0 463650.0 220800.0 464550.0 ;
      RECT  115500.0 482550.0 116400.0 483450.0 ;
      RECT  115500.0 484950.0 116400.0 485850.0 ;
      RECT  114150.0 482550.0 115950.0 483450.0 ;
      RECT  115500.0 483000.0 116400.0 485400.0 ;
      RECT  115950.0 484950.0 117900.0 485850.0 ;
      RECT  186900.0 482550.0 187800.0 483450.0 ;
      RECT  186900.0 487050.0 187800.0 487950.0 ;
      RECT  154050.0 482550.0 187350.0 483450.0 ;
      RECT  186900.0 483000.0 187800.0 487500.0 ;
      RECT  187350.0 487050.0 220800.0 487950.0 ;
      RECT  115500.0 495750.0 116400.0 496650.0 ;
      RECT  115500.0 493350.0 116400.0 494250.0 ;
      RECT  114150.0 495750.0 115950.0 496650.0 ;
      RECT  115500.0 493800.0 116400.0 496200.0 ;
      RECT  115950.0 493350.0 117900.0 494250.0 ;
      RECT  186900.0 495750.0 187800.0 496650.0 ;
      RECT  186900.0 491250.0 187800.0 492150.0 ;
      RECT  154050.0 495750.0 187350.0 496650.0 ;
      RECT  186900.0 491700.0 187800.0 496200.0 ;
      RECT  187350.0 491250.0 220800.0 492150.0 ;
      RECT  115500.0 510150.0 116400.0 511050.0 ;
      RECT  115500.0 512550.0 116400.0 513450.0 ;
      RECT  114150.0 510150.0 115950.0 511050.0 ;
      RECT  115500.0 510600.0 116400.0 513000.0 ;
      RECT  115950.0 512550.0 117900.0 513450.0 ;
      RECT  186900.0 510150.0 187800.0 511050.0 ;
      RECT  186900.0 514650.0 187800.0 515550.0 ;
      RECT  154050.0 510150.0 187350.0 511050.0 ;
      RECT  186900.0 510600.0 187800.0 515100.0 ;
      RECT  187350.0 514650.0 220800.0 515550.0 ;
      RECT  115500.0 523350.0 116400.0 524250.0 ;
      RECT  115500.0 520950.0 116400.0 521850.0 ;
      RECT  114150.0 523350.0 115950.0 524250.0 ;
      RECT  115500.0 521400.0 116400.0 523800.0 ;
      RECT  115950.0 520950.0 117900.0 521850.0 ;
      RECT  186900.0 523350.0 187800.0 524250.0 ;
      RECT  186900.0 518850.0 187800.0 519750.0 ;
      RECT  154050.0 523350.0 187350.0 524250.0 ;
      RECT  186900.0 519300.0 187800.0 523800.0 ;
      RECT  187350.0 518850.0 220800.0 519750.0 ;
      RECT  115500.0 537750.0 116400.0 538650.0 ;
      RECT  115500.0 540150.0 116400.0 541050.0 ;
      RECT  114150.0 537750.0 115950.0 538650.0 ;
      RECT  115500.0 538200.0 116400.0 540600.0 ;
      RECT  115950.0 540150.0 117900.0 541050.0 ;
      RECT  186900.0 537750.0 187800.0 538650.0 ;
      RECT  186900.0 542250.0 187800.0 543150.0 ;
      RECT  154050.0 537750.0 187350.0 538650.0 ;
      RECT  186900.0 538200.0 187800.0 542700.0 ;
      RECT  187350.0 542250.0 220800.0 543150.0 ;
      RECT  115500.0 550950.0 116400.0 551850.0 ;
      RECT  115500.0 548550.0 116400.0 549450.0 ;
      RECT  114150.0 550950.0 115950.0 551850.0 ;
      RECT  115500.0 549000.0 116400.0 551400.0 ;
      RECT  115950.0 548550.0 117900.0 549450.0 ;
      RECT  186900.0 550950.0 187800.0 551850.0 ;
      RECT  186900.0 546450.0 187800.0 547350.0 ;
      RECT  154050.0 550950.0 187350.0 551850.0 ;
      RECT  186900.0 546900.0 187800.0 551400.0 ;
      RECT  187350.0 546450.0 220800.0 547350.0 ;
      RECT  115500.0 565350.0 116400.0 566250.0 ;
      RECT  115500.0 567750.0 116400.0 568650.0 ;
      RECT  114150.0 565350.0 115950.0 566250.0 ;
      RECT  115500.0 565800.0 116400.0 568200.0 ;
      RECT  115950.0 567750.0 117900.0 568650.0 ;
      RECT  186900.0 565350.0 187800.0 566250.0 ;
      RECT  186900.0 569850.0 187800.0 570750.0 ;
      RECT  154050.0 565350.0 187350.0 566250.0 ;
      RECT  186900.0 565800.0 187800.0 570300.0 ;
      RECT  187350.0 569850.0 220800.0 570750.0 ;
      RECT  115500.0 578550.0 116400.0 579450.0 ;
      RECT  115500.0 576150.0 116400.0 577050.0 ;
      RECT  114150.0 578550.0 115950.0 579450.0 ;
      RECT  115500.0 576600.0 116400.0 579000.0 ;
      RECT  115950.0 576150.0 117900.0 577050.0 ;
      RECT  186900.0 578550.0 187800.0 579450.0 ;
      RECT  186900.0 574050.0 187800.0 574950.0 ;
      RECT  154050.0 578550.0 187350.0 579450.0 ;
      RECT  186900.0 574500.0 187800.0 579000.0 ;
      RECT  187350.0 574050.0 220800.0 574950.0 ;
      RECT  115500.0 592950.0 116400.0 593850.0 ;
      RECT  115500.0 595350.0 116400.0 596250.0 ;
      RECT  114150.0 592950.0 115950.0 593850.0 ;
      RECT  115500.0 593400.0 116400.0 595800.0 ;
      RECT  115950.0 595350.0 117900.0 596250.0 ;
      RECT  186900.0 592950.0 187800.0 593850.0 ;
      RECT  186900.0 597450.0 187800.0 598350.0 ;
      RECT  154050.0 592950.0 187350.0 593850.0 ;
      RECT  186900.0 593400.0 187800.0 597900.0 ;
      RECT  187350.0 597450.0 220800.0 598350.0 ;
      RECT  115500.0 606150.0 116400.0 607050.0 ;
      RECT  115500.0 603750.0 116400.0 604650.0 ;
      RECT  114150.0 606150.0 115950.0 607050.0 ;
      RECT  115500.0 604200.0 116400.0 606600.0 ;
      RECT  115950.0 603750.0 117900.0 604650.0 ;
      RECT  186900.0 606150.0 187800.0 607050.0 ;
      RECT  186900.0 601650.0 187800.0 602550.0 ;
      RECT  154050.0 606150.0 187350.0 607050.0 ;
      RECT  186900.0 602100.0 187800.0 606600.0 ;
      RECT  187350.0 601650.0 220800.0 602550.0 ;
      RECT  115500.0 620550.0 116400.0 621450.0 ;
      RECT  115500.0 622950.0 116400.0 623850.0 ;
      RECT  114150.0 620550.0 115950.0 621450.0 ;
      RECT  115500.0 621000.0 116400.0 623400.0 ;
      RECT  115950.0 622950.0 117900.0 623850.0 ;
      RECT  186900.0 620550.0 187800.0 621450.0 ;
      RECT  186900.0 625050.0 187800.0 625950.0 ;
      RECT  154050.0 620550.0 187350.0 621450.0 ;
      RECT  186900.0 621000.0 187800.0 625500.0 ;
      RECT  187350.0 625050.0 220800.0 625950.0 ;
      RECT  115500.0 633750.0 116400.0 634650.0 ;
      RECT  115500.0 631350.0 116400.0 632250.0 ;
      RECT  114150.0 633750.0 115950.0 634650.0 ;
      RECT  115500.0 631800.0 116400.0 634200.0 ;
      RECT  115950.0 631350.0 117900.0 632250.0 ;
      RECT  186900.0 633750.0 187800.0 634650.0 ;
      RECT  186900.0 629250.0 187800.0 630150.0 ;
      RECT  154050.0 633750.0 187350.0 634650.0 ;
      RECT  186900.0 629700.0 187800.0 634200.0 ;
      RECT  187350.0 629250.0 220800.0 630150.0 ;
      RECT  115500.0 648150.0 116400.0 649050.0 ;
      RECT  115500.0 650550.0 116400.0 651450.0 ;
      RECT  114150.0 648150.0 115950.0 649050.0 ;
      RECT  115500.0 648600.0 116400.0 651000.0 ;
      RECT  115950.0 650550.0 117900.0 651450.0 ;
      RECT  186900.0 648150.0 187800.0 649050.0 ;
      RECT  186900.0 652650.0 187800.0 653550.0 ;
      RECT  154050.0 648150.0 187350.0 649050.0 ;
      RECT  186900.0 648600.0 187800.0 653100.0 ;
      RECT  187350.0 652650.0 220800.0 653550.0 ;
      RECT  115500.0 661350.0 116400.0 662250.0 ;
      RECT  115500.0 658950.0 116400.0 659850.0 ;
      RECT  114150.0 661350.0 115950.0 662250.0 ;
      RECT  115500.0 659400.0 116400.0 661800.0 ;
      RECT  115950.0 658950.0 117900.0 659850.0 ;
      RECT  186900.0 661350.0 187800.0 662250.0 ;
      RECT  186900.0 656850.0 187800.0 657750.0 ;
      RECT  154050.0 661350.0 187350.0 662250.0 ;
      RECT  186900.0 657300.0 187800.0 661800.0 ;
      RECT  187350.0 656850.0 220800.0 657750.0 ;
      RECT  115500.0 675750.0 116400.0 676650.0 ;
      RECT  115500.0 678150.0 116400.0 679050.0 ;
      RECT  114150.0 675750.0 115950.0 676650.0 ;
      RECT  115500.0 676200.0 116400.0 678600.0 ;
      RECT  115950.0 678150.0 117900.0 679050.0 ;
      RECT  186900.0 675750.0 187800.0 676650.0 ;
      RECT  186900.0 680250.0 187800.0 681150.0 ;
      RECT  154050.0 675750.0 187350.0 676650.0 ;
      RECT  186900.0 676200.0 187800.0 680700.0 ;
      RECT  187350.0 680250.0 220800.0 681150.0 ;
      RECT  115500.0 688950.0 116400.0 689850.0 ;
      RECT  115500.0 686550.0 116400.0 687450.0 ;
      RECT  114150.0 688950.0 115950.0 689850.0 ;
      RECT  115500.0 687000.0 116400.0 689400.0 ;
      RECT  115950.0 686550.0 117900.0 687450.0 ;
      RECT  186900.0 688950.0 187800.0 689850.0 ;
      RECT  186900.0 684450.0 187800.0 685350.0 ;
      RECT  154050.0 688950.0 187350.0 689850.0 ;
      RECT  186900.0 684900.0 187800.0 689400.0 ;
      RECT  187350.0 684450.0 220800.0 685350.0 ;
      RECT  115500.0 703350.0 116400.0 704250.0 ;
      RECT  115500.0 705750.0 116400.0 706650.0 ;
      RECT  114150.0 703350.0 115950.0 704250.0 ;
      RECT  115500.0 703800.0 116400.0 706200.0 ;
      RECT  115950.0 705750.0 117900.0 706650.0 ;
      RECT  186900.0 703350.0 187800.0 704250.0 ;
      RECT  186900.0 707850.0 187800.0 708750.0 ;
      RECT  154050.0 703350.0 187350.0 704250.0 ;
      RECT  186900.0 703800.0 187800.0 708300.0 ;
      RECT  187350.0 707850.0 220800.0 708750.0 ;
      RECT  115500.0 716550.0 116400.0 717450.0 ;
      RECT  115500.0 714150.0 116400.0 715050.0 ;
      RECT  114150.0 716550.0 115950.0 717450.0 ;
      RECT  115500.0 714600.0 116400.0 717000.0 ;
      RECT  115950.0 714150.0 117900.0 715050.0 ;
      RECT  186900.0 716550.0 187800.0 717450.0 ;
      RECT  186900.0 712050.0 187800.0 712950.0 ;
      RECT  154050.0 716550.0 187350.0 717450.0 ;
      RECT  186900.0 712500.0 187800.0 717000.0 ;
      RECT  187350.0 712050.0 220800.0 712950.0 ;
      RECT  115500.0 730950.0 116400.0 731850.0 ;
      RECT  115500.0 733350.0 116400.0 734250.0 ;
      RECT  114150.0 730950.0 115950.0 731850.0 ;
      RECT  115500.0 731400.0 116400.0 733800.0 ;
      RECT  115950.0 733350.0 117900.0 734250.0 ;
      RECT  186900.0 730950.0 187800.0 731850.0 ;
      RECT  186900.0 735450.0 187800.0 736350.0 ;
      RECT  154050.0 730950.0 187350.0 731850.0 ;
      RECT  186900.0 731400.0 187800.0 735900.0 ;
      RECT  187350.0 735450.0 220800.0 736350.0 ;
      RECT  115500.0 744150.0 116400.0 745050.0 ;
      RECT  115500.0 741750.0 116400.0 742650.0 ;
      RECT  114150.0 744150.0 115950.0 745050.0 ;
      RECT  115500.0 742200.0 116400.0 744600.0 ;
      RECT  115950.0 741750.0 117900.0 742650.0 ;
      RECT  186900.0 744150.0 187800.0 745050.0 ;
      RECT  186900.0 739650.0 187800.0 740550.0 ;
      RECT  154050.0 744150.0 187350.0 745050.0 ;
      RECT  186900.0 740100.0 187800.0 744600.0 ;
      RECT  187350.0 739650.0 220800.0 740550.0 ;
      RECT  115500.0 758550.0 116400.0 759450.0 ;
      RECT  115500.0 760950.0 116400.0 761850.0 ;
      RECT  114150.0 758550.0 115950.0 759450.0 ;
      RECT  115500.0 759000.0 116400.0 761400.0 ;
      RECT  115950.0 760950.0 117900.0 761850.0 ;
      RECT  186900.0 758550.0 187800.0 759450.0 ;
      RECT  186900.0 763050.0 187800.0 763950.0 ;
      RECT  154050.0 758550.0 187350.0 759450.0 ;
      RECT  186900.0 759000.0 187800.0 763500.0 ;
      RECT  187350.0 763050.0 220800.0 763950.0 ;
      RECT  115500.0 771750.0 116400.0 772650.0 ;
      RECT  115500.0 769350.0 116400.0 770250.0 ;
      RECT  114150.0 771750.0 115950.0 772650.0 ;
      RECT  115500.0 769800.0 116400.0 772200.0 ;
      RECT  115950.0 769350.0 117900.0 770250.0 ;
      RECT  186900.0 771750.0 187800.0 772650.0 ;
      RECT  186900.0 767250.0 187800.0 768150.0 ;
      RECT  154050.0 771750.0 187350.0 772650.0 ;
      RECT  186900.0 767700.0 187800.0 772200.0 ;
      RECT  187350.0 767250.0 220800.0 768150.0 ;
      RECT  115500.0 786150.0 116400.0 787050.0 ;
      RECT  115500.0 788550.0 116400.0 789450.0 ;
      RECT  114150.0 786150.0 115950.0 787050.0 ;
      RECT  115500.0 786600.0 116400.0 789000.0 ;
      RECT  115950.0 788550.0 117900.0 789450.0 ;
      RECT  186900.0 786150.0 187800.0 787050.0 ;
      RECT  186900.0 790650.0 187800.0 791550.0 ;
      RECT  154050.0 786150.0 187350.0 787050.0 ;
      RECT  186900.0 786600.0 187800.0 791100.0 ;
      RECT  187350.0 790650.0 220800.0 791550.0 ;
      RECT  115500.0 799350.0 116400.0 800250.0 ;
      RECT  115500.0 796950.0 116400.0 797850.0 ;
      RECT  114150.0 799350.0 115950.0 800250.0 ;
      RECT  115500.0 797400.0 116400.0 799800.0 ;
      RECT  115950.0 796950.0 117900.0 797850.0 ;
      RECT  186900.0 799350.0 187800.0 800250.0 ;
      RECT  186900.0 794850.0 187800.0 795750.0 ;
      RECT  154050.0 799350.0 187350.0 800250.0 ;
      RECT  186900.0 795300.0 187800.0 799800.0 ;
      RECT  187350.0 794850.0 220800.0 795750.0 ;
      RECT  115500.0 813750.0 116400.0 814650.0 ;
      RECT  115500.0 816150.0 116400.0 817050.0 ;
      RECT  114150.0 813750.0 115950.0 814650.0 ;
      RECT  115500.0 814200.0 116400.0 816600.0 ;
      RECT  115950.0 816150.0 117900.0 817050.0 ;
      RECT  186900.0 813750.0 187800.0 814650.0 ;
      RECT  186900.0 818250.0 187800.0 819150.0 ;
      RECT  154050.0 813750.0 187350.0 814650.0 ;
      RECT  186900.0 814200.0 187800.0 818700.0 ;
      RECT  187350.0 818250.0 220800.0 819150.0 ;
      RECT  115500.0 826950.0 116400.0 827850.0 ;
      RECT  115500.0 824550.0 116400.0 825450.0 ;
      RECT  114150.0 826950.0 115950.0 827850.0 ;
      RECT  115500.0 825000.0 116400.0 827400.0 ;
      RECT  115950.0 824550.0 117900.0 825450.0 ;
      RECT  186900.0 826950.0 187800.0 827850.0 ;
      RECT  186900.0 822450.0 187800.0 823350.0 ;
      RECT  154050.0 826950.0 187350.0 827850.0 ;
      RECT  186900.0 822900.0 187800.0 827400.0 ;
      RECT  187350.0 822450.0 220800.0 823350.0 ;
      RECT  115500.0 841350.0 116400.0 842250.0 ;
      RECT  115500.0 843750.0 116400.0 844650.0 ;
      RECT  114150.0 841350.0 115950.0 842250.0 ;
      RECT  115500.0 841800.0 116400.0 844200.0 ;
      RECT  115950.0 843750.0 117900.0 844650.0 ;
      RECT  186900.0 841350.0 187800.0 842250.0 ;
      RECT  186900.0 845850.0 187800.0 846750.0 ;
      RECT  154050.0 841350.0 187350.0 842250.0 ;
      RECT  186900.0 841800.0 187800.0 846300.0 ;
      RECT  187350.0 845850.0 220800.0 846750.0 ;
      RECT  115500.0 854550.0 116400.0 855450.0 ;
      RECT  115500.0 852150.0 116400.0 853050.0 ;
      RECT  114150.0 854550.0 115950.0 855450.0 ;
      RECT  115500.0 852600.0 116400.0 855000.0 ;
      RECT  115950.0 852150.0 117900.0 853050.0 ;
      RECT  186900.0 854550.0 187800.0 855450.0 ;
      RECT  186900.0 850050.0 187800.0 850950.0 ;
      RECT  154050.0 854550.0 187350.0 855450.0 ;
      RECT  186900.0 850500.0 187800.0 855000.0 ;
      RECT  187350.0 850050.0 220800.0 850950.0 ;
      RECT  115500.0 868950.0 116400.0 869850.0 ;
      RECT  115500.0 871350.0 116400.0 872250.0 ;
      RECT  114150.0 868950.0 115950.0 869850.0 ;
      RECT  115500.0 869400.0 116400.0 871800.0 ;
      RECT  115950.0 871350.0 117900.0 872250.0 ;
      RECT  186900.0 868950.0 187800.0 869850.0 ;
      RECT  186900.0 873450.0 187800.0 874350.0 ;
      RECT  154050.0 868950.0 187350.0 869850.0 ;
      RECT  186900.0 869400.0 187800.0 873900.0 ;
      RECT  187350.0 873450.0 220800.0 874350.0 ;
      RECT  115500.0 882150.0 116400.0 883050.0 ;
      RECT  115500.0 879750.0 116400.0 880650.0 ;
      RECT  114150.0 882150.0 115950.0 883050.0 ;
      RECT  115500.0 880200.0 116400.0 882600.0 ;
      RECT  115950.0 879750.0 117900.0 880650.0 ;
      RECT  186900.0 882150.0 187800.0 883050.0 ;
      RECT  186900.0 877650.0 187800.0 878550.0 ;
      RECT  154050.0 882150.0 187350.0 883050.0 ;
      RECT  186900.0 878100.0 187800.0 882600.0 ;
      RECT  187350.0 877650.0 220800.0 878550.0 ;
      RECT  115500.0 896550.0 116400.0 897450.0 ;
      RECT  115500.0 898950.0 116400.0 899850.0 ;
      RECT  114150.0 896550.0 115950.0 897450.0 ;
      RECT  115500.0 897000.0 116400.0 899400.0 ;
      RECT  115950.0 898950.0 117900.0 899850.0 ;
      RECT  186900.0 896550.0 187800.0 897450.0 ;
      RECT  186900.0 901050.0 187800.0 901950.0 ;
      RECT  154050.0 896550.0 187350.0 897450.0 ;
      RECT  186900.0 897000.0 187800.0 901500.0 ;
      RECT  187350.0 901050.0 220800.0 901950.0 ;
      RECT  115500.0 909750.0 116400.0 910650.0 ;
      RECT  115500.0 907350.0 116400.0 908250.0 ;
      RECT  114150.0 909750.0 115950.0 910650.0 ;
      RECT  115500.0 907800.0 116400.0 910200.0 ;
      RECT  115950.0 907350.0 117900.0 908250.0 ;
      RECT  186900.0 909750.0 187800.0 910650.0 ;
      RECT  186900.0 905250.0 187800.0 906150.0 ;
      RECT  154050.0 909750.0 187350.0 910650.0 ;
      RECT  186900.0 905700.0 187800.0 910200.0 ;
      RECT  187350.0 905250.0 220800.0 906150.0 ;
      RECT  115500.0 924150.0 116400.0 925050.0 ;
      RECT  115500.0 926550.0 116400.0 927450.0 ;
      RECT  114150.0 924150.0 115950.0 925050.0 ;
      RECT  115500.0 924600.0 116400.0 927000.0 ;
      RECT  115950.0 926550.0 117900.0 927450.0 ;
      RECT  186900.0 924150.0 187800.0 925050.0 ;
      RECT  186900.0 928650.0 187800.0 929550.0 ;
      RECT  154050.0 924150.0 187350.0 925050.0 ;
      RECT  186900.0 924600.0 187800.0 929100.0 ;
      RECT  187350.0 928650.0 220800.0 929550.0 ;
      RECT  115500.0 937350.0 116400.0 938250.0 ;
      RECT  115500.0 934950.0 116400.0 935850.0 ;
      RECT  114150.0 937350.0 115950.0 938250.0 ;
      RECT  115500.0 935400.0 116400.0 937800.0 ;
      RECT  115950.0 934950.0 117900.0 935850.0 ;
      RECT  186900.0 937350.0 187800.0 938250.0 ;
      RECT  186900.0 932850.0 187800.0 933750.0 ;
      RECT  154050.0 937350.0 187350.0 938250.0 ;
      RECT  186900.0 933300.0 187800.0 937800.0 ;
      RECT  187350.0 932850.0 220800.0 933750.0 ;
      RECT  115500.0 951750.0 116400.0 952650.0 ;
      RECT  115500.0 954150.0 116400.0 955050.0 ;
      RECT  114150.0 951750.0 115950.0 952650.0 ;
      RECT  115500.0 952200.0 116400.0 954600.0 ;
      RECT  115950.0 954150.0 117900.0 955050.0 ;
      RECT  186900.0 951750.0 187800.0 952650.0 ;
      RECT  186900.0 956250.0 187800.0 957150.0 ;
      RECT  154050.0 951750.0 187350.0 952650.0 ;
      RECT  186900.0 952200.0 187800.0 956700.0 ;
      RECT  187350.0 956250.0 220800.0 957150.0 ;
      RECT  115500.0 964950.0 116400.0 965850.0 ;
      RECT  115500.0 962550.0 116400.0 963450.0 ;
      RECT  114150.0 964950.0 115950.0 965850.0 ;
      RECT  115500.0 963000.0 116400.0 965400.0 ;
      RECT  115950.0 962550.0 117900.0 963450.0 ;
      RECT  186900.0 964950.0 187800.0 965850.0 ;
      RECT  186900.0 960450.0 187800.0 961350.0 ;
      RECT  154050.0 964950.0 187350.0 965850.0 ;
      RECT  186900.0 960900.0 187800.0 965400.0 ;
      RECT  187350.0 960450.0 220800.0 961350.0 ;
      RECT  115500.0 979350.0 116400.0 980250.0 ;
      RECT  115500.0 981750.0 116400.0 982650.0 ;
      RECT  114150.0 979350.0 115950.0 980250.0 ;
      RECT  115500.0 979800.0 116400.0 982200.0 ;
      RECT  115950.0 981750.0 117900.0 982650.0 ;
      RECT  186900.0 979350.0 187800.0 980250.0 ;
      RECT  186900.0 983850.0 187800.0 984750.0 ;
      RECT  154050.0 979350.0 187350.0 980250.0 ;
      RECT  186900.0 979800.0 187800.0 984300.0 ;
      RECT  187350.0 983850.0 220800.0 984750.0 ;
      RECT  115500.0 992550.0 116400.0 993450.0 ;
      RECT  115500.0 990150.0 116400.0 991050.0 ;
      RECT  114150.0 992550.0 115950.0 993450.0 ;
      RECT  115500.0 990600.0 116400.0 993000.0 ;
      RECT  115950.0 990150.0 117900.0 991050.0 ;
      RECT  186900.0 992550.0 187800.0 993450.0 ;
      RECT  186900.0 988050.0 187800.0 988950.0 ;
      RECT  154050.0 992550.0 187350.0 993450.0 ;
      RECT  186900.0 988500.0 187800.0 993000.0 ;
      RECT  187350.0 988050.0 220800.0 988950.0 ;
      RECT  115500.0 1006950.0 116400.0 1007850.0 ;
      RECT  115500.0 1009350.0 116400.0 1010250.0 ;
      RECT  114150.0 1006950.0 115950.0 1007850.0 ;
      RECT  115500.0 1007400.0 116400.0 1009800.0 ;
      RECT  115950.0 1009350.0 117900.0 1010250.0 ;
      RECT  186900.0 1006950.0 187800.0 1007850.0 ;
      RECT  186900.0 1011450.0 187800.0 1012350.0 ;
      RECT  154050.0 1006950.0 187350.0 1007850.0 ;
      RECT  186900.0 1007400.0 187800.0 1011900.0 ;
      RECT  187350.0 1011450.0 220800.0 1012350.0 ;
      RECT  115500.0 1020150.0 116400.0 1021050.0 ;
      RECT  115500.0 1017750.0 116400.0 1018650.0 ;
      RECT  114150.0 1020150.0 115950.0 1021050.0 ;
      RECT  115500.0 1018200.0 116400.0 1020600.0 ;
      RECT  115950.0 1017750.0 117900.0 1018650.0 ;
      RECT  186900.0 1020150.0 187800.0 1021050.0 ;
      RECT  186900.0 1015650.0 187800.0 1016550.0 ;
      RECT  154050.0 1020150.0 187350.0 1021050.0 ;
      RECT  186900.0 1016100.0 187800.0 1020600.0 ;
      RECT  187350.0 1015650.0 220800.0 1016550.0 ;
      RECT  115500.0 1034550.0 116400.0 1035450.0 ;
      RECT  115500.0 1036950.0 116400.0 1037850.0 ;
      RECT  114150.0 1034550.0 115950.0 1035450.0 ;
      RECT  115500.0 1035000.0 116400.0 1037400.0 ;
      RECT  115950.0 1036950.0 117900.0 1037850.0 ;
      RECT  186900.0 1034550.0 187800.0 1035450.0 ;
      RECT  186900.0 1039050.0 187800.0 1039950.0 ;
      RECT  154050.0 1034550.0 187350.0 1035450.0 ;
      RECT  186900.0 1035000.0 187800.0 1039500.0 ;
      RECT  187350.0 1039050.0 220800.0 1039950.0 ;
      RECT  115500.0 1047750.0 116400.0 1048650.0 ;
      RECT  115500.0 1045350.0 116400.0 1046250.0 ;
      RECT  114150.0 1047750.0 115950.0 1048650.0 ;
      RECT  115500.0 1045800.0 116400.0 1048200.0 ;
      RECT  115950.0 1045350.0 117900.0 1046250.0 ;
      RECT  186900.0 1047750.0 187800.0 1048650.0 ;
      RECT  186900.0 1043250.0 187800.0 1044150.0 ;
      RECT  154050.0 1047750.0 187350.0 1048650.0 ;
      RECT  186900.0 1043700.0 187800.0 1048200.0 ;
      RECT  187350.0 1043250.0 220800.0 1044150.0 ;
      RECT  115500.0 1062150.0 116400.0 1063050.0 ;
      RECT  115500.0 1064550.0 116400.0 1065450.0 ;
      RECT  114150.0 1062150.0 115950.0 1063050.0 ;
      RECT  115500.0 1062600.0 116400.0 1065000.0 ;
      RECT  115950.0 1064550.0 117900.0 1065450.0 ;
      RECT  186900.0 1062150.0 187800.0 1063050.0 ;
      RECT  186900.0 1066650.0 187800.0 1067550.0 ;
      RECT  154050.0 1062150.0 187350.0 1063050.0 ;
      RECT  186900.0 1062600.0 187800.0 1067100.0 ;
      RECT  187350.0 1066650.0 220800.0 1067550.0 ;
      RECT  115500.0 1075350.0 116400.0 1076250.0 ;
      RECT  115500.0 1072950.0 116400.0 1073850.0 ;
      RECT  114150.0 1075350.0 115950.0 1076250.0 ;
      RECT  115500.0 1073400.0 116400.0 1075800.0 ;
      RECT  115950.0 1072950.0 117900.0 1073850.0 ;
      RECT  186900.0 1075350.0 187800.0 1076250.0 ;
      RECT  186900.0 1070850.0 187800.0 1071750.0 ;
      RECT  154050.0 1075350.0 187350.0 1076250.0 ;
      RECT  186900.0 1071300.0 187800.0 1075800.0 ;
      RECT  187350.0 1070850.0 220800.0 1071750.0 ;
      RECT  115500.0 1089750.0 116400.0 1090650.0 ;
      RECT  115500.0 1092150.0 116400.0 1093050.0 ;
      RECT  114150.0 1089750.0 115950.0 1090650.0 ;
      RECT  115500.0 1090200.0 116400.0 1092600.0 ;
      RECT  115950.0 1092150.0 117900.0 1093050.0 ;
      RECT  186900.0 1089750.0 187800.0 1090650.0 ;
      RECT  186900.0 1094250.0 187800.0 1095150.0 ;
      RECT  154050.0 1089750.0 187350.0 1090650.0 ;
      RECT  186900.0 1090200.0 187800.0 1094700.0 ;
      RECT  187350.0 1094250.0 220800.0 1095150.0 ;
      RECT  115500.0 1102950.0 116400.0 1103850.0 ;
      RECT  115500.0 1100550.0 116400.0 1101450.0 ;
      RECT  114150.0 1102950.0 115950.0 1103850.0 ;
      RECT  115500.0 1101000.0 116400.0 1103400.0 ;
      RECT  115950.0 1100550.0 117900.0 1101450.0 ;
      RECT  186900.0 1102950.0 187800.0 1103850.0 ;
      RECT  186900.0 1098450.0 187800.0 1099350.0 ;
      RECT  154050.0 1102950.0 187350.0 1103850.0 ;
      RECT  186900.0 1098900.0 187800.0 1103400.0 ;
      RECT  187350.0 1098450.0 220800.0 1099350.0 ;
      RECT  115500.0 1117350.0 116400.0 1118250.0 ;
      RECT  115500.0 1119750.0 116400.0 1120650.0 ;
      RECT  114150.0 1117350.0 115950.0 1118250.0 ;
      RECT  115500.0 1117800.0 116400.0 1120200.0 ;
      RECT  115950.0 1119750.0 117900.0 1120650.0 ;
      RECT  186900.0 1117350.0 187800.0 1118250.0 ;
      RECT  186900.0 1121850.0 187800.0 1122750.0 ;
      RECT  154050.0 1117350.0 187350.0 1118250.0 ;
      RECT  186900.0 1117800.0 187800.0 1122300.0 ;
      RECT  187350.0 1121850.0 220800.0 1122750.0 ;
      RECT  115500.0 1130550.0 116400.0 1131450.0 ;
      RECT  115500.0 1128150.0 116400.0 1129050.0 ;
      RECT  114150.0 1130550.0 115950.0 1131450.0 ;
      RECT  115500.0 1128600.0 116400.0 1131000.0 ;
      RECT  115950.0 1128150.0 117900.0 1129050.0 ;
      RECT  186900.0 1130550.0 187800.0 1131450.0 ;
      RECT  186900.0 1126050.0 187800.0 1126950.0 ;
      RECT  154050.0 1130550.0 187350.0 1131450.0 ;
      RECT  186900.0 1126500.0 187800.0 1131000.0 ;
      RECT  187350.0 1126050.0 220800.0 1126950.0 ;
      RECT  115500.0 1144950.0 116400.0 1145850.0 ;
      RECT  115500.0 1147350.0 116400.0 1148250.0 ;
      RECT  114150.0 1144950.0 115950.0 1145850.0 ;
      RECT  115500.0 1145400.0 116400.0 1147800.0 ;
      RECT  115950.0 1147350.0 117900.0 1148250.0 ;
      RECT  186900.0 1144950.0 187800.0 1145850.0 ;
      RECT  186900.0 1149450.0 187800.0 1150350.0 ;
      RECT  154050.0 1144950.0 187350.0 1145850.0 ;
      RECT  186900.0 1145400.0 187800.0 1149900.0 ;
      RECT  187350.0 1149450.0 220800.0 1150350.0 ;
      RECT  115500.0 1158150.0 116400.0 1159050.0 ;
      RECT  115500.0 1155750.0 116400.0 1156650.0 ;
      RECT  114150.0 1158150.0 115950.0 1159050.0 ;
      RECT  115500.0 1156200.0 116400.0 1158600.0 ;
      RECT  115950.0 1155750.0 117900.0 1156650.0 ;
      RECT  186900.0 1158150.0 187800.0 1159050.0 ;
      RECT  186900.0 1153650.0 187800.0 1154550.0 ;
      RECT  154050.0 1158150.0 187350.0 1159050.0 ;
      RECT  186900.0 1154100.0 187800.0 1158600.0 ;
      RECT  187350.0 1153650.0 220800.0 1154550.0 ;
      RECT  115500.0 1172550.0 116400.0 1173450.0 ;
      RECT  115500.0 1174950.0 116400.0 1175850.0 ;
      RECT  114150.0 1172550.0 115950.0 1173450.0 ;
      RECT  115500.0 1173000.0 116400.0 1175400.0 ;
      RECT  115950.0 1174950.0 117900.0 1175850.0 ;
      RECT  186900.0 1172550.0 187800.0 1173450.0 ;
      RECT  186900.0 1177050.0 187800.0 1177950.0 ;
      RECT  154050.0 1172550.0 187350.0 1173450.0 ;
      RECT  186900.0 1173000.0 187800.0 1177500.0 ;
      RECT  187350.0 1177050.0 220800.0 1177950.0 ;
      RECT  115500.0 1185750.0 116400.0 1186650.0 ;
      RECT  115500.0 1183350.0 116400.0 1184250.0 ;
      RECT  114150.0 1185750.0 115950.0 1186650.0 ;
      RECT  115500.0 1183800.0 116400.0 1186200.0 ;
      RECT  115950.0 1183350.0 117900.0 1184250.0 ;
      RECT  186900.0 1185750.0 187800.0 1186650.0 ;
      RECT  186900.0 1181250.0 187800.0 1182150.0 ;
      RECT  154050.0 1185750.0 187350.0 1186650.0 ;
      RECT  186900.0 1181700.0 187800.0 1186200.0 ;
      RECT  187350.0 1181250.0 220800.0 1182150.0 ;
      RECT  115500.0 1200150.0 116400.0 1201050.0 ;
      RECT  115500.0 1202550.0 116400.0 1203450.0 ;
      RECT  114150.0 1200150.0 115950.0 1201050.0 ;
      RECT  115500.0 1200600.0 116400.0 1203000.0 ;
      RECT  115950.0 1202550.0 117900.0 1203450.0 ;
      RECT  186900.0 1200150.0 187800.0 1201050.0 ;
      RECT  186900.0 1204650.0 187800.0 1205550.0 ;
      RECT  154050.0 1200150.0 187350.0 1201050.0 ;
      RECT  186900.0 1200600.0 187800.0 1205100.0 ;
      RECT  187350.0 1204650.0 220800.0 1205550.0 ;
      RECT  115500.0 1213350.0 116400.0 1214250.0 ;
      RECT  115500.0 1210950.0 116400.0 1211850.0 ;
      RECT  114150.0 1213350.0 115950.0 1214250.0 ;
      RECT  115500.0 1211400.0 116400.0 1213800.0 ;
      RECT  115950.0 1210950.0 117900.0 1211850.0 ;
      RECT  186900.0 1213350.0 187800.0 1214250.0 ;
      RECT  186900.0 1208850.0 187800.0 1209750.0 ;
      RECT  154050.0 1213350.0 187350.0 1214250.0 ;
      RECT  186900.0 1209300.0 187800.0 1213800.0 ;
      RECT  187350.0 1208850.0 220800.0 1209750.0 ;
      RECT  115500.0 1227750.0 116400.0 1228650.0 ;
      RECT  115500.0 1230150.0 116400.0 1231050.0 ;
      RECT  114150.0 1227750.0 115950.0 1228650.0 ;
      RECT  115500.0 1228200.0 116400.0 1230600.0 ;
      RECT  115950.0 1230150.0 117900.0 1231050.0 ;
      RECT  186900.0 1227750.0 187800.0 1228650.0 ;
      RECT  186900.0 1232250.0 187800.0 1233150.0 ;
      RECT  154050.0 1227750.0 187350.0 1228650.0 ;
      RECT  186900.0 1228200.0 187800.0 1232700.0 ;
      RECT  187350.0 1232250.0 220800.0 1233150.0 ;
      RECT  115500.0 1240950.0 116400.0 1241850.0 ;
      RECT  115500.0 1238550.0 116400.0 1239450.0 ;
      RECT  114150.0 1240950.0 115950.0 1241850.0 ;
      RECT  115500.0 1239000.0 116400.0 1241400.0 ;
      RECT  115950.0 1238550.0 117900.0 1239450.0 ;
      RECT  186900.0 1240950.0 187800.0 1241850.0 ;
      RECT  186900.0 1236450.0 187800.0 1237350.0 ;
      RECT  154050.0 1240950.0 187350.0 1241850.0 ;
      RECT  186900.0 1236900.0 187800.0 1241400.0 ;
      RECT  187350.0 1236450.0 220800.0 1237350.0 ;
      RECT  115500.0 1255350.0 116400.0 1256250.0 ;
      RECT  115500.0 1257750.0 116400.0 1258650.0 ;
      RECT  114150.0 1255350.0 115950.0 1256250.0 ;
      RECT  115500.0 1255800.0 116400.0 1258200.0 ;
      RECT  115950.0 1257750.0 117900.0 1258650.0 ;
      RECT  186900.0 1255350.0 187800.0 1256250.0 ;
      RECT  186900.0 1259850.0 187800.0 1260750.0 ;
      RECT  154050.0 1255350.0 187350.0 1256250.0 ;
      RECT  186900.0 1255800.0 187800.0 1260300.0 ;
      RECT  187350.0 1259850.0 220800.0 1260750.0 ;
      RECT  115500.0 1268550.0 116400.0 1269450.0 ;
      RECT  115500.0 1266150.0 116400.0 1267050.0 ;
      RECT  114150.0 1268550.0 115950.0 1269450.0 ;
      RECT  115500.0 1266600.0 116400.0 1269000.0 ;
      RECT  115950.0 1266150.0 117900.0 1267050.0 ;
      RECT  186900.0 1268550.0 187800.0 1269450.0 ;
      RECT  186900.0 1264050.0 187800.0 1264950.0 ;
      RECT  154050.0 1268550.0 187350.0 1269450.0 ;
      RECT  186900.0 1264500.0 187800.0 1269000.0 ;
      RECT  187350.0 1264050.0 220800.0 1264950.0 ;
      RECT  115500.0 1282950.0 116400.0 1283850.0 ;
      RECT  115500.0 1285350.0 116400.0 1286250.0 ;
      RECT  114150.0 1282950.0 115950.0 1283850.0 ;
      RECT  115500.0 1283400.0 116400.0 1285800.0 ;
      RECT  115950.0 1285350.0 117900.0 1286250.0 ;
      RECT  186900.0 1282950.0 187800.0 1283850.0 ;
      RECT  186900.0 1287450.0 187800.0 1288350.0 ;
      RECT  154050.0 1282950.0 187350.0 1283850.0 ;
      RECT  186900.0 1283400.0 187800.0 1287900.0 ;
      RECT  187350.0 1287450.0 220800.0 1288350.0 ;
      RECT  115500.0 1296150.0 116400.0 1297050.0 ;
      RECT  115500.0 1293750.0 116400.0 1294650.0 ;
      RECT  114150.0 1296150.0 115950.0 1297050.0 ;
      RECT  115500.0 1294200.0 116400.0 1296600.0 ;
      RECT  115950.0 1293750.0 117900.0 1294650.0 ;
      RECT  186900.0 1296150.0 187800.0 1297050.0 ;
      RECT  186900.0 1291650.0 187800.0 1292550.0 ;
      RECT  154050.0 1296150.0 187350.0 1297050.0 ;
      RECT  186900.0 1292100.0 187800.0 1296600.0 ;
      RECT  187350.0 1291650.0 220800.0 1292550.0 ;
      RECT  115500.0 1310550.0 116400.0 1311450.0 ;
      RECT  115500.0 1312950.0 116400.0 1313850.0 ;
      RECT  114150.0 1310550.0 115950.0 1311450.0 ;
      RECT  115500.0 1311000.0 116400.0 1313400.0 ;
      RECT  115950.0 1312950.0 117900.0 1313850.0 ;
      RECT  186900.0 1310550.0 187800.0 1311450.0 ;
      RECT  186900.0 1315050.0 187800.0 1315950.0 ;
      RECT  154050.0 1310550.0 187350.0 1311450.0 ;
      RECT  186900.0 1311000.0 187800.0 1315500.0 ;
      RECT  187350.0 1315050.0 220800.0 1315950.0 ;
      RECT  115500.0 1323750.0 116400.0 1324650.0 ;
      RECT  115500.0 1321350.0 116400.0 1322250.0 ;
      RECT  114150.0 1323750.0 115950.0 1324650.0 ;
      RECT  115500.0 1321800.0 116400.0 1324200.0 ;
      RECT  115950.0 1321350.0 117900.0 1322250.0 ;
      RECT  186900.0 1323750.0 187800.0 1324650.0 ;
      RECT  186900.0 1319250.0 187800.0 1320150.0 ;
      RECT  154050.0 1323750.0 187350.0 1324650.0 ;
      RECT  186900.0 1319700.0 187800.0 1324200.0 ;
      RECT  187350.0 1319250.0 220800.0 1320150.0 ;
      RECT  115500.0 1338150.0 116400.0 1339050.0 ;
      RECT  115500.0 1340550.0 116400.0 1341450.0 ;
      RECT  114150.0 1338150.0 115950.0 1339050.0 ;
      RECT  115500.0 1338600.0 116400.0 1341000.0 ;
      RECT  115950.0 1340550.0 117900.0 1341450.0 ;
      RECT  186900.0 1338150.0 187800.0 1339050.0 ;
      RECT  186900.0 1342650.0 187800.0 1343550.0 ;
      RECT  154050.0 1338150.0 187350.0 1339050.0 ;
      RECT  186900.0 1338600.0 187800.0 1343100.0 ;
      RECT  187350.0 1342650.0 220800.0 1343550.0 ;
      RECT  115500.0 1351350.0 116400.0 1352250.0 ;
      RECT  115500.0 1348950.0 116400.0 1349850.0 ;
      RECT  114150.0 1351350.0 115950.0 1352250.0 ;
      RECT  115500.0 1349400.0 116400.0 1351800.0 ;
      RECT  115950.0 1348950.0 117900.0 1349850.0 ;
      RECT  186900.0 1351350.0 187800.0 1352250.0 ;
      RECT  186900.0 1346850.0 187800.0 1347750.0 ;
      RECT  154050.0 1351350.0 187350.0 1352250.0 ;
      RECT  186900.0 1347300.0 187800.0 1351800.0 ;
      RECT  187350.0 1346850.0 220800.0 1347750.0 ;
      RECT  115500.0 1365750.0 116400.0 1366650.0 ;
      RECT  115500.0 1368150.0 116400.0 1369050.0 ;
      RECT  114150.0 1365750.0 115950.0 1366650.0 ;
      RECT  115500.0 1366200.0 116400.0 1368600.0 ;
      RECT  115950.0 1368150.0 117900.0 1369050.0 ;
      RECT  186900.0 1365750.0 187800.0 1366650.0 ;
      RECT  186900.0 1370250.0 187800.0 1371150.0 ;
      RECT  154050.0 1365750.0 187350.0 1366650.0 ;
      RECT  186900.0 1366200.0 187800.0 1370700.0 ;
      RECT  187350.0 1370250.0 220800.0 1371150.0 ;
      RECT  115500.0 1378950.0 116400.0 1379850.0 ;
      RECT  115500.0 1376550.0 116400.0 1377450.0 ;
      RECT  114150.0 1378950.0 115950.0 1379850.0 ;
      RECT  115500.0 1377000.0 116400.0 1379400.0 ;
      RECT  115950.0 1376550.0 117900.0 1377450.0 ;
      RECT  186900.0 1378950.0 187800.0 1379850.0 ;
      RECT  186900.0 1374450.0 187800.0 1375350.0 ;
      RECT  154050.0 1378950.0 187350.0 1379850.0 ;
      RECT  186900.0 1374900.0 187800.0 1379400.0 ;
      RECT  187350.0 1374450.0 220800.0 1375350.0 ;
      RECT  115500.0 1393350.0 116400.0 1394250.0 ;
      RECT  115500.0 1395750.0 116400.0 1396650.0 ;
      RECT  114150.0 1393350.0 115950.0 1394250.0 ;
      RECT  115500.0 1393800.0 116400.0 1396200.0 ;
      RECT  115950.0 1395750.0 117900.0 1396650.0 ;
      RECT  186900.0 1393350.0 187800.0 1394250.0 ;
      RECT  186900.0 1397850.0 187800.0 1398750.0 ;
      RECT  154050.0 1393350.0 187350.0 1394250.0 ;
      RECT  186900.0 1393800.0 187800.0 1398300.0 ;
      RECT  187350.0 1397850.0 220800.0 1398750.0 ;
      RECT  115500.0 1406550.0 116400.0 1407450.0 ;
      RECT  115500.0 1404150.0 116400.0 1405050.0 ;
      RECT  114150.0 1406550.0 115950.0 1407450.0 ;
      RECT  115500.0 1404600.0 116400.0 1407000.0 ;
      RECT  115950.0 1404150.0 117900.0 1405050.0 ;
      RECT  186900.0 1406550.0 187800.0 1407450.0 ;
      RECT  186900.0 1402050.0 187800.0 1402950.0 ;
      RECT  154050.0 1406550.0 187350.0 1407450.0 ;
      RECT  186900.0 1402500.0 187800.0 1407000.0 ;
      RECT  187350.0 1402050.0 220800.0 1402950.0 ;
      RECT  115500.0 1420950.0 116400.0 1421850.0 ;
      RECT  115500.0 1423350.0 116400.0 1424250.0 ;
      RECT  114150.0 1420950.0 115950.0 1421850.0 ;
      RECT  115500.0 1421400.0 116400.0 1423800.0 ;
      RECT  115950.0 1423350.0 117900.0 1424250.0 ;
      RECT  186900.0 1420950.0 187800.0 1421850.0 ;
      RECT  186900.0 1425450.0 187800.0 1426350.0 ;
      RECT  154050.0 1420950.0 187350.0 1421850.0 ;
      RECT  186900.0 1421400.0 187800.0 1425900.0 ;
      RECT  187350.0 1425450.0 220800.0 1426350.0 ;
      RECT  115500.0 1434150.0 116400.0 1435050.0 ;
      RECT  115500.0 1431750.0 116400.0 1432650.0 ;
      RECT  114150.0 1434150.0 115950.0 1435050.0 ;
      RECT  115500.0 1432200.0 116400.0 1434600.0 ;
      RECT  115950.0 1431750.0 117900.0 1432650.0 ;
      RECT  186900.0 1434150.0 187800.0 1435050.0 ;
      RECT  186900.0 1429650.0 187800.0 1430550.0 ;
      RECT  154050.0 1434150.0 187350.0 1435050.0 ;
      RECT  186900.0 1430100.0 187800.0 1434600.0 ;
      RECT  187350.0 1429650.0 220800.0 1430550.0 ;
      RECT  115500.0 1448550.0 116400.0 1449450.0 ;
      RECT  115500.0 1450950.0 116400.0 1451850.0 ;
      RECT  114150.0 1448550.0 115950.0 1449450.0 ;
      RECT  115500.0 1449000.0 116400.0 1451400.0 ;
      RECT  115950.0 1450950.0 117900.0 1451850.0 ;
      RECT  186900.0 1448550.0 187800.0 1449450.0 ;
      RECT  186900.0 1453050.0 187800.0 1453950.0 ;
      RECT  154050.0 1448550.0 187350.0 1449450.0 ;
      RECT  186900.0 1449000.0 187800.0 1453500.0 ;
      RECT  187350.0 1453050.0 220800.0 1453950.0 ;
      RECT  115500.0 1461750.0 116400.0 1462650.0 ;
      RECT  115500.0 1459350.0 116400.0 1460250.0 ;
      RECT  114150.0 1461750.0 115950.0 1462650.0 ;
      RECT  115500.0 1459800.0 116400.0 1462200.0 ;
      RECT  115950.0 1459350.0 117900.0 1460250.0 ;
      RECT  186900.0 1461750.0 187800.0 1462650.0 ;
      RECT  186900.0 1457250.0 187800.0 1458150.0 ;
      RECT  154050.0 1461750.0 187350.0 1462650.0 ;
      RECT  186900.0 1457700.0 187800.0 1462200.0 ;
      RECT  187350.0 1457250.0 220800.0 1458150.0 ;
      RECT  115500.0 1476150.0 116400.0 1477050.0 ;
      RECT  115500.0 1478550.0 116400.0 1479450.0 ;
      RECT  114150.0 1476150.0 115950.0 1477050.0 ;
      RECT  115500.0 1476600.0 116400.0 1479000.0 ;
      RECT  115950.0 1478550.0 117900.0 1479450.0 ;
      RECT  186900.0 1476150.0 187800.0 1477050.0 ;
      RECT  186900.0 1480650.0 187800.0 1481550.0 ;
      RECT  154050.0 1476150.0 187350.0 1477050.0 ;
      RECT  186900.0 1476600.0 187800.0 1481100.0 ;
      RECT  187350.0 1480650.0 220800.0 1481550.0 ;
      RECT  115500.0 1489350.0 116400.0 1490250.0 ;
      RECT  115500.0 1486950.0 116400.0 1487850.0 ;
      RECT  114150.0 1489350.0 115950.0 1490250.0 ;
      RECT  115500.0 1487400.0 116400.0 1489800.0 ;
      RECT  115950.0 1486950.0 117900.0 1487850.0 ;
      RECT  186900.0 1489350.0 187800.0 1490250.0 ;
      RECT  186900.0 1484850.0 187800.0 1485750.0 ;
      RECT  154050.0 1489350.0 187350.0 1490250.0 ;
      RECT  186900.0 1485300.0 187800.0 1489800.0 ;
      RECT  187350.0 1484850.0 220800.0 1485750.0 ;
      RECT  115500.0 1503750.0 116400.0 1504650.0 ;
      RECT  115500.0 1506150.0 116400.0 1507050.0 ;
      RECT  114150.0 1503750.0 115950.0 1504650.0 ;
      RECT  115500.0 1504200.0 116400.0 1506600.0 ;
      RECT  115950.0 1506150.0 117900.0 1507050.0 ;
      RECT  186900.0 1503750.0 187800.0 1504650.0 ;
      RECT  186900.0 1508250.0 187800.0 1509150.0 ;
      RECT  154050.0 1503750.0 187350.0 1504650.0 ;
      RECT  186900.0 1504200.0 187800.0 1508700.0 ;
      RECT  187350.0 1508250.0 220800.0 1509150.0 ;
      RECT  115500.0 1516950.0 116400.0 1517850.0 ;
      RECT  115500.0 1514550.0 116400.0 1515450.0 ;
      RECT  114150.0 1516950.0 115950.0 1517850.0 ;
      RECT  115500.0 1515000.0 116400.0 1517400.0 ;
      RECT  115950.0 1514550.0 117900.0 1515450.0 ;
      RECT  186900.0 1516950.0 187800.0 1517850.0 ;
      RECT  186900.0 1512450.0 187800.0 1513350.0 ;
      RECT  154050.0 1516950.0 187350.0 1517850.0 ;
      RECT  186900.0 1512900.0 187800.0 1517400.0 ;
      RECT  187350.0 1512450.0 220800.0 1513350.0 ;
      RECT  115500.0 1531350.0 116400.0 1532250.0 ;
      RECT  115500.0 1533750.0 116400.0 1534650.0 ;
      RECT  114150.0 1531350.0 115950.0 1532250.0 ;
      RECT  115500.0 1531800.0 116400.0 1534200.0 ;
      RECT  115950.0 1533750.0 117900.0 1534650.0 ;
      RECT  186900.0 1531350.0 187800.0 1532250.0 ;
      RECT  186900.0 1535850.0 187800.0 1536750.0 ;
      RECT  154050.0 1531350.0 187350.0 1532250.0 ;
      RECT  186900.0 1531800.0 187800.0 1536300.0 ;
      RECT  187350.0 1535850.0 220800.0 1536750.0 ;
      RECT  115500.0 1544550.0 116400.0 1545450.0 ;
      RECT  115500.0 1542150.0 116400.0 1543050.0 ;
      RECT  114150.0 1544550.0 115950.0 1545450.0 ;
      RECT  115500.0 1542600.0 116400.0 1545000.0 ;
      RECT  115950.0 1542150.0 117900.0 1543050.0 ;
      RECT  186900.0 1544550.0 187800.0 1545450.0 ;
      RECT  186900.0 1540050.0 187800.0 1540950.0 ;
      RECT  154050.0 1544550.0 187350.0 1545450.0 ;
      RECT  186900.0 1540500.0 187800.0 1545000.0 ;
      RECT  187350.0 1540050.0 220800.0 1540950.0 ;
      RECT  115500.0 1558950.0 116400.0 1559850.0 ;
      RECT  115500.0 1561350.0 116400.0 1562250.0 ;
      RECT  114150.0 1558950.0 115950.0 1559850.0 ;
      RECT  115500.0 1559400.0 116400.0 1561800.0 ;
      RECT  115950.0 1561350.0 117900.0 1562250.0 ;
      RECT  186900.0 1558950.0 187800.0 1559850.0 ;
      RECT  186900.0 1563450.0 187800.0 1564350.0 ;
      RECT  154050.0 1558950.0 187350.0 1559850.0 ;
      RECT  186900.0 1559400.0 187800.0 1563900.0 ;
      RECT  187350.0 1563450.0 220800.0 1564350.0 ;
      RECT  115500.0 1572150.0 116400.0 1573050.0 ;
      RECT  115500.0 1569750.0 116400.0 1570650.0 ;
      RECT  114150.0 1572150.0 115950.0 1573050.0 ;
      RECT  115500.0 1570200.0 116400.0 1572600.0 ;
      RECT  115950.0 1569750.0 117900.0 1570650.0 ;
      RECT  186900.0 1572150.0 187800.0 1573050.0 ;
      RECT  186900.0 1567650.0 187800.0 1568550.0 ;
      RECT  154050.0 1572150.0 187350.0 1573050.0 ;
      RECT  186900.0 1568100.0 187800.0 1572600.0 ;
      RECT  187350.0 1567650.0 220800.0 1568550.0 ;
      RECT  115500.0 1586550.0 116400.0 1587450.0 ;
      RECT  115500.0 1588950.0 116400.0 1589850.0 ;
      RECT  114150.0 1586550.0 115950.0 1587450.0 ;
      RECT  115500.0 1587000.0 116400.0 1589400.0 ;
      RECT  115950.0 1588950.0 117900.0 1589850.0 ;
      RECT  186900.0 1586550.0 187800.0 1587450.0 ;
      RECT  186900.0 1591050.0 187800.0 1591950.0 ;
      RECT  154050.0 1586550.0 187350.0 1587450.0 ;
      RECT  186900.0 1587000.0 187800.0 1591500.0 ;
      RECT  187350.0 1591050.0 220800.0 1591950.0 ;
      RECT  115500.0 1599750.0 116400.0 1600650.0 ;
      RECT  115500.0 1597350.0 116400.0 1598250.0 ;
      RECT  114150.0 1599750.0 115950.0 1600650.0 ;
      RECT  115500.0 1597800.0 116400.0 1600200.0 ;
      RECT  115950.0 1597350.0 117900.0 1598250.0 ;
      RECT  186900.0 1599750.0 187800.0 1600650.0 ;
      RECT  186900.0 1595250.0 187800.0 1596150.0 ;
      RECT  154050.0 1599750.0 187350.0 1600650.0 ;
      RECT  186900.0 1595700.0 187800.0 1600200.0 ;
      RECT  187350.0 1595250.0 220800.0 1596150.0 ;
      RECT  115500.0 1614150.0 116400.0 1615050.0 ;
      RECT  115500.0 1616550.0 116400.0 1617450.0 ;
      RECT  114150.0 1614150.0 115950.0 1615050.0 ;
      RECT  115500.0 1614600.0 116400.0 1617000.0 ;
      RECT  115950.0 1616550.0 117900.0 1617450.0 ;
      RECT  186900.0 1614150.0 187800.0 1615050.0 ;
      RECT  186900.0 1618650.0 187800.0 1619550.0 ;
      RECT  154050.0 1614150.0 187350.0 1615050.0 ;
      RECT  186900.0 1614600.0 187800.0 1619100.0 ;
      RECT  187350.0 1618650.0 220800.0 1619550.0 ;
      RECT  115500.0 1627350.0 116400.0 1628250.0 ;
      RECT  115500.0 1624950.0 116400.0 1625850.0 ;
      RECT  114150.0 1627350.0 115950.0 1628250.0 ;
      RECT  115500.0 1625400.0 116400.0 1627800.0 ;
      RECT  115950.0 1624950.0 117900.0 1625850.0 ;
      RECT  186900.0 1627350.0 187800.0 1628250.0 ;
      RECT  186900.0 1622850.0 187800.0 1623750.0 ;
      RECT  154050.0 1627350.0 187350.0 1628250.0 ;
      RECT  186900.0 1623300.0 187800.0 1627800.0 ;
      RECT  187350.0 1622850.0 220800.0 1623750.0 ;
      RECT  115500.0 1641750.0 116400.0 1642650.0 ;
      RECT  115500.0 1644150.0 116400.0 1645050.0 ;
      RECT  114150.0 1641750.0 115950.0 1642650.0 ;
      RECT  115500.0 1642200.0 116400.0 1644600.0 ;
      RECT  115950.0 1644150.0 117900.0 1645050.0 ;
      RECT  186900.0 1641750.0 187800.0 1642650.0 ;
      RECT  186900.0 1646250.0 187800.0 1647150.0 ;
      RECT  154050.0 1641750.0 187350.0 1642650.0 ;
      RECT  186900.0 1642200.0 187800.0 1646700.0 ;
      RECT  187350.0 1646250.0 220800.0 1647150.0 ;
      RECT  115500.0 1654950.0 116400.0 1655850.0 ;
      RECT  115500.0 1652550.0 116400.0 1653450.0 ;
      RECT  114150.0 1654950.0 115950.0 1655850.0 ;
      RECT  115500.0 1653000.0 116400.0 1655400.0 ;
      RECT  115950.0 1652550.0 117900.0 1653450.0 ;
      RECT  186900.0 1654950.0 187800.0 1655850.0 ;
      RECT  186900.0 1650450.0 187800.0 1651350.0 ;
      RECT  154050.0 1654950.0 187350.0 1655850.0 ;
      RECT  186900.0 1650900.0 187800.0 1655400.0 ;
      RECT  187350.0 1650450.0 220800.0 1651350.0 ;
      RECT  115500.0 1669350.0 116400.0 1670250.0 ;
      RECT  115500.0 1671750.0 116400.0 1672650.0 ;
      RECT  114150.0 1669350.0 115950.0 1670250.0 ;
      RECT  115500.0 1669800.0 116400.0 1672200.0 ;
      RECT  115950.0 1671750.0 117900.0 1672650.0 ;
      RECT  186900.0 1669350.0 187800.0 1670250.0 ;
      RECT  186900.0 1673850.0 187800.0 1674750.0 ;
      RECT  154050.0 1669350.0 187350.0 1670250.0 ;
      RECT  186900.0 1669800.0 187800.0 1674300.0 ;
      RECT  187350.0 1673850.0 220800.0 1674750.0 ;
      RECT  115500.0 1682550.0 116400.0 1683450.0 ;
      RECT  115500.0 1680150.0 116400.0 1681050.0 ;
      RECT  114150.0 1682550.0 115950.0 1683450.0 ;
      RECT  115500.0 1680600.0 116400.0 1683000.0 ;
      RECT  115950.0 1680150.0 117900.0 1681050.0 ;
      RECT  186900.0 1682550.0 187800.0 1683450.0 ;
      RECT  186900.0 1678050.0 187800.0 1678950.0 ;
      RECT  154050.0 1682550.0 187350.0 1683450.0 ;
      RECT  186900.0 1678500.0 187800.0 1683000.0 ;
      RECT  187350.0 1678050.0 220800.0 1678950.0 ;
      RECT  115500.0 1696950.0 116400.0 1697850.0 ;
      RECT  115500.0 1699350.0 116400.0 1700250.0 ;
      RECT  114150.0 1696950.0 115950.0 1697850.0 ;
      RECT  115500.0 1697400.0 116400.0 1699800.0 ;
      RECT  115950.0 1699350.0 117900.0 1700250.0 ;
      RECT  186900.0 1696950.0 187800.0 1697850.0 ;
      RECT  186900.0 1701450.0 187800.0 1702350.0 ;
      RECT  154050.0 1696950.0 187350.0 1697850.0 ;
      RECT  186900.0 1697400.0 187800.0 1701900.0 ;
      RECT  187350.0 1701450.0 220800.0 1702350.0 ;
      RECT  115500.0 1710150.0 116400.0 1711050.0 ;
      RECT  115500.0 1707750.0 116400.0 1708650.0 ;
      RECT  114150.0 1710150.0 115950.0 1711050.0 ;
      RECT  115500.0 1708200.0 116400.0 1710600.0 ;
      RECT  115950.0 1707750.0 117900.0 1708650.0 ;
      RECT  186900.0 1710150.0 187800.0 1711050.0 ;
      RECT  186900.0 1705650.0 187800.0 1706550.0 ;
      RECT  154050.0 1710150.0 187350.0 1711050.0 ;
      RECT  186900.0 1706100.0 187800.0 1710600.0 ;
      RECT  187350.0 1705650.0 220800.0 1706550.0 ;
      RECT  115500.0 1724550.0 116400.0 1725450.0 ;
      RECT  115500.0 1726950.0 116400.0 1727850.0 ;
      RECT  114150.0 1724550.0 115950.0 1725450.0 ;
      RECT  115500.0 1725000.0 116400.0 1727400.0 ;
      RECT  115950.0 1726950.0 117900.0 1727850.0 ;
      RECT  186900.0 1724550.0 187800.0 1725450.0 ;
      RECT  186900.0 1729050.0 187800.0 1729950.0 ;
      RECT  154050.0 1724550.0 187350.0 1725450.0 ;
      RECT  186900.0 1725000.0 187800.0 1729500.0 ;
      RECT  187350.0 1729050.0 220800.0 1729950.0 ;
      RECT  115500.0 1737750.0 116400.0 1738650.0 ;
      RECT  115500.0 1735350.0 116400.0 1736250.0 ;
      RECT  114150.0 1737750.0 115950.0 1738650.0 ;
      RECT  115500.0 1735800.0 116400.0 1738200.0 ;
      RECT  115950.0 1735350.0 117900.0 1736250.0 ;
      RECT  186900.0 1737750.0 187800.0 1738650.0 ;
      RECT  186900.0 1733250.0 187800.0 1734150.0 ;
      RECT  154050.0 1737750.0 187350.0 1738650.0 ;
      RECT  186900.0 1733700.0 187800.0 1738200.0 ;
      RECT  187350.0 1733250.0 220800.0 1734150.0 ;
      RECT  115500.0 1752150.0 116400.0 1753050.0 ;
      RECT  115500.0 1754550.0 116400.0 1755450.0 ;
      RECT  114150.0 1752150.0 115950.0 1753050.0 ;
      RECT  115500.0 1752600.0 116400.0 1755000.0 ;
      RECT  115950.0 1754550.0 117900.0 1755450.0 ;
      RECT  186900.0 1752150.0 187800.0 1753050.0 ;
      RECT  186900.0 1756650.0 187800.0 1757550.0 ;
      RECT  154050.0 1752150.0 187350.0 1753050.0 ;
      RECT  186900.0 1752600.0 187800.0 1757100.0 ;
      RECT  187350.0 1756650.0 220800.0 1757550.0 ;
      RECT  115500.0 1765350.0 116400.0 1766250.0 ;
      RECT  115500.0 1762950.0 116400.0 1763850.0 ;
      RECT  114150.0 1765350.0 115950.0 1766250.0 ;
      RECT  115500.0 1763400.0 116400.0 1765800.0 ;
      RECT  115950.0 1762950.0 117900.0 1763850.0 ;
      RECT  186900.0 1765350.0 187800.0 1766250.0 ;
      RECT  186900.0 1760850.0 187800.0 1761750.0 ;
      RECT  154050.0 1765350.0 187350.0 1766250.0 ;
      RECT  186900.0 1761300.0 187800.0 1765800.0 ;
      RECT  187350.0 1760850.0 220800.0 1761750.0 ;
      RECT  115500.0 1779750.0 116400.0 1780650.0 ;
      RECT  115500.0 1782150.0 116400.0 1783050.0 ;
      RECT  114150.0 1779750.0 115950.0 1780650.0 ;
      RECT  115500.0 1780200.0 116400.0 1782600.0 ;
      RECT  115950.0 1782150.0 117900.0 1783050.0 ;
      RECT  186900.0 1779750.0 187800.0 1780650.0 ;
      RECT  186900.0 1784250.0 187800.0 1785150.0 ;
      RECT  154050.0 1779750.0 187350.0 1780650.0 ;
      RECT  186900.0 1780200.0 187800.0 1784700.0 ;
      RECT  187350.0 1784250.0 220800.0 1785150.0 ;
      RECT  115500.0 1792950.0 116400.0 1793850.0 ;
      RECT  115500.0 1790550.0 116400.0 1791450.0 ;
      RECT  114150.0 1792950.0 115950.0 1793850.0 ;
      RECT  115500.0 1791000.0 116400.0 1793400.0 ;
      RECT  115950.0 1790550.0 117900.0 1791450.0 ;
      RECT  186900.0 1792950.0 187800.0 1793850.0 ;
      RECT  186900.0 1788450.0 187800.0 1789350.0 ;
      RECT  154050.0 1792950.0 187350.0 1793850.0 ;
      RECT  186900.0 1788900.0 187800.0 1793400.0 ;
      RECT  187350.0 1788450.0 220800.0 1789350.0 ;
      RECT  115500.0 1807350.0 116400.0 1808250.0 ;
      RECT  115500.0 1809750.0 116400.0 1810650.0 ;
      RECT  114150.0 1807350.0 115950.0 1808250.0 ;
      RECT  115500.0 1807800.0 116400.0 1810200.0 ;
      RECT  115950.0 1809750.0 117900.0 1810650.0 ;
      RECT  186900.0 1807350.0 187800.0 1808250.0 ;
      RECT  186900.0 1811850.0 187800.0 1812750.0 ;
      RECT  154050.0 1807350.0 187350.0 1808250.0 ;
      RECT  186900.0 1807800.0 187800.0 1812300.0 ;
      RECT  187350.0 1811850.0 220800.0 1812750.0 ;
      RECT  115500.0 1820550.0 116400.0 1821450.0 ;
      RECT  115500.0 1818150.0 116400.0 1819050.0 ;
      RECT  114150.0 1820550.0 115950.0 1821450.0 ;
      RECT  115500.0 1818600.0 116400.0 1821000.0 ;
      RECT  115950.0 1818150.0 117900.0 1819050.0 ;
      RECT  186900.0 1820550.0 187800.0 1821450.0 ;
      RECT  186900.0 1816050.0 187800.0 1816950.0 ;
      RECT  154050.0 1820550.0 187350.0 1821450.0 ;
      RECT  186900.0 1816500.0 187800.0 1821000.0 ;
      RECT  187350.0 1816050.0 220800.0 1816950.0 ;
      RECT  115500.0 1834950.0 116400.0 1835850.0 ;
      RECT  115500.0 1837350.0 116400.0 1838250.0 ;
      RECT  114150.0 1834950.0 115950.0 1835850.0 ;
      RECT  115500.0 1835400.0 116400.0 1837800.0 ;
      RECT  115950.0 1837350.0 117900.0 1838250.0 ;
      RECT  186900.0 1834950.0 187800.0 1835850.0 ;
      RECT  186900.0 1839450.0 187800.0 1840350.0 ;
      RECT  154050.0 1834950.0 187350.0 1835850.0 ;
      RECT  186900.0 1835400.0 187800.0 1839900.0 ;
      RECT  187350.0 1839450.0 220800.0 1840350.0 ;
      RECT  115500.0 1848150.0 116400.0 1849050.0 ;
      RECT  115500.0 1845750.0 116400.0 1846650.0 ;
      RECT  114150.0 1848150.0 115950.0 1849050.0 ;
      RECT  115500.0 1846200.0 116400.0 1848600.0 ;
      RECT  115950.0 1845750.0 117900.0 1846650.0 ;
      RECT  186900.0 1848150.0 187800.0 1849050.0 ;
      RECT  186900.0 1843650.0 187800.0 1844550.0 ;
      RECT  154050.0 1848150.0 187350.0 1849050.0 ;
      RECT  186900.0 1844100.0 187800.0 1848600.0 ;
      RECT  187350.0 1843650.0 220800.0 1844550.0 ;
      RECT  115500.0 1862550.0 116400.0 1863450.0 ;
      RECT  115500.0 1864950.0 116400.0 1865850.0 ;
      RECT  114150.0 1862550.0 115950.0 1863450.0 ;
      RECT  115500.0 1863000.0 116400.0 1865400.0 ;
      RECT  115950.0 1864950.0 117900.0 1865850.0 ;
      RECT  186900.0 1862550.0 187800.0 1863450.0 ;
      RECT  186900.0 1867050.0 187800.0 1867950.0 ;
      RECT  154050.0 1862550.0 187350.0 1863450.0 ;
      RECT  186900.0 1863000.0 187800.0 1867500.0 ;
      RECT  187350.0 1867050.0 220800.0 1867950.0 ;
      RECT  115500.0 1875750.0 116400.0 1876650.0 ;
      RECT  115500.0 1873350.0 116400.0 1874250.0 ;
      RECT  114150.0 1875750.0 115950.0 1876650.0 ;
      RECT  115500.0 1873800.0 116400.0 1876200.0 ;
      RECT  115950.0 1873350.0 117900.0 1874250.0 ;
      RECT  186900.0 1875750.0 187800.0 1876650.0 ;
      RECT  186900.0 1871250.0 187800.0 1872150.0 ;
      RECT  154050.0 1875750.0 187350.0 1876650.0 ;
      RECT  186900.0 1871700.0 187800.0 1876200.0 ;
      RECT  187350.0 1871250.0 220800.0 1872150.0 ;
      RECT  115500.0 1890150.0 116400.0 1891050.0 ;
      RECT  115500.0 1892550.0 116400.0 1893450.0 ;
      RECT  114150.0 1890150.0 115950.0 1891050.0 ;
      RECT  115500.0 1890600.0 116400.0 1893000.0 ;
      RECT  115950.0 1892550.0 117900.0 1893450.0 ;
      RECT  186900.0 1890150.0 187800.0 1891050.0 ;
      RECT  186900.0 1894650.0 187800.0 1895550.0 ;
      RECT  154050.0 1890150.0 187350.0 1891050.0 ;
      RECT  186900.0 1890600.0 187800.0 1895100.0 ;
      RECT  187350.0 1894650.0 220800.0 1895550.0 ;
      RECT  115500.0 1903350.0 116400.0 1904250.0 ;
      RECT  115500.0 1900950.0 116400.0 1901850.0 ;
      RECT  114150.0 1903350.0 115950.0 1904250.0 ;
      RECT  115500.0 1901400.0 116400.0 1903800.0 ;
      RECT  115950.0 1900950.0 117900.0 1901850.0 ;
      RECT  186900.0 1903350.0 187800.0 1904250.0 ;
      RECT  186900.0 1898850.0 187800.0 1899750.0 ;
      RECT  154050.0 1903350.0 187350.0 1904250.0 ;
      RECT  186900.0 1899300.0 187800.0 1903800.0 ;
      RECT  187350.0 1898850.0 220800.0 1899750.0 ;
      RECT  115500.0 1917750.0 116400.0 1918650.0 ;
      RECT  115500.0 1920150.0 116400.0 1921050.0 ;
      RECT  114150.0 1917750.0 115950.0 1918650.0 ;
      RECT  115500.0 1918200.0 116400.0 1920600.0 ;
      RECT  115950.0 1920150.0 117900.0 1921050.0 ;
      RECT  186900.0 1917750.0 187800.0 1918650.0 ;
      RECT  186900.0 1922250.0 187800.0 1923150.0 ;
      RECT  154050.0 1917750.0 187350.0 1918650.0 ;
      RECT  186900.0 1918200.0 187800.0 1922700.0 ;
      RECT  187350.0 1922250.0 220800.0 1923150.0 ;
      RECT  115500.0 1930950.0 116400.0 1931850.0 ;
      RECT  115500.0 1928550.0 116400.0 1929450.0 ;
      RECT  114150.0 1930950.0 115950.0 1931850.0 ;
      RECT  115500.0 1929000.0 116400.0 1931400.0 ;
      RECT  115950.0 1928550.0 117900.0 1929450.0 ;
      RECT  186900.0 1930950.0 187800.0 1931850.0 ;
      RECT  186900.0 1926450.0 187800.0 1927350.0 ;
      RECT  154050.0 1930950.0 187350.0 1931850.0 ;
      RECT  186900.0 1926900.0 187800.0 1931400.0 ;
      RECT  187350.0 1926450.0 220800.0 1927350.0 ;
      RECT  115500.0 1945350.0 116400.0 1946250.0 ;
      RECT  115500.0 1947750.0 116400.0 1948650.0 ;
      RECT  114150.0 1945350.0 115950.0 1946250.0 ;
      RECT  115500.0 1945800.0 116400.0 1948200.0 ;
      RECT  115950.0 1947750.0 117900.0 1948650.0 ;
      RECT  186900.0 1945350.0 187800.0 1946250.0 ;
      RECT  186900.0 1949850.0 187800.0 1950750.0 ;
      RECT  154050.0 1945350.0 187350.0 1946250.0 ;
      RECT  186900.0 1945800.0 187800.0 1950300.0 ;
      RECT  187350.0 1949850.0 220800.0 1950750.0 ;
      RECT  115500.0 1958550.0 116400.0 1959450.0 ;
      RECT  115500.0 1956150.0 116400.0 1957050.0 ;
      RECT  114150.0 1958550.0 115950.0 1959450.0 ;
      RECT  115500.0 1956600.0 116400.0 1959000.0 ;
      RECT  115950.0 1956150.0 117900.0 1957050.0 ;
      RECT  186900.0 1958550.0 187800.0 1959450.0 ;
      RECT  186900.0 1954050.0 187800.0 1954950.0 ;
      RECT  154050.0 1958550.0 187350.0 1959450.0 ;
      RECT  186900.0 1954500.0 187800.0 1959000.0 ;
      RECT  187350.0 1954050.0 220800.0 1954950.0 ;
      RECT  115500.0 1972950.0 116400.0 1973850.0 ;
      RECT  115500.0 1975350.0 116400.0 1976250.0 ;
      RECT  114150.0 1972950.0 115950.0 1973850.0 ;
      RECT  115500.0 1973400.0 116400.0 1975800.0 ;
      RECT  115950.0 1975350.0 117900.0 1976250.0 ;
      RECT  186900.0 1972950.0 187800.0 1973850.0 ;
      RECT  186900.0 1977450.0 187800.0 1978350.0 ;
      RECT  154050.0 1972950.0 187350.0 1973850.0 ;
      RECT  186900.0 1973400.0 187800.0 1977900.0 ;
      RECT  187350.0 1977450.0 220800.0 1978350.0 ;
      RECT  115500.0 1986150.0 116400.0 1987050.0 ;
      RECT  115500.0 1983750.0 116400.0 1984650.0 ;
      RECT  114150.0 1986150.0 115950.0 1987050.0 ;
      RECT  115500.0 1984200.0 116400.0 1986600.0 ;
      RECT  115950.0 1983750.0 117900.0 1984650.0 ;
      RECT  186900.0 1986150.0 187800.0 1987050.0 ;
      RECT  186900.0 1981650.0 187800.0 1982550.0 ;
      RECT  154050.0 1986150.0 187350.0 1987050.0 ;
      RECT  186900.0 1982100.0 187800.0 1986600.0 ;
      RECT  187350.0 1981650.0 220800.0 1982550.0 ;
      RECT  115500.0 2000550.0 116400.0 2001450.0 ;
      RECT  115500.0 2002950.0 116400.0 2003850.0 ;
      RECT  114150.0 2000550.0 115950.0 2001450.0 ;
      RECT  115500.0 2001000.0 116400.0 2003400.0 ;
      RECT  115950.0 2002950.0 117900.0 2003850.0 ;
      RECT  186900.0 2000550.0 187800.0 2001450.0 ;
      RECT  186900.0 2005050.0 187800.0 2005950.0 ;
      RECT  154050.0 2000550.0 187350.0 2001450.0 ;
      RECT  186900.0 2001000.0 187800.0 2005500.0 ;
      RECT  187350.0 2005050.0 220800.0 2005950.0 ;
      RECT  115500.0 2013750.0 116400.0 2014650.0 ;
      RECT  115500.0 2011350.0 116400.0 2012250.0 ;
      RECT  114150.0 2013750.0 115950.0 2014650.0 ;
      RECT  115500.0 2011800.0 116400.0 2014200.0 ;
      RECT  115950.0 2011350.0 117900.0 2012250.0 ;
      RECT  186900.0 2013750.0 187800.0 2014650.0 ;
      RECT  186900.0 2009250.0 187800.0 2010150.0 ;
      RECT  154050.0 2013750.0 187350.0 2014650.0 ;
      RECT  186900.0 2009700.0 187800.0 2014200.0 ;
      RECT  187350.0 2009250.0 220800.0 2010150.0 ;
      RECT  115500.0 2028150.0 116400.0 2029050.0 ;
      RECT  115500.0 2030550.0 116400.0 2031450.0 ;
      RECT  114150.0 2028150.0 115950.0 2029050.0 ;
      RECT  115500.0 2028600.0 116400.0 2031000.0 ;
      RECT  115950.0 2030550.0 117900.0 2031450.0 ;
      RECT  186900.0 2028150.0 187800.0 2029050.0 ;
      RECT  186900.0 2032650.0 187800.0 2033550.0 ;
      RECT  154050.0 2028150.0 187350.0 2029050.0 ;
      RECT  186900.0 2028600.0 187800.0 2033100.0 ;
      RECT  187350.0 2032650.0 220800.0 2033550.0 ;
      RECT  115500.0 2041350.0 116400.0 2042250.0 ;
      RECT  115500.0 2038950.0 116400.0 2039850.0 ;
      RECT  114150.0 2041350.0 115950.0 2042250.0 ;
      RECT  115500.0 2039400.0 116400.0 2041800.0 ;
      RECT  115950.0 2038950.0 117900.0 2039850.0 ;
      RECT  186900.0 2041350.0 187800.0 2042250.0 ;
      RECT  186900.0 2036850.0 187800.0 2037750.0 ;
      RECT  154050.0 2041350.0 187350.0 2042250.0 ;
      RECT  186900.0 2037300.0 187800.0 2041800.0 ;
      RECT  187350.0 2036850.0 220800.0 2037750.0 ;
      RECT  115500.0 2055750.0 116400.0 2056650.0 ;
      RECT  115500.0 2058150.0 116400.0 2059050.0 ;
      RECT  114150.0 2055750.0 115950.0 2056650.0 ;
      RECT  115500.0 2056200.0 116400.0 2058600.0 ;
      RECT  115950.0 2058150.0 117900.0 2059050.0 ;
      RECT  186900.0 2055750.0 187800.0 2056650.0 ;
      RECT  186900.0 2060250.0 187800.0 2061150.0 ;
      RECT  154050.0 2055750.0 187350.0 2056650.0 ;
      RECT  186900.0 2056200.0 187800.0 2060700.0 ;
      RECT  187350.0 2060250.0 220800.0 2061150.0 ;
      RECT  115500.0 2068950.0 116400.0 2069850.0 ;
      RECT  115500.0 2066550.0 116400.0 2067450.0 ;
      RECT  114150.0 2068950.0 115950.0 2069850.0 ;
      RECT  115500.0 2067000.0 116400.0 2069400.0 ;
      RECT  115950.0 2066550.0 117900.0 2067450.0 ;
      RECT  186900.0 2068950.0 187800.0 2069850.0 ;
      RECT  186900.0 2064450.0 187800.0 2065350.0 ;
      RECT  154050.0 2068950.0 187350.0 2069850.0 ;
      RECT  186900.0 2064900.0 187800.0 2069400.0 ;
      RECT  187350.0 2064450.0 220800.0 2065350.0 ;
      RECT  115500.0 2083350.0 116400.0 2084250.0 ;
      RECT  115500.0 2085750.0 116400.0 2086650.0 ;
      RECT  114150.0 2083350.0 115950.0 2084250.0 ;
      RECT  115500.0 2083800.0 116400.0 2086200.0 ;
      RECT  115950.0 2085750.0 117900.0 2086650.0 ;
      RECT  186900.0 2083350.0 187800.0 2084250.0 ;
      RECT  186900.0 2087850.0 187800.0 2088750.0 ;
      RECT  154050.0 2083350.0 187350.0 2084250.0 ;
      RECT  186900.0 2083800.0 187800.0 2088300.0 ;
      RECT  187350.0 2087850.0 220800.0 2088750.0 ;
      RECT  115500.0 2096550.0 116400.0 2097450.0 ;
      RECT  115500.0 2094150.0 116400.0 2095050.0 ;
      RECT  114150.0 2096550.0 115950.0 2097450.0 ;
      RECT  115500.0 2094600.0 116400.0 2097000.0 ;
      RECT  115950.0 2094150.0 117900.0 2095050.0 ;
      RECT  186900.0 2096550.0 187800.0 2097450.0 ;
      RECT  186900.0 2092050.0 187800.0 2092950.0 ;
      RECT  154050.0 2096550.0 187350.0 2097450.0 ;
      RECT  186900.0 2092500.0 187800.0 2097000.0 ;
      RECT  187350.0 2092050.0 220800.0 2092950.0 ;
      RECT  115500.0 2110950.0 116400.0 2111850.0 ;
      RECT  115500.0 2113350.0 116400.0 2114250.0 ;
      RECT  114150.0 2110950.0 115950.0 2111850.0 ;
      RECT  115500.0 2111400.0 116400.0 2113800.0 ;
      RECT  115950.0 2113350.0 117900.0 2114250.0 ;
      RECT  186900.0 2110950.0 187800.0 2111850.0 ;
      RECT  186900.0 2115450.0 187800.0 2116350.0 ;
      RECT  154050.0 2110950.0 187350.0 2111850.0 ;
      RECT  186900.0 2111400.0 187800.0 2115900.0 ;
      RECT  187350.0 2115450.0 220800.0 2116350.0 ;
      RECT  115500.0 2124150.0 116400.0 2125050.0 ;
      RECT  115500.0 2121750.0 116400.0 2122650.0 ;
      RECT  114150.0 2124150.0 115950.0 2125050.0 ;
      RECT  115500.0 2122200.0 116400.0 2124600.0 ;
      RECT  115950.0 2121750.0 117900.0 2122650.0 ;
      RECT  186900.0 2124150.0 187800.0 2125050.0 ;
      RECT  186900.0 2119650.0 187800.0 2120550.0 ;
      RECT  154050.0 2124150.0 187350.0 2125050.0 ;
      RECT  186900.0 2120100.0 187800.0 2124600.0 ;
      RECT  187350.0 2119650.0 220800.0 2120550.0 ;
      RECT  115500.0 2138550.0 116400.0 2139450.0 ;
      RECT  115500.0 2140950.0 116400.0 2141850.0 ;
      RECT  114150.0 2138550.0 115950.0 2139450.0 ;
      RECT  115500.0 2139000.0 116400.0 2141400.0 ;
      RECT  115950.0 2140950.0 117900.0 2141850.0 ;
      RECT  186900.0 2138550.0 187800.0 2139450.0 ;
      RECT  186900.0 2143050.0 187800.0 2143950.0 ;
      RECT  154050.0 2138550.0 187350.0 2139450.0 ;
      RECT  186900.0 2139000.0 187800.0 2143500.0 ;
      RECT  187350.0 2143050.0 220800.0 2143950.0 ;
      RECT  124200.0 378750.0 221400.0 379650.0 ;
      RECT  124200.0 406350.0 221400.0 407250.0 ;
      RECT  124200.0 433950.0 221400.0 434850.0 ;
      RECT  124200.0 461550.0 221400.0 462450.0 ;
      RECT  124200.0 489150.0 221400.0 490050.0 ;
      RECT  124200.0 516750.0 221400.0 517650.0 ;
      RECT  124200.0 544350.0 221400.0 545250.0 ;
      RECT  124200.0 571950.0 221400.0 572850.0 ;
      RECT  124200.0 599550.0 221400.0 600450.0 ;
      RECT  124200.0 627150.0 221400.0 628050.0 ;
      RECT  124200.0 654750.0 221400.0 655650.0 ;
      RECT  124200.0 682350.0 221400.0 683250.0 ;
      RECT  124200.0 709950.0 221400.0 710850.0 ;
      RECT  124200.0 737550.0 221400.0 738450.0 ;
      RECT  124200.0 765150.0 221400.0 766050.0 ;
      RECT  124200.0 792750.0 221400.0 793650.0 ;
      RECT  124200.0 820350.0 221400.0 821250.0 ;
      RECT  124200.0 847950.0 221400.0 848850.0 ;
      RECT  124200.0 875550.0 221400.0 876450.0 ;
      RECT  124200.0 903150.0 221400.0 904050.0 ;
      RECT  124200.0 930750.0 221400.0 931650.0 ;
      RECT  124200.0 958350.0 221400.0 959250.0 ;
      RECT  124200.0 985950.0 221400.0 986850.0 ;
      RECT  124200.0 1013550.0 221400.0 1014450.0 ;
      RECT  124200.0 1041150.0 221400.0 1042050.0 ;
      RECT  124200.0 1068750.0 221400.0 1069650.0 ;
      RECT  124200.0 1096350.0 221400.0 1097250.0 ;
      RECT  124200.0 1123950.0 221400.0 1124850.0 ;
      RECT  124200.0 1151550.0 221400.0 1152450.0 ;
      RECT  124200.0 1179150.0 221400.0 1180050.0 ;
      RECT  124200.0 1206750.0 221400.0 1207650.0 ;
      RECT  124200.0 1234350.0 221400.0 1235250.0 ;
      RECT  124200.0 1261950.0 221400.0 1262850.0 ;
      RECT  124200.0 1289550.0 221400.0 1290450.0 ;
      RECT  124200.0 1317150.0 221400.0 1318050.0 ;
      RECT  124200.0 1344750.0 221400.0 1345650.0 ;
      RECT  124200.0 1372350.0 221400.0 1373250.0 ;
      RECT  124200.0 1399950.0 221400.0 1400850.0 ;
      RECT  124200.0 1427550.0 221400.0 1428450.0 ;
      RECT  124200.0 1455150.0 221400.0 1456050.0 ;
      RECT  124200.0 1482750.0 221400.0 1483650.0 ;
      RECT  124200.0 1510350.0 221400.0 1511250.0 ;
      RECT  124200.0 1537950.0 221400.0 1538850.0 ;
      RECT  124200.0 1565550.0 221400.0 1566450.0 ;
      RECT  124200.0 1593150.0 221400.0 1594050.0 ;
      RECT  124200.0 1620750.0 221400.0 1621650.0 ;
      RECT  124200.0 1648350.0 221400.0 1649250.0 ;
      RECT  124200.0 1675950.0 221400.0 1676850.0 ;
      RECT  124200.0 1703550.0 221400.0 1704450.0 ;
      RECT  124200.0 1731150.0 221400.0 1732050.0 ;
      RECT  124200.0 1758750.0 221400.0 1759650.0 ;
      RECT  124200.0 1786350.0 221400.0 1787250.0 ;
      RECT  124200.0 1813950.0 221400.0 1814850.0 ;
      RECT  124200.0 1841550.0 221400.0 1842450.0 ;
      RECT  124200.0 1869150.0 221400.0 1870050.0 ;
      RECT  124200.0 1896750.0 221400.0 1897650.0 ;
      RECT  124200.0 1924350.0 221400.0 1925250.0 ;
      RECT  124200.0 1951950.0 221400.0 1952850.0 ;
      RECT  124200.0 1979550.0 221400.0 1980450.0 ;
      RECT  124200.0 2007150.0 221400.0 2008050.0 ;
      RECT  124200.0 2034750.0 221400.0 2035650.0 ;
      RECT  124200.0 2062350.0 221400.0 2063250.0 ;
      RECT  124200.0 2089950.0 221400.0 2090850.0 ;
      RECT  124200.0 2117550.0 221400.0 2118450.0 ;
      RECT  124200.0 2145150.0 221400.0 2146050.0 ;
      RECT  52800.0 392550.0 1534200.0 393450.0 ;
      RECT  52800.0 420150.0 1534200.0 421050.0 ;
      RECT  52800.0 447750.0 1534200.0 448650.0 ;
      RECT  52800.0 475350.0 1534200.0 476250.0 ;
      RECT  52800.0 502950.0 1534200.0 503850.0 ;
      RECT  52800.0 530550.0 1534200.0 531450.0 ;
      RECT  52800.0 558150.0 1534200.0 559050.0 ;
      RECT  52800.0 585750.0 1534200.0 586650.0 ;
      RECT  52800.0 613350.0 1534200.0 614250.0 ;
      RECT  52800.0 640950.0 1534200.0 641850.0 ;
      RECT  52800.0 668550.0 1534200.0 669450.0 ;
      RECT  52800.0 696150.0 1534200.0 697050.0 ;
      RECT  52800.0 723750.0 1534200.0 724650.0 ;
      RECT  52800.0 751350.0 1534200.0 752250.0 ;
      RECT  52800.0 778950.0 1534200.0 779850.0 ;
      RECT  52800.0 806550.0 1534200.0 807450.0 ;
      RECT  52800.0 834150.0 1534200.0 835050.0 ;
      RECT  52800.0 861750.0 1534200.0 862650.0 ;
      RECT  52800.0 889350.0 1534200.0 890250.0 ;
      RECT  52800.0 916950.0 1534200.0 917850.0 ;
      RECT  52800.0 944550.0 1534200.0 945450.0 ;
      RECT  52800.0 972150.0 1534200.0 973050.0 ;
      RECT  52800.0 999750.0 1534200.0 1000650.0 ;
      RECT  52800.0 1027350.0 1534200.0 1028250.0 ;
      RECT  52800.0 1054950.0 1534200.0 1055850.0 ;
      RECT  52800.0 1082550.0 1534200.0 1083450.0 ;
      RECT  52800.0 1110150.0 1534200.0 1111050.0 ;
      RECT  52800.0 1137750.0 1534200.0 1138650.0 ;
      RECT  52800.0 1165350.0 1534200.0 1166250.0 ;
      RECT  52800.0 1192950.0 1534200.0 1193850.0 ;
      RECT  52800.0 1220550.0 1534200.0 1221450.0 ;
      RECT  52800.0 1248150.0 1534200.0 1249050.0 ;
      RECT  52800.0 1275750.0 1534200.0 1276650.0 ;
      RECT  52800.0 1303350.0 1534200.0 1304250.0 ;
      RECT  52800.0 1330950.0 1534200.0 1331850.0 ;
      RECT  52800.0 1358550.0 1534200.0 1359450.0 ;
      RECT  52800.0 1386150.0 1534200.0 1387050.0 ;
      RECT  52800.0 1413750.0 1534200.0 1414650.0 ;
      RECT  52800.0 1441350.0 1534200.0 1442250.0 ;
      RECT  52800.0 1468950.0 1534200.0 1469850.0 ;
      RECT  52800.0 1496550.0 1534200.0 1497450.0 ;
      RECT  52800.0 1524150.0 1534200.0 1525050.0 ;
      RECT  52800.0 1551750.0 1534200.0 1552650.0 ;
      RECT  52800.0 1579350.0 1534200.0 1580250.0 ;
      RECT  52800.0 1606950.0 1534200.0 1607850.0 ;
      RECT  52800.0 1634550.0 1534200.0 1635450.0 ;
      RECT  52800.0 1662150.0 1534200.0 1663050.0 ;
      RECT  52800.0 1689750.0 1534200.0 1690650.0 ;
      RECT  52800.0 1717350.0 1534200.0 1718250.0 ;
      RECT  52800.0 1744950.0 1534200.0 1745850.0 ;
      RECT  52800.0 1772550.0 1534200.0 1773450.0 ;
      RECT  52800.0 1800150.0 1534200.0 1801050.0 ;
      RECT  52800.0 1827750.0 1534200.0 1828650.0 ;
      RECT  52800.0 1855350.0 1534200.0 1856250.0 ;
      RECT  52800.0 1882950.0 1534200.0 1883850.0 ;
      RECT  52800.0 1910550.0 1534200.0 1911450.0 ;
      RECT  52800.0 1938150.0 1534200.0 1939050.0 ;
      RECT  52800.0 1965750.0 1534200.0 1966650.0 ;
      RECT  52800.0 1993350.0 1534200.0 1994250.0 ;
      RECT  52800.0 2020950.0 1534200.0 2021850.0 ;
      RECT  52800.0 2048550.0 1534200.0 2049450.0 ;
      RECT  52800.0 2076150.0 1534200.0 2077050.0 ;
      RECT  52800.0 2103750.0 1534200.0 2104650.0 ;
      RECT  52800.0 2131350.0 1534200.0 2132250.0 ;
      RECT  147300.0 160650.0 162000.0 161550.0 ;
      RECT  144300.0 174450.0 164700.0 175350.0 ;
      RECT  147300.0 215850.0 167400.0 216750.0 ;
      RECT  144300.0 229650.0 170100.0 230550.0 ;
      RECT  157500.0 271050.0 172800.0 271950.0 ;
      RECT  154500.0 284850.0 175500.0 285750.0 ;
      RECT  151500.0 298650.0 178200.0 299550.0 ;
      RECT  157500.0 157950.0 159000.0 158850.0 ;
      RECT  157500.0 185550.0 159000.0 186450.0 ;
      RECT  157500.0 213150.0 159000.0 214050.0 ;
      RECT  157500.0 240750.0 159000.0 241650.0 ;
      RECT  157500.0 268350.0 159000.0 269250.0 ;
      RECT  157500.0 295950.0 159000.0 296850.0 ;
      RECT  157500.0 323550.0 159000.0 324450.0 ;
      RECT  157500.0 351150.0 159000.0 352050.0 ;
      RECT  52800.0 171750.0 157500.0 172650.0 ;
      RECT  52800.0 199350.0 157500.0 200250.0 ;
      RECT  52800.0 226950.0 157500.0 227850.0 ;
      RECT  52800.0 254550.0 157500.0 255450.0 ;
      RECT  52800.0 282150.0 157500.0 283050.0 ;
      RECT  52800.0 309750.0 157500.0 310650.0 ;
      RECT  52800.0 337350.0 157500.0 338250.0 ;
      RECT  52800.0 364950.0 157500.0 365850.0 ;
      RECT  180900.0 351300.0 221400.0 352200.0 ;
      RECT  183600.0 349200.0 221400.0 350100.0 ;
      RECT  186300.0 347100.0 221400.0 348000.0 ;
      RECT  189000.0 345000.0 221400.0 345900.0 ;
      RECT  152100.0 6750.0 180900.0 7650.0 ;
      RECT  152100.0 21150.0 183600.0 22050.0 ;
      RECT  152100.0 34350.0 186300.0 35250.0 ;
      RECT  152100.0 48750.0 189000.0 49650.0 ;
      RECT  152100.0 150.0 193950.0 1050.0 ;
      RECT  152100.0 27750.0 193950.0 28650.0 ;
      RECT  152100.0 55350.0 193950.0 56250.0 ;
      RECT  52800.0 13950.0 193950.0 14850.0 ;
      RECT  52800.0 41550.0 193950.0 42450.0 ;
      RECT  117900.0 146700.0 162000.0 147600.0 ;
      RECT  117900.0 138000.0 164700.0 138900.0 ;
      RECT  117900.0 126300.0 167400.0 127200.0 ;
      RECT  117900.0 117600.0 170100.0 118500.0 ;
      RECT  117900.0 105900.0 172800.0 106800.0 ;
      RECT  117900.0 97200.0 175500.0 98100.0 ;
      RECT  117900.0 85500.0 178200.0 86400.0 ;
      RECT  119100.0 142350.0 195150.0 143250.0 ;
      RECT  119100.0 121950.0 195150.0 122850.0 ;
      RECT  119100.0 101550.0 195150.0 102450.0 ;
      RECT  119100.0 81150.0 195150.0 82050.0 ;
      RECT  119100.0 60750.0 195150.0 61650.0 ;
      RECT  115500.0 58650.0 116400.0 59550.0 ;
      RECT  115500.0 59100.0 116400.0 61200.0 ;
      RECT  52800.0 58650.0 115950.0 59550.0 ;
      RECT  209700.0 171450.0 221400.0 172350.0 ;
      RECT  204300.0 166950.0 221400.0 167850.0 ;
      RECT  207000.0 164550.0 221400.0 165450.0 ;
      RECT  209700.0 2154000.0 221400.0 2154900.0 ;
      RECT  212400.0 236250.0 221400.0 237150.0 ;
      RECT  215100.0 334350.0 221400.0 335250.0 ;
      RECT  61500.0 154650.0 62400.0 155550.0 ;
      RECT  61500.0 153000.0 62400.0 155100.0 ;
      RECT  61950.0 154650.0 201600.0 155550.0 ;
      RECT  121050.0 2147250.0 202500.0 2148150.0 ;
      RECT  221400.0 2165100.0 1529700.0 2166000.0 ;
      RECT  221400.0 307050.0 1529700.0 307950.0 ;
      RECT  221400.0 238350.0 1529700.0 239250.0 ;
      RECT  221400.0 225450.0 1529700.0 226350.0 ;
      RECT  221400.0 148650.0 1529700.0 149550.0 ;
      RECT  198450.0 162450.0 221400.0 163350.0 ;
      RECT  198450.0 332250.0 221400.0 333150.0 ;
      RECT  198450.0 234150.0 221400.0 235050.0 ;
      RECT  221400.0 379200.0 231600.0 393000.0 ;
      RECT  221400.0 406800.0 231600.0 393000.0 ;
      RECT  221400.0 406800.0 231600.0 420600.0 ;
      RECT  221400.0 434400.0 231600.0 420600.0 ;
      RECT  221400.0 434400.0 231600.0 448200.0 ;
      RECT  221400.0 462000.0 231600.0 448200.0 ;
      RECT  221400.0 462000.0 231600.0 475800.0 ;
      RECT  221400.0 489600.0 231600.0 475800.0 ;
      RECT  221400.0 489600.0 231600.0 503400.0 ;
      RECT  221400.0 517200.0 231600.0 503400.0 ;
      RECT  221400.0 517200.0 231600.0 531000.0 ;
      RECT  221400.0 544800.0 231600.0 531000.0 ;
      RECT  221400.0 544800.0 231600.0 558600.0 ;
      RECT  221400.0 572400.0 231600.0 558600.0 ;
      RECT  221400.0 572400.0 231600.0 586200.0 ;
      RECT  221400.0 600000.0 231600.0 586200.0 ;
      RECT  221400.0 600000.0 231600.0 613800.0 ;
      RECT  221400.0 627600.0 231600.0 613800.0 ;
      RECT  221400.0 627600.0 231600.0 641400.0 ;
      RECT  221400.0 655200.0 231600.0 641400.0 ;
      RECT  221400.0 655200.0 231600.0 669000.0 ;
      RECT  221400.0 682800.0 231600.0 669000.0 ;
      RECT  221400.0 682800.0 231600.0 696600.0 ;
      RECT  221400.0 710400.0 231600.0 696600.0 ;
      RECT  221400.0 710400.0 231600.0 724200.0 ;
      RECT  221400.0 738000.0 231600.0 724200.0 ;
      RECT  221400.0 738000.0 231600.0 751800.0 ;
      RECT  221400.0 765600.0 231600.0 751800.0 ;
      RECT  221400.0 765600.0 231600.0 779400.0 ;
      RECT  221400.0 793200.0 231600.0 779400.0 ;
      RECT  221400.0 793200.0 231600.0 807000.0 ;
      RECT  221400.0 820800.0 231600.0 807000.0 ;
      RECT  221400.0 820800.0 231600.0 834600.0 ;
      RECT  221400.0 848400.0 231600.0 834600.0 ;
      RECT  221400.0 848400.0 231600.0 862200.0 ;
      RECT  221400.0 876000.0 231600.0 862200.0 ;
      RECT  221400.0 876000.0 231600.0 889800.0 ;
      RECT  221400.0 903600.0 231600.0 889800.0 ;
      RECT  221400.0 903600.0 231600.0 917400.0 ;
      RECT  221400.0 931200.0 231600.0 917400.0 ;
      RECT  221400.0 931200.0 231600.0 945000.0 ;
      RECT  221400.0 958800.0 231600.0 945000.0 ;
      RECT  221400.0 958800.0 231600.0 972600.0 ;
      RECT  221400.0 986400.0 231600.0 972600.0 ;
      RECT  221400.0 986400.0 231600.0 1000200.0 ;
      RECT  221400.0 1014000.0 231600.0 1000200.0 ;
      RECT  221400.0 1014000.0 231600.0 1027800.0 ;
      RECT  221400.0 1041600.0 231600.0 1027800.0 ;
      RECT  221400.0 1041600.0 231600.0 1055400.0 ;
      RECT  221400.0 1069200.0 231600.0 1055400.0 ;
      RECT  221400.0 1069200.0 231600.0 1083000.0 ;
      RECT  221400.0 1096800.0 231600.0 1083000.0 ;
      RECT  221400.0 1096800.0 231600.0 1110600.0 ;
      RECT  221400.0 1124400.0 231600.0 1110600.0 ;
      RECT  221400.0 1124400.0 231600.0 1138200.0 ;
      RECT  221400.0 1152000.0 231600.0 1138200.0 ;
      RECT  221400.0 1152000.0 231600.0 1165800.0 ;
      RECT  221400.0 1179600.0 231600.0 1165800.0 ;
      RECT  221400.0 1179600.0 231600.0 1193400.0 ;
      RECT  221400.0 1207200.0 231600.0 1193400.0 ;
      RECT  221400.0 1207200.0 231600.0 1221000.0 ;
      RECT  221400.0 1234800.0 231600.0 1221000.0 ;
      RECT  221400.0 1234800.0 231600.0 1248600.0 ;
      RECT  221400.0 1262400.0 231600.0 1248600.0 ;
      RECT  221400.0 1262400.0 231600.0 1276200.0 ;
      RECT  221400.0 1290000.0 231600.0 1276200.0 ;
      RECT  221400.0 1290000.0 231600.0 1303800.0 ;
      RECT  221400.0 1317600.0 231600.0 1303800.0 ;
      RECT  221400.0 1317600.0 231600.0 1331400.0 ;
      RECT  221400.0 1345200.0 231600.0 1331400.0 ;
      RECT  221400.0 1345200.0 231600.0 1359000.0 ;
      RECT  221400.0 1372800.0 231600.0 1359000.0 ;
      RECT  221400.0 1372800.0 231600.0 1386600.0 ;
      RECT  221400.0 1400400.0 231600.0 1386600.0 ;
      RECT  221400.0 1400400.0 231600.0 1414200.0 ;
      RECT  221400.0 1428000.0 231600.0 1414200.0 ;
      RECT  221400.0 1428000.0 231600.0 1441800.0 ;
      RECT  221400.0 1455600.0 231600.0 1441800.0 ;
      RECT  221400.0 1455600.0 231600.0 1469400.0 ;
      RECT  221400.0 1483200.0 231600.0 1469400.0 ;
      RECT  221400.0 1483200.0 231600.0 1497000.0 ;
      RECT  221400.0 1510800.0 231600.0 1497000.0 ;
      RECT  221400.0 1510800.0 231600.0 1524600.0 ;
      RECT  221400.0 1538400.0 231600.0 1524600.0 ;
      RECT  221400.0 1538400.0 231600.0 1552200.0 ;
      RECT  221400.0 1566000.0 231600.0 1552200.0 ;
      RECT  221400.0 1566000.0 231600.0 1579800.0 ;
      RECT  221400.0 1593600.0 231600.0 1579800.0 ;
      RECT  221400.0 1593600.0 231600.0 1607400.0 ;
      RECT  221400.0 1621200.0 231600.0 1607400.0 ;
      RECT  221400.0 1621200.0 231600.0 1635000.0 ;
      RECT  221400.0 1648800.0 231600.0 1635000.0 ;
      RECT  221400.0 1648800.0 231600.0 1662600.0 ;
      RECT  221400.0 1676400.0 231600.0 1662600.0 ;
      RECT  221400.0 1676400.0 231600.0 1690200.0 ;
      RECT  221400.0 1704000.0 231600.0 1690200.0 ;
      RECT  221400.0 1704000.0 231600.0 1717800.0 ;
      RECT  221400.0 1731600.0 231600.0 1717800.0 ;
      RECT  221400.0 1731600.0 231600.0 1745400.0 ;
      RECT  221400.0 1759200.0 231600.0 1745400.0 ;
      RECT  221400.0 1759200.0 231600.0 1773000.0 ;
      RECT  221400.0 1786800.0 231600.0 1773000.0 ;
      RECT  221400.0 1786800.0 231600.0 1800600.0 ;
      RECT  221400.0 1814400.0 231600.0 1800600.0 ;
      RECT  221400.0 1814400.0 231600.0 1828200.0 ;
      RECT  221400.0 1842000.0 231600.0 1828200.0 ;
      RECT  221400.0 1842000.0 231600.0 1855800.0 ;
      RECT  221400.0 1869600.0 231600.0 1855800.0 ;
      RECT  221400.0 1869600.0 231600.0 1883400.0 ;
      RECT  221400.0 1897200.0 231600.0 1883400.0 ;
      RECT  221400.0 1897200.0 231600.0 1911000.0 ;
      RECT  221400.0 1924800.0 231600.0 1911000.0 ;
      RECT  221400.0 1924800.0 231600.0 1938600.0 ;
      RECT  221400.0 1952400.0 231600.0 1938600.0 ;
      RECT  221400.0 1952400.0 231600.0 1966200.0 ;
      RECT  221400.0 1980000.0 231600.0 1966200.0 ;
      RECT  221400.0 1980000.0 231600.0 1993800.0 ;
      RECT  221400.0 2007600.0 231600.0 1993800.0 ;
      RECT  221400.0 2007600.0 231600.0 2021400.0 ;
      RECT  221400.0 2035200.0 231600.0 2021400.0 ;
      RECT  221400.0 2035200.0 231600.0 2049000.0 ;
      RECT  221400.0 2062800.0 231600.0 2049000.0 ;
      RECT  221400.0 2062800.0 231600.0 2076600.0 ;
      RECT  221400.0 2090400.0 231600.0 2076600.0 ;
      RECT  221400.0 2090400.0 231600.0 2104200.0 ;
      RECT  221400.0 2118000.0 231600.0 2104200.0 ;
      RECT  221400.0 2118000.0 231600.0 2131800.0 ;
      RECT  221400.0 2145600.0 231600.0 2131800.0 ;
      RECT  231600.0 379200.0 241800.0 393000.0 ;
      RECT  231600.0 406800.0 241800.0 393000.0 ;
      RECT  231600.0 406800.0 241800.0 420600.0 ;
      RECT  231600.0 434400.0 241800.0 420600.0 ;
      RECT  231600.0 434400.0 241800.0 448200.0 ;
      RECT  231600.0 462000.0 241800.0 448200.0 ;
      RECT  231600.0 462000.0 241800.0 475800.0 ;
      RECT  231600.0 489600.0 241800.0 475800.0 ;
      RECT  231600.0 489600.0 241800.0 503400.0 ;
      RECT  231600.0 517200.0 241800.0 503400.0 ;
      RECT  231600.0 517200.0 241800.0 531000.0 ;
      RECT  231600.0 544800.0 241800.0 531000.0 ;
      RECT  231600.0 544800.0 241800.0 558600.0 ;
      RECT  231600.0 572400.0 241800.0 558600.0 ;
      RECT  231600.0 572400.0 241800.0 586200.0 ;
      RECT  231600.0 600000.0 241800.0 586200.0 ;
      RECT  231600.0 600000.0 241800.0 613800.0 ;
      RECT  231600.0 627600.0 241800.0 613800.0 ;
      RECT  231600.0 627600.0 241800.0 641400.0 ;
      RECT  231600.0 655200.0 241800.0 641400.0 ;
      RECT  231600.0 655200.0 241800.0 669000.0 ;
      RECT  231600.0 682800.0 241800.0 669000.0 ;
      RECT  231600.0 682800.0 241800.0 696600.0 ;
      RECT  231600.0 710400.0 241800.0 696600.0 ;
      RECT  231600.0 710400.0 241800.0 724200.0 ;
      RECT  231600.0 738000.0 241800.0 724200.0 ;
      RECT  231600.0 738000.0 241800.0 751800.0 ;
      RECT  231600.0 765600.0 241800.0 751800.0 ;
      RECT  231600.0 765600.0 241800.0 779400.0 ;
      RECT  231600.0 793200.0 241800.0 779400.0 ;
      RECT  231600.0 793200.0 241800.0 807000.0 ;
      RECT  231600.0 820800.0 241800.0 807000.0 ;
      RECT  231600.0 820800.0 241800.0 834600.0 ;
      RECT  231600.0 848400.0 241800.0 834600.0 ;
      RECT  231600.0 848400.0 241800.0 862200.0 ;
      RECT  231600.0 876000.0 241800.0 862200.0 ;
      RECT  231600.0 876000.0 241800.0 889800.0 ;
      RECT  231600.0 903600.0 241800.0 889800.0 ;
      RECT  231600.0 903600.0 241800.0 917400.0 ;
      RECT  231600.0 931200.0 241800.0 917400.0 ;
      RECT  231600.0 931200.0 241800.0 945000.0 ;
      RECT  231600.0 958800.0 241800.0 945000.0 ;
      RECT  231600.0 958800.0 241800.0 972600.0 ;
      RECT  231600.0 986400.0 241800.0 972600.0 ;
      RECT  231600.0 986400.0 241800.0 1000200.0 ;
      RECT  231600.0 1014000.0 241800.0 1000200.0 ;
      RECT  231600.0 1014000.0 241800.0 1027800.0 ;
      RECT  231600.0 1041600.0 241800.0 1027800.0 ;
      RECT  231600.0 1041600.0 241800.0 1055400.0 ;
      RECT  231600.0 1069200.0 241800.0 1055400.0 ;
      RECT  231600.0 1069200.0 241800.0 1083000.0 ;
      RECT  231600.0 1096800.0 241800.0 1083000.0 ;
      RECT  231600.0 1096800.0 241800.0 1110600.0 ;
      RECT  231600.0 1124400.0 241800.0 1110600.0 ;
      RECT  231600.0 1124400.0 241800.0 1138200.0 ;
      RECT  231600.0 1152000.0 241800.0 1138200.0 ;
      RECT  231600.0 1152000.0 241800.0 1165800.0 ;
      RECT  231600.0 1179600.0 241800.0 1165800.0 ;
      RECT  231600.0 1179600.0 241800.0 1193400.0 ;
      RECT  231600.0 1207200.0 241800.0 1193400.0 ;
      RECT  231600.0 1207200.0 241800.0 1221000.0 ;
      RECT  231600.0 1234800.0 241800.0 1221000.0 ;
      RECT  231600.0 1234800.0 241800.0 1248600.0 ;
      RECT  231600.0 1262400.0 241800.0 1248600.0 ;
      RECT  231600.0 1262400.0 241800.0 1276200.0 ;
      RECT  231600.0 1290000.0 241800.0 1276200.0 ;
      RECT  231600.0 1290000.0 241800.0 1303800.0 ;
      RECT  231600.0 1317600.0 241800.0 1303800.0 ;
      RECT  231600.0 1317600.0 241800.0 1331400.0 ;
      RECT  231600.0 1345200.0 241800.0 1331400.0 ;
      RECT  231600.0 1345200.0 241800.0 1359000.0 ;
      RECT  231600.0 1372800.0 241800.0 1359000.0 ;
      RECT  231600.0 1372800.0 241800.0 1386600.0 ;
      RECT  231600.0 1400400.0 241800.0 1386600.0 ;
      RECT  231600.0 1400400.0 241800.0 1414200.0 ;
      RECT  231600.0 1428000.0 241800.0 1414200.0 ;
      RECT  231600.0 1428000.0 241800.0 1441800.0 ;
      RECT  231600.0 1455600.0 241800.0 1441800.0 ;
      RECT  231600.0 1455600.0 241800.0 1469400.0 ;
      RECT  231600.0 1483200.0 241800.0 1469400.0 ;
      RECT  231600.0 1483200.0 241800.0 1497000.0 ;
      RECT  231600.0 1510800.0 241800.0 1497000.0 ;
      RECT  231600.0 1510800.0 241800.0 1524600.0 ;
      RECT  231600.0 1538400.0 241800.0 1524600.0 ;
      RECT  231600.0 1538400.0 241800.0 1552200.0 ;
      RECT  231600.0 1566000.0 241800.0 1552200.0 ;
      RECT  231600.0 1566000.0 241800.0 1579800.0 ;
      RECT  231600.0 1593600.0 241800.0 1579800.0 ;
      RECT  231600.0 1593600.0 241800.0 1607400.0 ;
      RECT  231600.0 1621200.0 241800.0 1607400.0 ;
      RECT  231600.0 1621200.0 241800.0 1635000.0 ;
      RECT  231600.0 1648800.0 241800.0 1635000.0 ;
      RECT  231600.0 1648800.0 241800.0 1662600.0 ;
      RECT  231600.0 1676400.0 241800.0 1662600.0 ;
      RECT  231600.0 1676400.0 241800.0 1690200.0 ;
      RECT  231600.0 1704000.0 241800.0 1690200.0 ;
      RECT  231600.0 1704000.0 241800.0 1717800.0 ;
      RECT  231600.0 1731600.0 241800.0 1717800.0 ;
      RECT  231600.0 1731600.0 241800.0 1745400.0 ;
      RECT  231600.0 1759200.0 241800.0 1745400.0 ;
      RECT  231600.0 1759200.0 241800.0 1773000.0 ;
      RECT  231600.0 1786800.0 241800.0 1773000.0 ;
      RECT  231600.0 1786800.0 241800.0 1800600.0 ;
      RECT  231600.0 1814400.0 241800.0 1800600.0 ;
      RECT  231600.0 1814400.0 241800.0 1828200.0 ;
      RECT  231600.0 1842000.0 241800.0 1828200.0 ;
      RECT  231600.0 1842000.0 241800.0 1855800.0 ;
      RECT  231600.0 1869600.0 241800.0 1855800.0 ;
      RECT  231600.0 1869600.0 241800.0 1883400.0 ;
      RECT  231600.0 1897200.0 241800.0 1883400.0 ;
      RECT  231600.0 1897200.0 241800.0 1911000.0 ;
      RECT  231600.0 1924800.0 241800.0 1911000.0 ;
      RECT  231600.0 1924800.0 241800.0 1938600.0 ;
      RECT  231600.0 1952400.0 241800.0 1938600.0 ;
      RECT  231600.0 1952400.0 241800.0 1966200.0 ;
      RECT  231600.0 1980000.0 241800.0 1966200.0 ;
      RECT  231600.0 1980000.0 241800.0 1993800.0 ;
      RECT  231600.0 2007600.0 241800.0 1993800.0 ;
      RECT  231600.0 2007600.0 241800.0 2021400.0 ;
      RECT  231600.0 2035200.0 241800.0 2021400.0 ;
      RECT  231600.0 2035200.0 241800.0 2049000.0 ;
      RECT  231600.0 2062800.0 241800.0 2049000.0 ;
      RECT  231600.0 2062800.0 241800.0 2076600.0 ;
      RECT  231600.0 2090400.0 241800.0 2076600.0 ;
      RECT  231600.0 2090400.0 241800.0 2104200.0 ;
      RECT  231600.0 2118000.0 241800.0 2104200.0 ;
      RECT  231600.0 2118000.0 241800.0 2131800.0 ;
      RECT  231600.0 2145600.0 241800.0 2131800.0 ;
      RECT  241800.0 379200.0 252000.0 393000.0 ;
      RECT  241800.0 406800.0 252000.0 393000.0 ;
      RECT  241800.0 406800.0 252000.0 420600.0 ;
      RECT  241800.0 434400.0 252000.0 420600.0 ;
      RECT  241800.0 434400.0 252000.0 448200.0 ;
      RECT  241800.0 462000.0 252000.0 448200.0 ;
      RECT  241800.0 462000.0 252000.0 475800.0 ;
      RECT  241800.0 489600.0 252000.0 475800.0 ;
      RECT  241800.0 489600.0 252000.0 503400.0 ;
      RECT  241800.0 517200.0 252000.0 503400.0 ;
      RECT  241800.0 517200.0 252000.0 531000.0 ;
      RECT  241800.0 544800.0 252000.0 531000.0 ;
      RECT  241800.0 544800.0 252000.0 558600.0 ;
      RECT  241800.0 572400.0 252000.0 558600.0 ;
      RECT  241800.0 572400.0 252000.0 586200.0 ;
      RECT  241800.0 600000.0 252000.0 586200.0 ;
      RECT  241800.0 600000.0 252000.0 613800.0 ;
      RECT  241800.0 627600.0 252000.0 613800.0 ;
      RECT  241800.0 627600.0 252000.0 641400.0 ;
      RECT  241800.0 655200.0 252000.0 641400.0 ;
      RECT  241800.0 655200.0 252000.0 669000.0 ;
      RECT  241800.0 682800.0 252000.0 669000.0 ;
      RECT  241800.0 682800.0 252000.0 696600.0 ;
      RECT  241800.0 710400.0 252000.0 696600.0 ;
      RECT  241800.0 710400.0 252000.0 724200.0 ;
      RECT  241800.0 738000.0 252000.0 724200.0 ;
      RECT  241800.0 738000.0 252000.0 751800.0 ;
      RECT  241800.0 765600.0 252000.0 751800.0 ;
      RECT  241800.0 765600.0 252000.0 779400.0 ;
      RECT  241800.0 793200.0 252000.0 779400.0 ;
      RECT  241800.0 793200.0 252000.0 807000.0 ;
      RECT  241800.0 820800.0 252000.0 807000.0 ;
      RECT  241800.0 820800.0 252000.0 834600.0 ;
      RECT  241800.0 848400.0 252000.0 834600.0 ;
      RECT  241800.0 848400.0 252000.0 862200.0 ;
      RECT  241800.0 876000.0 252000.0 862200.0 ;
      RECT  241800.0 876000.0 252000.0 889800.0 ;
      RECT  241800.0 903600.0 252000.0 889800.0 ;
      RECT  241800.0 903600.0 252000.0 917400.0 ;
      RECT  241800.0 931200.0 252000.0 917400.0 ;
      RECT  241800.0 931200.0 252000.0 945000.0 ;
      RECT  241800.0 958800.0 252000.0 945000.0 ;
      RECT  241800.0 958800.0 252000.0 972600.0 ;
      RECT  241800.0 986400.0 252000.0 972600.0 ;
      RECT  241800.0 986400.0 252000.0 1000200.0 ;
      RECT  241800.0 1014000.0 252000.0 1000200.0 ;
      RECT  241800.0 1014000.0 252000.0 1027800.0 ;
      RECT  241800.0 1041600.0 252000.0 1027800.0 ;
      RECT  241800.0 1041600.0 252000.0 1055400.0 ;
      RECT  241800.0 1069200.0 252000.0 1055400.0 ;
      RECT  241800.0 1069200.0 252000.0 1083000.0 ;
      RECT  241800.0 1096800.0 252000.0 1083000.0 ;
      RECT  241800.0 1096800.0 252000.0 1110600.0 ;
      RECT  241800.0 1124400.0 252000.0 1110600.0 ;
      RECT  241800.0 1124400.0 252000.0 1138200.0 ;
      RECT  241800.0 1152000.0 252000.0 1138200.0 ;
      RECT  241800.0 1152000.0 252000.0 1165800.0 ;
      RECT  241800.0 1179600.0 252000.0 1165800.0 ;
      RECT  241800.0 1179600.0 252000.0 1193400.0 ;
      RECT  241800.0 1207200.0 252000.0 1193400.0 ;
      RECT  241800.0 1207200.0 252000.0 1221000.0 ;
      RECT  241800.0 1234800.0 252000.0 1221000.0 ;
      RECT  241800.0 1234800.0 252000.0 1248600.0 ;
      RECT  241800.0 1262400.0 252000.0 1248600.0 ;
      RECT  241800.0 1262400.0 252000.0 1276200.0 ;
      RECT  241800.0 1290000.0 252000.0 1276200.0 ;
      RECT  241800.0 1290000.0 252000.0 1303800.0 ;
      RECT  241800.0 1317600.0 252000.0 1303800.0 ;
      RECT  241800.0 1317600.0 252000.0 1331400.0 ;
      RECT  241800.0 1345200.0 252000.0 1331400.0 ;
      RECT  241800.0 1345200.0 252000.0 1359000.0 ;
      RECT  241800.0 1372800.0 252000.0 1359000.0 ;
      RECT  241800.0 1372800.0 252000.0 1386600.0 ;
      RECT  241800.0 1400400.0 252000.0 1386600.0 ;
      RECT  241800.0 1400400.0 252000.0 1414200.0 ;
      RECT  241800.0 1428000.0 252000.0 1414200.0 ;
      RECT  241800.0 1428000.0 252000.0 1441800.0 ;
      RECT  241800.0 1455600.0 252000.0 1441800.0 ;
      RECT  241800.0 1455600.0 252000.0 1469400.0 ;
      RECT  241800.0 1483200.0 252000.0 1469400.0 ;
      RECT  241800.0 1483200.0 252000.0 1497000.0 ;
      RECT  241800.0 1510800.0 252000.0 1497000.0 ;
      RECT  241800.0 1510800.0 252000.0 1524600.0 ;
      RECT  241800.0 1538400.0 252000.0 1524600.0 ;
      RECT  241800.0 1538400.0 252000.0 1552200.0 ;
      RECT  241800.0 1566000.0 252000.0 1552200.0 ;
      RECT  241800.0 1566000.0 252000.0 1579800.0 ;
      RECT  241800.0 1593600.0 252000.0 1579800.0 ;
      RECT  241800.0 1593600.0 252000.0 1607400.0 ;
      RECT  241800.0 1621200.0 252000.0 1607400.0 ;
      RECT  241800.0 1621200.0 252000.0 1635000.0 ;
      RECT  241800.0 1648800.0 252000.0 1635000.0 ;
      RECT  241800.0 1648800.0 252000.0 1662600.0 ;
      RECT  241800.0 1676400.0 252000.0 1662600.0 ;
      RECT  241800.0 1676400.0 252000.0 1690200.0 ;
      RECT  241800.0 1704000.0 252000.0 1690200.0 ;
      RECT  241800.0 1704000.0 252000.0 1717800.0 ;
      RECT  241800.0 1731600.0 252000.0 1717800.0 ;
      RECT  241800.0 1731600.0 252000.0 1745400.0 ;
      RECT  241800.0 1759200.0 252000.0 1745400.0 ;
      RECT  241800.0 1759200.0 252000.0 1773000.0 ;
      RECT  241800.0 1786800.0 252000.0 1773000.0 ;
      RECT  241800.0 1786800.0 252000.0 1800600.0 ;
      RECT  241800.0 1814400.0 252000.0 1800600.0 ;
      RECT  241800.0 1814400.0 252000.0 1828200.0 ;
      RECT  241800.0 1842000.0 252000.0 1828200.0 ;
      RECT  241800.0 1842000.0 252000.0 1855800.0 ;
      RECT  241800.0 1869600.0 252000.0 1855800.0 ;
      RECT  241800.0 1869600.0 252000.0 1883400.0 ;
      RECT  241800.0 1897200.0 252000.0 1883400.0 ;
      RECT  241800.0 1897200.0 252000.0 1911000.0 ;
      RECT  241800.0 1924800.0 252000.0 1911000.0 ;
      RECT  241800.0 1924800.0 252000.0 1938600.0 ;
      RECT  241800.0 1952400.0 252000.0 1938600.0 ;
      RECT  241800.0 1952400.0 252000.0 1966200.0 ;
      RECT  241800.0 1980000.0 252000.0 1966200.0 ;
      RECT  241800.0 1980000.0 252000.0 1993800.0 ;
      RECT  241800.0 2007600.0 252000.0 1993800.0 ;
      RECT  241800.0 2007600.0 252000.0 2021400.0 ;
      RECT  241800.0 2035200.0 252000.0 2021400.0 ;
      RECT  241800.0 2035200.0 252000.0 2049000.0 ;
      RECT  241800.0 2062800.0 252000.0 2049000.0 ;
      RECT  241800.0 2062800.0 252000.0 2076600.0 ;
      RECT  241800.0 2090400.0 252000.0 2076600.0 ;
      RECT  241800.0 2090400.0 252000.0 2104200.0 ;
      RECT  241800.0 2118000.0 252000.0 2104200.0 ;
      RECT  241800.0 2118000.0 252000.0 2131800.0 ;
      RECT  241800.0 2145600.0 252000.0 2131800.0 ;
      RECT  252000.0 379200.0 262200.0 393000.0 ;
      RECT  252000.0 406800.0 262200.0 393000.0 ;
      RECT  252000.0 406800.0 262200.0 420600.0 ;
      RECT  252000.0 434400.0 262200.0 420600.0 ;
      RECT  252000.0 434400.0 262200.0 448200.0 ;
      RECT  252000.0 462000.0 262200.0 448200.0 ;
      RECT  252000.0 462000.0 262200.0 475800.0 ;
      RECT  252000.0 489600.0 262200.0 475800.0 ;
      RECT  252000.0 489600.0 262200.0 503400.0 ;
      RECT  252000.0 517200.0 262200.0 503400.0 ;
      RECT  252000.0 517200.0 262200.0 531000.0 ;
      RECT  252000.0 544800.0 262200.0 531000.0 ;
      RECT  252000.0 544800.0 262200.0 558600.0 ;
      RECT  252000.0 572400.0 262200.0 558600.0 ;
      RECT  252000.0 572400.0 262200.0 586200.0 ;
      RECT  252000.0 600000.0 262200.0 586200.0 ;
      RECT  252000.0 600000.0 262200.0 613800.0 ;
      RECT  252000.0 627600.0 262200.0 613800.0 ;
      RECT  252000.0 627600.0 262200.0 641400.0 ;
      RECT  252000.0 655200.0 262200.0 641400.0 ;
      RECT  252000.0 655200.0 262200.0 669000.0 ;
      RECT  252000.0 682800.0 262200.0 669000.0 ;
      RECT  252000.0 682800.0 262200.0 696600.0 ;
      RECT  252000.0 710400.0 262200.0 696600.0 ;
      RECT  252000.0 710400.0 262200.0 724200.0 ;
      RECT  252000.0 738000.0 262200.0 724200.0 ;
      RECT  252000.0 738000.0 262200.0 751800.0 ;
      RECT  252000.0 765600.0 262200.0 751800.0 ;
      RECT  252000.0 765600.0 262200.0 779400.0 ;
      RECT  252000.0 793200.0 262200.0 779400.0 ;
      RECT  252000.0 793200.0 262200.0 807000.0 ;
      RECT  252000.0 820800.0 262200.0 807000.0 ;
      RECT  252000.0 820800.0 262200.0 834600.0 ;
      RECT  252000.0 848400.0 262200.0 834600.0 ;
      RECT  252000.0 848400.0 262200.0 862200.0 ;
      RECT  252000.0 876000.0 262200.0 862200.0 ;
      RECT  252000.0 876000.0 262200.0 889800.0 ;
      RECT  252000.0 903600.0 262200.0 889800.0 ;
      RECT  252000.0 903600.0 262200.0 917400.0 ;
      RECT  252000.0 931200.0 262200.0 917400.0 ;
      RECT  252000.0 931200.0 262200.0 945000.0 ;
      RECT  252000.0 958800.0 262200.0 945000.0 ;
      RECT  252000.0 958800.0 262200.0 972600.0 ;
      RECT  252000.0 986400.0 262200.0 972600.0 ;
      RECT  252000.0 986400.0 262200.0 1000200.0 ;
      RECT  252000.0 1014000.0 262200.0 1000200.0 ;
      RECT  252000.0 1014000.0 262200.0 1027800.0 ;
      RECT  252000.0 1041600.0 262200.0 1027800.0 ;
      RECT  252000.0 1041600.0 262200.0 1055400.0 ;
      RECT  252000.0 1069200.0 262200.0 1055400.0 ;
      RECT  252000.0 1069200.0 262200.0 1083000.0 ;
      RECT  252000.0 1096800.0 262200.0 1083000.0 ;
      RECT  252000.0 1096800.0 262200.0 1110600.0 ;
      RECT  252000.0 1124400.0 262200.0 1110600.0 ;
      RECT  252000.0 1124400.0 262200.0 1138200.0 ;
      RECT  252000.0 1152000.0 262200.0 1138200.0 ;
      RECT  252000.0 1152000.0 262200.0 1165800.0 ;
      RECT  252000.0 1179600.0 262200.0 1165800.0 ;
      RECT  252000.0 1179600.0 262200.0 1193400.0 ;
      RECT  252000.0 1207200.0 262200.0 1193400.0 ;
      RECT  252000.0 1207200.0 262200.0 1221000.0 ;
      RECT  252000.0 1234800.0 262200.0 1221000.0 ;
      RECT  252000.0 1234800.0 262200.0 1248600.0 ;
      RECT  252000.0 1262400.0 262200.0 1248600.0 ;
      RECT  252000.0 1262400.0 262200.0 1276200.0 ;
      RECT  252000.0 1290000.0 262200.0 1276200.0 ;
      RECT  252000.0 1290000.0 262200.0 1303800.0 ;
      RECT  252000.0 1317600.0 262200.0 1303800.0 ;
      RECT  252000.0 1317600.0 262200.0 1331400.0 ;
      RECT  252000.0 1345200.0 262200.0 1331400.0 ;
      RECT  252000.0 1345200.0 262200.0 1359000.0 ;
      RECT  252000.0 1372800.0 262200.0 1359000.0 ;
      RECT  252000.0 1372800.0 262200.0 1386600.0 ;
      RECT  252000.0 1400400.0 262200.0 1386600.0 ;
      RECT  252000.0 1400400.0 262200.0 1414200.0 ;
      RECT  252000.0 1428000.0 262200.0 1414200.0 ;
      RECT  252000.0 1428000.0 262200.0 1441800.0 ;
      RECT  252000.0 1455600.0 262200.0 1441800.0 ;
      RECT  252000.0 1455600.0 262200.0 1469400.0 ;
      RECT  252000.0 1483200.0 262200.0 1469400.0 ;
      RECT  252000.0 1483200.0 262200.0 1497000.0 ;
      RECT  252000.0 1510800.0 262200.0 1497000.0 ;
      RECT  252000.0 1510800.0 262200.0 1524600.0 ;
      RECT  252000.0 1538400.0 262200.0 1524600.0 ;
      RECT  252000.0 1538400.0 262200.0 1552200.0 ;
      RECT  252000.0 1566000.0 262200.0 1552200.0 ;
      RECT  252000.0 1566000.0 262200.0 1579800.0 ;
      RECT  252000.0 1593600.0 262200.0 1579800.0 ;
      RECT  252000.0 1593600.0 262200.0 1607400.0 ;
      RECT  252000.0 1621200.0 262200.0 1607400.0 ;
      RECT  252000.0 1621200.0 262200.0 1635000.0 ;
      RECT  252000.0 1648800.0 262200.0 1635000.0 ;
      RECT  252000.0 1648800.0 262200.0 1662600.0 ;
      RECT  252000.0 1676400.0 262200.0 1662600.0 ;
      RECT  252000.0 1676400.0 262200.0 1690200.0 ;
      RECT  252000.0 1704000.0 262200.0 1690200.0 ;
      RECT  252000.0 1704000.0 262200.0 1717800.0 ;
      RECT  252000.0 1731600.0 262200.0 1717800.0 ;
      RECT  252000.0 1731600.0 262200.0 1745400.0 ;
      RECT  252000.0 1759200.0 262200.0 1745400.0 ;
      RECT  252000.0 1759200.0 262200.0 1773000.0 ;
      RECT  252000.0 1786800.0 262200.0 1773000.0 ;
      RECT  252000.0 1786800.0 262200.0 1800600.0 ;
      RECT  252000.0 1814400.0 262200.0 1800600.0 ;
      RECT  252000.0 1814400.0 262200.0 1828200.0 ;
      RECT  252000.0 1842000.0 262200.0 1828200.0 ;
      RECT  252000.0 1842000.0 262200.0 1855800.0 ;
      RECT  252000.0 1869600.0 262200.0 1855800.0 ;
      RECT  252000.0 1869600.0 262200.0 1883400.0 ;
      RECT  252000.0 1897200.0 262200.0 1883400.0 ;
      RECT  252000.0 1897200.0 262200.0 1911000.0 ;
      RECT  252000.0 1924800.0 262200.0 1911000.0 ;
      RECT  252000.0 1924800.0 262200.0 1938600.0 ;
      RECT  252000.0 1952400.0 262200.0 1938600.0 ;
      RECT  252000.0 1952400.0 262200.0 1966200.0 ;
      RECT  252000.0 1980000.0 262200.0 1966200.0 ;
      RECT  252000.0 1980000.0 262200.0 1993800.0 ;
      RECT  252000.0 2007600.0 262200.0 1993800.0 ;
      RECT  252000.0 2007600.0 262200.0 2021400.0 ;
      RECT  252000.0 2035200.0 262200.0 2021400.0 ;
      RECT  252000.0 2035200.0 262200.0 2049000.0 ;
      RECT  252000.0 2062800.0 262200.0 2049000.0 ;
      RECT  252000.0 2062800.0 262200.0 2076600.0 ;
      RECT  252000.0 2090400.0 262200.0 2076600.0 ;
      RECT  252000.0 2090400.0 262200.0 2104200.0 ;
      RECT  252000.0 2118000.0 262200.0 2104200.0 ;
      RECT  252000.0 2118000.0 262200.0 2131800.0 ;
      RECT  252000.0 2145600.0 262200.0 2131800.0 ;
      RECT  262200.0 379200.0 272400.0 393000.0 ;
      RECT  262200.0 406800.0 272400.0 393000.0 ;
      RECT  262200.0 406800.0 272400.0 420600.0 ;
      RECT  262200.0 434400.0 272400.0 420600.0 ;
      RECT  262200.0 434400.0 272400.0 448200.0 ;
      RECT  262200.0 462000.0 272400.0 448200.0 ;
      RECT  262200.0 462000.0 272400.0 475800.0 ;
      RECT  262200.0 489600.0 272400.0 475800.0 ;
      RECT  262200.0 489600.0 272400.0 503400.0 ;
      RECT  262200.0 517200.0 272400.0 503400.0 ;
      RECT  262200.0 517200.0 272400.0 531000.0 ;
      RECT  262200.0 544800.0 272400.0 531000.0 ;
      RECT  262200.0 544800.0 272400.0 558600.0 ;
      RECT  262200.0 572400.0 272400.0 558600.0 ;
      RECT  262200.0 572400.0 272400.0 586200.0 ;
      RECT  262200.0 600000.0 272400.0 586200.0 ;
      RECT  262200.0 600000.0 272400.0 613800.0 ;
      RECT  262200.0 627600.0 272400.0 613800.0 ;
      RECT  262200.0 627600.0 272400.0 641400.0 ;
      RECT  262200.0 655200.0 272400.0 641400.0 ;
      RECT  262200.0 655200.0 272400.0 669000.0 ;
      RECT  262200.0 682800.0 272400.0 669000.0 ;
      RECT  262200.0 682800.0 272400.0 696600.0 ;
      RECT  262200.0 710400.0 272400.0 696600.0 ;
      RECT  262200.0 710400.0 272400.0 724200.0 ;
      RECT  262200.0 738000.0 272400.0 724200.0 ;
      RECT  262200.0 738000.0 272400.0 751800.0 ;
      RECT  262200.0 765600.0 272400.0 751800.0 ;
      RECT  262200.0 765600.0 272400.0 779400.0 ;
      RECT  262200.0 793200.0 272400.0 779400.0 ;
      RECT  262200.0 793200.0 272400.0 807000.0 ;
      RECT  262200.0 820800.0 272400.0 807000.0 ;
      RECT  262200.0 820800.0 272400.0 834600.0 ;
      RECT  262200.0 848400.0 272400.0 834600.0 ;
      RECT  262200.0 848400.0 272400.0 862200.0 ;
      RECT  262200.0 876000.0 272400.0 862200.0 ;
      RECT  262200.0 876000.0 272400.0 889800.0 ;
      RECT  262200.0 903600.0 272400.0 889800.0 ;
      RECT  262200.0 903600.0 272400.0 917400.0 ;
      RECT  262200.0 931200.0 272400.0 917400.0 ;
      RECT  262200.0 931200.0 272400.0 945000.0 ;
      RECT  262200.0 958800.0 272400.0 945000.0 ;
      RECT  262200.0 958800.0 272400.0 972600.0 ;
      RECT  262200.0 986400.0 272400.0 972600.0 ;
      RECT  262200.0 986400.0 272400.0 1000200.0 ;
      RECT  262200.0 1014000.0 272400.0 1000200.0 ;
      RECT  262200.0 1014000.0 272400.0 1027800.0 ;
      RECT  262200.0 1041600.0 272400.0 1027800.0 ;
      RECT  262200.0 1041600.0 272400.0 1055400.0 ;
      RECT  262200.0 1069200.0 272400.0 1055400.0 ;
      RECT  262200.0 1069200.0 272400.0 1083000.0 ;
      RECT  262200.0 1096800.0 272400.0 1083000.0 ;
      RECT  262200.0 1096800.0 272400.0 1110600.0 ;
      RECT  262200.0 1124400.0 272400.0 1110600.0 ;
      RECT  262200.0 1124400.0 272400.0 1138200.0 ;
      RECT  262200.0 1152000.0 272400.0 1138200.0 ;
      RECT  262200.0 1152000.0 272400.0 1165800.0 ;
      RECT  262200.0 1179600.0 272400.0 1165800.0 ;
      RECT  262200.0 1179600.0 272400.0 1193400.0 ;
      RECT  262200.0 1207200.0 272400.0 1193400.0 ;
      RECT  262200.0 1207200.0 272400.0 1221000.0 ;
      RECT  262200.0 1234800.0 272400.0 1221000.0 ;
      RECT  262200.0 1234800.0 272400.0 1248600.0 ;
      RECT  262200.0 1262400.0 272400.0 1248600.0 ;
      RECT  262200.0 1262400.0 272400.0 1276200.0 ;
      RECT  262200.0 1290000.0 272400.0 1276200.0 ;
      RECT  262200.0 1290000.0 272400.0 1303800.0 ;
      RECT  262200.0 1317600.0 272400.0 1303800.0 ;
      RECT  262200.0 1317600.0 272400.0 1331400.0 ;
      RECT  262200.0 1345200.0 272400.0 1331400.0 ;
      RECT  262200.0 1345200.0 272400.0 1359000.0 ;
      RECT  262200.0 1372800.0 272400.0 1359000.0 ;
      RECT  262200.0 1372800.0 272400.0 1386600.0 ;
      RECT  262200.0 1400400.0 272400.0 1386600.0 ;
      RECT  262200.0 1400400.0 272400.0 1414200.0 ;
      RECT  262200.0 1428000.0 272400.0 1414200.0 ;
      RECT  262200.0 1428000.0 272400.0 1441800.0 ;
      RECT  262200.0 1455600.0 272400.0 1441800.0 ;
      RECT  262200.0 1455600.0 272400.0 1469400.0 ;
      RECT  262200.0 1483200.0 272400.0 1469400.0 ;
      RECT  262200.0 1483200.0 272400.0 1497000.0 ;
      RECT  262200.0 1510800.0 272400.0 1497000.0 ;
      RECT  262200.0 1510800.0 272400.0 1524600.0 ;
      RECT  262200.0 1538400.0 272400.0 1524600.0 ;
      RECT  262200.0 1538400.0 272400.0 1552200.0 ;
      RECT  262200.0 1566000.0 272400.0 1552200.0 ;
      RECT  262200.0 1566000.0 272400.0 1579800.0 ;
      RECT  262200.0 1593600.0 272400.0 1579800.0 ;
      RECT  262200.0 1593600.0 272400.0 1607400.0 ;
      RECT  262200.0 1621200.0 272400.0 1607400.0 ;
      RECT  262200.0 1621200.0 272400.0 1635000.0 ;
      RECT  262200.0 1648800.0 272400.0 1635000.0 ;
      RECT  262200.0 1648800.0 272400.0 1662600.0 ;
      RECT  262200.0 1676400.0 272400.0 1662600.0 ;
      RECT  262200.0 1676400.0 272400.0 1690200.0 ;
      RECT  262200.0 1704000.0 272400.0 1690200.0 ;
      RECT  262200.0 1704000.0 272400.0 1717800.0 ;
      RECT  262200.0 1731600.0 272400.0 1717800.0 ;
      RECT  262200.0 1731600.0 272400.0 1745400.0 ;
      RECT  262200.0 1759200.0 272400.0 1745400.0 ;
      RECT  262200.0 1759200.0 272400.0 1773000.0 ;
      RECT  262200.0 1786800.0 272400.0 1773000.0 ;
      RECT  262200.0 1786800.0 272400.0 1800600.0 ;
      RECT  262200.0 1814400.0 272400.0 1800600.0 ;
      RECT  262200.0 1814400.0 272400.0 1828200.0 ;
      RECT  262200.0 1842000.0 272400.0 1828200.0 ;
      RECT  262200.0 1842000.0 272400.0 1855800.0 ;
      RECT  262200.0 1869600.0 272400.0 1855800.0 ;
      RECT  262200.0 1869600.0 272400.0 1883400.0 ;
      RECT  262200.0 1897200.0 272400.0 1883400.0 ;
      RECT  262200.0 1897200.0 272400.0 1911000.0 ;
      RECT  262200.0 1924800.0 272400.0 1911000.0 ;
      RECT  262200.0 1924800.0 272400.0 1938600.0 ;
      RECT  262200.0 1952400.0 272400.0 1938600.0 ;
      RECT  262200.0 1952400.0 272400.0 1966200.0 ;
      RECT  262200.0 1980000.0 272400.0 1966200.0 ;
      RECT  262200.0 1980000.0 272400.0 1993800.0 ;
      RECT  262200.0 2007600.0 272400.0 1993800.0 ;
      RECT  262200.0 2007600.0 272400.0 2021400.0 ;
      RECT  262200.0 2035200.0 272400.0 2021400.0 ;
      RECT  262200.0 2035200.0 272400.0 2049000.0 ;
      RECT  262200.0 2062800.0 272400.0 2049000.0 ;
      RECT  262200.0 2062800.0 272400.0 2076600.0 ;
      RECT  262200.0 2090400.0 272400.0 2076600.0 ;
      RECT  262200.0 2090400.0 272400.0 2104200.0 ;
      RECT  262200.0 2118000.0 272400.0 2104200.0 ;
      RECT  262200.0 2118000.0 272400.0 2131800.0 ;
      RECT  262200.0 2145600.0 272400.0 2131800.0 ;
      RECT  272400.0 379200.0 282600.0 393000.0 ;
      RECT  272400.0 406800.0 282600.0 393000.0 ;
      RECT  272400.0 406800.0 282600.0 420600.0 ;
      RECT  272400.0 434400.0 282600.0 420600.0 ;
      RECT  272400.0 434400.0 282600.0 448200.0 ;
      RECT  272400.0 462000.0 282600.0 448200.0 ;
      RECT  272400.0 462000.0 282600.0 475800.0 ;
      RECT  272400.0 489600.0 282600.0 475800.0 ;
      RECT  272400.0 489600.0 282600.0 503400.0 ;
      RECT  272400.0 517200.0 282600.0 503400.0 ;
      RECT  272400.0 517200.0 282600.0 531000.0 ;
      RECT  272400.0 544800.0 282600.0 531000.0 ;
      RECT  272400.0 544800.0 282600.0 558600.0 ;
      RECT  272400.0 572400.0 282600.0 558600.0 ;
      RECT  272400.0 572400.0 282600.0 586200.0 ;
      RECT  272400.0 600000.0 282600.0 586200.0 ;
      RECT  272400.0 600000.0 282600.0 613800.0 ;
      RECT  272400.0 627600.0 282600.0 613800.0 ;
      RECT  272400.0 627600.0 282600.0 641400.0 ;
      RECT  272400.0 655200.0 282600.0 641400.0 ;
      RECT  272400.0 655200.0 282600.0 669000.0 ;
      RECT  272400.0 682800.0 282600.0 669000.0 ;
      RECT  272400.0 682800.0 282600.0 696600.0 ;
      RECT  272400.0 710400.0 282600.0 696600.0 ;
      RECT  272400.0 710400.0 282600.0 724200.0 ;
      RECT  272400.0 738000.0 282600.0 724200.0 ;
      RECT  272400.0 738000.0 282600.0 751800.0 ;
      RECT  272400.0 765600.0 282600.0 751800.0 ;
      RECT  272400.0 765600.0 282600.0 779400.0 ;
      RECT  272400.0 793200.0 282600.0 779400.0 ;
      RECT  272400.0 793200.0 282600.0 807000.0 ;
      RECT  272400.0 820800.0 282600.0 807000.0 ;
      RECT  272400.0 820800.0 282600.0 834600.0 ;
      RECT  272400.0 848400.0 282600.0 834600.0 ;
      RECT  272400.0 848400.0 282600.0 862200.0 ;
      RECT  272400.0 876000.0 282600.0 862200.0 ;
      RECT  272400.0 876000.0 282600.0 889800.0 ;
      RECT  272400.0 903600.0 282600.0 889800.0 ;
      RECT  272400.0 903600.0 282600.0 917400.0 ;
      RECT  272400.0 931200.0 282600.0 917400.0 ;
      RECT  272400.0 931200.0 282600.0 945000.0 ;
      RECT  272400.0 958800.0 282600.0 945000.0 ;
      RECT  272400.0 958800.0 282600.0 972600.0 ;
      RECT  272400.0 986400.0 282600.0 972600.0 ;
      RECT  272400.0 986400.0 282600.0 1000200.0 ;
      RECT  272400.0 1014000.0 282600.0 1000200.0 ;
      RECT  272400.0 1014000.0 282600.0 1027800.0 ;
      RECT  272400.0 1041600.0 282600.0 1027800.0 ;
      RECT  272400.0 1041600.0 282600.0 1055400.0 ;
      RECT  272400.0 1069200.0 282600.0 1055400.0 ;
      RECT  272400.0 1069200.0 282600.0 1083000.0 ;
      RECT  272400.0 1096800.0 282600.0 1083000.0 ;
      RECT  272400.0 1096800.0 282600.0 1110600.0 ;
      RECT  272400.0 1124400.0 282600.0 1110600.0 ;
      RECT  272400.0 1124400.0 282600.0 1138200.0 ;
      RECT  272400.0 1152000.0 282600.0 1138200.0 ;
      RECT  272400.0 1152000.0 282600.0 1165800.0 ;
      RECT  272400.0 1179600.0 282600.0 1165800.0 ;
      RECT  272400.0 1179600.0 282600.0 1193400.0 ;
      RECT  272400.0 1207200.0 282600.0 1193400.0 ;
      RECT  272400.0 1207200.0 282600.0 1221000.0 ;
      RECT  272400.0 1234800.0 282600.0 1221000.0 ;
      RECT  272400.0 1234800.0 282600.0 1248600.0 ;
      RECT  272400.0 1262400.0 282600.0 1248600.0 ;
      RECT  272400.0 1262400.0 282600.0 1276200.0 ;
      RECT  272400.0 1290000.0 282600.0 1276200.0 ;
      RECT  272400.0 1290000.0 282600.0 1303800.0 ;
      RECT  272400.0 1317600.0 282600.0 1303800.0 ;
      RECT  272400.0 1317600.0 282600.0 1331400.0 ;
      RECT  272400.0 1345200.0 282600.0 1331400.0 ;
      RECT  272400.0 1345200.0 282600.0 1359000.0 ;
      RECT  272400.0 1372800.0 282600.0 1359000.0 ;
      RECT  272400.0 1372800.0 282600.0 1386600.0 ;
      RECT  272400.0 1400400.0 282600.0 1386600.0 ;
      RECT  272400.0 1400400.0 282600.0 1414200.0 ;
      RECT  272400.0 1428000.0 282600.0 1414200.0 ;
      RECT  272400.0 1428000.0 282600.0 1441800.0 ;
      RECT  272400.0 1455600.0 282600.0 1441800.0 ;
      RECT  272400.0 1455600.0 282600.0 1469400.0 ;
      RECT  272400.0 1483200.0 282600.0 1469400.0 ;
      RECT  272400.0 1483200.0 282600.0 1497000.0 ;
      RECT  272400.0 1510800.0 282600.0 1497000.0 ;
      RECT  272400.0 1510800.0 282600.0 1524600.0 ;
      RECT  272400.0 1538400.0 282600.0 1524600.0 ;
      RECT  272400.0 1538400.0 282600.0 1552200.0 ;
      RECT  272400.0 1566000.0 282600.0 1552200.0 ;
      RECT  272400.0 1566000.0 282600.0 1579800.0 ;
      RECT  272400.0 1593600.0 282600.0 1579800.0 ;
      RECT  272400.0 1593600.0 282600.0 1607400.0 ;
      RECT  272400.0 1621200.0 282600.0 1607400.0 ;
      RECT  272400.0 1621200.0 282600.0 1635000.0 ;
      RECT  272400.0 1648800.0 282600.0 1635000.0 ;
      RECT  272400.0 1648800.0 282600.0 1662600.0 ;
      RECT  272400.0 1676400.0 282600.0 1662600.0 ;
      RECT  272400.0 1676400.0 282600.0 1690200.0 ;
      RECT  272400.0 1704000.0 282600.0 1690200.0 ;
      RECT  272400.0 1704000.0 282600.0 1717800.0 ;
      RECT  272400.0 1731600.0 282600.0 1717800.0 ;
      RECT  272400.0 1731600.0 282600.0 1745400.0 ;
      RECT  272400.0 1759200.0 282600.0 1745400.0 ;
      RECT  272400.0 1759200.0 282600.0 1773000.0 ;
      RECT  272400.0 1786800.0 282600.0 1773000.0 ;
      RECT  272400.0 1786800.0 282600.0 1800600.0 ;
      RECT  272400.0 1814400.0 282600.0 1800600.0 ;
      RECT  272400.0 1814400.0 282600.0 1828200.0 ;
      RECT  272400.0 1842000.0 282600.0 1828200.0 ;
      RECT  272400.0 1842000.0 282600.0 1855800.0 ;
      RECT  272400.0 1869600.0 282600.0 1855800.0 ;
      RECT  272400.0 1869600.0 282600.0 1883400.0 ;
      RECT  272400.0 1897200.0 282600.0 1883400.0 ;
      RECT  272400.0 1897200.0 282600.0 1911000.0 ;
      RECT  272400.0 1924800.0 282600.0 1911000.0 ;
      RECT  272400.0 1924800.0 282600.0 1938600.0 ;
      RECT  272400.0 1952400.0 282600.0 1938600.0 ;
      RECT  272400.0 1952400.0 282600.0 1966200.0 ;
      RECT  272400.0 1980000.0 282600.0 1966200.0 ;
      RECT  272400.0 1980000.0 282600.0 1993800.0 ;
      RECT  272400.0 2007600.0 282600.0 1993800.0 ;
      RECT  272400.0 2007600.0 282600.0 2021400.0 ;
      RECT  272400.0 2035200.0 282600.0 2021400.0 ;
      RECT  272400.0 2035200.0 282600.0 2049000.0 ;
      RECT  272400.0 2062800.0 282600.0 2049000.0 ;
      RECT  272400.0 2062800.0 282600.0 2076600.0 ;
      RECT  272400.0 2090400.0 282600.0 2076600.0 ;
      RECT  272400.0 2090400.0 282600.0 2104200.0 ;
      RECT  272400.0 2118000.0 282600.0 2104200.0 ;
      RECT  272400.0 2118000.0 282600.0 2131800.0 ;
      RECT  272400.0 2145600.0 282600.0 2131800.0 ;
      RECT  282600.0 379200.0 292800.0 393000.0 ;
      RECT  282600.0 406800.0 292800.0 393000.0 ;
      RECT  282600.0 406800.0 292800.0 420600.0 ;
      RECT  282600.0 434400.0 292800.0 420600.0 ;
      RECT  282600.0 434400.0 292800.0 448200.0 ;
      RECT  282600.0 462000.0 292800.0 448200.0 ;
      RECT  282600.0 462000.0 292800.0 475800.0 ;
      RECT  282600.0 489600.0 292800.0 475800.0 ;
      RECT  282600.0 489600.0 292800.0 503400.0 ;
      RECT  282600.0 517200.0 292800.0 503400.0 ;
      RECT  282600.0 517200.0 292800.0 531000.0 ;
      RECT  282600.0 544800.0 292800.0 531000.0 ;
      RECT  282600.0 544800.0 292800.0 558600.0 ;
      RECT  282600.0 572400.0 292800.0 558600.0 ;
      RECT  282600.0 572400.0 292800.0 586200.0 ;
      RECT  282600.0 600000.0 292800.0 586200.0 ;
      RECT  282600.0 600000.0 292800.0 613800.0 ;
      RECT  282600.0 627600.0 292800.0 613800.0 ;
      RECT  282600.0 627600.0 292800.0 641400.0 ;
      RECT  282600.0 655200.0 292800.0 641400.0 ;
      RECT  282600.0 655200.0 292800.0 669000.0 ;
      RECT  282600.0 682800.0 292800.0 669000.0 ;
      RECT  282600.0 682800.0 292800.0 696600.0 ;
      RECT  282600.0 710400.0 292800.0 696600.0 ;
      RECT  282600.0 710400.0 292800.0 724200.0 ;
      RECT  282600.0 738000.0 292800.0 724200.0 ;
      RECT  282600.0 738000.0 292800.0 751800.0 ;
      RECT  282600.0 765600.0 292800.0 751800.0 ;
      RECT  282600.0 765600.0 292800.0 779400.0 ;
      RECT  282600.0 793200.0 292800.0 779400.0 ;
      RECT  282600.0 793200.0 292800.0 807000.0 ;
      RECT  282600.0 820800.0 292800.0 807000.0 ;
      RECT  282600.0 820800.0 292800.0 834600.0 ;
      RECT  282600.0 848400.0 292800.0 834600.0 ;
      RECT  282600.0 848400.0 292800.0 862200.0 ;
      RECT  282600.0 876000.0 292800.0 862200.0 ;
      RECT  282600.0 876000.0 292800.0 889800.0 ;
      RECT  282600.0 903600.0 292800.0 889800.0 ;
      RECT  282600.0 903600.0 292800.0 917400.0 ;
      RECT  282600.0 931200.0 292800.0 917400.0 ;
      RECT  282600.0 931200.0 292800.0 945000.0 ;
      RECT  282600.0 958800.0 292800.0 945000.0 ;
      RECT  282600.0 958800.0 292800.0 972600.0 ;
      RECT  282600.0 986400.0 292800.0 972600.0 ;
      RECT  282600.0 986400.0 292800.0 1000200.0 ;
      RECT  282600.0 1014000.0 292800.0 1000200.0 ;
      RECT  282600.0 1014000.0 292800.0 1027800.0 ;
      RECT  282600.0 1041600.0 292800.0 1027800.0 ;
      RECT  282600.0 1041600.0 292800.0 1055400.0 ;
      RECT  282600.0 1069200.0 292800.0 1055400.0 ;
      RECT  282600.0 1069200.0 292800.0 1083000.0 ;
      RECT  282600.0 1096800.0 292800.0 1083000.0 ;
      RECT  282600.0 1096800.0 292800.0 1110600.0 ;
      RECT  282600.0 1124400.0 292800.0 1110600.0 ;
      RECT  282600.0 1124400.0 292800.0 1138200.0 ;
      RECT  282600.0 1152000.0 292800.0 1138200.0 ;
      RECT  282600.0 1152000.0 292800.0 1165800.0 ;
      RECT  282600.0 1179600.0 292800.0 1165800.0 ;
      RECT  282600.0 1179600.0 292800.0 1193400.0 ;
      RECT  282600.0 1207200.0 292800.0 1193400.0 ;
      RECT  282600.0 1207200.0 292800.0 1221000.0 ;
      RECT  282600.0 1234800.0 292800.0 1221000.0 ;
      RECT  282600.0 1234800.0 292800.0 1248600.0 ;
      RECT  282600.0 1262400.0 292800.0 1248600.0 ;
      RECT  282600.0 1262400.0 292800.0 1276200.0 ;
      RECT  282600.0 1290000.0 292800.0 1276200.0 ;
      RECT  282600.0 1290000.0 292800.0 1303800.0 ;
      RECT  282600.0 1317600.0 292800.0 1303800.0 ;
      RECT  282600.0 1317600.0 292800.0 1331400.0 ;
      RECT  282600.0 1345200.0 292800.0 1331400.0 ;
      RECT  282600.0 1345200.0 292800.0 1359000.0 ;
      RECT  282600.0 1372800.0 292800.0 1359000.0 ;
      RECT  282600.0 1372800.0 292800.0 1386600.0 ;
      RECT  282600.0 1400400.0 292800.0 1386600.0 ;
      RECT  282600.0 1400400.0 292800.0 1414200.0 ;
      RECT  282600.0 1428000.0 292800.0 1414200.0 ;
      RECT  282600.0 1428000.0 292800.0 1441800.0 ;
      RECT  282600.0 1455600.0 292800.0 1441800.0 ;
      RECT  282600.0 1455600.0 292800.0 1469400.0 ;
      RECT  282600.0 1483200.0 292800.0 1469400.0 ;
      RECT  282600.0 1483200.0 292800.0 1497000.0 ;
      RECT  282600.0 1510800.0 292800.0 1497000.0 ;
      RECT  282600.0 1510800.0 292800.0 1524600.0 ;
      RECT  282600.0 1538400.0 292800.0 1524600.0 ;
      RECT  282600.0 1538400.0 292800.0 1552200.0 ;
      RECT  282600.0 1566000.0 292800.0 1552200.0 ;
      RECT  282600.0 1566000.0 292800.0 1579800.0 ;
      RECT  282600.0 1593600.0 292800.0 1579800.0 ;
      RECT  282600.0 1593600.0 292800.0 1607400.0 ;
      RECT  282600.0 1621200.0 292800.0 1607400.0 ;
      RECT  282600.0 1621200.0 292800.0 1635000.0 ;
      RECT  282600.0 1648800.0 292800.0 1635000.0 ;
      RECT  282600.0 1648800.0 292800.0 1662600.0 ;
      RECT  282600.0 1676400.0 292800.0 1662600.0 ;
      RECT  282600.0 1676400.0 292800.0 1690200.0 ;
      RECT  282600.0 1704000.0 292800.0 1690200.0 ;
      RECT  282600.0 1704000.0 292800.0 1717800.0 ;
      RECT  282600.0 1731600.0 292800.0 1717800.0 ;
      RECT  282600.0 1731600.0 292800.0 1745400.0 ;
      RECT  282600.0 1759200.0 292800.0 1745400.0 ;
      RECT  282600.0 1759200.0 292800.0 1773000.0 ;
      RECT  282600.0 1786800.0 292800.0 1773000.0 ;
      RECT  282600.0 1786800.0 292800.0 1800600.0 ;
      RECT  282600.0 1814400.0 292800.0 1800600.0 ;
      RECT  282600.0 1814400.0 292800.0 1828200.0 ;
      RECT  282600.0 1842000.0 292800.0 1828200.0 ;
      RECT  282600.0 1842000.0 292800.0 1855800.0 ;
      RECT  282600.0 1869600.0 292800.0 1855800.0 ;
      RECT  282600.0 1869600.0 292800.0 1883400.0 ;
      RECT  282600.0 1897200.0 292800.0 1883400.0 ;
      RECT  282600.0 1897200.0 292800.0 1911000.0 ;
      RECT  282600.0 1924800.0 292800.0 1911000.0 ;
      RECT  282600.0 1924800.0 292800.0 1938600.0 ;
      RECT  282600.0 1952400.0 292800.0 1938600.0 ;
      RECT  282600.0 1952400.0 292800.0 1966200.0 ;
      RECT  282600.0 1980000.0 292800.0 1966200.0 ;
      RECT  282600.0 1980000.0 292800.0 1993800.0 ;
      RECT  282600.0 2007600.0 292800.0 1993800.0 ;
      RECT  282600.0 2007600.0 292800.0 2021400.0 ;
      RECT  282600.0 2035200.0 292800.0 2021400.0 ;
      RECT  282600.0 2035200.0 292800.0 2049000.0 ;
      RECT  282600.0 2062800.0 292800.0 2049000.0 ;
      RECT  282600.0 2062800.0 292800.0 2076600.0 ;
      RECT  282600.0 2090400.0 292800.0 2076600.0 ;
      RECT  282600.0 2090400.0 292800.0 2104200.0 ;
      RECT  282600.0 2118000.0 292800.0 2104200.0 ;
      RECT  282600.0 2118000.0 292800.0 2131800.0 ;
      RECT  282600.0 2145600.0 292800.0 2131800.0 ;
      RECT  292800.0 379200.0 303000.0 393000.0 ;
      RECT  292800.0 406800.0 303000.0 393000.0 ;
      RECT  292800.0 406800.0 303000.0 420600.0 ;
      RECT  292800.0 434400.0 303000.0 420600.0 ;
      RECT  292800.0 434400.0 303000.0 448200.0 ;
      RECT  292800.0 462000.0 303000.0 448200.0 ;
      RECT  292800.0 462000.0 303000.0 475800.0 ;
      RECT  292800.0 489600.0 303000.0 475800.0 ;
      RECT  292800.0 489600.0 303000.0 503400.0 ;
      RECT  292800.0 517200.0 303000.0 503400.0 ;
      RECT  292800.0 517200.0 303000.0 531000.0 ;
      RECT  292800.0 544800.0 303000.0 531000.0 ;
      RECT  292800.0 544800.0 303000.0 558600.0 ;
      RECT  292800.0 572400.0 303000.0 558600.0 ;
      RECT  292800.0 572400.0 303000.0 586200.0 ;
      RECT  292800.0 600000.0 303000.0 586200.0 ;
      RECT  292800.0 600000.0 303000.0 613800.0 ;
      RECT  292800.0 627600.0 303000.0 613800.0 ;
      RECT  292800.0 627600.0 303000.0 641400.0 ;
      RECT  292800.0 655200.0 303000.0 641400.0 ;
      RECT  292800.0 655200.0 303000.0 669000.0 ;
      RECT  292800.0 682800.0 303000.0 669000.0 ;
      RECT  292800.0 682800.0 303000.0 696600.0 ;
      RECT  292800.0 710400.0 303000.0 696600.0 ;
      RECT  292800.0 710400.0 303000.0 724200.0 ;
      RECT  292800.0 738000.0 303000.0 724200.0 ;
      RECT  292800.0 738000.0 303000.0 751800.0 ;
      RECT  292800.0 765600.0 303000.0 751800.0 ;
      RECT  292800.0 765600.0 303000.0 779400.0 ;
      RECT  292800.0 793200.0 303000.0 779400.0 ;
      RECT  292800.0 793200.0 303000.0 807000.0 ;
      RECT  292800.0 820800.0 303000.0 807000.0 ;
      RECT  292800.0 820800.0 303000.0 834600.0 ;
      RECT  292800.0 848400.0 303000.0 834600.0 ;
      RECT  292800.0 848400.0 303000.0 862200.0 ;
      RECT  292800.0 876000.0 303000.0 862200.0 ;
      RECT  292800.0 876000.0 303000.0 889800.0 ;
      RECT  292800.0 903600.0 303000.0 889800.0 ;
      RECT  292800.0 903600.0 303000.0 917400.0 ;
      RECT  292800.0 931200.0 303000.0 917400.0 ;
      RECT  292800.0 931200.0 303000.0 945000.0 ;
      RECT  292800.0 958800.0 303000.0 945000.0 ;
      RECT  292800.0 958800.0 303000.0 972600.0 ;
      RECT  292800.0 986400.0 303000.0 972600.0 ;
      RECT  292800.0 986400.0 303000.0 1000200.0 ;
      RECT  292800.0 1014000.0 303000.0 1000200.0 ;
      RECT  292800.0 1014000.0 303000.0 1027800.0 ;
      RECT  292800.0 1041600.0 303000.0 1027800.0 ;
      RECT  292800.0 1041600.0 303000.0 1055400.0 ;
      RECT  292800.0 1069200.0 303000.0 1055400.0 ;
      RECT  292800.0 1069200.0 303000.0 1083000.0 ;
      RECT  292800.0 1096800.0 303000.0 1083000.0 ;
      RECT  292800.0 1096800.0 303000.0 1110600.0 ;
      RECT  292800.0 1124400.0 303000.0 1110600.0 ;
      RECT  292800.0 1124400.0 303000.0 1138200.0 ;
      RECT  292800.0 1152000.0 303000.0 1138200.0 ;
      RECT  292800.0 1152000.0 303000.0 1165800.0 ;
      RECT  292800.0 1179600.0 303000.0 1165800.0 ;
      RECT  292800.0 1179600.0 303000.0 1193400.0 ;
      RECT  292800.0 1207200.0 303000.0 1193400.0 ;
      RECT  292800.0 1207200.0 303000.0 1221000.0 ;
      RECT  292800.0 1234800.0 303000.0 1221000.0 ;
      RECT  292800.0 1234800.0 303000.0 1248600.0 ;
      RECT  292800.0 1262400.0 303000.0 1248600.0 ;
      RECT  292800.0 1262400.0 303000.0 1276200.0 ;
      RECT  292800.0 1290000.0 303000.0 1276200.0 ;
      RECT  292800.0 1290000.0 303000.0 1303800.0 ;
      RECT  292800.0 1317600.0 303000.0 1303800.0 ;
      RECT  292800.0 1317600.0 303000.0 1331400.0 ;
      RECT  292800.0 1345200.0 303000.0 1331400.0 ;
      RECT  292800.0 1345200.0 303000.0 1359000.0 ;
      RECT  292800.0 1372800.0 303000.0 1359000.0 ;
      RECT  292800.0 1372800.0 303000.0 1386600.0 ;
      RECT  292800.0 1400400.0 303000.0 1386600.0 ;
      RECT  292800.0 1400400.0 303000.0 1414200.0 ;
      RECT  292800.0 1428000.0 303000.0 1414200.0 ;
      RECT  292800.0 1428000.0 303000.0 1441800.0 ;
      RECT  292800.0 1455600.0 303000.0 1441800.0 ;
      RECT  292800.0 1455600.0 303000.0 1469400.0 ;
      RECT  292800.0 1483200.0 303000.0 1469400.0 ;
      RECT  292800.0 1483200.0 303000.0 1497000.0 ;
      RECT  292800.0 1510800.0 303000.0 1497000.0 ;
      RECT  292800.0 1510800.0 303000.0 1524600.0 ;
      RECT  292800.0 1538400.0 303000.0 1524600.0 ;
      RECT  292800.0 1538400.0 303000.0 1552200.0 ;
      RECT  292800.0 1566000.0 303000.0 1552200.0 ;
      RECT  292800.0 1566000.0 303000.0 1579800.0 ;
      RECT  292800.0 1593600.0 303000.0 1579800.0 ;
      RECT  292800.0 1593600.0 303000.0 1607400.0 ;
      RECT  292800.0 1621200.0 303000.0 1607400.0 ;
      RECT  292800.0 1621200.0 303000.0 1635000.0 ;
      RECT  292800.0 1648800.0 303000.0 1635000.0 ;
      RECT  292800.0 1648800.0 303000.0 1662600.0 ;
      RECT  292800.0 1676400.0 303000.0 1662600.0 ;
      RECT  292800.0 1676400.0 303000.0 1690200.0 ;
      RECT  292800.0 1704000.0 303000.0 1690200.0 ;
      RECT  292800.0 1704000.0 303000.0 1717800.0 ;
      RECT  292800.0 1731600.0 303000.0 1717800.0 ;
      RECT  292800.0 1731600.0 303000.0 1745400.0 ;
      RECT  292800.0 1759200.0 303000.0 1745400.0 ;
      RECT  292800.0 1759200.0 303000.0 1773000.0 ;
      RECT  292800.0 1786800.0 303000.0 1773000.0 ;
      RECT  292800.0 1786800.0 303000.0 1800600.0 ;
      RECT  292800.0 1814400.0 303000.0 1800600.0 ;
      RECT  292800.0 1814400.0 303000.0 1828200.0 ;
      RECT  292800.0 1842000.0 303000.0 1828200.0 ;
      RECT  292800.0 1842000.0 303000.0 1855800.0 ;
      RECT  292800.0 1869600.0 303000.0 1855800.0 ;
      RECT  292800.0 1869600.0 303000.0 1883400.0 ;
      RECT  292800.0 1897200.0 303000.0 1883400.0 ;
      RECT  292800.0 1897200.0 303000.0 1911000.0 ;
      RECT  292800.0 1924800.0 303000.0 1911000.0 ;
      RECT  292800.0 1924800.0 303000.0 1938600.0 ;
      RECT  292800.0 1952400.0 303000.0 1938600.0 ;
      RECT  292800.0 1952400.0 303000.0 1966200.0 ;
      RECT  292800.0 1980000.0 303000.0 1966200.0 ;
      RECT  292800.0 1980000.0 303000.0 1993800.0 ;
      RECT  292800.0 2007600.0 303000.0 1993800.0 ;
      RECT  292800.0 2007600.0 303000.0 2021400.0 ;
      RECT  292800.0 2035200.0 303000.0 2021400.0 ;
      RECT  292800.0 2035200.0 303000.0 2049000.0 ;
      RECT  292800.0 2062800.0 303000.0 2049000.0 ;
      RECT  292800.0 2062800.0 303000.0 2076600.0 ;
      RECT  292800.0 2090400.0 303000.0 2076600.0 ;
      RECT  292800.0 2090400.0 303000.0 2104200.0 ;
      RECT  292800.0 2118000.0 303000.0 2104200.0 ;
      RECT  292800.0 2118000.0 303000.0 2131800.0 ;
      RECT  292800.0 2145600.0 303000.0 2131800.0 ;
      RECT  303000.0 379200.0 313200.0 393000.0 ;
      RECT  303000.0 406800.0 313200.0 393000.0 ;
      RECT  303000.0 406800.0 313200.0 420600.0 ;
      RECT  303000.0 434400.0 313200.0 420600.0 ;
      RECT  303000.0 434400.0 313200.0 448200.0 ;
      RECT  303000.0 462000.0 313200.0 448200.0 ;
      RECT  303000.0 462000.0 313200.0 475800.0 ;
      RECT  303000.0 489600.0 313200.0 475800.0 ;
      RECT  303000.0 489600.0 313200.0 503400.0 ;
      RECT  303000.0 517200.0 313200.0 503400.0 ;
      RECT  303000.0 517200.0 313200.0 531000.0 ;
      RECT  303000.0 544800.0 313200.0 531000.0 ;
      RECT  303000.0 544800.0 313200.0 558600.0 ;
      RECT  303000.0 572400.0 313200.0 558600.0 ;
      RECT  303000.0 572400.0 313200.0 586200.0 ;
      RECT  303000.0 600000.0 313200.0 586200.0 ;
      RECT  303000.0 600000.0 313200.0 613800.0 ;
      RECT  303000.0 627600.0 313200.0 613800.0 ;
      RECT  303000.0 627600.0 313200.0 641400.0 ;
      RECT  303000.0 655200.0 313200.0 641400.0 ;
      RECT  303000.0 655200.0 313200.0 669000.0 ;
      RECT  303000.0 682800.0 313200.0 669000.0 ;
      RECT  303000.0 682800.0 313200.0 696600.0 ;
      RECT  303000.0 710400.0 313200.0 696600.0 ;
      RECT  303000.0 710400.0 313200.0 724200.0 ;
      RECT  303000.0 738000.0 313200.0 724200.0 ;
      RECT  303000.0 738000.0 313200.0 751800.0 ;
      RECT  303000.0 765600.0 313200.0 751800.0 ;
      RECT  303000.0 765600.0 313200.0 779400.0 ;
      RECT  303000.0 793200.0 313200.0 779400.0 ;
      RECT  303000.0 793200.0 313200.0 807000.0 ;
      RECT  303000.0 820800.0 313200.0 807000.0 ;
      RECT  303000.0 820800.0 313200.0 834600.0 ;
      RECT  303000.0 848400.0 313200.0 834600.0 ;
      RECT  303000.0 848400.0 313200.0 862200.0 ;
      RECT  303000.0 876000.0 313200.0 862200.0 ;
      RECT  303000.0 876000.0 313200.0 889800.0 ;
      RECT  303000.0 903600.0 313200.0 889800.0 ;
      RECT  303000.0 903600.0 313200.0 917400.0 ;
      RECT  303000.0 931200.0 313200.0 917400.0 ;
      RECT  303000.0 931200.0 313200.0 945000.0 ;
      RECT  303000.0 958800.0 313200.0 945000.0 ;
      RECT  303000.0 958800.0 313200.0 972600.0 ;
      RECT  303000.0 986400.0 313200.0 972600.0 ;
      RECT  303000.0 986400.0 313200.0 1000200.0 ;
      RECT  303000.0 1014000.0 313200.0 1000200.0 ;
      RECT  303000.0 1014000.0 313200.0 1027800.0 ;
      RECT  303000.0 1041600.0 313200.0 1027800.0 ;
      RECT  303000.0 1041600.0 313200.0 1055400.0 ;
      RECT  303000.0 1069200.0 313200.0 1055400.0 ;
      RECT  303000.0 1069200.0 313200.0 1083000.0 ;
      RECT  303000.0 1096800.0 313200.0 1083000.0 ;
      RECT  303000.0 1096800.0 313200.0 1110600.0 ;
      RECT  303000.0 1124400.0 313200.0 1110600.0 ;
      RECT  303000.0 1124400.0 313200.0 1138200.0 ;
      RECT  303000.0 1152000.0 313200.0 1138200.0 ;
      RECT  303000.0 1152000.0 313200.0 1165800.0 ;
      RECT  303000.0 1179600.0 313200.0 1165800.0 ;
      RECT  303000.0 1179600.0 313200.0 1193400.0 ;
      RECT  303000.0 1207200.0 313200.0 1193400.0 ;
      RECT  303000.0 1207200.0 313200.0 1221000.0 ;
      RECT  303000.0 1234800.0 313200.0 1221000.0 ;
      RECT  303000.0 1234800.0 313200.0 1248600.0 ;
      RECT  303000.0 1262400.0 313200.0 1248600.0 ;
      RECT  303000.0 1262400.0 313200.0 1276200.0 ;
      RECT  303000.0 1290000.0 313200.0 1276200.0 ;
      RECT  303000.0 1290000.0 313200.0 1303800.0 ;
      RECT  303000.0 1317600.0 313200.0 1303800.0 ;
      RECT  303000.0 1317600.0 313200.0 1331400.0 ;
      RECT  303000.0 1345200.0 313200.0 1331400.0 ;
      RECT  303000.0 1345200.0 313200.0 1359000.0 ;
      RECT  303000.0 1372800.0 313200.0 1359000.0 ;
      RECT  303000.0 1372800.0 313200.0 1386600.0 ;
      RECT  303000.0 1400400.0 313200.0 1386600.0 ;
      RECT  303000.0 1400400.0 313200.0 1414200.0 ;
      RECT  303000.0 1428000.0 313200.0 1414200.0 ;
      RECT  303000.0 1428000.0 313200.0 1441800.0 ;
      RECT  303000.0 1455600.0 313200.0 1441800.0 ;
      RECT  303000.0 1455600.0 313200.0 1469400.0 ;
      RECT  303000.0 1483200.0 313200.0 1469400.0 ;
      RECT  303000.0 1483200.0 313200.0 1497000.0 ;
      RECT  303000.0 1510800.0 313200.0 1497000.0 ;
      RECT  303000.0 1510800.0 313200.0 1524600.0 ;
      RECT  303000.0 1538400.0 313200.0 1524600.0 ;
      RECT  303000.0 1538400.0 313200.0 1552200.0 ;
      RECT  303000.0 1566000.0 313200.0 1552200.0 ;
      RECT  303000.0 1566000.0 313200.0 1579800.0 ;
      RECT  303000.0 1593600.0 313200.0 1579800.0 ;
      RECT  303000.0 1593600.0 313200.0 1607400.0 ;
      RECT  303000.0 1621200.0 313200.0 1607400.0 ;
      RECT  303000.0 1621200.0 313200.0 1635000.0 ;
      RECT  303000.0 1648800.0 313200.0 1635000.0 ;
      RECT  303000.0 1648800.0 313200.0 1662600.0 ;
      RECT  303000.0 1676400.0 313200.0 1662600.0 ;
      RECT  303000.0 1676400.0 313200.0 1690200.0 ;
      RECT  303000.0 1704000.0 313200.0 1690200.0 ;
      RECT  303000.0 1704000.0 313200.0 1717800.0 ;
      RECT  303000.0 1731600.0 313200.0 1717800.0 ;
      RECT  303000.0 1731600.0 313200.0 1745400.0 ;
      RECT  303000.0 1759200.0 313200.0 1745400.0 ;
      RECT  303000.0 1759200.0 313200.0 1773000.0 ;
      RECT  303000.0 1786800.0 313200.0 1773000.0 ;
      RECT  303000.0 1786800.0 313200.0 1800600.0 ;
      RECT  303000.0 1814400.0 313200.0 1800600.0 ;
      RECT  303000.0 1814400.0 313200.0 1828200.0 ;
      RECT  303000.0 1842000.0 313200.0 1828200.0 ;
      RECT  303000.0 1842000.0 313200.0 1855800.0 ;
      RECT  303000.0 1869600.0 313200.0 1855800.0 ;
      RECT  303000.0 1869600.0 313200.0 1883400.0 ;
      RECT  303000.0 1897200.0 313200.0 1883400.0 ;
      RECT  303000.0 1897200.0 313200.0 1911000.0 ;
      RECT  303000.0 1924800.0 313200.0 1911000.0 ;
      RECT  303000.0 1924800.0 313200.0 1938600.0 ;
      RECT  303000.0 1952400.0 313200.0 1938600.0 ;
      RECT  303000.0 1952400.0 313200.0 1966200.0 ;
      RECT  303000.0 1980000.0 313200.0 1966200.0 ;
      RECT  303000.0 1980000.0 313200.0 1993800.0 ;
      RECT  303000.0 2007600.0 313200.0 1993800.0 ;
      RECT  303000.0 2007600.0 313200.0 2021400.0 ;
      RECT  303000.0 2035200.0 313200.0 2021400.0 ;
      RECT  303000.0 2035200.0 313200.0 2049000.0 ;
      RECT  303000.0 2062800.0 313200.0 2049000.0 ;
      RECT  303000.0 2062800.0 313200.0 2076600.0 ;
      RECT  303000.0 2090400.0 313200.0 2076600.0 ;
      RECT  303000.0 2090400.0 313200.0 2104200.0 ;
      RECT  303000.0 2118000.0 313200.0 2104200.0 ;
      RECT  303000.0 2118000.0 313200.0 2131800.0 ;
      RECT  303000.0 2145600.0 313200.0 2131800.0 ;
      RECT  313200.0 379200.0 323400.0 393000.0 ;
      RECT  313200.0 406800.0 323400.0 393000.0 ;
      RECT  313200.0 406800.0 323400.0 420600.0 ;
      RECT  313200.0 434400.0 323400.0 420600.0 ;
      RECT  313200.0 434400.0 323400.0 448200.0 ;
      RECT  313200.0 462000.0 323400.0 448200.0 ;
      RECT  313200.0 462000.0 323400.0 475800.0 ;
      RECT  313200.0 489600.0 323400.0 475800.0 ;
      RECT  313200.0 489600.0 323400.0 503400.0 ;
      RECT  313200.0 517200.0 323400.0 503400.0 ;
      RECT  313200.0 517200.0 323400.0 531000.0 ;
      RECT  313200.0 544800.0 323400.0 531000.0 ;
      RECT  313200.0 544800.0 323400.0 558600.0 ;
      RECT  313200.0 572400.0 323400.0 558600.0 ;
      RECT  313200.0 572400.0 323400.0 586200.0 ;
      RECT  313200.0 600000.0 323400.0 586200.0 ;
      RECT  313200.0 600000.0 323400.0 613800.0 ;
      RECT  313200.0 627600.0 323400.0 613800.0 ;
      RECT  313200.0 627600.0 323400.0 641400.0 ;
      RECT  313200.0 655200.0 323400.0 641400.0 ;
      RECT  313200.0 655200.0 323400.0 669000.0 ;
      RECT  313200.0 682800.0 323400.0 669000.0 ;
      RECT  313200.0 682800.0 323400.0 696600.0 ;
      RECT  313200.0 710400.0 323400.0 696600.0 ;
      RECT  313200.0 710400.0 323400.0 724200.0 ;
      RECT  313200.0 738000.0 323400.0 724200.0 ;
      RECT  313200.0 738000.0 323400.0 751800.0 ;
      RECT  313200.0 765600.0 323400.0 751800.0 ;
      RECT  313200.0 765600.0 323400.0 779400.0 ;
      RECT  313200.0 793200.0 323400.0 779400.0 ;
      RECT  313200.0 793200.0 323400.0 807000.0 ;
      RECT  313200.0 820800.0 323400.0 807000.0 ;
      RECT  313200.0 820800.0 323400.0 834600.0 ;
      RECT  313200.0 848400.0 323400.0 834600.0 ;
      RECT  313200.0 848400.0 323400.0 862200.0 ;
      RECT  313200.0 876000.0 323400.0 862200.0 ;
      RECT  313200.0 876000.0 323400.0 889800.0 ;
      RECT  313200.0 903600.0 323400.0 889800.0 ;
      RECT  313200.0 903600.0 323400.0 917400.0 ;
      RECT  313200.0 931200.0 323400.0 917400.0 ;
      RECT  313200.0 931200.0 323400.0 945000.0 ;
      RECT  313200.0 958800.0 323400.0 945000.0 ;
      RECT  313200.0 958800.0 323400.0 972600.0 ;
      RECT  313200.0 986400.0 323400.0 972600.0 ;
      RECT  313200.0 986400.0 323400.0 1000200.0 ;
      RECT  313200.0 1014000.0 323400.0 1000200.0 ;
      RECT  313200.0 1014000.0 323400.0 1027800.0 ;
      RECT  313200.0 1041600.0 323400.0 1027800.0 ;
      RECT  313200.0 1041600.0 323400.0 1055400.0 ;
      RECT  313200.0 1069200.0 323400.0 1055400.0 ;
      RECT  313200.0 1069200.0 323400.0 1083000.0 ;
      RECT  313200.0 1096800.0 323400.0 1083000.0 ;
      RECT  313200.0 1096800.0 323400.0 1110600.0 ;
      RECT  313200.0 1124400.0 323400.0 1110600.0 ;
      RECT  313200.0 1124400.0 323400.0 1138200.0 ;
      RECT  313200.0 1152000.0 323400.0 1138200.0 ;
      RECT  313200.0 1152000.0 323400.0 1165800.0 ;
      RECT  313200.0 1179600.0 323400.0 1165800.0 ;
      RECT  313200.0 1179600.0 323400.0 1193400.0 ;
      RECT  313200.0 1207200.0 323400.0 1193400.0 ;
      RECT  313200.0 1207200.0 323400.0 1221000.0 ;
      RECT  313200.0 1234800.0 323400.0 1221000.0 ;
      RECT  313200.0 1234800.0 323400.0 1248600.0 ;
      RECT  313200.0 1262400.0 323400.0 1248600.0 ;
      RECT  313200.0 1262400.0 323400.0 1276200.0 ;
      RECT  313200.0 1290000.0 323400.0 1276200.0 ;
      RECT  313200.0 1290000.0 323400.0 1303800.0 ;
      RECT  313200.0 1317600.0 323400.0 1303800.0 ;
      RECT  313200.0 1317600.0 323400.0 1331400.0 ;
      RECT  313200.0 1345200.0 323400.0 1331400.0 ;
      RECT  313200.0 1345200.0 323400.0 1359000.0 ;
      RECT  313200.0 1372800.0 323400.0 1359000.0 ;
      RECT  313200.0 1372800.0 323400.0 1386600.0 ;
      RECT  313200.0 1400400.0 323400.0 1386600.0 ;
      RECT  313200.0 1400400.0 323400.0 1414200.0 ;
      RECT  313200.0 1428000.0 323400.0 1414200.0 ;
      RECT  313200.0 1428000.0 323400.0 1441800.0 ;
      RECT  313200.0 1455600.0 323400.0 1441800.0 ;
      RECT  313200.0 1455600.0 323400.0 1469400.0 ;
      RECT  313200.0 1483200.0 323400.0 1469400.0 ;
      RECT  313200.0 1483200.0 323400.0 1497000.0 ;
      RECT  313200.0 1510800.0 323400.0 1497000.0 ;
      RECT  313200.0 1510800.0 323400.0 1524600.0 ;
      RECT  313200.0 1538400.0 323400.0 1524600.0 ;
      RECT  313200.0 1538400.0 323400.0 1552200.0 ;
      RECT  313200.0 1566000.0 323400.0 1552200.0 ;
      RECT  313200.0 1566000.0 323400.0 1579800.0 ;
      RECT  313200.0 1593600.0 323400.0 1579800.0 ;
      RECT  313200.0 1593600.0 323400.0 1607400.0 ;
      RECT  313200.0 1621200.0 323400.0 1607400.0 ;
      RECT  313200.0 1621200.0 323400.0 1635000.0 ;
      RECT  313200.0 1648800.0 323400.0 1635000.0 ;
      RECT  313200.0 1648800.0 323400.0 1662600.0 ;
      RECT  313200.0 1676400.0 323400.0 1662600.0 ;
      RECT  313200.0 1676400.0 323400.0 1690200.0 ;
      RECT  313200.0 1704000.0 323400.0 1690200.0 ;
      RECT  313200.0 1704000.0 323400.0 1717800.0 ;
      RECT  313200.0 1731600.0 323400.0 1717800.0 ;
      RECT  313200.0 1731600.0 323400.0 1745400.0 ;
      RECT  313200.0 1759200.0 323400.0 1745400.0 ;
      RECT  313200.0 1759200.0 323400.0 1773000.0 ;
      RECT  313200.0 1786800.0 323400.0 1773000.0 ;
      RECT  313200.0 1786800.0 323400.0 1800600.0 ;
      RECT  313200.0 1814400.0 323400.0 1800600.0 ;
      RECT  313200.0 1814400.0 323400.0 1828200.0 ;
      RECT  313200.0 1842000.0 323400.0 1828200.0 ;
      RECT  313200.0 1842000.0 323400.0 1855800.0 ;
      RECT  313200.0 1869600.0 323400.0 1855800.0 ;
      RECT  313200.0 1869600.0 323400.0 1883400.0 ;
      RECT  313200.0 1897200.0 323400.0 1883400.0 ;
      RECT  313200.0 1897200.0 323400.0 1911000.0 ;
      RECT  313200.0 1924800.0 323400.0 1911000.0 ;
      RECT  313200.0 1924800.0 323400.0 1938600.0 ;
      RECT  313200.0 1952400.0 323400.0 1938600.0 ;
      RECT  313200.0 1952400.0 323400.0 1966200.0 ;
      RECT  313200.0 1980000.0 323400.0 1966200.0 ;
      RECT  313200.0 1980000.0 323400.0 1993800.0 ;
      RECT  313200.0 2007600.0 323400.0 1993800.0 ;
      RECT  313200.0 2007600.0 323400.0 2021400.0 ;
      RECT  313200.0 2035200.0 323400.0 2021400.0 ;
      RECT  313200.0 2035200.0 323400.0 2049000.0 ;
      RECT  313200.0 2062800.0 323400.0 2049000.0 ;
      RECT  313200.0 2062800.0 323400.0 2076600.0 ;
      RECT  313200.0 2090400.0 323400.0 2076600.0 ;
      RECT  313200.0 2090400.0 323400.0 2104200.0 ;
      RECT  313200.0 2118000.0 323400.0 2104200.0 ;
      RECT  313200.0 2118000.0 323400.0 2131800.0 ;
      RECT  313200.0 2145600.0 323400.0 2131800.0 ;
      RECT  323400.0 379200.0 333600.0 393000.0 ;
      RECT  323400.0 406800.0 333600.0 393000.0 ;
      RECT  323400.0 406800.0 333600.0 420600.0 ;
      RECT  323400.0 434400.0 333600.0 420600.0 ;
      RECT  323400.0 434400.0 333600.0 448200.0 ;
      RECT  323400.0 462000.0 333600.0 448200.0 ;
      RECT  323400.0 462000.0 333600.0 475800.0 ;
      RECT  323400.0 489600.0 333600.0 475800.0 ;
      RECT  323400.0 489600.0 333600.0 503400.0 ;
      RECT  323400.0 517200.0 333600.0 503400.0 ;
      RECT  323400.0 517200.0 333600.0 531000.0 ;
      RECT  323400.0 544800.0 333600.0 531000.0 ;
      RECT  323400.0 544800.0 333600.0 558600.0 ;
      RECT  323400.0 572400.0 333600.0 558600.0 ;
      RECT  323400.0 572400.0 333600.0 586200.0 ;
      RECT  323400.0 600000.0 333600.0 586200.0 ;
      RECT  323400.0 600000.0 333600.0 613800.0 ;
      RECT  323400.0 627600.0 333600.0 613800.0 ;
      RECT  323400.0 627600.0 333600.0 641400.0 ;
      RECT  323400.0 655200.0 333600.0 641400.0 ;
      RECT  323400.0 655200.0 333600.0 669000.0 ;
      RECT  323400.0 682800.0 333600.0 669000.0 ;
      RECT  323400.0 682800.0 333600.0 696600.0 ;
      RECT  323400.0 710400.0 333600.0 696600.0 ;
      RECT  323400.0 710400.0 333600.0 724200.0 ;
      RECT  323400.0 738000.0 333600.0 724200.0 ;
      RECT  323400.0 738000.0 333600.0 751800.0 ;
      RECT  323400.0 765600.0 333600.0 751800.0 ;
      RECT  323400.0 765600.0 333600.0 779400.0 ;
      RECT  323400.0 793200.0 333600.0 779400.0 ;
      RECT  323400.0 793200.0 333600.0 807000.0 ;
      RECT  323400.0 820800.0 333600.0 807000.0 ;
      RECT  323400.0 820800.0 333600.0 834600.0 ;
      RECT  323400.0 848400.0 333600.0 834600.0 ;
      RECT  323400.0 848400.0 333600.0 862200.0 ;
      RECT  323400.0 876000.0 333600.0 862200.0 ;
      RECT  323400.0 876000.0 333600.0 889800.0 ;
      RECT  323400.0 903600.0 333600.0 889800.0 ;
      RECT  323400.0 903600.0 333600.0 917400.0 ;
      RECT  323400.0 931200.0 333600.0 917400.0 ;
      RECT  323400.0 931200.0 333600.0 945000.0 ;
      RECT  323400.0 958800.0 333600.0 945000.0 ;
      RECT  323400.0 958800.0 333600.0 972600.0 ;
      RECT  323400.0 986400.0 333600.0 972600.0 ;
      RECT  323400.0 986400.0 333600.0 1000200.0 ;
      RECT  323400.0 1014000.0 333600.0 1000200.0 ;
      RECT  323400.0 1014000.0 333600.0 1027800.0 ;
      RECT  323400.0 1041600.0 333600.0 1027800.0 ;
      RECT  323400.0 1041600.0 333600.0 1055400.0 ;
      RECT  323400.0 1069200.0 333600.0 1055400.0 ;
      RECT  323400.0 1069200.0 333600.0 1083000.0 ;
      RECT  323400.0 1096800.0 333600.0 1083000.0 ;
      RECT  323400.0 1096800.0 333600.0 1110600.0 ;
      RECT  323400.0 1124400.0 333600.0 1110600.0 ;
      RECT  323400.0 1124400.0 333600.0 1138200.0 ;
      RECT  323400.0 1152000.0 333600.0 1138200.0 ;
      RECT  323400.0 1152000.0 333600.0 1165800.0 ;
      RECT  323400.0 1179600.0 333600.0 1165800.0 ;
      RECT  323400.0 1179600.0 333600.0 1193400.0 ;
      RECT  323400.0 1207200.0 333600.0 1193400.0 ;
      RECT  323400.0 1207200.0 333600.0 1221000.0 ;
      RECT  323400.0 1234800.0 333600.0 1221000.0 ;
      RECT  323400.0 1234800.0 333600.0 1248600.0 ;
      RECT  323400.0 1262400.0 333600.0 1248600.0 ;
      RECT  323400.0 1262400.0 333600.0 1276200.0 ;
      RECT  323400.0 1290000.0 333600.0 1276200.0 ;
      RECT  323400.0 1290000.0 333600.0 1303800.0 ;
      RECT  323400.0 1317600.0 333600.0 1303800.0 ;
      RECT  323400.0 1317600.0 333600.0 1331400.0 ;
      RECT  323400.0 1345200.0 333600.0 1331400.0 ;
      RECT  323400.0 1345200.0 333600.0 1359000.0 ;
      RECT  323400.0 1372800.0 333600.0 1359000.0 ;
      RECT  323400.0 1372800.0 333600.0 1386600.0 ;
      RECT  323400.0 1400400.0 333600.0 1386600.0 ;
      RECT  323400.0 1400400.0 333600.0 1414200.0 ;
      RECT  323400.0 1428000.0 333600.0 1414200.0 ;
      RECT  323400.0 1428000.0 333600.0 1441800.0 ;
      RECT  323400.0 1455600.0 333600.0 1441800.0 ;
      RECT  323400.0 1455600.0 333600.0 1469400.0 ;
      RECT  323400.0 1483200.0 333600.0 1469400.0 ;
      RECT  323400.0 1483200.0 333600.0 1497000.0 ;
      RECT  323400.0 1510800.0 333600.0 1497000.0 ;
      RECT  323400.0 1510800.0 333600.0 1524600.0 ;
      RECT  323400.0 1538400.0 333600.0 1524600.0 ;
      RECT  323400.0 1538400.0 333600.0 1552200.0 ;
      RECT  323400.0 1566000.0 333600.0 1552200.0 ;
      RECT  323400.0 1566000.0 333600.0 1579800.0 ;
      RECT  323400.0 1593600.0 333600.0 1579800.0 ;
      RECT  323400.0 1593600.0 333600.0 1607400.0 ;
      RECT  323400.0 1621200.0 333600.0 1607400.0 ;
      RECT  323400.0 1621200.0 333600.0 1635000.0 ;
      RECT  323400.0 1648800.0 333600.0 1635000.0 ;
      RECT  323400.0 1648800.0 333600.0 1662600.0 ;
      RECT  323400.0 1676400.0 333600.0 1662600.0 ;
      RECT  323400.0 1676400.0 333600.0 1690200.0 ;
      RECT  323400.0 1704000.0 333600.0 1690200.0 ;
      RECT  323400.0 1704000.0 333600.0 1717800.0 ;
      RECT  323400.0 1731600.0 333600.0 1717800.0 ;
      RECT  323400.0 1731600.0 333600.0 1745400.0 ;
      RECT  323400.0 1759200.0 333600.0 1745400.0 ;
      RECT  323400.0 1759200.0 333600.0 1773000.0 ;
      RECT  323400.0 1786800.0 333600.0 1773000.0 ;
      RECT  323400.0 1786800.0 333600.0 1800600.0 ;
      RECT  323400.0 1814400.0 333600.0 1800600.0 ;
      RECT  323400.0 1814400.0 333600.0 1828200.0 ;
      RECT  323400.0 1842000.0 333600.0 1828200.0 ;
      RECT  323400.0 1842000.0 333600.0 1855800.0 ;
      RECT  323400.0 1869600.0 333600.0 1855800.0 ;
      RECT  323400.0 1869600.0 333600.0 1883400.0 ;
      RECT  323400.0 1897200.0 333600.0 1883400.0 ;
      RECT  323400.0 1897200.0 333600.0 1911000.0 ;
      RECT  323400.0 1924800.0 333600.0 1911000.0 ;
      RECT  323400.0 1924800.0 333600.0 1938600.0 ;
      RECT  323400.0 1952400.0 333600.0 1938600.0 ;
      RECT  323400.0 1952400.0 333600.0 1966200.0 ;
      RECT  323400.0 1980000.0 333600.0 1966200.0 ;
      RECT  323400.0 1980000.0 333600.0 1993800.0 ;
      RECT  323400.0 2007600.0 333600.0 1993800.0 ;
      RECT  323400.0 2007600.0 333600.0 2021400.0 ;
      RECT  323400.0 2035200.0 333600.0 2021400.0 ;
      RECT  323400.0 2035200.0 333600.0 2049000.0 ;
      RECT  323400.0 2062800.0 333600.0 2049000.0 ;
      RECT  323400.0 2062800.0 333600.0 2076600.0 ;
      RECT  323400.0 2090400.0 333600.0 2076600.0 ;
      RECT  323400.0 2090400.0 333600.0 2104200.0 ;
      RECT  323400.0 2118000.0 333600.0 2104200.0 ;
      RECT  323400.0 2118000.0 333600.0 2131800.0 ;
      RECT  323400.0 2145600.0 333600.0 2131800.0 ;
      RECT  333600.0 379200.0 343800.0 393000.0 ;
      RECT  333600.0 406800.0 343800.0 393000.0 ;
      RECT  333600.0 406800.0 343800.0 420600.0 ;
      RECT  333600.0 434400.0 343800.0 420600.0 ;
      RECT  333600.0 434400.0 343800.0 448200.0 ;
      RECT  333600.0 462000.0 343800.0 448200.0 ;
      RECT  333600.0 462000.0 343800.0 475800.0 ;
      RECT  333600.0 489600.0 343800.0 475800.0 ;
      RECT  333600.0 489600.0 343800.0 503400.0 ;
      RECT  333600.0 517200.0 343800.0 503400.0 ;
      RECT  333600.0 517200.0 343800.0 531000.0 ;
      RECT  333600.0 544800.0 343800.0 531000.0 ;
      RECT  333600.0 544800.0 343800.0 558600.0 ;
      RECT  333600.0 572400.0 343800.0 558600.0 ;
      RECT  333600.0 572400.0 343800.0 586200.0 ;
      RECT  333600.0 600000.0 343800.0 586200.0 ;
      RECT  333600.0 600000.0 343800.0 613800.0 ;
      RECT  333600.0 627600.0 343800.0 613800.0 ;
      RECT  333600.0 627600.0 343800.0 641400.0 ;
      RECT  333600.0 655200.0 343800.0 641400.0 ;
      RECT  333600.0 655200.0 343800.0 669000.0 ;
      RECT  333600.0 682800.0 343800.0 669000.0 ;
      RECT  333600.0 682800.0 343800.0 696600.0 ;
      RECT  333600.0 710400.0 343800.0 696600.0 ;
      RECT  333600.0 710400.0 343800.0 724200.0 ;
      RECT  333600.0 738000.0 343800.0 724200.0 ;
      RECT  333600.0 738000.0 343800.0 751800.0 ;
      RECT  333600.0 765600.0 343800.0 751800.0 ;
      RECT  333600.0 765600.0 343800.0 779400.0 ;
      RECT  333600.0 793200.0 343800.0 779400.0 ;
      RECT  333600.0 793200.0 343800.0 807000.0 ;
      RECT  333600.0 820800.0 343800.0 807000.0 ;
      RECT  333600.0 820800.0 343800.0 834600.0 ;
      RECT  333600.0 848400.0 343800.0 834600.0 ;
      RECT  333600.0 848400.0 343800.0 862200.0 ;
      RECT  333600.0 876000.0 343800.0 862200.0 ;
      RECT  333600.0 876000.0 343800.0 889800.0 ;
      RECT  333600.0 903600.0 343800.0 889800.0 ;
      RECT  333600.0 903600.0 343800.0 917400.0 ;
      RECT  333600.0 931200.0 343800.0 917400.0 ;
      RECT  333600.0 931200.0 343800.0 945000.0 ;
      RECT  333600.0 958800.0 343800.0 945000.0 ;
      RECT  333600.0 958800.0 343800.0 972600.0 ;
      RECT  333600.0 986400.0 343800.0 972600.0 ;
      RECT  333600.0 986400.0 343800.0 1000200.0 ;
      RECT  333600.0 1014000.0 343800.0 1000200.0 ;
      RECT  333600.0 1014000.0 343800.0 1027800.0 ;
      RECT  333600.0 1041600.0 343800.0 1027800.0 ;
      RECT  333600.0 1041600.0 343800.0 1055400.0 ;
      RECT  333600.0 1069200.0 343800.0 1055400.0 ;
      RECT  333600.0 1069200.0 343800.0 1083000.0 ;
      RECT  333600.0 1096800.0 343800.0 1083000.0 ;
      RECT  333600.0 1096800.0 343800.0 1110600.0 ;
      RECT  333600.0 1124400.0 343800.0 1110600.0 ;
      RECT  333600.0 1124400.0 343800.0 1138200.0 ;
      RECT  333600.0 1152000.0 343800.0 1138200.0 ;
      RECT  333600.0 1152000.0 343800.0 1165800.0 ;
      RECT  333600.0 1179600.0 343800.0 1165800.0 ;
      RECT  333600.0 1179600.0 343800.0 1193400.0 ;
      RECT  333600.0 1207200.0 343800.0 1193400.0 ;
      RECT  333600.0 1207200.0 343800.0 1221000.0 ;
      RECT  333600.0 1234800.0 343800.0 1221000.0 ;
      RECT  333600.0 1234800.0 343800.0 1248600.0 ;
      RECT  333600.0 1262400.0 343800.0 1248600.0 ;
      RECT  333600.0 1262400.0 343800.0 1276200.0 ;
      RECT  333600.0 1290000.0 343800.0 1276200.0 ;
      RECT  333600.0 1290000.0 343800.0 1303800.0 ;
      RECT  333600.0 1317600.0 343800.0 1303800.0 ;
      RECT  333600.0 1317600.0 343800.0 1331400.0 ;
      RECT  333600.0 1345200.0 343800.0 1331400.0 ;
      RECT  333600.0 1345200.0 343800.0 1359000.0 ;
      RECT  333600.0 1372800.0 343800.0 1359000.0 ;
      RECT  333600.0 1372800.0 343800.0 1386600.0 ;
      RECT  333600.0 1400400.0 343800.0 1386600.0 ;
      RECT  333600.0 1400400.0 343800.0 1414200.0 ;
      RECT  333600.0 1428000.0 343800.0 1414200.0 ;
      RECT  333600.0 1428000.0 343800.0 1441800.0 ;
      RECT  333600.0 1455600.0 343800.0 1441800.0 ;
      RECT  333600.0 1455600.0 343800.0 1469400.0 ;
      RECT  333600.0 1483200.0 343800.0 1469400.0 ;
      RECT  333600.0 1483200.0 343800.0 1497000.0 ;
      RECT  333600.0 1510800.0 343800.0 1497000.0 ;
      RECT  333600.0 1510800.0 343800.0 1524600.0 ;
      RECT  333600.0 1538400.0 343800.0 1524600.0 ;
      RECT  333600.0 1538400.0 343800.0 1552200.0 ;
      RECT  333600.0 1566000.0 343800.0 1552200.0 ;
      RECT  333600.0 1566000.0 343800.0 1579800.0 ;
      RECT  333600.0 1593600.0 343800.0 1579800.0 ;
      RECT  333600.0 1593600.0 343800.0 1607400.0 ;
      RECT  333600.0 1621200.0 343800.0 1607400.0 ;
      RECT  333600.0 1621200.0 343800.0 1635000.0 ;
      RECT  333600.0 1648800.0 343800.0 1635000.0 ;
      RECT  333600.0 1648800.0 343800.0 1662600.0 ;
      RECT  333600.0 1676400.0 343800.0 1662600.0 ;
      RECT  333600.0 1676400.0 343800.0 1690200.0 ;
      RECT  333600.0 1704000.0 343800.0 1690200.0 ;
      RECT  333600.0 1704000.0 343800.0 1717800.0 ;
      RECT  333600.0 1731600.0 343800.0 1717800.0 ;
      RECT  333600.0 1731600.0 343800.0 1745400.0 ;
      RECT  333600.0 1759200.0 343800.0 1745400.0 ;
      RECT  333600.0 1759200.0 343800.0 1773000.0 ;
      RECT  333600.0 1786800.0 343800.0 1773000.0 ;
      RECT  333600.0 1786800.0 343800.0 1800600.0 ;
      RECT  333600.0 1814400.0 343800.0 1800600.0 ;
      RECT  333600.0 1814400.0 343800.0 1828200.0 ;
      RECT  333600.0 1842000.0 343800.0 1828200.0 ;
      RECT  333600.0 1842000.0 343800.0 1855800.0 ;
      RECT  333600.0 1869600.0 343800.0 1855800.0 ;
      RECT  333600.0 1869600.0 343800.0 1883400.0 ;
      RECT  333600.0 1897200.0 343800.0 1883400.0 ;
      RECT  333600.0 1897200.0 343800.0 1911000.0 ;
      RECT  333600.0 1924800.0 343800.0 1911000.0 ;
      RECT  333600.0 1924800.0 343800.0 1938600.0 ;
      RECT  333600.0 1952400.0 343800.0 1938600.0 ;
      RECT  333600.0 1952400.0 343800.0 1966200.0 ;
      RECT  333600.0 1980000.0 343800.0 1966200.0 ;
      RECT  333600.0 1980000.0 343800.0 1993800.0 ;
      RECT  333600.0 2007600.0 343800.0 1993800.0 ;
      RECT  333600.0 2007600.0 343800.0 2021400.0 ;
      RECT  333600.0 2035200.0 343800.0 2021400.0 ;
      RECT  333600.0 2035200.0 343800.0 2049000.0 ;
      RECT  333600.0 2062800.0 343800.0 2049000.0 ;
      RECT  333600.0 2062800.0 343800.0 2076600.0 ;
      RECT  333600.0 2090400.0 343800.0 2076600.0 ;
      RECT  333600.0 2090400.0 343800.0 2104200.0 ;
      RECT  333600.0 2118000.0 343800.0 2104200.0 ;
      RECT  333600.0 2118000.0 343800.0 2131800.0 ;
      RECT  333600.0 2145600.0 343800.0 2131800.0 ;
      RECT  343800.0 379200.0 354000.0 393000.0 ;
      RECT  343800.0 406800.0 354000.0 393000.0 ;
      RECT  343800.0 406800.0 354000.0 420600.0 ;
      RECT  343800.0 434400.0 354000.0 420600.0 ;
      RECT  343800.0 434400.0 354000.0 448200.0 ;
      RECT  343800.0 462000.0 354000.0 448200.0 ;
      RECT  343800.0 462000.0 354000.0 475800.0 ;
      RECT  343800.0 489600.0 354000.0 475800.0 ;
      RECT  343800.0 489600.0 354000.0 503400.0 ;
      RECT  343800.0 517200.0 354000.0 503400.0 ;
      RECT  343800.0 517200.0 354000.0 531000.0 ;
      RECT  343800.0 544800.0 354000.0 531000.0 ;
      RECT  343800.0 544800.0 354000.0 558600.0 ;
      RECT  343800.0 572400.0 354000.0 558600.0 ;
      RECT  343800.0 572400.0 354000.0 586200.0 ;
      RECT  343800.0 600000.0 354000.0 586200.0 ;
      RECT  343800.0 600000.0 354000.0 613800.0 ;
      RECT  343800.0 627600.0 354000.0 613800.0 ;
      RECT  343800.0 627600.0 354000.0 641400.0 ;
      RECT  343800.0 655200.0 354000.0 641400.0 ;
      RECT  343800.0 655200.0 354000.0 669000.0 ;
      RECT  343800.0 682800.0 354000.0 669000.0 ;
      RECT  343800.0 682800.0 354000.0 696600.0 ;
      RECT  343800.0 710400.0 354000.0 696600.0 ;
      RECT  343800.0 710400.0 354000.0 724200.0 ;
      RECT  343800.0 738000.0 354000.0 724200.0 ;
      RECT  343800.0 738000.0 354000.0 751800.0 ;
      RECT  343800.0 765600.0 354000.0 751800.0 ;
      RECT  343800.0 765600.0 354000.0 779400.0 ;
      RECT  343800.0 793200.0 354000.0 779400.0 ;
      RECT  343800.0 793200.0 354000.0 807000.0 ;
      RECT  343800.0 820800.0 354000.0 807000.0 ;
      RECT  343800.0 820800.0 354000.0 834600.0 ;
      RECT  343800.0 848400.0 354000.0 834600.0 ;
      RECT  343800.0 848400.0 354000.0 862200.0 ;
      RECT  343800.0 876000.0 354000.0 862200.0 ;
      RECT  343800.0 876000.0 354000.0 889800.0 ;
      RECT  343800.0 903600.0 354000.0 889800.0 ;
      RECT  343800.0 903600.0 354000.0 917400.0 ;
      RECT  343800.0 931200.0 354000.0 917400.0 ;
      RECT  343800.0 931200.0 354000.0 945000.0 ;
      RECT  343800.0 958800.0 354000.0 945000.0 ;
      RECT  343800.0 958800.0 354000.0 972600.0 ;
      RECT  343800.0 986400.0 354000.0 972600.0 ;
      RECT  343800.0 986400.0 354000.0 1000200.0 ;
      RECT  343800.0 1014000.0 354000.0 1000200.0 ;
      RECT  343800.0 1014000.0 354000.0 1027800.0 ;
      RECT  343800.0 1041600.0 354000.0 1027800.0 ;
      RECT  343800.0 1041600.0 354000.0 1055400.0 ;
      RECT  343800.0 1069200.0 354000.0 1055400.0 ;
      RECT  343800.0 1069200.0 354000.0 1083000.0 ;
      RECT  343800.0 1096800.0 354000.0 1083000.0 ;
      RECT  343800.0 1096800.0 354000.0 1110600.0 ;
      RECT  343800.0 1124400.0 354000.0 1110600.0 ;
      RECT  343800.0 1124400.0 354000.0 1138200.0 ;
      RECT  343800.0 1152000.0 354000.0 1138200.0 ;
      RECT  343800.0 1152000.0 354000.0 1165800.0 ;
      RECT  343800.0 1179600.0 354000.0 1165800.0 ;
      RECT  343800.0 1179600.0 354000.0 1193400.0 ;
      RECT  343800.0 1207200.0 354000.0 1193400.0 ;
      RECT  343800.0 1207200.0 354000.0 1221000.0 ;
      RECT  343800.0 1234800.0 354000.0 1221000.0 ;
      RECT  343800.0 1234800.0 354000.0 1248600.0 ;
      RECT  343800.0 1262400.0 354000.0 1248600.0 ;
      RECT  343800.0 1262400.0 354000.0 1276200.0 ;
      RECT  343800.0 1290000.0 354000.0 1276200.0 ;
      RECT  343800.0 1290000.0 354000.0 1303800.0 ;
      RECT  343800.0 1317600.0 354000.0 1303800.0 ;
      RECT  343800.0 1317600.0 354000.0 1331400.0 ;
      RECT  343800.0 1345200.0 354000.0 1331400.0 ;
      RECT  343800.0 1345200.0 354000.0 1359000.0 ;
      RECT  343800.0 1372800.0 354000.0 1359000.0 ;
      RECT  343800.0 1372800.0 354000.0 1386600.0 ;
      RECT  343800.0 1400400.0 354000.0 1386600.0 ;
      RECT  343800.0 1400400.0 354000.0 1414200.0 ;
      RECT  343800.0 1428000.0 354000.0 1414200.0 ;
      RECT  343800.0 1428000.0 354000.0 1441800.0 ;
      RECT  343800.0 1455600.0 354000.0 1441800.0 ;
      RECT  343800.0 1455600.0 354000.0 1469400.0 ;
      RECT  343800.0 1483200.0 354000.0 1469400.0 ;
      RECT  343800.0 1483200.0 354000.0 1497000.0 ;
      RECT  343800.0 1510800.0 354000.0 1497000.0 ;
      RECT  343800.0 1510800.0 354000.0 1524600.0 ;
      RECT  343800.0 1538400.0 354000.0 1524600.0 ;
      RECT  343800.0 1538400.0 354000.0 1552200.0 ;
      RECT  343800.0 1566000.0 354000.0 1552200.0 ;
      RECT  343800.0 1566000.0 354000.0 1579800.0 ;
      RECT  343800.0 1593600.0 354000.0 1579800.0 ;
      RECT  343800.0 1593600.0 354000.0 1607400.0 ;
      RECT  343800.0 1621200.0 354000.0 1607400.0 ;
      RECT  343800.0 1621200.0 354000.0 1635000.0 ;
      RECT  343800.0 1648800.0 354000.0 1635000.0 ;
      RECT  343800.0 1648800.0 354000.0 1662600.0 ;
      RECT  343800.0 1676400.0 354000.0 1662600.0 ;
      RECT  343800.0 1676400.0 354000.0 1690200.0 ;
      RECT  343800.0 1704000.0 354000.0 1690200.0 ;
      RECT  343800.0 1704000.0 354000.0 1717800.0 ;
      RECT  343800.0 1731600.0 354000.0 1717800.0 ;
      RECT  343800.0 1731600.0 354000.0 1745400.0 ;
      RECT  343800.0 1759200.0 354000.0 1745400.0 ;
      RECT  343800.0 1759200.0 354000.0 1773000.0 ;
      RECT  343800.0 1786800.0 354000.0 1773000.0 ;
      RECT  343800.0 1786800.0 354000.0 1800600.0 ;
      RECT  343800.0 1814400.0 354000.0 1800600.0 ;
      RECT  343800.0 1814400.0 354000.0 1828200.0 ;
      RECT  343800.0 1842000.0 354000.0 1828200.0 ;
      RECT  343800.0 1842000.0 354000.0 1855800.0 ;
      RECT  343800.0 1869600.0 354000.0 1855800.0 ;
      RECT  343800.0 1869600.0 354000.0 1883400.0 ;
      RECT  343800.0 1897200.0 354000.0 1883400.0 ;
      RECT  343800.0 1897200.0 354000.0 1911000.0 ;
      RECT  343800.0 1924800.0 354000.0 1911000.0 ;
      RECT  343800.0 1924800.0 354000.0 1938600.0 ;
      RECT  343800.0 1952400.0 354000.0 1938600.0 ;
      RECT  343800.0 1952400.0 354000.0 1966200.0 ;
      RECT  343800.0 1980000.0 354000.0 1966200.0 ;
      RECT  343800.0 1980000.0 354000.0 1993800.0 ;
      RECT  343800.0 2007600.0 354000.0 1993800.0 ;
      RECT  343800.0 2007600.0 354000.0 2021400.0 ;
      RECT  343800.0 2035200.0 354000.0 2021400.0 ;
      RECT  343800.0 2035200.0 354000.0 2049000.0 ;
      RECT  343800.0 2062800.0 354000.0 2049000.0 ;
      RECT  343800.0 2062800.0 354000.0 2076600.0 ;
      RECT  343800.0 2090400.0 354000.0 2076600.0 ;
      RECT  343800.0 2090400.0 354000.0 2104200.0 ;
      RECT  343800.0 2118000.0 354000.0 2104200.0 ;
      RECT  343800.0 2118000.0 354000.0 2131800.0 ;
      RECT  343800.0 2145600.0 354000.0 2131800.0 ;
      RECT  354000.0 379200.0 364200.0 393000.0 ;
      RECT  354000.0 406800.0 364200.0 393000.0 ;
      RECT  354000.0 406800.0 364200.0 420600.0 ;
      RECT  354000.0 434400.0 364200.0 420600.0 ;
      RECT  354000.0 434400.0 364200.0 448200.0 ;
      RECT  354000.0 462000.0 364200.0 448200.0 ;
      RECT  354000.0 462000.0 364200.0 475800.0 ;
      RECT  354000.0 489600.0 364200.0 475800.0 ;
      RECT  354000.0 489600.0 364200.0 503400.0 ;
      RECT  354000.0 517200.0 364200.0 503400.0 ;
      RECT  354000.0 517200.0 364200.0 531000.0 ;
      RECT  354000.0 544800.0 364200.0 531000.0 ;
      RECT  354000.0 544800.0 364200.0 558600.0 ;
      RECT  354000.0 572400.0 364200.0 558600.0 ;
      RECT  354000.0 572400.0 364200.0 586200.0 ;
      RECT  354000.0 600000.0 364200.0 586200.0 ;
      RECT  354000.0 600000.0 364200.0 613800.0 ;
      RECT  354000.0 627600.0 364200.0 613800.0 ;
      RECT  354000.0 627600.0 364200.0 641400.0 ;
      RECT  354000.0 655200.0 364200.0 641400.0 ;
      RECT  354000.0 655200.0 364200.0 669000.0 ;
      RECT  354000.0 682800.0 364200.0 669000.0 ;
      RECT  354000.0 682800.0 364200.0 696600.0 ;
      RECT  354000.0 710400.0 364200.0 696600.0 ;
      RECT  354000.0 710400.0 364200.0 724200.0 ;
      RECT  354000.0 738000.0 364200.0 724200.0 ;
      RECT  354000.0 738000.0 364200.0 751800.0 ;
      RECT  354000.0 765600.0 364200.0 751800.0 ;
      RECT  354000.0 765600.0 364200.0 779400.0 ;
      RECT  354000.0 793200.0 364200.0 779400.0 ;
      RECT  354000.0 793200.0 364200.0 807000.0 ;
      RECT  354000.0 820800.0 364200.0 807000.0 ;
      RECT  354000.0 820800.0 364200.0 834600.0 ;
      RECT  354000.0 848400.0 364200.0 834600.0 ;
      RECT  354000.0 848400.0 364200.0 862200.0 ;
      RECT  354000.0 876000.0 364200.0 862200.0 ;
      RECT  354000.0 876000.0 364200.0 889800.0 ;
      RECT  354000.0 903600.0 364200.0 889800.0 ;
      RECT  354000.0 903600.0 364200.0 917400.0 ;
      RECT  354000.0 931200.0 364200.0 917400.0 ;
      RECT  354000.0 931200.0 364200.0 945000.0 ;
      RECT  354000.0 958800.0 364200.0 945000.0 ;
      RECT  354000.0 958800.0 364200.0 972600.0 ;
      RECT  354000.0 986400.0 364200.0 972600.0 ;
      RECT  354000.0 986400.0 364200.0 1000200.0 ;
      RECT  354000.0 1014000.0 364200.0 1000200.0 ;
      RECT  354000.0 1014000.0 364200.0 1027800.0 ;
      RECT  354000.0 1041600.0 364200.0 1027800.0 ;
      RECT  354000.0 1041600.0 364200.0 1055400.0 ;
      RECT  354000.0 1069200.0 364200.0 1055400.0 ;
      RECT  354000.0 1069200.0 364200.0 1083000.0 ;
      RECT  354000.0 1096800.0 364200.0 1083000.0 ;
      RECT  354000.0 1096800.0 364200.0 1110600.0 ;
      RECT  354000.0 1124400.0 364200.0 1110600.0 ;
      RECT  354000.0 1124400.0 364200.0 1138200.0 ;
      RECT  354000.0 1152000.0 364200.0 1138200.0 ;
      RECT  354000.0 1152000.0 364200.0 1165800.0 ;
      RECT  354000.0 1179600.0 364200.0 1165800.0 ;
      RECT  354000.0 1179600.0 364200.0 1193400.0 ;
      RECT  354000.0 1207200.0 364200.0 1193400.0 ;
      RECT  354000.0 1207200.0 364200.0 1221000.0 ;
      RECT  354000.0 1234800.0 364200.0 1221000.0 ;
      RECT  354000.0 1234800.0 364200.0 1248600.0 ;
      RECT  354000.0 1262400.0 364200.0 1248600.0 ;
      RECT  354000.0 1262400.0 364200.0 1276200.0 ;
      RECT  354000.0 1290000.0 364200.0 1276200.0 ;
      RECT  354000.0 1290000.0 364200.0 1303800.0 ;
      RECT  354000.0 1317600.0 364200.0 1303800.0 ;
      RECT  354000.0 1317600.0 364200.0 1331400.0 ;
      RECT  354000.0 1345200.0 364200.0 1331400.0 ;
      RECT  354000.0 1345200.0 364200.0 1359000.0 ;
      RECT  354000.0 1372800.0 364200.0 1359000.0 ;
      RECT  354000.0 1372800.0 364200.0 1386600.0 ;
      RECT  354000.0 1400400.0 364200.0 1386600.0 ;
      RECT  354000.0 1400400.0 364200.0 1414200.0 ;
      RECT  354000.0 1428000.0 364200.0 1414200.0 ;
      RECT  354000.0 1428000.0 364200.0 1441800.0 ;
      RECT  354000.0 1455600.0 364200.0 1441800.0 ;
      RECT  354000.0 1455600.0 364200.0 1469400.0 ;
      RECT  354000.0 1483200.0 364200.0 1469400.0 ;
      RECT  354000.0 1483200.0 364200.0 1497000.0 ;
      RECT  354000.0 1510800.0 364200.0 1497000.0 ;
      RECT  354000.0 1510800.0 364200.0 1524600.0 ;
      RECT  354000.0 1538400.0 364200.0 1524600.0 ;
      RECT  354000.0 1538400.0 364200.0 1552200.0 ;
      RECT  354000.0 1566000.0 364200.0 1552200.0 ;
      RECT  354000.0 1566000.0 364200.0 1579800.0 ;
      RECT  354000.0 1593600.0 364200.0 1579800.0 ;
      RECT  354000.0 1593600.0 364200.0 1607400.0 ;
      RECT  354000.0 1621200.0 364200.0 1607400.0 ;
      RECT  354000.0 1621200.0 364200.0 1635000.0 ;
      RECT  354000.0 1648800.0 364200.0 1635000.0 ;
      RECT  354000.0 1648800.0 364200.0 1662600.0 ;
      RECT  354000.0 1676400.0 364200.0 1662600.0 ;
      RECT  354000.0 1676400.0 364200.0 1690200.0 ;
      RECT  354000.0 1704000.0 364200.0 1690200.0 ;
      RECT  354000.0 1704000.0 364200.0 1717800.0 ;
      RECT  354000.0 1731600.0 364200.0 1717800.0 ;
      RECT  354000.0 1731600.0 364200.0 1745400.0 ;
      RECT  354000.0 1759200.0 364200.0 1745400.0 ;
      RECT  354000.0 1759200.0 364200.0 1773000.0 ;
      RECT  354000.0 1786800.0 364200.0 1773000.0 ;
      RECT  354000.0 1786800.0 364200.0 1800600.0 ;
      RECT  354000.0 1814400.0 364200.0 1800600.0 ;
      RECT  354000.0 1814400.0 364200.0 1828200.0 ;
      RECT  354000.0 1842000.0 364200.0 1828200.0 ;
      RECT  354000.0 1842000.0 364200.0 1855800.0 ;
      RECT  354000.0 1869600.0 364200.0 1855800.0 ;
      RECT  354000.0 1869600.0 364200.0 1883400.0 ;
      RECT  354000.0 1897200.0 364200.0 1883400.0 ;
      RECT  354000.0 1897200.0 364200.0 1911000.0 ;
      RECT  354000.0 1924800.0 364200.0 1911000.0 ;
      RECT  354000.0 1924800.0 364200.0 1938600.0 ;
      RECT  354000.0 1952400.0 364200.0 1938600.0 ;
      RECT  354000.0 1952400.0 364200.0 1966200.0 ;
      RECT  354000.0 1980000.0 364200.0 1966200.0 ;
      RECT  354000.0 1980000.0 364200.0 1993800.0 ;
      RECT  354000.0 2007600.0 364200.0 1993800.0 ;
      RECT  354000.0 2007600.0 364200.0 2021400.0 ;
      RECT  354000.0 2035200.0 364200.0 2021400.0 ;
      RECT  354000.0 2035200.0 364200.0 2049000.0 ;
      RECT  354000.0 2062800.0 364200.0 2049000.0 ;
      RECT  354000.0 2062800.0 364200.0 2076600.0 ;
      RECT  354000.0 2090400.0 364200.0 2076600.0 ;
      RECT  354000.0 2090400.0 364200.0 2104200.0 ;
      RECT  354000.0 2118000.0 364200.0 2104200.0 ;
      RECT  354000.0 2118000.0 364200.0 2131800.0 ;
      RECT  354000.0 2145600.0 364200.0 2131800.0 ;
      RECT  364200.0 379200.0 374400.0 393000.0 ;
      RECT  364200.0 406800.0 374400.0 393000.0 ;
      RECT  364200.0 406800.0 374400.0 420600.0 ;
      RECT  364200.0 434400.0 374400.0 420600.0 ;
      RECT  364200.0 434400.0 374400.0 448200.0 ;
      RECT  364200.0 462000.0 374400.0 448200.0 ;
      RECT  364200.0 462000.0 374400.0 475800.0 ;
      RECT  364200.0 489600.0 374400.0 475800.0 ;
      RECT  364200.0 489600.0 374400.0 503400.0 ;
      RECT  364200.0 517200.0 374400.0 503400.0 ;
      RECT  364200.0 517200.0 374400.0 531000.0 ;
      RECT  364200.0 544800.0 374400.0 531000.0 ;
      RECT  364200.0 544800.0 374400.0 558600.0 ;
      RECT  364200.0 572400.0 374400.0 558600.0 ;
      RECT  364200.0 572400.0 374400.0 586200.0 ;
      RECT  364200.0 600000.0 374400.0 586200.0 ;
      RECT  364200.0 600000.0 374400.0 613800.0 ;
      RECT  364200.0 627600.0 374400.0 613800.0 ;
      RECT  364200.0 627600.0 374400.0 641400.0 ;
      RECT  364200.0 655200.0 374400.0 641400.0 ;
      RECT  364200.0 655200.0 374400.0 669000.0 ;
      RECT  364200.0 682800.0 374400.0 669000.0 ;
      RECT  364200.0 682800.0 374400.0 696600.0 ;
      RECT  364200.0 710400.0 374400.0 696600.0 ;
      RECT  364200.0 710400.0 374400.0 724200.0 ;
      RECT  364200.0 738000.0 374400.0 724200.0 ;
      RECT  364200.0 738000.0 374400.0 751800.0 ;
      RECT  364200.0 765600.0 374400.0 751800.0 ;
      RECT  364200.0 765600.0 374400.0 779400.0 ;
      RECT  364200.0 793200.0 374400.0 779400.0 ;
      RECT  364200.0 793200.0 374400.0 807000.0 ;
      RECT  364200.0 820800.0 374400.0 807000.0 ;
      RECT  364200.0 820800.0 374400.0 834600.0 ;
      RECT  364200.0 848400.0 374400.0 834600.0 ;
      RECT  364200.0 848400.0 374400.0 862200.0 ;
      RECT  364200.0 876000.0 374400.0 862200.0 ;
      RECT  364200.0 876000.0 374400.0 889800.0 ;
      RECT  364200.0 903600.0 374400.0 889800.0 ;
      RECT  364200.0 903600.0 374400.0 917400.0 ;
      RECT  364200.0 931200.0 374400.0 917400.0 ;
      RECT  364200.0 931200.0 374400.0 945000.0 ;
      RECT  364200.0 958800.0 374400.0 945000.0 ;
      RECT  364200.0 958800.0 374400.0 972600.0 ;
      RECT  364200.0 986400.0 374400.0 972600.0 ;
      RECT  364200.0 986400.0 374400.0 1000200.0 ;
      RECT  364200.0 1014000.0 374400.0 1000200.0 ;
      RECT  364200.0 1014000.0 374400.0 1027800.0 ;
      RECT  364200.0 1041600.0 374400.0 1027800.0 ;
      RECT  364200.0 1041600.0 374400.0 1055400.0 ;
      RECT  364200.0 1069200.0 374400.0 1055400.0 ;
      RECT  364200.0 1069200.0 374400.0 1083000.0 ;
      RECT  364200.0 1096800.0 374400.0 1083000.0 ;
      RECT  364200.0 1096800.0 374400.0 1110600.0 ;
      RECT  364200.0 1124400.0 374400.0 1110600.0 ;
      RECT  364200.0 1124400.0 374400.0 1138200.0 ;
      RECT  364200.0 1152000.0 374400.0 1138200.0 ;
      RECT  364200.0 1152000.0 374400.0 1165800.0 ;
      RECT  364200.0 1179600.0 374400.0 1165800.0 ;
      RECT  364200.0 1179600.0 374400.0 1193400.0 ;
      RECT  364200.0 1207200.0 374400.0 1193400.0 ;
      RECT  364200.0 1207200.0 374400.0 1221000.0 ;
      RECT  364200.0 1234800.0 374400.0 1221000.0 ;
      RECT  364200.0 1234800.0 374400.0 1248600.0 ;
      RECT  364200.0 1262400.0 374400.0 1248600.0 ;
      RECT  364200.0 1262400.0 374400.0 1276200.0 ;
      RECT  364200.0 1290000.0 374400.0 1276200.0 ;
      RECT  364200.0 1290000.0 374400.0 1303800.0 ;
      RECT  364200.0 1317600.0 374400.0 1303800.0 ;
      RECT  364200.0 1317600.0 374400.0 1331400.0 ;
      RECT  364200.0 1345200.0 374400.0 1331400.0 ;
      RECT  364200.0 1345200.0 374400.0 1359000.0 ;
      RECT  364200.0 1372800.0 374400.0 1359000.0 ;
      RECT  364200.0 1372800.0 374400.0 1386600.0 ;
      RECT  364200.0 1400400.0 374400.0 1386600.0 ;
      RECT  364200.0 1400400.0 374400.0 1414200.0 ;
      RECT  364200.0 1428000.0 374400.0 1414200.0 ;
      RECT  364200.0 1428000.0 374400.0 1441800.0 ;
      RECT  364200.0 1455600.0 374400.0 1441800.0 ;
      RECT  364200.0 1455600.0 374400.0 1469400.0 ;
      RECT  364200.0 1483200.0 374400.0 1469400.0 ;
      RECT  364200.0 1483200.0 374400.0 1497000.0 ;
      RECT  364200.0 1510800.0 374400.0 1497000.0 ;
      RECT  364200.0 1510800.0 374400.0 1524600.0 ;
      RECT  364200.0 1538400.0 374400.0 1524600.0 ;
      RECT  364200.0 1538400.0 374400.0 1552200.0 ;
      RECT  364200.0 1566000.0 374400.0 1552200.0 ;
      RECT  364200.0 1566000.0 374400.0 1579800.0 ;
      RECT  364200.0 1593600.0 374400.0 1579800.0 ;
      RECT  364200.0 1593600.0 374400.0 1607400.0 ;
      RECT  364200.0 1621200.0 374400.0 1607400.0 ;
      RECT  364200.0 1621200.0 374400.0 1635000.0 ;
      RECT  364200.0 1648800.0 374400.0 1635000.0 ;
      RECT  364200.0 1648800.0 374400.0 1662600.0 ;
      RECT  364200.0 1676400.0 374400.0 1662600.0 ;
      RECT  364200.0 1676400.0 374400.0 1690200.0 ;
      RECT  364200.0 1704000.0 374400.0 1690200.0 ;
      RECT  364200.0 1704000.0 374400.0 1717800.0 ;
      RECT  364200.0 1731600.0 374400.0 1717800.0 ;
      RECT  364200.0 1731600.0 374400.0 1745400.0 ;
      RECT  364200.0 1759200.0 374400.0 1745400.0 ;
      RECT  364200.0 1759200.0 374400.0 1773000.0 ;
      RECT  364200.0 1786800.0 374400.0 1773000.0 ;
      RECT  364200.0 1786800.0 374400.0 1800600.0 ;
      RECT  364200.0 1814400.0 374400.0 1800600.0 ;
      RECT  364200.0 1814400.0 374400.0 1828200.0 ;
      RECT  364200.0 1842000.0 374400.0 1828200.0 ;
      RECT  364200.0 1842000.0 374400.0 1855800.0 ;
      RECT  364200.0 1869600.0 374400.0 1855800.0 ;
      RECT  364200.0 1869600.0 374400.0 1883400.0 ;
      RECT  364200.0 1897200.0 374400.0 1883400.0 ;
      RECT  364200.0 1897200.0 374400.0 1911000.0 ;
      RECT  364200.0 1924800.0 374400.0 1911000.0 ;
      RECT  364200.0 1924800.0 374400.0 1938600.0 ;
      RECT  364200.0 1952400.0 374400.0 1938600.0 ;
      RECT  364200.0 1952400.0 374400.0 1966200.0 ;
      RECT  364200.0 1980000.0 374400.0 1966200.0 ;
      RECT  364200.0 1980000.0 374400.0 1993800.0 ;
      RECT  364200.0 2007600.0 374400.0 1993800.0 ;
      RECT  364200.0 2007600.0 374400.0 2021400.0 ;
      RECT  364200.0 2035200.0 374400.0 2021400.0 ;
      RECT  364200.0 2035200.0 374400.0 2049000.0 ;
      RECT  364200.0 2062800.0 374400.0 2049000.0 ;
      RECT  364200.0 2062800.0 374400.0 2076600.0 ;
      RECT  364200.0 2090400.0 374400.0 2076600.0 ;
      RECT  364200.0 2090400.0 374400.0 2104200.0 ;
      RECT  364200.0 2118000.0 374400.0 2104200.0 ;
      RECT  364200.0 2118000.0 374400.0 2131800.0 ;
      RECT  364200.0 2145600.0 374400.0 2131800.0 ;
      RECT  374400.0 379200.0 384600.0 393000.0 ;
      RECT  374400.0 406800.0 384600.0 393000.0 ;
      RECT  374400.0 406800.0 384600.0 420600.0 ;
      RECT  374400.0 434400.0 384600.0 420600.0 ;
      RECT  374400.0 434400.0 384600.0 448200.0 ;
      RECT  374400.0 462000.0 384600.0 448200.0 ;
      RECT  374400.0 462000.0 384600.0 475800.0 ;
      RECT  374400.0 489600.0 384600.0 475800.0 ;
      RECT  374400.0 489600.0 384600.0 503400.0 ;
      RECT  374400.0 517200.0 384600.0 503400.0 ;
      RECT  374400.0 517200.0 384600.0 531000.0 ;
      RECT  374400.0 544800.0 384600.0 531000.0 ;
      RECT  374400.0 544800.0 384600.0 558600.0 ;
      RECT  374400.0 572400.0 384600.0 558600.0 ;
      RECT  374400.0 572400.0 384600.0 586200.0 ;
      RECT  374400.0 600000.0 384600.0 586200.0 ;
      RECT  374400.0 600000.0 384600.0 613800.0 ;
      RECT  374400.0 627600.0 384600.0 613800.0 ;
      RECT  374400.0 627600.0 384600.0 641400.0 ;
      RECT  374400.0 655200.0 384600.0 641400.0 ;
      RECT  374400.0 655200.0 384600.0 669000.0 ;
      RECT  374400.0 682800.0 384600.0 669000.0 ;
      RECT  374400.0 682800.0 384600.0 696600.0 ;
      RECT  374400.0 710400.0 384600.0 696600.0 ;
      RECT  374400.0 710400.0 384600.0 724200.0 ;
      RECT  374400.0 738000.0 384600.0 724200.0 ;
      RECT  374400.0 738000.0 384600.0 751800.0 ;
      RECT  374400.0 765600.0 384600.0 751800.0 ;
      RECT  374400.0 765600.0 384600.0 779400.0 ;
      RECT  374400.0 793200.0 384600.0 779400.0 ;
      RECT  374400.0 793200.0 384600.0 807000.0 ;
      RECT  374400.0 820800.0 384600.0 807000.0 ;
      RECT  374400.0 820800.0 384600.0 834600.0 ;
      RECT  374400.0 848400.0 384600.0 834600.0 ;
      RECT  374400.0 848400.0 384600.0 862200.0 ;
      RECT  374400.0 876000.0 384600.0 862200.0 ;
      RECT  374400.0 876000.0 384600.0 889800.0 ;
      RECT  374400.0 903600.0 384600.0 889800.0 ;
      RECT  374400.0 903600.0 384600.0 917400.0 ;
      RECT  374400.0 931200.0 384600.0 917400.0 ;
      RECT  374400.0 931200.0 384600.0 945000.0 ;
      RECT  374400.0 958800.0 384600.0 945000.0 ;
      RECT  374400.0 958800.0 384600.0 972600.0 ;
      RECT  374400.0 986400.0 384600.0 972600.0 ;
      RECT  374400.0 986400.0 384600.0 1000200.0 ;
      RECT  374400.0 1014000.0 384600.0 1000200.0 ;
      RECT  374400.0 1014000.0 384600.0 1027800.0 ;
      RECT  374400.0 1041600.0 384600.0 1027800.0 ;
      RECT  374400.0 1041600.0 384600.0 1055400.0 ;
      RECT  374400.0 1069200.0 384600.0 1055400.0 ;
      RECT  374400.0 1069200.0 384600.0 1083000.0 ;
      RECT  374400.0 1096800.0 384600.0 1083000.0 ;
      RECT  374400.0 1096800.0 384600.0 1110600.0 ;
      RECT  374400.0 1124400.0 384600.0 1110600.0 ;
      RECT  374400.0 1124400.0 384600.0 1138200.0 ;
      RECT  374400.0 1152000.0 384600.0 1138200.0 ;
      RECT  374400.0 1152000.0 384600.0 1165800.0 ;
      RECT  374400.0 1179600.0 384600.0 1165800.0 ;
      RECT  374400.0 1179600.0 384600.0 1193400.0 ;
      RECT  374400.0 1207200.0 384600.0 1193400.0 ;
      RECT  374400.0 1207200.0 384600.0 1221000.0 ;
      RECT  374400.0 1234800.0 384600.0 1221000.0 ;
      RECT  374400.0 1234800.0 384600.0 1248600.0 ;
      RECT  374400.0 1262400.0 384600.0 1248600.0 ;
      RECT  374400.0 1262400.0 384600.0 1276200.0 ;
      RECT  374400.0 1290000.0 384600.0 1276200.0 ;
      RECT  374400.0 1290000.0 384600.0 1303800.0 ;
      RECT  374400.0 1317600.0 384600.0 1303800.0 ;
      RECT  374400.0 1317600.0 384600.0 1331400.0 ;
      RECT  374400.0 1345200.0 384600.0 1331400.0 ;
      RECT  374400.0 1345200.0 384600.0 1359000.0 ;
      RECT  374400.0 1372800.0 384600.0 1359000.0 ;
      RECT  374400.0 1372800.0 384600.0 1386600.0 ;
      RECT  374400.0 1400400.0 384600.0 1386600.0 ;
      RECT  374400.0 1400400.0 384600.0 1414200.0 ;
      RECT  374400.0 1428000.0 384600.0 1414200.0 ;
      RECT  374400.0 1428000.0 384600.0 1441800.0 ;
      RECT  374400.0 1455600.0 384600.0 1441800.0 ;
      RECT  374400.0 1455600.0 384600.0 1469400.0 ;
      RECT  374400.0 1483200.0 384600.0 1469400.0 ;
      RECT  374400.0 1483200.0 384600.0 1497000.0 ;
      RECT  374400.0 1510800.0 384600.0 1497000.0 ;
      RECT  374400.0 1510800.0 384600.0 1524600.0 ;
      RECT  374400.0 1538400.0 384600.0 1524600.0 ;
      RECT  374400.0 1538400.0 384600.0 1552200.0 ;
      RECT  374400.0 1566000.0 384600.0 1552200.0 ;
      RECT  374400.0 1566000.0 384600.0 1579800.0 ;
      RECT  374400.0 1593600.0 384600.0 1579800.0 ;
      RECT  374400.0 1593600.0 384600.0 1607400.0 ;
      RECT  374400.0 1621200.0 384600.0 1607400.0 ;
      RECT  374400.0 1621200.0 384600.0 1635000.0 ;
      RECT  374400.0 1648800.0 384600.0 1635000.0 ;
      RECT  374400.0 1648800.0 384600.0 1662600.0 ;
      RECT  374400.0 1676400.0 384600.0 1662600.0 ;
      RECT  374400.0 1676400.0 384600.0 1690200.0 ;
      RECT  374400.0 1704000.0 384600.0 1690200.0 ;
      RECT  374400.0 1704000.0 384600.0 1717800.0 ;
      RECT  374400.0 1731600.0 384600.0 1717800.0 ;
      RECT  374400.0 1731600.0 384600.0 1745400.0 ;
      RECT  374400.0 1759200.0 384600.0 1745400.0 ;
      RECT  374400.0 1759200.0 384600.0 1773000.0 ;
      RECT  374400.0 1786800.0 384600.0 1773000.0 ;
      RECT  374400.0 1786800.0 384600.0 1800600.0 ;
      RECT  374400.0 1814400.0 384600.0 1800600.0 ;
      RECT  374400.0 1814400.0 384600.0 1828200.0 ;
      RECT  374400.0 1842000.0 384600.0 1828200.0 ;
      RECT  374400.0 1842000.0 384600.0 1855800.0 ;
      RECT  374400.0 1869600.0 384600.0 1855800.0 ;
      RECT  374400.0 1869600.0 384600.0 1883400.0 ;
      RECT  374400.0 1897200.0 384600.0 1883400.0 ;
      RECT  374400.0 1897200.0 384600.0 1911000.0 ;
      RECT  374400.0 1924800.0 384600.0 1911000.0 ;
      RECT  374400.0 1924800.0 384600.0 1938600.0 ;
      RECT  374400.0 1952400.0 384600.0 1938600.0 ;
      RECT  374400.0 1952400.0 384600.0 1966200.0 ;
      RECT  374400.0 1980000.0 384600.0 1966200.0 ;
      RECT  374400.0 1980000.0 384600.0 1993800.0 ;
      RECT  374400.0 2007600.0 384600.0 1993800.0 ;
      RECT  374400.0 2007600.0 384600.0 2021400.0 ;
      RECT  374400.0 2035200.0 384600.0 2021400.0 ;
      RECT  374400.0 2035200.0 384600.0 2049000.0 ;
      RECT  374400.0 2062800.0 384600.0 2049000.0 ;
      RECT  374400.0 2062800.0 384600.0 2076600.0 ;
      RECT  374400.0 2090400.0 384600.0 2076600.0 ;
      RECT  374400.0 2090400.0 384600.0 2104200.0 ;
      RECT  374400.0 2118000.0 384600.0 2104200.0 ;
      RECT  374400.0 2118000.0 384600.0 2131800.0 ;
      RECT  374400.0 2145600.0 384600.0 2131800.0 ;
      RECT  384600.0 379200.0 394800.0 393000.0 ;
      RECT  384600.0 406800.0 394800.0 393000.0 ;
      RECT  384600.0 406800.0 394800.0 420600.0 ;
      RECT  384600.0 434400.0 394800.0 420600.0 ;
      RECT  384600.0 434400.0 394800.0 448200.0 ;
      RECT  384600.0 462000.0 394800.0 448200.0 ;
      RECT  384600.0 462000.0 394800.0 475800.0 ;
      RECT  384600.0 489600.0 394800.0 475800.0 ;
      RECT  384600.0 489600.0 394800.0 503400.0 ;
      RECT  384600.0 517200.0 394800.0 503400.0 ;
      RECT  384600.0 517200.0 394800.0 531000.0 ;
      RECT  384600.0 544800.0 394800.0 531000.0 ;
      RECT  384600.0 544800.0 394800.0 558600.0 ;
      RECT  384600.0 572400.0 394800.0 558600.0 ;
      RECT  384600.0 572400.0 394800.0 586200.0 ;
      RECT  384600.0 600000.0 394800.0 586200.0 ;
      RECT  384600.0 600000.0 394800.0 613800.0 ;
      RECT  384600.0 627600.0 394800.0 613800.0 ;
      RECT  384600.0 627600.0 394800.0 641400.0 ;
      RECT  384600.0 655200.0 394800.0 641400.0 ;
      RECT  384600.0 655200.0 394800.0 669000.0 ;
      RECT  384600.0 682800.0 394800.0 669000.0 ;
      RECT  384600.0 682800.0 394800.0 696600.0 ;
      RECT  384600.0 710400.0 394800.0 696600.0 ;
      RECT  384600.0 710400.0 394800.0 724200.0 ;
      RECT  384600.0 738000.0 394800.0 724200.0 ;
      RECT  384600.0 738000.0 394800.0 751800.0 ;
      RECT  384600.0 765600.0 394800.0 751800.0 ;
      RECT  384600.0 765600.0 394800.0 779400.0 ;
      RECT  384600.0 793200.0 394800.0 779400.0 ;
      RECT  384600.0 793200.0 394800.0 807000.0 ;
      RECT  384600.0 820800.0 394800.0 807000.0 ;
      RECT  384600.0 820800.0 394800.0 834600.0 ;
      RECT  384600.0 848400.0 394800.0 834600.0 ;
      RECT  384600.0 848400.0 394800.0 862200.0 ;
      RECT  384600.0 876000.0 394800.0 862200.0 ;
      RECT  384600.0 876000.0 394800.0 889800.0 ;
      RECT  384600.0 903600.0 394800.0 889800.0 ;
      RECT  384600.0 903600.0 394800.0 917400.0 ;
      RECT  384600.0 931200.0 394800.0 917400.0 ;
      RECT  384600.0 931200.0 394800.0 945000.0 ;
      RECT  384600.0 958800.0 394800.0 945000.0 ;
      RECT  384600.0 958800.0 394800.0 972600.0 ;
      RECT  384600.0 986400.0 394800.0 972600.0 ;
      RECT  384600.0 986400.0 394800.0 1000200.0 ;
      RECT  384600.0 1014000.0 394800.0 1000200.0 ;
      RECT  384600.0 1014000.0 394800.0 1027800.0 ;
      RECT  384600.0 1041600.0 394800.0 1027800.0 ;
      RECT  384600.0 1041600.0 394800.0 1055400.0 ;
      RECT  384600.0 1069200.0 394800.0 1055400.0 ;
      RECT  384600.0 1069200.0 394800.0 1083000.0 ;
      RECT  384600.0 1096800.0 394800.0 1083000.0 ;
      RECT  384600.0 1096800.0 394800.0 1110600.0 ;
      RECT  384600.0 1124400.0 394800.0 1110600.0 ;
      RECT  384600.0 1124400.0 394800.0 1138200.0 ;
      RECT  384600.0 1152000.0 394800.0 1138200.0 ;
      RECT  384600.0 1152000.0 394800.0 1165800.0 ;
      RECT  384600.0 1179600.0 394800.0 1165800.0 ;
      RECT  384600.0 1179600.0 394800.0 1193400.0 ;
      RECT  384600.0 1207200.0 394800.0 1193400.0 ;
      RECT  384600.0 1207200.0 394800.0 1221000.0 ;
      RECT  384600.0 1234800.0 394800.0 1221000.0 ;
      RECT  384600.0 1234800.0 394800.0 1248600.0 ;
      RECT  384600.0 1262400.0 394800.0 1248600.0 ;
      RECT  384600.0 1262400.0 394800.0 1276200.0 ;
      RECT  384600.0 1290000.0 394800.0 1276200.0 ;
      RECT  384600.0 1290000.0 394800.0 1303800.0 ;
      RECT  384600.0 1317600.0 394800.0 1303800.0 ;
      RECT  384600.0 1317600.0 394800.0 1331400.0 ;
      RECT  384600.0 1345200.0 394800.0 1331400.0 ;
      RECT  384600.0 1345200.0 394800.0 1359000.0 ;
      RECT  384600.0 1372800.0 394800.0 1359000.0 ;
      RECT  384600.0 1372800.0 394800.0 1386600.0 ;
      RECT  384600.0 1400400.0 394800.0 1386600.0 ;
      RECT  384600.0 1400400.0 394800.0 1414200.0 ;
      RECT  384600.0 1428000.0 394800.0 1414200.0 ;
      RECT  384600.0 1428000.0 394800.0 1441800.0 ;
      RECT  384600.0 1455600.0 394800.0 1441800.0 ;
      RECT  384600.0 1455600.0 394800.0 1469400.0 ;
      RECT  384600.0 1483200.0 394800.0 1469400.0 ;
      RECT  384600.0 1483200.0 394800.0 1497000.0 ;
      RECT  384600.0 1510800.0 394800.0 1497000.0 ;
      RECT  384600.0 1510800.0 394800.0 1524600.0 ;
      RECT  384600.0 1538400.0 394800.0 1524600.0 ;
      RECT  384600.0 1538400.0 394800.0 1552200.0 ;
      RECT  384600.0 1566000.0 394800.0 1552200.0 ;
      RECT  384600.0 1566000.0 394800.0 1579800.0 ;
      RECT  384600.0 1593600.0 394800.0 1579800.0 ;
      RECT  384600.0 1593600.0 394800.0 1607400.0 ;
      RECT  384600.0 1621200.0 394800.0 1607400.0 ;
      RECT  384600.0 1621200.0 394800.0 1635000.0 ;
      RECT  384600.0 1648800.0 394800.0 1635000.0 ;
      RECT  384600.0 1648800.0 394800.0 1662600.0 ;
      RECT  384600.0 1676400.0 394800.0 1662600.0 ;
      RECT  384600.0 1676400.0 394800.0 1690200.0 ;
      RECT  384600.0 1704000.0 394800.0 1690200.0 ;
      RECT  384600.0 1704000.0 394800.0 1717800.0 ;
      RECT  384600.0 1731600.0 394800.0 1717800.0 ;
      RECT  384600.0 1731600.0 394800.0 1745400.0 ;
      RECT  384600.0 1759200.0 394800.0 1745400.0 ;
      RECT  384600.0 1759200.0 394800.0 1773000.0 ;
      RECT  384600.0 1786800.0 394800.0 1773000.0 ;
      RECT  384600.0 1786800.0 394800.0 1800600.0 ;
      RECT  384600.0 1814400.0 394800.0 1800600.0 ;
      RECT  384600.0 1814400.0 394800.0 1828200.0 ;
      RECT  384600.0 1842000.0 394800.0 1828200.0 ;
      RECT  384600.0 1842000.0 394800.0 1855800.0 ;
      RECT  384600.0 1869600.0 394800.0 1855800.0 ;
      RECT  384600.0 1869600.0 394800.0 1883400.0 ;
      RECT  384600.0 1897200.0 394800.0 1883400.0 ;
      RECT  384600.0 1897200.0 394800.0 1911000.0 ;
      RECT  384600.0 1924800.0 394800.0 1911000.0 ;
      RECT  384600.0 1924800.0 394800.0 1938600.0 ;
      RECT  384600.0 1952400.0 394800.0 1938600.0 ;
      RECT  384600.0 1952400.0 394800.0 1966200.0 ;
      RECT  384600.0 1980000.0 394800.0 1966200.0 ;
      RECT  384600.0 1980000.0 394800.0 1993800.0 ;
      RECT  384600.0 2007600.0 394800.0 1993800.0 ;
      RECT  384600.0 2007600.0 394800.0 2021400.0 ;
      RECT  384600.0 2035200.0 394800.0 2021400.0 ;
      RECT  384600.0 2035200.0 394800.0 2049000.0 ;
      RECT  384600.0 2062800.0 394800.0 2049000.0 ;
      RECT  384600.0 2062800.0 394800.0 2076600.0 ;
      RECT  384600.0 2090400.0 394800.0 2076600.0 ;
      RECT  384600.0 2090400.0 394800.0 2104200.0 ;
      RECT  384600.0 2118000.0 394800.0 2104200.0 ;
      RECT  384600.0 2118000.0 394800.0 2131800.0 ;
      RECT  384600.0 2145600.0 394800.0 2131800.0 ;
      RECT  394800.0 379200.0 405000.0 393000.0 ;
      RECT  394800.0 406800.0 405000.0 393000.0 ;
      RECT  394800.0 406800.0 405000.0 420600.0 ;
      RECT  394800.0 434400.0 405000.0 420600.0 ;
      RECT  394800.0 434400.0 405000.0 448200.0 ;
      RECT  394800.0 462000.0 405000.0 448200.0 ;
      RECT  394800.0 462000.0 405000.0 475800.0 ;
      RECT  394800.0 489600.0 405000.0 475800.0 ;
      RECT  394800.0 489600.0 405000.0 503400.0 ;
      RECT  394800.0 517200.0 405000.0 503400.0 ;
      RECT  394800.0 517200.0 405000.0 531000.0 ;
      RECT  394800.0 544800.0 405000.0 531000.0 ;
      RECT  394800.0 544800.0 405000.0 558600.0 ;
      RECT  394800.0 572400.0 405000.0 558600.0 ;
      RECT  394800.0 572400.0 405000.0 586200.0 ;
      RECT  394800.0 600000.0 405000.0 586200.0 ;
      RECT  394800.0 600000.0 405000.0 613800.0 ;
      RECT  394800.0 627600.0 405000.0 613800.0 ;
      RECT  394800.0 627600.0 405000.0 641400.0 ;
      RECT  394800.0 655200.0 405000.0 641400.0 ;
      RECT  394800.0 655200.0 405000.0 669000.0 ;
      RECT  394800.0 682800.0 405000.0 669000.0 ;
      RECT  394800.0 682800.0 405000.0 696600.0 ;
      RECT  394800.0 710400.0 405000.0 696600.0 ;
      RECT  394800.0 710400.0 405000.0 724200.0 ;
      RECT  394800.0 738000.0 405000.0 724200.0 ;
      RECT  394800.0 738000.0 405000.0 751800.0 ;
      RECT  394800.0 765600.0 405000.0 751800.0 ;
      RECT  394800.0 765600.0 405000.0 779400.0 ;
      RECT  394800.0 793200.0 405000.0 779400.0 ;
      RECT  394800.0 793200.0 405000.0 807000.0 ;
      RECT  394800.0 820800.0 405000.0 807000.0 ;
      RECT  394800.0 820800.0 405000.0 834600.0 ;
      RECT  394800.0 848400.0 405000.0 834600.0 ;
      RECT  394800.0 848400.0 405000.0 862200.0 ;
      RECT  394800.0 876000.0 405000.0 862200.0 ;
      RECT  394800.0 876000.0 405000.0 889800.0 ;
      RECT  394800.0 903600.0 405000.0 889800.0 ;
      RECT  394800.0 903600.0 405000.0 917400.0 ;
      RECT  394800.0 931200.0 405000.0 917400.0 ;
      RECT  394800.0 931200.0 405000.0 945000.0 ;
      RECT  394800.0 958800.0 405000.0 945000.0 ;
      RECT  394800.0 958800.0 405000.0 972600.0 ;
      RECT  394800.0 986400.0 405000.0 972600.0 ;
      RECT  394800.0 986400.0 405000.0 1000200.0 ;
      RECT  394800.0 1014000.0 405000.0 1000200.0 ;
      RECT  394800.0 1014000.0 405000.0 1027800.0 ;
      RECT  394800.0 1041600.0 405000.0 1027800.0 ;
      RECT  394800.0 1041600.0 405000.0 1055400.0 ;
      RECT  394800.0 1069200.0 405000.0 1055400.0 ;
      RECT  394800.0 1069200.0 405000.0 1083000.0 ;
      RECT  394800.0 1096800.0 405000.0 1083000.0 ;
      RECT  394800.0 1096800.0 405000.0 1110600.0 ;
      RECT  394800.0 1124400.0 405000.0 1110600.0 ;
      RECT  394800.0 1124400.0 405000.0 1138200.0 ;
      RECT  394800.0 1152000.0 405000.0 1138200.0 ;
      RECT  394800.0 1152000.0 405000.0 1165800.0 ;
      RECT  394800.0 1179600.0 405000.0 1165800.0 ;
      RECT  394800.0 1179600.0 405000.0 1193400.0 ;
      RECT  394800.0 1207200.0 405000.0 1193400.0 ;
      RECT  394800.0 1207200.0 405000.0 1221000.0 ;
      RECT  394800.0 1234800.0 405000.0 1221000.0 ;
      RECT  394800.0 1234800.0 405000.0 1248600.0 ;
      RECT  394800.0 1262400.0 405000.0 1248600.0 ;
      RECT  394800.0 1262400.0 405000.0 1276200.0 ;
      RECT  394800.0 1290000.0 405000.0 1276200.0 ;
      RECT  394800.0 1290000.0 405000.0 1303800.0 ;
      RECT  394800.0 1317600.0 405000.0 1303800.0 ;
      RECT  394800.0 1317600.0 405000.0 1331400.0 ;
      RECT  394800.0 1345200.0 405000.0 1331400.0 ;
      RECT  394800.0 1345200.0 405000.0 1359000.0 ;
      RECT  394800.0 1372800.0 405000.0 1359000.0 ;
      RECT  394800.0 1372800.0 405000.0 1386600.0 ;
      RECT  394800.0 1400400.0 405000.0 1386600.0 ;
      RECT  394800.0 1400400.0 405000.0 1414200.0 ;
      RECT  394800.0 1428000.0 405000.0 1414200.0 ;
      RECT  394800.0 1428000.0 405000.0 1441800.0 ;
      RECT  394800.0 1455600.0 405000.0 1441800.0 ;
      RECT  394800.0 1455600.0 405000.0 1469400.0 ;
      RECT  394800.0 1483200.0 405000.0 1469400.0 ;
      RECT  394800.0 1483200.0 405000.0 1497000.0 ;
      RECT  394800.0 1510800.0 405000.0 1497000.0 ;
      RECT  394800.0 1510800.0 405000.0 1524600.0 ;
      RECT  394800.0 1538400.0 405000.0 1524600.0 ;
      RECT  394800.0 1538400.0 405000.0 1552200.0 ;
      RECT  394800.0 1566000.0 405000.0 1552200.0 ;
      RECT  394800.0 1566000.0 405000.0 1579800.0 ;
      RECT  394800.0 1593600.0 405000.0 1579800.0 ;
      RECT  394800.0 1593600.0 405000.0 1607400.0 ;
      RECT  394800.0 1621200.0 405000.0 1607400.0 ;
      RECT  394800.0 1621200.0 405000.0 1635000.0 ;
      RECT  394800.0 1648800.0 405000.0 1635000.0 ;
      RECT  394800.0 1648800.0 405000.0 1662600.0 ;
      RECT  394800.0 1676400.0 405000.0 1662600.0 ;
      RECT  394800.0 1676400.0 405000.0 1690200.0 ;
      RECT  394800.0 1704000.0 405000.0 1690200.0 ;
      RECT  394800.0 1704000.0 405000.0 1717800.0 ;
      RECT  394800.0 1731600.0 405000.0 1717800.0 ;
      RECT  394800.0 1731600.0 405000.0 1745400.0 ;
      RECT  394800.0 1759200.0 405000.0 1745400.0 ;
      RECT  394800.0 1759200.0 405000.0 1773000.0 ;
      RECT  394800.0 1786800.0 405000.0 1773000.0 ;
      RECT  394800.0 1786800.0 405000.0 1800600.0 ;
      RECT  394800.0 1814400.0 405000.0 1800600.0 ;
      RECT  394800.0 1814400.0 405000.0 1828200.0 ;
      RECT  394800.0 1842000.0 405000.0 1828200.0 ;
      RECT  394800.0 1842000.0 405000.0 1855800.0 ;
      RECT  394800.0 1869600.0 405000.0 1855800.0 ;
      RECT  394800.0 1869600.0 405000.0 1883400.0 ;
      RECT  394800.0 1897200.0 405000.0 1883400.0 ;
      RECT  394800.0 1897200.0 405000.0 1911000.0 ;
      RECT  394800.0 1924800.0 405000.0 1911000.0 ;
      RECT  394800.0 1924800.0 405000.0 1938600.0 ;
      RECT  394800.0 1952400.0 405000.0 1938600.0 ;
      RECT  394800.0 1952400.0 405000.0 1966200.0 ;
      RECT  394800.0 1980000.0 405000.0 1966200.0 ;
      RECT  394800.0 1980000.0 405000.0 1993800.0 ;
      RECT  394800.0 2007600.0 405000.0 1993800.0 ;
      RECT  394800.0 2007600.0 405000.0 2021400.0 ;
      RECT  394800.0 2035200.0 405000.0 2021400.0 ;
      RECT  394800.0 2035200.0 405000.0 2049000.0 ;
      RECT  394800.0 2062800.0 405000.0 2049000.0 ;
      RECT  394800.0 2062800.0 405000.0 2076600.0 ;
      RECT  394800.0 2090400.0 405000.0 2076600.0 ;
      RECT  394800.0 2090400.0 405000.0 2104200.0 ;
      RECT  394800.0 2118000.0 405000.0 2104200.0 ;
      RECT  394800.0 2118000.0 405000.0 2131800.0 ;
      RECT  394800.0 2145600.0 405000.0 2131800.0 ;
      RECT  405000.0 379200.0 415200.0 393000.0 ;
      RECT  405000.0 406800.0 415200.0 393000.0 ;
      RECT  405000.0 406800.0 415200.0 420600.0 ;
      RECT  405000.0 434400.0 415200.0 420600.0 ;
      RECT  405000.0 434400.0 415200.0 448200.0 ;
      RECT  405000.0 462000.0 415200.0 448200.0 ;
      RECT  405000.0 462000.0 415200.0 475800.0 ;
      RECT  405000.0 489600.0 415200.0 475800.0 ;
      RECT  405000.0 489600.0 415200.0 503400.0 ;
      RECT  405000.0 517200.0 415200.0 503400.0 ;
      RECT  405000.0 517200.0 415200.0 531000.0 ;
      RECT  405000.0 544800.0 415200.0 531000.0 ;
      RECT  405000.0 544800.0 415200.0 558600.0 ;
      RECT  405000.0 572400.0 415200.0 558600.0 ;
      RECT  405000.0 572400.0 415200.0 586200.0 ;
      RECT  405000.0 600000.0 415200.0 586200.0 ;
      RECT  405000.0 600000.0 415200.0 613800.0 ;
      RECT  405000.0 627600.0 415200.0 613800.0 ;
      RECT  405000.0 627600.0 415200.0 641400.0 ;
      RECT  405000.0 655200.0 415200.0 641400.0 ;
      RECT  405000.0 655200.0 415200.0 669000.0 ;
      RECT  405000.0 682800.0 415200.0 669000.0 ;
      RECT  405000.0 682800.0 415200.0 696600.0 ;
      RECT  405000.0 710400.0 415200.0 696600.0 ;
      RECT  405000.0 710400.0 415200.0 724200.0 ;
      RECT  405000.0 738000.0 415200.0 724200.0 ;
      RECT  405000.0 738000.0 415200.0 751800.0 ;
      RECT  405000.0 765600.0 415200.0 751800.0 ;
      RECT  405000.0 765600.0 415200.0 779400.0 ;
      RECT  405000.0 793200.0 415200.0 779400.0 ;
      RECT  405000.0 793200.0 415200.0 807000.0 ;
      RECT  405000.0 820800.0 415200.0 807000.0 ;
      RECT  405000.0 820800.0 415200.0 834600.0 ;
      RECT  405000.0 848400.0 415200.0 834600.0 ;
      RECT  405000.0 848400.0 415200.0 862200.0 ;
      RECT  405000.0 876000.0 415200.0 862200.0 ;
      RECT  405000.0 876000.0 415200.0 889800.0 ;
      RECT  405000.0 903600.0 415200.0 889800.0 ;
      RECT  405000.0 903600.0 415200.0 917400.0 ;
      RECT  405000.0 931200.0 415200.0 917400.0 ;
      RECT  405000.0 931200.0 415200.0 945000.0 ;
      RECT  405000.0 958800.0 415200.0 945000.0 ;
      RECT  405000.0 958800.0 415200.0 972600.0 ;
      RECT  405000.0 986400.0 415200.0 972600.0 ;
      RECT  405000.0 986400.0 415200.0 1000200.0 ;
      RECT  405000.0 1014000.0 415200.0 1000200.0 ;
      RECT  405000.0 1014000.0 415200.0 1027800.0 ;
      RECT  405000.0 1041600.0 415200.0 1027800.0 ;
      RECT  405000.0 1041600.0 415200.0 1055400.0 ;
      RECT  405000.0 1069200.0 415200.0 1055400.0 ;
      RECT  405000.0 1069200.0 415200.0 1083000.0 ;
      RECT  405000.0 1096800.0 415200.0 1083000.0 ;
      RECT  405000.0 1096800.0 415200.0 1110600.0 ;
      RECT  405000.0 1124400.0 415200.0 1110600.0 ;
      RECT  405000.0 1124400.0 415200.0 1138200.0 ;
      RECT  405000.0 1152000.0 415200.0 1138200.0 ;
      RECT  405000.0 1152000.0 415200.0 1165800.0 ;
      RECT  405000.0 1179600.0 415200.0 1165800.0 ;
      RECT  405000.0 1179600.0 415200.0 1193400.0 ;
      RECT  405000.0 1207200.0 415200.0 1193400.0 ;
      RECT  405000.0 1207200.0 415200.0 1221000.0 ;
      RECT  405000.0 1234800.0 415200.0 1221000.0 ;
      RECT  405000.0 1234800.0 415200.0 1248600.0 ;
      RECT  405000.0 1262400.0 415200.0 1248600.0 ;
      RECT  405000.0 1262400.0 415200.0 1276200.0 ;
      RECT  405000.0 1290000.0 415200.0 1276200.0 ;
      RECT  405000.0 1290000.0 415200.0 1303800.0 ;
      RECT  405000.0 1317600.0 415200.0 1303800.0 ;
      RECT  405000.0 1317600.0 415200.0 1331400.0 ;
      RECT  405000.0 1345200.0 415200.0 1331400.0 ;
      RECT  405000.0 1345200.0 415200.0 1359000.0 ;
      RECT  405000.0 1372800.0 415200.0 1359000.0 ;
      RECT  405000.0 1372800.0 415200.0 1386600.0 ;
      RECT  405000.0 1400400.0 415200.0 1386600.0 ;
      RECT  405000.0 1400400.0 415200.0 1414200.0 ;
      RECT  405000.0 1428000.0 415200.0 1414200.0 ;
      RECT  405000.0 1428000.0 415200.0 1441800.0 ;
      RECT  405000.0 1455600.0 415200.0 1441800.0 ;
      RECT  405000.0 1455600.0 415200.0 1469400.0 ;
      RECT  405000.0 1483200.0 415200.0 1469400.0 ;
      RECT  405000.0 1483200.0 415200.0 1497000.0 ;
      RECT  405000.0 1510800.0 415200.0 1497000.0 ;
      RECT  405000.0 1510800.0 415200.0 1524600.0 ;
      RECT  405000.0 1538400.0 415200.0 1524600.0 ;
      RECT  405000.0 1538400.0 415200.0 1552200.0 ;
      RECT  405000.0 1566000.0 415200.0 1552200.0 ;
      RECT  405000.0 1566000.0 415200.0 1579800.0 ;
      RECT  405000.0 1593600.0 415200.0 1579800.0 ;
      RECT  405000.0 1593600.0 415200.0 1607400.0 ;
      RECT  405000.0 1621200.0 415200.0 1607400.0 ;
      RECT  405000.0 1621200.0 415200.0 1635000.0 ;
      RECT  405000.0 1648800.0 415200.0 1635000.0 ;
      RECT  405000.0 1648800.0 415200.0 1662600.0 ;
      RECT  405000.0 1676400.0 415200.0 1662600.0 ;
      RECT  405000.0 1676400.0 415200.0 1690200.0 ;
      RECT  405000.0 1704000.0 415200.0 1690200.0 ;
      RECT  405000.0 1704000.0 415200.0 1717800.0 ;
      RECT  405000.0 1731600.0 415200.0 1717800.0 ;
      RECT  405000.0 1731600.0 415200.0 1745400.0 ;
      RECT  405000.0 1759200.0 415200.0 1745400.0 ;
      RECT  405000.0 1759200.0 415200.0 1773000.0 ;
      RECT  405000.0 1786800.0 415200.0 1773000.0 ;
      RECT  405000.0 1786800.0 415200.0 1800600.0 ;
      RECT  405000.0 1814400.0 415200.0 1800600.0 ;
      RECT  405000.0 1814400.0 415200.0 1828200.0 ;
      RECT  405000.0 1842000.0 415200.0 1828200.0 ;
      RECT  405000.0 1842000.0 415200.0 1855800.0 ;
      RECT  405000.0 1869600.0 415200.0 1855800.0 ;
      RECT  405000.0 1869600.0 415200.0 1883400.0 ;
      RECT  405000.0 1897200.0 415200.0 1883400.0 ;
      RECT  405000.0 1897200.0 415200.0 1911000.0 ;
      RECT  405000.0 1924800.0 415200.0 1911000.0 ;
      RECT  405000.0 1924800.0 415200.0 1938600.0 ;
      RECT  405000.0 1952400.0 415200.0 1938600.0 ;
      RECT  405000.0 1952400.0 415200.0 1966200.0 ;
      RECT  405000.0 1980000.0 415200.0 1966200.0 ;
      RECT  405000.0 1980000.0 415200.0 1993800.0 ;
      RECT  405000.0 2007600.0 415200.0 1993800.0 ;
      RECT  405000.0 2007600.0 415200.0 2021400.0 ;
      RECT  405000.0 2035200.0 415200.0 2021400.0 ;
      RECT  405000.0 2035200.0 415200.0 2049000.0 ;
      RECT  405000.0 2062800.0 415200.0 2049000.0 ;
      RECT  405000.0 2062800.0 415200.0 2076600.0 ;
      RECT  405000.0 2090400.0 415200.0 2076600.0 ;
      RECT  405000.0 2090400.0 415200.0 2104200.0 ;
      RECT  405000.0 2118000.0 415200.0 2104200.0 ;
      RECT  405000.0 2118000.0 415200.0 2131800.0 ;
      RECT  405000.0 2145600.0 415200.0 2131800.0 ;
      RECT  415200.0 379200.0 425400.0 393000.0 ;
      RECT  415200.0 406800.0 425400.0 393000.0 ;
      RECT  415200.0 406800.0 425400.0 420600.0 ;
      RECT  415200.0 434400.0 425400.0 420600.0 ;
      RECT  415200.0 434400.0 425400.0 448200.0 ;
      RECT  415200.0 462000.0 425400.0 448200.0 ;
      RECT  415200.0 462000.0 425400.0 475800.0 ;
      RECT  415200.0 489600.0 425400.0 475800.0 ;
      RECT  415200.0 489600.0 425400.0 503400.0 ;
      RECT  415200.0 517200.0 425400.0 503400.0 ;
      RECT  415200.0 517200.0 425400.0 531000.0 ;
      RECT  415200.0 544800.0 425400.0 531000.0 ;
      RECT  415200.0 544800.0 425400.0 558600.0 ;
      RECT  415200.0 572400.0 425400.0 558600.0 ;
      RECT  415200.0 572400.0 425400.0 586200.0 ;
      RECT  415200.0 600000.0 425400.0 586200.0 ;
      RECT  415200.0 600000.0 425400.0 613800.0 ;
      RECT  415200.0 627600.0 425400.0 613800.0 ;
      RECT  415200.0 627600.0 425400.0 641400.0 ;
      RECT  415200.0 655200.0 425400.0 641400.0 ;
      RECT  415200.0 655200.0 425400.0 669000.0 ;
      RECT  415200.0 682800.0 425400.0 669000.0 ;
      RECT  415200.0 682800.0 425400.0 696600.0 ;
      RECT  415200.0 710400.0 425400.0 696600.0 ;
      RECT  415200.0 710400.0 425400.0 724200.0 ;
      RECT  415200.0 738000.0 425400.0 724200.0 ;
      RECT  415200.0 738000.0 425400.0 751800.0 ;
      RECT  415200.0 765600.0 425400.0 751800.0 ;
      RECT  415200.0 765600.0 425400.0 779400.0 ;
      RECT  415200.0 793200.0 425400.0 779400.0 ;
      RECT  415200.0 793200.0 425400.0 807000.0 ;
      RECT  415200.0 820800.0 425400.0 807000.0 ;
      RECT  415200.0 820800.0 425400.0 834600.0 ;
      RECT  415200.0 848400.0 425400.0 834600.0 ;
      RECT  415200.0 848400.0 425400.0 862200.0 ;
      RECT  415200.0 876000.0 425400.0 862200.0 ;
      RECT  415200.0 876000.0 425400.0 889800.0 ;
      RECT  415200.0 903600.0 425400.0 889800.0 ;
      RECT  415200.0 903600.0 425400.0 917400.0 ;
      RECT  415200.0 931200.0 425400.0 917400.0 ;
      RECT  415200.0 931200.0 425400.0 945000.0 ;
      RECT  415200.0 958800.0 425400.0 945000.0 ;
      RECT  415200.0 958800.0 425400.0 972600.0 ;
      RECT  415200.0 986400.0 425400.0 972600.0 ;
      RECT  415200.0 986400.0 425400.0 1000200.0 ;
      RECT  415200.0 1014000.0 425400.0 1000200.0 ;
      RECT  415200.0 1014000.0 425400.0 1027800.0 ;
      RECT  415200.0 1041600.0 425400.0 1027800.0 ;
      RECT  415200.0 1041600.0 425400.0 1055400.0 ;
      RECT  415200.0 1069200.0 425400.0 1055400.0 ;
      RECT  415200.0 1069200.0 425400.0 1083000.0 ;
      RECT  415200.0 1096800.0 425400.0 1083000.0 ;
      RECT  415200.0 1096800.0 425400.0 1110600.0 ;
      RECT  415200.0 1124400.0 425400.0 1110600.0 ;
      RECT  415200.0 1124400.0 425400.0 1138200.0 ;
      RECT  415200.0 1152000.0 425400.0 1138200.0 ;
      RECT  415200.0 1152000.0 425400.0 1165800.0 ;
      RECT  415200.0 1179600.0 425400.0 1165800.0 ;
      RECT  415200.0 1179600.0 425400.0 1193400.0 ;
      RECT  415200.0 1207200.0 425400.0 1193400.0 ;
      RECT  415200.0 1207200.0 425400.0 1221000.0 ;
      RECT  415200.0 1234800.0 425400.0 1221000.0 ;
      RECT  415200.0 1234800.0 425400.0 1248600.0 ;
      RECT  415200.0 1262400.0 425400.0 1248600.0 ;
      RECT  415200.0 1262400.0 425400.0 1276200.0 ;
      RECT  415200.0 1290000.0 425400.0 1276200.0 ;
      RECT  415200.0 1290000.0 425400.0 1303800.0 ;
      RECT  415200.0 1317600.0 425400.0 1303800.0 ;
      RECT  415200.0 1317600.0 425400.0 1331400.0 ;
      RECT  415200.0 1345200.0 425400.0 1331400.0 ;
      RECT  415200.0 1345200.0 425400.0 1359000.0 ;
      RECT  415200.0 1372800.0 425400.0 1359000.0 ;
      RECT  415200.0 1372800.0 425400.0 1386600.0 ;
      RECT  415200.0 1400400.0 425400.0 1386600.0 ;
      RECT  415200.0 1400400.0 425400.0 1414200.0 ;
      RECT  415200.0 1428000.0 425400.0 1414200.0 ;
      RECT  415200.0 1428000.0 425400.0 1441800.0 ;
      RECT  415200.0 1455600.0 425400.0 1441800.0 ;
      RECT  415200.0 1455600.0 425400.0 1469400.0 ;
      RECT  415200.0 1483200.0 425400.0 1469400.0 ;
      RECT  415200.0 1483200.0 425400.0 1497000.0 ;
      RECT  415200.0 1510800.0 425400.0 1497000.0 ;
      RECT  415200.0 1510800.0 425400.0 1524600.0 ;
      RECT  415200.0 1538400.0 425400.0 1524600.0 ;
      RECT  415200.0 1538400.0 425400.0 1552200.0 ;
      RECT  415200.0 1566000.0 425400.0 1552200.0 ;
      RECT  415200.0 1566000.0 425400.0 1579800.0 ;
      RECT  415200.0 1593600.0 425400.0 1579800.0 ;
      RECT  415200.0 1593600.0 425400.0 1607400.0 ;
      RECT  415200.0 1621200.0 425400.0 1607400.0 ;
      RECT  415200.0 1621200.0 425400.0 1635000.0 ;
      RECT  415200.0 1648800.0 425400.0 1635000.0 ;
      RECT  415200.0 1648800.0 425400.0 1662600.0 ;
      RECT  415200.0 1676400.0 425400.0 1662600.0 ;
      RECT  415200.0 1676400.0 425400.0 1690200.0 ;
      RECT  415200.0 1704000.0 425400.0 1690200.0 ;
      RECT  415200.0 1704000.0 425400.0 1717800.0 ;
      RECT  415200.0 1731600.0 425400.0 1717800.0 ;
      RECT  415200.0 1731600.0 425400.0 1745400.0 ;
      RECT  415200.0 1759200.0 425400.0 1745400.0 ;
      RECT  415200.0 1759200.0 425400.0 1773000.0 ;
      RECT  415200.0 1786800.0 425400.0 1773000.0 ;
      RECT  415200.0 1786800.0 425400.0 1800600.0 ;
      RECT  415200.0 1814400.0 425400.0 1800600.0 ;
      RECT  415200.0 1814400.0 425400.0 1828200.0 ;
      RECT  415200.0 1842000.0 425400.0 1828200.0 ;
      RECT  415200.0 1842000.0 425400.0 1855800.0 ;
      RECT  415200.0 1869600.0 425400.0 1855800.0 ;
      RECT  415200.0 1869600.0 425400.0 1883400.0 ;
      RECT  415200.0 1897200.0 425400.0 1883400.0 ;
      RECT  415200.0 1897200.0 425400.0 1911000.0 ;
      RECT  415200.0 1924800.0 425400.0 1911000.0 ;
      RECT  415200.0 1924800.0 425400.0 1938600.0 ;
      RECT  415200.0 1952400.0 425400.0 1938600.0 ;
      RECT  415200.0 1952400.0 425400.0 1966200.0 ;
      RECT  415200.0 1980000.0 425400.0 1966200.0 ;
      RECT  415200.0 1980000.0 425400.0 1993800.0 ;
      RECT  415200.0 2007600.0 425400.0 1993800.0 ;
      RECT  415200.0 2007600.0 425400.0 2021400.0 ;
      RECT  415200.0 2035200.0 425400.0 2021400.0 ;
      RECT  415200.0 2035200.0 425400.0 2049000.0 ;
      RECT  415200.0 2062800.0 425400.0 2049000.0 ;
      RECT  415200.0 2062800.0 425400.0 2076600.0 ;
      RECT  415200.0 2090400.0 425400.0 2076600.0 ;
      RECT  415200.0 2090400.0 425400.0 2104200.0 ;
      RECT  415200.0 2118000.0 425400.0 2104200.0 ;
      RECT  415200.0 2118000.0 425400.0 2131800.0 ;
      RECT  415200.0 2145600.0 425400.0 2131800.0 ;
      RECT  425400.0 379200.0 435600.0 393000.0 ;
      RECT  425400.0 406800.0 435600.0 393000.0 ;
      RECT  425400.0 406800.0 435600.0 420600.0 ;
      RECT  425400.0 434400.0 435600.0 420600.0 ;
      RECT  425400.0 434400.0 435600.0 448200.0 ;
      RECT  425400.0 462000.0 435600.0 448200.0 ;
      RECT  425400.0 462000.0 435600.0 475800.0 ;
      RECT  425400.0 489600.0 435600.0 475800.0 ;
      RECT  425400.0 489600.0 435600.0 503400.0 ;
      RECT  425400.0 517200.0 435600.0 503400.0 ;
      RECT  425400.0 517200.0 435600.0 531000.0 ;
      RECT  425400.0 544800.0 435600.0 531000.0 ;
      RECT  425400.0 544800.0 435600.0 558600.0 ;
      RECT  425400.0 572400.0 435600.0 558600.0 ;
      RECT  425400.0 572400.0 435600.0 586200.0 ;
      RECT  425400.0 600000.0 435600.0 586200.0 ;
      RECT  425400.0 600000.0 435600.0 613800.0 ;
      RECT  425400.0 627600.0 435600.0 613800.0 ;
      RECT  425400.0 627600.0 435600.0 641400.0 ;
      RECT  425400.0 655200.0 435600.0 641400.0 ;
      RECT  425400.0 655200.0 435600.0 669000.0 ;
      RECT  425400.0 682800.0 435600.0 669000.0 ;
      RECT  425400.0 682800.0 435600.0 696600.0 ;
      RECT  425400.0 710400.0 435600.0 696600.0 ;
      RECT  425400.0 710400.0 435600.0 724200.0 ;
      RECT  425400.0 738000.0 435600.0 724200.0 ;
      RECT  425400.0 738000.0 435600.0 751800.0 ;
      RECT  425400.0 765600.0 435600.0 751800.0 ;
      RECT  425400.0 765600.0 435600.0 779400.0 ;
      RECT  425400.0 793200.0 435600.0 779400.0 ;
      RECT  425400.0 793200.0 435600.0 807000.0 ;
      RECT  425400.0 820800.0 435600.0 807000.0 ;
      RECT  425400.0 820800.0 435600.0 834600.0 ;
      RECT  425400.0 848400.0 435600.0 834600.0 ;
      RECT  425400.0 848400.0 435600.0 862200.0 ;
      RECT  425400.0 876000.0 435600.0 862200.0 ;
      RECT  425400.0 876000.0 435600.0 889800.0 ;
      RECT  425400.0 903600.0 435600.0 889800.0 ;
      RECT  425400.0 903600.0 435600.0 917400.0 ;
      RECT  425400.0 931200.0 435600.0 917400.0 ;
      RECT  425400.0 931200.0 435600.0 945000.0 ;
      RECT  425400.0 958800.0 435600.0 945000.0 ;
      RECT  425400.0 958800.0 435600.0 972600.0 ;
      RECT  425400.0 986400.0 435600.0 972600.0 ;
      RECT  425400.0 986400.0 435600.0 1000200.0 ;
      RECT  425400.0 1014000.0 435600.0 1000200.0 ;
      RECT  425400.0 1014000.0 435600.0 1027800.0 ;
      RECT  425400.0 1041600.0 435600.0 1027800.0 ;
      RECT  425400.0 1041600.0 435600.0 1055400.0 ;
      RECT  425400.0 1069200.0 435600.0 1055400.0 ;
      RECT  425400.0 1069200.0 435600.0 1083000.0 ;
      RECT  425400.0 1096800.0 435600.0 1083000.0 ;
      RECT  425400.0 1096800.0 435600.0 1110600.0 ;
      RECT  425400.0 1124400.0 435600.0 1110600.0 ;
      RECT  425400.0 1124400.0 435600.0 1138200.0 ;
      RECT  425400.0 1152000.0 435600.0 1138200.0 ;
      RECT  425400.0 1152000.0 435600.0 1165800.0 ;
      RECT  425400.0 1179600.0 435600.0 1165800.0 ;
      RECT  425400.0 1179600.0 435600.0 1193400.0 ;
      RECT  425400.0 1207200.0 435600.0 1193400.0 ;
      RECT  425400.0 1207200.0 435600.0 1221000.0 ;
      RECT  425400.0 1234800.0 435600.0 1221000.0 ;
      RECT  425400.0 1234800.0 435600.0 1248600.0 ;
      RECT  425400.0 1262400.0 435600.0 1248600.0 ;
      RECT  425400.0 1262400.0 435600.0 1276200.0 ;
      RECT  425400.0 1290000.0 435600.0 1276200.0 ;
      RECT  425400.0 1290000.0 435600.0 1303800.0 ;
      RECT  425400.0 1317600.0 435600.0 1303800.0 ;
      RECT  425400.0 1317600.0 435600.0 1331400.0 ;
      RECT  425400.0 1345200.0 435600.0 1331400.0 ;
      RECT  425400.0 1345200.0 435600.0 1359000.0 ;
      RECT  425400.0 1372800.0 435600.0 1359000.0 ;
      RECT  425400.0 1372800.0 435600.0 1386600.0 ;
      RECT  425400.0 1400400.0 435600.0 1386600.0 ;
      RECT  425400.0 1400400.0 435600.0 1414200.0 ;
      RECT  425400.0 1428000.0 435600.0 1414200.0 ;
      RECT  425400.0 1428000.0 435600.0 1441800.0 ;
      RECT  425400.0 1455600.0 435600.0 1441800.0 ;
      RECT  425400.0 1455600.0 435600.0 1469400.0 ;
      RECT  425400.0 1483200.0 435600.0 1469400.0 ;
      RECT  425400.0 1483200.0 435600.0 1497000.0 ;
      RECT  425400.0 1510800.0 435600.0 1497000.0 ;
      RECT  425400.0 1510800.0 435600.0 1524600.0 ;
      RECT  425400.0 1538400.0 435600.0 1524600.0 ;
      RECT  425400.0 1538400.0 435600.0 1552200.0 ;
      RECT  425400.0 1566000.0 435600.0 1552200.0 ;
      RECT  425400.0 1566000.0 435600.0 1579800.0 ;
      RECT  425400.0 1593600.0 435600.0 1579800.0 ;
      RECT  425400.0 1593600.0 435600.0 1607400.0 ;
      RECT  425400.0 1621200.0 435600.0 1607400.0 ;
      RECT  425400.0 1621200.0 435600.0 1635000.0 ;
      RECT  425400.0 1648800.0 435600.0 1635000.0 ;
      RECT  425400.0 1648800.0 435600.0 1662600.0 ;
      RECT  425400.0 1676400.0 435600.0 1662600.0 ;
      RECT  425400.0 1676400.0 435600.0 1690200.0 ;
      RECT  425400.0 1704000.0 435600.0 1690200.0 ;
      RECT  425400.0 1704000.0 435600.0 1717800.0 ;
      RECT  425400.0 1731600.0 435600.0 1717800.0 ;
      RECT  425400.0 1731600.0 435600.0 1745400.0 ;
      RECT  425400.0 1759200.0 435600.0 1745400.0 ;
      RECT  425400.0 1759200.0 435600.0 1773000.0 ;
      RECT  425400.0 1786800.0 435600.0 1773000.0 ;
      RECT  425400.0 1786800.0 435600.0 1800600.0 ;
      RECT  425400.0 1814400.0 435600.0 1800600.0 ;
      RECT  425400.0 1814400.0 435600.0 1828200.0 ;
      RECT  425400.0 1842000.0 435600.0 1828200.0 ;
      RECT  425400.0 1842000.0 435600.0 1855800.0 ;
      RECT  425400.0 1869600.0 435600.0 1855800.0 ;
      RECT  425400.0 1869600.0 435600.0 1883400.0 ;
      RECT  425400.0 1897200.0 435600.0 1883400.0 ;
      RECT  425400.0 1897200.0 435600.0 1911000.0 ;
      RECT  425400.0 1924800.0 435600.0 1911000.0 ;
      RECT  425400.0 1924800.0 435600.0 1938600.0 ;
      RECT  425400.0 1952400.0 435600.0 1938600.0 ;
      RECT  425400.0 1952400.0 435600.0 1966200.0 ;
      RECT  425400.0 1980000.0 435600.0 1966200.0 ;
      RECT  425400.0 1980000.0 435600.0 1993800.0 ;
      RECT  425400.0 2007600.0 435600.0 1993800.0 ;
      RECT  425400.0 2007600.0 435600.0 2021400.0 ;
      RECT  425400.0 2035200.0 435600.0 2021400.0 ;
      RECT  425400.0 2035200.0 435600.0 2049000.0 ;
      RECT  425400.0 2062800.0 435600.0 2049000.0 ;
      RECT  425400.0 2062800.0 435600.0 2076600.0 ;
      RECT  425400.0 2090400.0 435600.0 2076600.0 ;
      RECT  425400.0 2090400.0 435600.0 2104200.0 ;
      RECT  425400.0 2118000.0 435600.0 2104200.0 ;
      RECT  425400.0 2118000.0 435600.0 2131800.0 ;
      RECT  425400.0 2145600.0 435600.0 2131800.0 ;
      RECT  435600.0 379200.0 445800.0 393000.0 ;
      RECT  435600.0 406800.0 445800.0 393000.0 ;
      RECT  435600.0 406800.0 445800.0 420600.0 ;
      RECT  435600.0 434400.0 445800.0 420600.0 ;
      RECT  435600.0 434400.0 445800.0 448200.0 ;
      RECT  435600.0 462000.0 445800.0 448200.0 ;
      RECT  435600.0 462000.0 445800.0 475800.0 ;
      RECT  435600.0 489600.0 445800.0 475800.0 ;
      RECT  435600.0 489600.0 445800.0 503400.0 ;
      RECT  435600.0 517200.0 445800.0 503400.0 ;
      RECT  435600.0 517200.0 445800.0 531000.0 ;
      RECT  435600.0 544800.0 445800.0 531000.0 ;
      RECT  435600.0 544800.0 445800.0 558600.0 ;
      RECT  435600.0 572400.0 445800.0 558600.0 ;
      RECT  435600.0 572400.0 445800.0 586200.0 ;
      RECT  435600.0 600000.0 445800.0 586200.0 ;
      RECT  435600.0 600000.0 445800.0 613800.0 ;
      RECT  435600.0 627600.0 445800.0 613800.0 ;
      RECT  435600.0 627600.0 445800.0 641400.0 ;
      RECT  435600.0 655200.0 445800.0 641400.0 ;
      RECT  435600.0 655200.0 445800.0 669000.0 ;
      RECT  435600.0 682800.0 445800.0 669000.0 ;
      RECT  435600.0 682800.0 445800.0 696600.0 ;
      RECT  435600.0 710400.0 445800.0 696600.0 ;
      RECT  435600.0 710400.0 445800.0 724200.0 ;
      RECT  435600.0 738000.0 445800.0 724200.0 ;
      RECT  435600.0 738000.0 445800.0 751800.0 ;
      RECT  435600.0 765600.0 445800.0 751800.0 ;
      RECT  435600.0 765600.0 445800.0 779400.0 ;
      RECT  435600.0 793200.0 445800.0 779400.0 ;
      RECT  435600.0 793200.0 445800.0 807000.0 ;
      RECT  435600.0 820800.0 445800.0 807000.0 ;
      RECT  435600.0 820800.0 445800.0 834600.0 ;
      RECT  435600.0 848400.0 445800.0 834600.0 ;
      RECT  435600.0 848400.0 445800.0 862200.0 ;
      RECT  435600.0 876000.0 445800.0 862200.0 ;
      RECT  435600.0 876000.0 445800.0 889800.0 ;
      RECT  435600.0 903600.0 445800.0 889800.0 ;
      RECT  435600.0 903600.0 445800.0 917400.0 ;
      RECT  435600.0 931200.0 445800.0 917400.0 ;
      RECT  435600.0 931200.0 445800.0 945000.0 ;
      RECT  435600.0 958800.0 445800.0 945000.0 ;
      RECT  435600.0 958800.0 445800.0 972600.0 ;
      RECT  435600.0 986400.0 445800.0 972600.0 ;
      RECT  435600.0 986400.0 445800.0 1000200.0 ;
      RECT  435600.0 1014000.0 445800.0 1000200.0 ;
      RECT  435600.0 1014000.0 445800.0 1027800.0 ;
      RECT  435600.0 1041600.0 445800.0 1027800.0 ;
      RECT  435600.0 1041600.0 445800.0 1055400.0 ;
      RECT  435600.0 1069200.0 445800.0 1055400.0 ;
      RECT  435600.0 1069200.0 445800.0 1083000.0 ;
      RECT  435600.0 1096800.0 445800.0 1083000.0 ;
      RECT  435600.0 1096800.0 445800.0 1110600.0 ;
      RECT  435600.0 1124400.0 445800.0 1110600.0 ;
      RECT  435600.0 1124400.0 445800.0 1138200.0 ;
      RECT  435600.0 1152000.0 445800.0 1138200.0 ;
      RECT  435600.0 1152000.0 445800.0 1165800.0 ;
      RECT  435600.0 1179600.0 445800.0 1165800.0 ;
      RECT  435600.0 1179600.0 445800.0 1193400.0 ;
      RECT  435600.0 1207200.0 445800.0 1193400.0 ;
      RECT  435600.0 1207200.0 445800.0 1221000.0 ;
      RECT  435600.0 1234800.0 445800.0 1221000.0 ;
      RECT  435600.0 1234800.0 445800.0 1248600.0 ;
      RECT  435600.0 1262400.0 445800.0 1248600.0 ;
      RECT  435600.0 1262400.0 445800.0 1276200.0 ;
      RECT  435600.0 1290000.0 445800.0 1276200.0 ;
      RECT  435600.0 1290000.0 445800.0 1303800.0 ;
      RECT  435600.0 1317600.0 445800.0 1303800.0 ;
      RECT  435600.0 1317600.0 445800.0 1331400.0 ;
      RECT  435600.0 1345200.0 445800.0 1331400.0 ;
      RECT  435600.0 1345200.0 445800.0 1359000.0 ;
      RECT  435600.0 1372800.0 445800.0 1359000.0 ;
      RECT  435600.0 1372800.0 445800.0 1386600.0 ;
      RECT  435600.0 1400400.0 445800.0 1386600.0 ;
      RECT  435600.0 1400400.0 445800.0 1414200.0 ;
      RECT  435600.0 1428000.0 445800.0 1414200.0 ;
      RECT  435600.0 1428000.0 445800.0 1441800.0 ;
      RECT  435600.0 1455600.0 445800.0 1441800.0 ;
      RECT  435600.0 1455600.0 445800.0 1469400.0 ;
      RECT  435600.0 1483200.0 445800.0 1469400.0 ;
      RECT  435600.0 1483200.0 445800.0 1497000.0 ;
      RECT  435600.0 1510800.0 445800.0 1497000.0 ;
      RECT  435600.0 1510800.0 445800.0 1524600.0 ;
      RECT  435600.0 1538400.0 445800.0 1524600.0 ;
      RECT  435600.0 1538400.0 445800.0 1552200.0 ;
      RECT  435600.0 1566000.0 445800.0 1552200.0 ;
      RECT  435600.0 1566000.0 445800.0 1579800.0 ;
      RECT  435600.0 1593600.0 445800.0 1579800.0 ;
      RECT  435600.0 1593600.0 445800.0 1607400.0 ;
      RECT  435600.0 1621200.0 445800.0 1607400.0 ;
      RECT  435600.0 1621200.0 445800.0 1635000.0 ;
      RECT  435600.0 1648800.0 445800.0 1635000.0 ;
      RECT  435600.0 1648800.0 445800.0 1662600.0 ;
      RECT  435600.0 1676400.0 445800.0 1662600.0 ;
      RECT  435600.0 1676400.0 445800.0 1690200.0 ;
      RECT  435600.0 1704000.0 445800.0 1690200.0 ;
      RECT  435600.0 1704000.0 445800.0 1717800.0 ;
      RECT  435600.0 1731600.0 445800.0 1717800.0 ;
      RECT  435600.0 1731600.0 445800.0 1745400.0 ;
      RECT  435600.0 1759200.0 445800.0 1745400.0 ;
      RECT  435600.0 1759200.0 445800.0 1773000.0 ;
      RECT  435600.0 1786800.0 445800.0 1773000.0 ;
      RECT  435600.0 1786800.0 445800.0 1800600.0 ;
      RECT  435600.0 1814400.0 445800.0 1800600.0 ;
      RECT  435600.0 1814400.0 445800.0 1828200.0 ;
      RECT  435600.0 1842000.0 445800.0 1828200.0 ;
      RECT  435600.0 1842000.0 445800.0 1855800.0 ;
      RECT  435600.0 1869600.0 445800.0 1855800.0 ;
      RECT  435600.0 1869600.0 445800.0 1883400.0 ;
      RECT  435600.0 1897200.0 445800.0 1883400.0 ;
      RECT  435600.0 1897200.0 445800.0 1911000.0 ;
      RECT  435600.0 1924800.0 445800.0 1911000.0 ;
      RECT  435600.0 1924800.0 445800.0 1938600.0 ;
      RECT  435600.0 1952400.0 445800.0 1938600.0 ;
      RECT  435600.0 1952400.0 445800.0 1966200.0 ;
      RECT  435600.0 1980000.0 445800.0 1966200.0 ;
      RECT  435600.0 1980000.0 445800.0 1993800.0 ;
      RECT  435600.0 2007600.0 445800.0 1993800.0 ;
      RECT  435600.0 2007600.0 445800.0 2021400.0 ;
      RECT  435600.0 2035200.0 445800.0 2021400.0 ;
      RECT  435600.0 2035200.0 445800.0 2049000.0 ;
      RECT  435600.0 2062800.0 445800.0 2049000.0 ;
      RECT  435600.0 2062800.0 445800.0 2076600.0 ;
      RECT  435600.0 2090400.0 445800.0 2076600.0 ;
      RECT  435600.0 2090400.0 445800.0 2104200.0 ;
      RECT  435600.0 2118000.0 445800.0 2104200.0 ;
      RECT  435600.0 2118000.0 445800.0 2131800.0 ;
      RECT  435600.0 2145600.0 445800.0 2131800.0 ;
      RECT  445800.0 379200.0 456000.0 393000.0 ;
      RECT  445800.0 406800.0 456000.0 393000.0 ;
      RECT  445800.0 406800.0 456000.0 420600.0 ;
      RECT  445800.0 434400.0 456000.0 420600.0 ;
      RECT  445800.0 434400.0 456000.0 448200.0 ;
      RECT  445800.0 462000.0 456000.0 448200.0 ;
      RECT  445800.0 462000.0 456000.0 475800.0 ;
      RECT  445800.0 489600.0 456000.0 475800.0 ;
      RECT  445800.0 489600.0 456000.0 503400.0 ;
      RECT  445800.0 517200.0 456000.0 503400.0 ;
      RECT  445800.0 517200.0 456000.0 531000.0 ;
      RECT  445800.0 544800.0 456000.0 531000.0 ;
      RECT  445800.0 544800.0 456000.0 558600.0 ;
      RECT  445800.0 572400.0 456000.0 558600.0 ;
      RECT  445800.0 572400.0 456000.0 586200.0 ;
      RECT  445800.0 600000.0 456000.0 586200.0 ;
      RECT  445800.0 600000.0 456000.0 613800.0 ;
      RECT  445800.0 627600.0 456000.0 613800.0 ;
      RECT  445800.0 627600.0 456000.0 641400.0 ;
      RECT  445800.0 655200.0 456000.0 641400.0 ;
      RECT  445800.0 655200.0 456000.0 669000.0 ;
      RECT  445800.0 682800.0 456000.0 669000.0 ;
      RECT  445800.0 682800.0 456000.0 696600.0 ;
      RECT  445800.0 710400.0 456000.0 696600.0 ;
      RECT  445800.0 710400.0 456000.0 724200.0 ;
      RECT  445800.0 738000.0 456000.0 724200.0 ;
      RECT  445800.0 738000.0 456000.0 751800.0 ;
      RECT  445800.0 765600.0 456000.0 751800.0 ;
      RECT  445800.0 765600.0 456000.0 779400.0 ;
      RECT  445800.0 793200.0 456000.0 779400.0 ;
      RECT  445800.0 793200.0 456000.0 807000.0 ;
      RECT  445800.0 820800.0 456000.0 807000.0 ;
      RECT  445800.0 820800.0 456000.0 834600.0 ;
      RECT  445800.0 848400.0 456000.0 834600.0 ;
      RECT  445800.0 848400.0 456000.0 862200.0 ;
      RECT  445800.0 876000.0 456000.0 862200.0 ;
      RECT  445800.0 876000.0 456000.0 889800.0 ;
      RECT  445800.0 903600.0 456000.0 889800.0 ;
      RECT  445800.0 903600.0 456000.0 917400.0 ;
      RECT  445800.0 931200.0 456000.0 917400.0 ;
      RECT  445800.0 931200.0 456000.0 945000.0 ;
      RECT  445800.0 958800.0 456000.0 945000.0 ;
      RECT  445800.0 958800.0 456000.0 972600.0 ;
      RECT  445800.0 986400.0 456000.0 972600.0 ;
      RECT  445800.0 986400.0 456000.0 1000200.0 ;
      RECT  445800.0 1014000.0 456000.0 1000200.0 ;
      RECT  445800.0 1014000.0 456000.0 1027800.0 ;
      RECT  445800.0 1041600.0 456000.0 1027800.0 ;
      RECT  445800.0 1041600.0 456000.0 1055400.0 ;
      RECT  445800.0 1069200.0 456000.0 1055400.0 ;
      RECT  445800.0 1069200.0 456000.0 1083000.0 ;
      RECT  445800.0 1096800.0 456000.0 1083000.0 ;
      RECT  445800.0 1096800.0 456000.0 1110600.0 ;
      RECT  445800.0 1124400.0 456000.0 1110600.0 ;
      RECT  445800.0 1124400.0 456000.0 1138200.0 ;
      RECT  445800.0 1152000.0 456000.0 1138200.0 ;
      RECT  445800.0 1152000.0 456000.0 1165800.0 ;
      RECT  445800.0 1179600.0 456000.0 1165800.0 ;
      RECT  445800.0 1179600.0 456000.0 1193400.0 ;
      RECT  445800.0 1207200.0 456000.0 1193400.0 ;
      RECT  445800.0 1207200.0 456000.0 1221000.0 ;
      RECT  445800.0 1234800.0 456000.0 1221000.0 ;
      RECT  445800.0 1234800.0 456000.0 1248600.0 ;
      RECT  445800.0 1262400.0 456000.0 1248600.0 ;
      RECT  445800.0 1262400.0 456000.0 1276200.0 ;
      RECT  445800.0 1290000.0 456000.0 1276200.0 ;
      RECT  445800.0 1290000.0 456000.0 1303800.0 ;
      RECT  445800.0 1317600.0 456000.0 1303800.0 ;
      RECT  445800.0 1317600.0 456000.0 1331400.0 ;
      RECT  445800.0 1345200.0 456000.0 1331400.0 ;
      RECT  445800.0 1345200.0 456000.0 1359000.0 ;
      RECT  445800.0 1372800.0 456000.0 1359000.0 ;
      RECT  445800.0 1372800.0 456000.0 1386600.0 ;
      RECT  445800.0 1400400.0 456000.0 1386600.0 ;
      RECT  445800.0 1400400.0 456000.0 1414200.0 ;
      RECT  445800.0 1428000.0 456000.0 1414200.0 ;
      RECT  445800.0 1428000.0 456000.0 1441800.0 ;
      RECT  445800.0 1455600.0 456000.0 1441800.0 ;
      RECT  445800.0 1455600.0 456000.0 1469400.0 ;
      RECT  445800.0 1483200.0 456000.0 1469400.0 ;
      RECT  445800.0 1483200.0 456000.0 1497000.0 ;
      RECT  445800.0 1510800.0 456000.0 1497000.0 ;
      RECT  445800.0 1510800.0 456000.0 1524600.0 ;
      RECT  445800.0 1538400.0 456000.0 1524600.0 ;
      RECT  445800.0 1538400.0 456000.0 1552200.0 ;
      RECT  445800.0 1566000.0 456000.0 1552200.0 ;
      RECT  445800.0 1566000.0 456000.0 1579800.0 ;
      RECT  445800.0 1593600.0 456000.0 1579800.0 ;
      RECT  445800.0 1593600.0 456000.0 1607400.0 ;
      RECT  445800.0 1621200.0 456000.0 1607400.0 ;
      RECT  445800.0 1621200.0 456000.0 1635000.0 ;
      RECT  445800.0 1648800.0 456000.0 1635000.0 ;
      RECT  445800.0 1648800.0 456000.0 1662600.0 ;
      RECT  445800.0 1676400.0 456000.0 1662600.0 ;
      RECT  445800.0 1676400.0 456000.0 1690200.0 ;
      RECT  445800.0 1704000.0 456000.0 1690200.0 ;
      RECT  445800.0 1704000.0 456000.0 1717800.0 ;
      RECT  445800.0 1731600.0 456000.0 1717800.0 ;
      RECT  445800.0 1731600.0 456000.0 1745400.0 ;
      RECT  445800.0 1759200.0 456000.0 1745400.0 ;
      RECT  445800.0 1759200.0 456000.0 1773000.0 ;
      RECT  445800.0 1786800.0 456000.0 1773000.0 ;
      RECT  445800.0 1786800.0 456000.0 1800600.0 ;
      RECT  445800.0 1814400.0 456000.0 1800600.0 ;
      RECT  445800.0 1814400.0 456000.0 1828200.0 ;
      RECT  445800.0 1842000.0 456000.0 1828200.0 ;
      RECT  445800.0 1842000.0 456000.0 1855800.0 ;
      RECT  445800.0 1869600.0 456000.0 1855800.0 ;
      RECT  445800.0 1869600.0 456000.0 1883400.0 ;
      RECT  445800.0 1897200.0 456000.0 1883400.0 ;
      RECT  445800.0 1897200.0 456000.0 1911000.0 ;
      RECT  445800.0 1924800.0 456000.0 1911000.0 ;
      RECT  445800.0 1924800.0 456000.0 1938600.0 ;
      RECT  445800.0 1952400.0 456000.0 1938600.0 ;
      RECT  445800.0 1952400.0 456000.0 1966200.0 ;
      RECT  445800.0 1980000.0 456000.0 1966200.0 ;
      RECT  445800.0 1980000.0 456000.0 1993800.0 ;
      RECT  445800.0 2007600.0 456000.0 1993800.0 ;
      RECT  445800.0 2007600.0 456000.0 2021400.0 ;
      RECT  445800.0 2035200.0 456000.0 2021400.0 ;
      RECT  445800.0 2035200.0 456000.0 2049000.0 ;
      RECT  445800.0 2062800.0 456000.0 2049000.0 ;
      RECT  445800.0 2062800.0 456000.0 2076600.0 ;
      RECT  445800.0 2090400.0 456000.0 2076600.0 ;
      RECT  445800.0 2090400.0 456000.0 2104200.0 ;
      RECT  445800.0 2118000.0 456000.0 2104200.0 ;
      RECT  445800.0 2118000.0 456000.0 2131800.0 ;
      RECT  445800.0 2145600.0 456000.0 2131800.0 ;
      RECT  456000.0 379200.0 466200.0 393000.0 ;
      RECT  456000.0 406800.0 466200.0 393000.0 ;
      RECT  456000.0 406800.0 466200.0 420600.0 ;
      RECT  456000.0 434400.0 466200.0 420600.0 ;
      RECT  456000.0 434400.0 466200.0 448200.0 ;
      RECT  456000.0 462000.0 466200.0 448200.0 ;
      RECT  456000.0 462000.0 466200.0 475800.0 ;
      RECT  456000.0 489600.0 466200.0 475800.0 ;
      RECT  456000.0 489600.0 466200.0 503400.0 ;
      RECT  456000.0 517200.0 466200.0 503400.0 ;
      RECT  456000.0 517200.0 466200.0 531000.0 ;
      RECT  456000.0 544800.0 466200.0 531000.0 ;
      RECT  456000.0 544800.0 466200.0 558600.0 ;
      RECT  456000.0 572400.0 466200.0 558600.0 ;
      RECT  456000.0 572400.0 466200.0 586200.0 ;
      RECT  456000.0 600000.0 466200.0 586200.0 ;
      RECT  456000.0 600000.0 466200.0 613800.0 ;
      RECT  456000.0 627600.0 466200.0 613800.0 ;
      RECT  456000.0 627600.0 466200.0 641400.0 ;
      RECT  456000.0 655200.0 466200.0 641400.0 ;
      RECT  456000.0 655200.0 466200.0 669000.0 ;
      RECT  456000.0 682800.0 466200.0 669000.0 ;
      RECT  456000.0 682800.0 466200.0 696600.0 ;
      RECT  456000.0 710400.0 466200.0 696600.0 ;
      RECT  456000.0 710400.0 466200.0 724200.0 ;
      RECT  456000.0 738000.0 466200.0 724200.0 ;
      RECT  456000.0 738000.0 466200.0 751800.0 ;
      RECT  456000.0 765600.0 466200.0 751800.0 ;
      RECT  456000.0 765600.0 466200.0 779400.0 ;
      RECT  456000.0 793200.0 466200.0 779400.0 ;
      RECT  456000.0 793200.0 466200.0 807000.0 ;
      RECT  456000.0 820800.0 466200.0 807000.0 ;
      RECT  456000.0 820800.0 466200.0 834600.0 ;
      RECT  456000.0 848400.0 466200.0 834600.0 ;
      RECT  456000.0 848400.0 466200.0 862200.0 ;
      RECT  456000.0 876000.0 466200.0 862200.0 ;
      RECT  456000.0 876000.0 466200.0 889800.0 ;
      RECT  456000.0 903600.0 466200.0 889800.0 ;
      RECT  456000.0 903600.0 466200.0 917400.0 ;
      RECT  456000.0 931200.0 466200.0 917400.0 ;
      RECT  456000.0 931200.0 466200.0 945000.0 ;
      RECT  456000.0 958800.0 466200.0 945000.0 ;
      RECT  456000.0 958800.0 466200.0 972600.0 ;
      RECT  456000.0 986400.0 466200.0 972600.0 ;
      RECT  456000.0 986400.0 466200.0 1000200.0 ;
      RECT  456000.0 1014000.0 466200.0 1000200.0 ;
      RECT  456000.0 1014000.0 466200.0 1027800.0 ;
      RECT  456000.0 1041600.0 466200.0 1027800.0 ;
      RECT  456000.0 1041600.0 466200.0 1055400.0 ;
      RECT  456000.0 1069200.0 466200.0 1055400.0 ;
      RECT  456000.0 1069200.0 466200.0 1083000.0 ;
      RECT  456000.0 1096800.0 466200.0 1083000.0 ;
      RECT  456000.0 1096800.0 466200.0 1110600.0 ;
      RECT  456000.0 1124400.0 466200.0 1110600.0 ;
      RECT  456000.0 1124400.0 466200.0 1138200.0 ;
      RECT  456000.0 1152000.0 466200.0 1138200.0 ;
      RECT  456000.0 1152000.0 466200.0 1165800.0 ;
      RECT  456000.0 1179600.0 466200.0 1165800.0 ;
      RECT  456000.0 1179600.0 466200.0 1193400.0 ;
      RECT  456000.0 1207200.0 466200.0 1193400.0 ;
      RECT  456000.0 1207200.0 466200.0 1221000.0 ;
      RECT  456000.0 1234800.0 466200.0 1221000.0 ;
      RECT  456000.0 1234800.0 466200.0 1248600.0 ;
      RECT  456000.0 1262400.0 466200.0 1248600.0 ;
      RECT  456000.0 1262400.0 466200.0 1276200.0 ;
      RECT  456000.0 1290000.0 466200.0 1276200.0 ;
      RECT  456000.0 1290000.0 466200.0 1303800.0 ;
      RECT  456000.0 1317600.0 466200.0 1303800.0 ;
      RECT  456000.0 1317600.0 466200.0 1331400.0 ;
      RECT  456000.0 1345200.0 466200.0 1331400.0 ;
      RECT  456000.0 1345200.0 466200.0 1359000.0 ;
      RECT  456000.0 1372800.0 466200.0 1359000.0 ;
      RECT  456000.0 1372800.0 466200.0 1386600.0 ;
      RECT  456000.0 1400400.0 466200.0 1386600.0 ;
      RECT  456000.0 1400400.0 466200.0 1414200.0 ;
      RECT  456000.0 1428000.0 466200.0 1414200.0 ;
      RECT  456000.0 1428000.0 466200.0 1441800.0 ;
      RECT  456000.0 1455600.0 466200.0 1441800.0 ;
      RECT  456000.0 1455600.0 466200.0 1469400.0 ;
      RECT  456000.0 1483200.0 466200.0 1469400.0 ;
      RECT  456000.0 1483200.0 466200.0 1497000.0 ;
      RECT  456000.0 1510800.0 466200.0 1497000.0 ;
      RECT  456000.0 1510800.0 466200.0 1524600.0 ;
      RECT  456000.0 1538400.0 466200.0 1524600.0 ;
      RECT  456000.0 1538400.0 466200.0 1552200.0 ;
      RECT  456000.0 1566000.0 466200.0 1552200.0 ;
      RECT  456000.0 1566000.0 466200.0 1579800.0 ;
      RECT  456000.0 1593600.0 466200.0 1579800.0 ;
      RECT  456000.0 1593600.0 466200.0 1607400.0 ;
      RECT  456000.0 1621200.0 466200.0 1607400.0 ;
      RECT  456000.0 1621200.0 466200.0 1635000.0 ;
      RECT  456000.0 1648800.0 466200.0 1635000.0 ;
      RECT  456000.0 1648800.0 466200.0 1662600.0 ;
      RECT  456000.0 1676400.0 466200.0 1662600.0 ;
      RECT  456000.0 1676400.0 466200.0 1690200.0 ;
      RECT  456000.0 1704000.0 466200.0 1690200.0 ;
      RECT  456000.0 1704000.0 466200.0 1717800.0 ;
      RECT  456000.0 1731600.0 466200.0 1717800.0 ;
      RECT  456000.0 1731600.0 466200.0 1745400.0 ;
      RECT  456000.0 1759200.0 466200.0 1745400.0 ;
      RECT  456000.0 1759200.0 466200.0 1773000.0 ;
      RECT  456000.0 1786800.0 466200.0 1773000.0 ;
      RECT  456000.0 1786800.0 466200.0 1800600.0 ;
      RECT  456000.0 1814400.0 466200.0 1800600.0 ;
      RECT  456000.0 1814400.0 466200.0 1828200.0 ;
      RECT  456000.0 1842000.0 466200.0 1828200.0 ;
      RECT  456000.0 1842000.0 466200.0 1855800.0 ;
      RECT  456000.0 1869600.0 466200.0 1855800.0 ;
      RECT  456000.0 1869600.0 466200.0 1883400.0 ;
      RECT  456000.0 1897200.0 466200.0 1883400.0 ;
      RECT  456000.0 1897200.0 466200.0 1911000.0 ;
      RECT  456000.0 1924800.0 466200.0 1911000.0 ;
      RECT  456000.0 1924800.0 466200.0 1938600.0 ;
      RECT  456000.0 1952400.0 466200.0 1938600.0 ;
      RECT  456000.0 1952400.0 466200.0 1966200.0 ;
      RECT  456000.0 1980000.0 466200.0 1966200.0 ;
      RECT  456000.0 1980000.0 466200.0 1993800.0 ;
      RECT  456000.0 2007600.0 466200.0 1993800.0 ;
      RECT  456000.0 2007600.0 466200.0 2021400.0 ;
      RECT  456000.0 2035200.0 466200.0 2021400.0 ;
      RECT  456000.0 2035200.0 466200.0 2049000.0 ;
      RECT  456000.0 2062800.0 466200.0 2049000.0 ;
      RECT  456000.0 2062800.0 466200.0 2076600.0 ;
      RECT  456000.0 2090400.0 466200.0 2076600.0 ;
      RECT  456000.0 2090400.0 466200.0 2104200.0 ;
      RECT  456000.0 2118000.0 466200.0 2104200.0 ;
      RECT  456000.0 2118000.0 466200.0 2131800.0 ;
      RECT  456000.0 2145600.0 466200.0 2131800.0 ;
      RECT  466200.0 379200.0 476400.0 393000.0 ;
      RECT  466200.0 406800.0 476400.0 393000.0 ;
      RECT  466200.0 406800.0 476400.0 420600.0 ;
      RECT  466200.0 434400.0 476400.0 420600.0 ;
      RECT  466200.0 434400.0 476400.0 448200.0 ;
      RECT  466200.0 462000.0 476400.0 448200.0 ;
      RECT  466200.0 462000.0 476400.0 475800.0 ;
      RECT  466200.0 489600.0 476400.0 475800.0 ;
      RECT  466200.0 489600.0 476400.0 503400.0 ;
      RECT  466200.0 517200.0 476400.0 503400.0 ;
      RECT  466200.0 517200.0 476400.0 531000.0 ;
      RECT  466200.0 544800.0 476400.0 531000.0 ;
      RECT  466200.0 544800.0 476400.0 558600.0 ;
      RECT  466200.0 572400.0 476400.0 558600.0 ;
      RECT  466200.0 572400.0 476400.0 586200.0 ;
      RECT  466200.0 600000.0 476400.0 586200.0 ;
      RECT  466200.0 600000.0 476400.0 613800.0 ;
      RECT  466200.0 627600.0 476400.0 613800.0 ;
      RECT  466200.0 627600.0 476400.0 641400.0 ;
      RECT  466200.0 655200.0 476400.0 641400.0 ;
      RECT  466200.0 655200.0 476400.0 669000.0 ;
      RECT  466200.0 682800.0 476400.0 669000.0 ;
      RECT  466200.0 682800.0 476400.0 696600.0 ;
      RECT  466200.0 710400.0 476400.0 696600.0 ;
      RECT  466200.0 710400.0 476400.0 724200.0 ;
      RECT  466200.0 738000.0 476400.0 724200.0 ;
      RECT  466200.0 738000.0 476400.0 751800.0 ;
      RECT  466200.0 765600.0 476400.0 751800.0 ;
      RECT  466200.0 765600.0 476400.0 779400.0 ;
      RECT  466200.0 793200.0 476400.0 779400.0 ;
      RECT  466200.0 793200.0 476400.0 807000.0 ;
      RECT  466200.0 820800.0 476400.0 807000.0 ;
      RECT  466200.0 820800.0 476400.0 834600.0 ;
      RECT  466200.0 848400.0 476400.0 834600.0 ;
      RECT  466200.0 848400.0 476400.0 862200.0 ;
      RECT  466200.0 876000.0 476400.0 862200.0 ;
      RECT  466200.0 876000.0 476400.0 889800.0 ;
      RECT  466200.0 903600.0 476400.0 889800.0 ;
      RECT  466200.0 903600.0 476400.0 917400.0 ;
      RECT  466200.0 931200.0 476400.0 917400.0 ;
      RECT  466200.0 931200.0 476400.0 945000.0 ;
      RECT  466200.0 958800.0 476400.0 945000.0 ;
      RECT  466200.0 958800.0 476400.0 972600.0 ;
      RECT  466200.0 986400.0 476400.0 972600.0 ;
      RECT  466200.0 986400.0 476400.0 1000200.0 ;
      RECT  466200.0 1014000.0 476400.0 1000200.0 ;
      RECT  466200.0 1014000.0 476400.0 1027800.0 ;
      RECT  466200.0 1041600.0 476400.0 1027800.0 ;
      RECT  466200.0 1041600.0 476400.0 1055400.0 ;
      RECT  466200.0 1069200.0 476400.0 1055400.0 ;
      RECT  466200.0 1069200.0 476400.0 1083000.0 ;
      RECT  466200.0 1096800.0 476400.0 1083000.0 ;
      RECT  466200.0 1096800.0 476400.0 1110600.0 ;
      RECT  466200.0 1124400.0 476400.0 1110600.0 ;
      RECT  466200.0 1124400.0 476400.0 1138200.0 ;
      RECT  466200.0 1152000.0 476400.0 1138200.0 ;
      RECT  466200.0 1152000.0 476400.0 1165800.0 ;
      RECT  466200.0 1179600.0 476400.0 1165800.0 ;
      RECT  466200.0 1179600.0 476400.0 1193400.0 ;
      RECT  466200.0 1207200.0 476400.0 1193400.0 ;
      RECT  466200.0 1207200.0 476400.0 1221000.0 ;
      RECT  466200.0 1234800.0 476400.0 1221000.0 ;
      RECT  466200.0 1234800.0 476400.0 1248600.0 ;
      RECT  466200.0 1262400.0 476400.0 1248600.0 ;
      RECT  466200.0 1262400.0 476400.0 1276200.0 ;
      RECT  466200.0 1290000.0 476400.0 1276200.0 ;
      RECT  466200.0 1290000.0 476400.0 1303800.0 ;
      RECT  466200.0 1317600.0 476400.0 1303800.0 ;
      RECT  466200.0 1317600.0 476400.0 1331400.0 ;
      RECT  466200.0 1345200.0 476400.0 1331400.0 ;
      RECT  466200.0 1345200.0 476400.0 1359000.0 ;
      RECT  466200.0 1372800.0 476400.0 1359000.0 ;
      RECT  466200.0 1372800.0 476400.0 1386600.0 ;
      RECT  466200.0 1400400.0 476400.0 1386600.0 ;
      RECT  466200.0 1400400.0 476400.0 1414200.0 ;
      RECT  466200.0 1428000.0 476400.0 1414200.0 ;
      RECT  466200.0 1428000.0 476400.0 1441800.0 ;
      RECT  466200.0 1455600.0 476400.0 1441800.0 ;
      RECT  466200.0 1455600.0 476400.0 1469400.0 ;
      RECT  466200.0 1483200.0 476400.0 1469400.0 ;
      RECT  466200.0 1483200.0 476400.0 1497000.0 ;
      RECT  466200.0 1510800.0 476400.0 1497000.0 ;
      RECT  466200.0 1510800.0 476400.0 1524600.0 ;
      RECT  466200.0 1538400.0 476400.0 1524600.0 ;
      RECT  466200.0 1538400.0 476400.0 1552200.0 ;
      RECT  466200.0 1566000.0 476400.0 1552200.0 ;
      RECT  466200.0 1566000.0 476400.0 1579800.0 ;
      RECT  466200.0 1593600.0 476400.0 1579800.0 ;
      RECT  466200.0 1593600.0 476400.0 1607400.0 ;
      RECT  466200.0 1621200.0 476400.0 1607400.0 ;
      RECT  466200.0 1621200.0 476400.0 1635000.0 ;
      RECT  466200.0 1648800.0 476400.0 1635000.0 ;
      RECT  466200.0 1648800.0 476400.0 1662600.0 ;
      RECT  466200.0 1676400.0 476400.0 1662600.0 ;
      RECT  466200.0 1676400.0 476400.0 1690200.0 ;
      RECT  466200.0 1704000.0 476400.0 1690200.0 ;
      RECT  466200.0 1704000.0 476400.0 1717800.0 ;
      RECT  466200.0 1731600.0 476400.0 1717800.0 ;
      RECT  466200.0 1731600.0 476400.0 1745400.0 ;
      RECT  466200.0 1759200.0 476400.0 1745400.0 ;
      RECT  466200.0 1759200.0 476400.0 1773000.0 ;
      RECT  466200.0 1786800.0 476400.0 1773000.0 ;
      RECT  466200.0 1786800.0 476400.0 1800600.0 ;
      RECT  466200.0 1814400.0 476400.0 1800600.0 ;
      RECT  466200.0 1814400.0 476400.0 1828200.0 ;
      RECT  466200.0 1842000.0 476400.0 1828200.0 ;
      RECT  466200.0 1842000.0 476400.0 1855800.0 ;
      RECT  466200.0 1869600.0 476400.0 1855800.0 ;
      RECT  466200.0 1869600.0 476400.0 1883400.0 ;
      RECT  466200.0 1897200.0 476400.0 1883400.0 ;
      RECT  466200.0 1897200.0 476400.0 1911000.0 ;
      RECT  466200.0 1924800.0 476400.0 1911000.0 ;
      RECT  466200.0 1924800.0 476400.0 1938600.0 ;
      RECT  466200.0 1952400.0 476400.0 1938600.0 ;
      RECT  466200.0 1952400.0 476400.0 1966200.0 ;
      RECT  466200.0 1980000.0 476400.0 1966200.0 ;
      RECT  466200.0 1980000.0 476400.0 1993800.0 ;
      RECT  466200.0 2007600.0 476400.0 1993800.0 ;
      RECT  466200.0 2007600.0 476400.0 2021400.0 ;
      RECT  466200.0 2035200.0 476400.0 2021400.0 ;
      RECT  466200.0 2035200.0 476400.0 2049000.0 ;
      RECT  466200.0 2062800.0 476400.0 2049000.0 ;
      RECT  466200.0 2062800.0 476400.0 2076600.0 ;
      RECT  466200.0 2090400.0 476400.0 2076600.0 ;
      RECT  466200.0 2090400.0 476400.0 2104200.0 ;
      RECT  466200.0 2118000.0 476400.0 2104200.0 ;
      RECT  466200.0 2118000.0 476400.0 2131800.0 ;
      RECT  466200.0 2145600.0 476400.0 2131800.0 ;
      RECT  476400.0 379200.0 486600.0 393000.0 ;
      RECT  476400.0 406800.0 486600.0 393000.0 ;
      RECT  476400.0 406800.0 486600.0 420600.0 ;
      RECT  476400.0 434400.0 486600.0 420600.0 ;
      RECT  476400.0 434400.0 486600.0 448200.0 ;
      RECT  476400.0 462000.0 486600.0 448200.0 ;
      RECT  476400.0 462000.0 486600.0 475800.0 ;
      RECT  476400.0 489600.0 486600.0 475800.0 ;
      RECT  476400.0 489600.0 486600.0 503400.0 ;
      RECT  476400.0 517200.0 486600.0 503400.0 ;
      RECT  476400.0 517200.0 486600.0 531000.0 ;
      RECT  476400.0 544800.0 486600.0 531000.0 ;
      RECT  476400.0 544800.0 486600.0 558600.0 ;
      RECT  476400.0 572400.0 486600.0 558600.0 ;
      RECT  476400.0 572400.0 486600.0 586200.0 ;
      RECT  476400.0 600000.0 486600.0 586200.0 ;
      RECT  476400.0 600000.0 486600.0 613800.0 ;
      RECT  476400.0 627600.0 486600.0 613800.0 ;
      RECT  476400.0 627600.0 486600.0 641400.0 ;
      RECT  476400.0 655200.0 486600.0 641400.0 ;
      RECT  476400.0 655200.0 486600.0 669000.0 ;
      RECT  476400.0 682800.0 486600.0 669000.0 ;
      RECT  476400.0 682800.0 486600.0 696600.0 ;
      RECT  476400.0 710400.0 486600.0 696600.0 ;
      RECT  476400.0 710400.0 486600.0 724200.0 ;
      RECT  476400.0 738000.0 486600.0 724200.0 ;
      RECT  476400.0 738000.0 486600.0 751800.0 ;
      RECT  476400.0 765600.0 486600.0 751800.0 ;
      RECT  476400.0 765600.0 486600.0 779400.0 ;
      RECT  476400.0 793200.0 486600.0 779400.0 ;
      RECT  476400.0 793200.0 486600.0 807000.0 ;
      RECT  476400.0 820800.0 486600.0 807000.0 ;
      RECT  476400.0 820800.0 486600.0 834600.0 ;
      RECT  476400.0 848400.0 486600.0 834600.0 ;
      RECT  476400.0 848400.0 486600.0 862200.0 ;
      RECT  476400.0 876000.0 486600.0 862200.0 ;
      RECT  476400.0 876000.0 486600.0 889800.0 ;
      RECT  476400.0 903600.0 486600.0 889800.0 ;
      RECT  476400.0 903600.0 486600.0 917400.0 ;
      RECT  476400.0 931200.0 486600.0 917400.0 ;
      RECT  476400.0 931200.0 486600.0 945000.0 ;
      RECT  476400.0 958800.0 486600.0 945000.0 ;
      RECT  476400.0 958800.0 486600.0 972600.0 ;
      RECT  476400.0 986400.0 486600.0 972600.0 ;
      RECT  476400.0 986400.0 486600.0 1000200.0 ;
      RECT  476400.0 1014000.0 486600.0 1000200.0 ;
      RECT  476400.0 1014000.0 486600.0 1027800.0 ;
      RECT  476400.0 1041600.0 486600.0 1027800.0 ;
      RECT  476400.0 1041600.0 486600.0 1055400.0 ;
      RECT  476400.0 1069200.0 486600.0 1055400.0 ;
      RECT  476400.0 1069200.0 486600.0 1083000.0 ;
      RECT  476400.0 1096800.0 486600.0 1083000.0 ;
      RECT  476400.0 1096800.0 486600.0 1110600.0 ;
      RECT  476400.0 1124400.0 486600.0 1110600.0 ;
      RECT  476400.0 1124400.0 486600.0 1138200.0 ;
      RECT  476400.0 1152000.0 486600.0 1138200.0 ;
      RECT  476400.0 1152000.0 486600.0 1165800.0 ;
      RECT  476400.0 1179600.0 486600.0 1165800.0 ;
      RECT  476400.0 1179600.0 486600.0 1193400.0 ;
      RECT  476400.0 1207200.0 486600.0 1193400.0 ;
      RECT  476400.0 1207200.0 486600.0 1221000.0 ;
      RECT  476400.0 1234800.0 486600.0 1221000.0 ;
      RECT  476400.0 1234800.0 486600.0 1248600.0 ;
      RECT  476400.0 1262400.0 486600.0 1248600.0 ;
      RECT  476400.0 1262400.0 486600.0 1276200.0 ;
      RECT  476400.0 1290000.0 486600.0 1276200.0 ;
      RECT  476400.0 1290000.0 486600.0 1303800.0 ;
      RECT  476400.0 1317600.0 486600.0 1303800.0 ;
      RECT  476400.0 1317600.0 486600.0 1331400.0 ;
      RECT  476400.0 1345200.0 486600.0 1331400.0 ;
      RECT  476400.0 1345200.0 486600.0 1359000.0 ;
      RECT  476400.0 1372800.0 486600.0 1359000.0 ;
      RECT  476400.0 1372800.0 486600.0 1386600.0 ;
      RECT  476400.0 1400400.0 486600.0 1386600.0 ;
      RECT  476400.0 1400400.0 486600.0 1414200.0 ;
      RECT  476400.0 1428000.0 486600.0 1414200.0 ;
      RECT  476400.0 1428000.0 486600.0 1441800.0 ;
      RECT  476400.0 1455600.0 486600.0 1441800.0 ;
      RECT  476400.0 1455600.0 486600.0 1469400.0 ;
      RECT  476400.0 1483200.0 486600.0 1469400.0 ;
      RECT  476400.0 1483200.0 486600.0 1497000.0 ;
      RECT  476400.0 1510800.0 486600.0 1497000.0 ;
      RECT  476400.0 1510800.0 486600.0 1524600.0 ;
      RECT  476400.0 1538400.0 486600.0 1524600.0 ;
      RECT  476400.0 1538400.0 486600.0 1552200.0 ;
      RECT  476400.0 1566000.0 486600.0 1552200.0 ;
      RECT  476400.0 1566000.0 486600.0 1579800.0 ;
      RECT  476400.0 1593600.0 486600.0 1579800.0 ;
      RECT  476400.0 1593600.0 486600.0 1607400.0 ;
      RECT  476400.0 1621200.0 486600.0 1607400.0 ;
      RECT  476400.0 1621200.0 486600.0 1635000.0 ;
      RECT  476400.0 1648800.0 486600.0 1635000.0 ;
      RECT  476400.0 1648800.0 486600.0 1662600.0 ;
      RECT  476400.0 1676400.0 486600.0 1662600.0 ;
      RECT  476400.0 1676400.0 486600.0 1690200.0 ;
      RECT  476400.0 1704000.0 486600.0 1690200.0 ;
      RECT  476400.0 1704000.0 486600.0 1717800.0 ;
      RECT  476400.0 1731600.0 486600.0 1717800.0 ;
      RECT  476400.0 1731600.0 486600.0 1745400.0 ;
      RECT  476400.0 1759200.0 486600.0 1745400.0 ;
      RECT  476400.0 1759200.0 486600.0 1773000.0 ;
      RECT  476400.0 1786800.0 486600.0 1773000.0 ;
      RECT  476400.0 1786800.0 486600.0 1800600.0 ;
      RECT  476400.0 1814400.0 486600.0 1800600.0 ;
      RECT  476400.0 1814400.0 486600.0 1828200.0 ;
      RECT  476400.0 1842000.0 486600.0 1828200.0 ;
      RECT  476400.0 1842000.0 486600.0 1855800.0 ;
      RECT  476400.0 1869600.0 486600.0 1855800.0 ;
      RECT  476400.0 1869600.0 486600.0 1883400.0 ;
      RECT  476400.0 1897200.0 486600.0 1883400.0 ;
      RECT  476400.0 1897200.0 486600.0 1911000.0 ;
      RECT  476400.0 1924800.0 486600.0 1911000.0 ;
      RECT  476400.0 1924800.0 486600.0 1938600.0 ;
      RECT  476400.0 1952400.0 486600.0 1938600.0 ;
      RECT  476400.0 1952400.0 486600.0 1966200.0 ;
      RECT  476400.0 1980000.0 486600.0 1966200.0 ;
      RECT  476400.0 1980000.0 486600.0 1993800.0 ;
      RECT  476400.0 2007600.0 486600.0 1993800.0 ;
      RECT  476400.0 2007600.0 486600.0 2021400.0 ;
      RECT  476400.0 2035200.0 486600.0 2021400.0 ;
      RECT  476400.0 2035200.0 486600.0 2049000.0 ;
      RECT  476400.0 2062800.0 486600.0 2049000.0 ;
      RECT  476400.0 2062800.0 486600.0 2076600.0 ;
      RECT  476400.0 2090400.0 486600.0 2076600.0 ;
      RECT  476400.0 2090400.0 486600.0 2104200.0 ;
      RECT  476400.0 2118000.0 486600.0 2104200.0 ;
      RECT  476400.0 2118000.0 486600.0 2131800.0 ;
      RECT  476400.0 2145600.0 486600.0 2131800.0 ;
      RECT  486600.0 379200.0 496800.0 393000.0 ;
      RECT  486600.0 406800.0 496800.0 393000.0 ;
      RECT  486600.0 406800.0 496800.0 420600.0 ;
      RECT  486600.0 434400.0 496800.0 420600.0 ;
      RECT  486600.0 434400.0 496800.0 448200.0 ;
      RECT  486600.0 462000.0 496800.0 448200.0 ;
      RECT  486600.0 462000.0 496800.0 475800.0 ;
      RECT  486600.0 489600.0 496800.0 475800.0 ;
      RECT  486600.0 489600.0 496800.0 503400.0 ;
      RECT  486600.0 517200.0 496800.0 503400.0 ;
      RECT  486600.0 517200.0 496800.0 531000.0 ;
      RECT  486600.0 544800.0 496800.0 531000.0 ;
      RECT  486600.0 544800.0 496800.0 558600.0 ;
      RECT  486600.0 572400.0 496800.0 558600.0 ;
      RECT  486600.0 572400.0 496800.0 586200.0 ;
      RECT  486600.0 600000.0 496800.0 586200.0 ;
      RECT  486600.0 600000.0 496800.0 613800.0 ;
      RECT  486600.0 627600.0 496800.0 613800.0 ;
      RECT  486600.0 627600.0 496800.0 641400.0 ;
      RECT  486600.0 655200.0 496800.0 641400.0 ;
      RECT  486600.0 655200.0 496800.0 669000.0 ;
      RECT  486600.0 682800.0 496800.0 669000.0 ;
      RECT  486600.0 682800.0 496800.0 696600.0 ;
      RECT  486600.0 710400.0 496800.0 696600.0 ;
      RECT  486600.0 710400.0 496800.0 724200.0 ;
      RECT  486600.0 738000.0 496800.0 724200.0 ;
      RECT  486600.0 738000.0 496800.0 751800.0 ;
      RECT  486600.0 765600.0 496800.0 751800.0 ;
      RECT  486600.0 765600.0 496800.0 779400.0 ;
      RECT  486600.0 793200.0 496800.0 779400.0 ;
      RECT  486600.0 793200.0 496800.0 807000.0 ;
      RECT  486600.0 820800.0 496800.0 807000.0 ;
      RECT  486600.0 820800.0 496800.0 834600.0 ;
      RECT  486600.0 848400.0 496800.0 834600.0 ;
      RECT  486600.0 848400.0 496800.0 862200.0 ;
      RECT  486600.0 876000.0 496800.0 862200.0 ;
      RECT  486600.0 876000.0 496800.0 889800.0 ;
      RECT  486600.0 903600.0 496800.0 889800.0 ;
      RECT  486600.0 903600.0 496800.0 917400.0 ;
      RECT  486600.0 931200.0 496800.0 917400.0 ;
      RECT  486600.0 931200.0 496800.0 945000.0 ;
      RECT  486600.0 958800.0 496800.0 945000.0 ;
      RECT  486600.0 958800.0 496800.0 972600.0 ;
      RECT  486600.0 986400.0 496800.0 972600.0 ;
      RECT  486600.0 986400.0 496800.0 1000200.0 ;
      RECT  486600.0 1014000.0 496800.0 1000200.0 ;
      RECT  486600.0 1014000.0 496800.0 1027800.0 ;
      RECT  486600.0 1041600.0 496800.0 1027800.0 ;
      RECT  486600.0 1041600.0 496800.0 1055400.0 ;
      RECT  486600.0 1069200.0 496800.0 1055400.0 ;
      RECT  486600.0 1069200.0 496800.0 1083000.0 ;
      RECT  486600.0 1096800.0 496800.0 1083000.0 ;
      RECT  486600.0 1096800.0 496800.0 1110600.0 ;
      RECT  486600.0 1124400.0 496800.0 1110600.0 ;
      RECT  486600.0 1124400.0 496800.0 1138200.0 ;
      RECT  486600.0 1152000.0 496800.0 1138200.0 ;
      RECT  486600.0 1152000.0 496800.0 1165800.0 ;
      RECT  486600.0 1179600.0 496800.0 1165800.0 ;
      RECT  486600.0 1179600.0 496800.0 1193400.0 ;
      RECT  486600.0 1207200.0 496800.0 1193400.0 ;
      RECT  486600.0 1207200.0 496800.0 1221000.0 ;
      RECT  486600.0 1234800.0 496800.0 1221000.0 ;
      RECT  486600.0 1234800.0 496800.0 1248600.0 ;
      RECT  486600.0 1262400.0 496800.0 1248600.0 ;
      RECT  486600.0 1262400.0 496800.0 1276200.0 ;
      RECT  486600.0 1290000.0 496800.0 1276200.0 ;
      RECT  486600.0 1290000.0 496800.0 1303800.0 ;
      RECT  486600.0 1317600.0 496800.0 1303800.0 ;
      RECT  486600.0 1317600.0 496800.0 1331400.0 ;
      RECT  486600.0 1345200.0 496800.0 1331400.0 ;
      RECT  486600.0 1345200.0 496800.0 1359000.0 ;
      RECT  486600.0 1372800.0 496800.0 1359000.0 ;
      RECT  486600.0 1372800.0 496800.0 1386600.0 ;
      RECT  486600.0 1400400.0 496800.0 1386600.0 ;
      RECT  486600.0 1400400.0 496800.0 1414200.0 ;
      RECT  486600.0 1428000.0 496800.0 1414200.0 ;
      RECT  486600.0 1428000.0 496800.0 1441800.0 ;
      RECT  486600.0 1455600.0 496800.0 1441800.0 ;
      RECT  486600.0 1455600.0 496800.0 1469400.0 ;
      RECT  486600.0 1483200.0 496800.0 1469400.0 ;
      RECT  486600.0 1483200.0 496800.0 1497000.0 ;
      RECT  486600.0 1510800.0 496800.0 1497000.0 ;
      RECT  486600.0 1510800.0 496800.0 1524600.0 ;
      RECT  486600.0 1538400.0 496800.0 1524600.0 ;
      RECT  486600.0 1538400.0 496800.0 1552200.0 ;
      RECT  486600.0 1566000.0 496800.0 1552200.0 ;
      RECT  486600.0 1566000.0 496800.0 1579800.0 ;
      RECT  486600.0 1593600.0 496800.0 1579800.0 ;
      RECT  486600.0 1593600.0 496800.0 1607400.0 ;
      RECT  486600.0 1621200.0 496800.0 1607400.0 ;
      RECT  486600.0 1621200.0 496800.0 1635000.0 ;
      RECT  486600.0 1648800.0 496800.0 1635000.0 ;
      RECT  486600.0 1648800.0 496800.0 1662600.0 ;
      RECT  486600.0 1676400.0 496800.0 1662600.0 ;
      RECT  486600.0 1676400.0 496800.0 1690200.0 ;
      RECT  486600.0 1704000.0 496800.0 1690200.0 ;
      RECT  486600.0 1704000.0 496800.0 1717800.0 ;
      RECT  486600.0 1731600.0 496800.0 1717800.0 ;
      RECT  486600.0 1731600.0 496800.0 1745400.0 ;
      RECT  486600.0 1759200.0 496800.0 1745400.0 ;
      RECT  486600.0 1759200.0 496800.0 1773000.0 ;
      RECT  486600.0 1786800.0 496800.0 1773000.0 ;
      RECT  486600.0 1786800.0 496800.0 1800600.0 ;
      RECT  486600.0 1814400.0 496800.0 1800600.0 ;
      RECT  486600.0 1814400.0 496800.0 1828200.0 ;
      RECT  486600.0 1842000.0 496800.0 1828200.0 ;
      RECT  486600.0 1842000.0 496800.0 1855800.0 ;
      RECT  486600.0 1869600.0 496800.0 1855800.0 ;
      RECT  486600.0 1869600.0 496800.0 1883400.0 ;
      RECT  486600.0 1897200.0 496800.0 1883400.0 ;
      RECT  486600.0 1897200.0 496800.0 1911000.0 ;
      RECT  486600.0 1924800.0 496800.0 1911000.0 ;
      RECT  486600.0 1924800.0 496800.0 1938600.0 ;
      RECT  486600.0 1952400.0 496800.0 1938600.0 ;
      RECT  486600.0 1952400.0 496800.0 1966200.0 ;
      RECT  486600.0 1980000.0 496800.0 1966200.0 ;
      RECT  486600.0 1980000.0 496800.0 1993800.0 ;
      RECT  486600.0 2007600.0 496800.0 1993800.0 ;
      RECT  486600.0 2007600.0 496800.0 2021400.0 ;
      RECT  486600.0 2035200.0 496800.0 2021400.0 ;
      RECT  486600.0 2035200.0 496800.0 2049000.0 ;
      RECT  486600.0 2062800.0 496800.0 2049000.0 ;
      RECT  486600.0 2062800.0 496800.0 2076600.0 ;
      RECT  486600.0 2090400.0 496800.0 2076600.0 ;
      RECT  486600.0 2090400.0 496800.0 2104200.0 ;
      RECT  486600.0 2118000.0 496800.0 2104200.0 ;
      RECT  486600.0 2118000.0 496800.0 2131800.0 ;
      RECT  486600.0 2145600.0 496800.0 2131800.0 ;
      RECT  496800.0 379200.0 507000.0 393000.0 ;
      RECT  496800.0 406800.0 507000.0 393000.0 ;
      RECT  496800.0 406800.0 507000.0 420600.0 ;
      RECT  496800.0 434400.0 507000.0 420600.0 ;
      RECT  496800.0 434400.0 507000.0 448200.0 ;
      RECT  496800.0 462000.0 507000.0 448200.0 ;
      RECT  496800.0 462000.0 507000.0 475800.0 ;
      RECT  496800.0 489600.0 507000.0 475800.0 ;
      RECT  496800.0 489600.0 507000.0 503400.0 ;
      RECT  496800.0 517200.0 507000.0 503400.0 ;
      RECT  496800.0 517200.0 507000.0 531000.0 ;
      RECT  496800.0 544800.0 507000.0 531000.0 ;
      RECT  496800.0 544800.0 507000.0 558600.0 ;
      RECT  496800.0 572400.0 507000.0 558600.0 ;
      RECT  496800.0 572400.0 507000.0 586200.0 ;
      RECT  496800.0 600000.0 507000.0 586200.0 ;
      RECT  496800.0 600000.0 507000.0 613800.0 ;
      RECT  496800.0 627600.0 507000.0 613800.0 ;
      RECT  496800.0 627600.0 507000.0 641400.0 ;
      RECT  496800.0 655200.0 507000.0 641400.0 ;
      RECT  496800.0 655200.0 507000.0 669000.0 ;
      RECT  496800.0 682800.0 507000.0 669000.0 ;
      RECT  496800.0 682800.0 507000.0 696600.0 ;
      RECT  496800.0 710400.0 507000.0 696600.0 ;
      RECT  496800.0 710400.0 507000.0 724200.0 ;
      RECT  496800.0 738000.0 507000.0 724200.0 ;
      RECT  496800.0 738000.0 507000.0 751800.0 ;
      RECT  496800.0 765600.0 507000.0 751800.0 ;
      RECT  496800.0 765600.0 507000.0 779400.0 ;
      RECT  496800.0 793200.0 507000.0 779400.0 ;
      RECT  496800.0 793200.0 507000.0 807000.0 ;
      RECT  496800.0 820800.0 507000.0 807000.0 ;
      RECT  496800.0 820800.0 507000.0 834600.0 ;
      RECT  496800.0 848400.0 507000.0 834600.0 ;
      RECT  496800.0 848400.0 507000.0 862200.0 ;
      RECT  496800.0 876000.0 507000.0 862200.0 ;
      RECT  496800.0 876000.0 507000.0 889800.0 ;
      RECT  496800.0 903600.0 507000.0 889800.0 ;
      RECT  496800.0 903600.0 507000.0 917400.0 ;
      RECT  496800.0 931200.0 507000.0 917400.0 ;
      RECT  496800.0 931200.0 507000.0 945000.0 ;
      RECT  496800.0 958800.0 507000.0 945000.0 ;
      RECT  496800.0 958800.0 507000.0 972600.0 ;
      RECT  496800.0 986400.0 507000.0 972600.0 ;
      RECT  496800.0 986400.0 507000.0 1000200.0 ;
      RECT  496800.0 1014000.0 507000.0 1000200.0 ;
      RECT  496800.0 1014000.0 507000.0 1027800.0 ;
      RECT  496800.0 1041600.0 507000.0 1027800.0 ;
      RECT  496800.0 1041600.0 507000.0 1055400.0 ;
      RECT  496800.0 1069200.0 507000.0 1055400.0 ;
      RECT  496800.0 1069200.0 507000.0 1083000.0 ;
      RECT  496800.0 1096800.0 507000.0 1083000.0 ;
      RECT  496800.0 1096800.0 507000.0 1110600.0 ;
      RECT  496800.0 1124400.0 507000.0 1110600.0 ;
      RECT  496800.0 1124400.0 507000.0 1138200.0 ;
      RECT  496800.0 1152000.0 507000.0 1138200.0 ;
      RECT  496800.0 1152000.0 507000.0 1165800.0 ;
      RECT  496800.0 1179600.0 507000.0 1165800.0 ;
      RECT  496800.0 1179600.0 507000.0 1193400.0 ;
      RECT  496800.0 1207200.0 507000.0 1193400.0 ;
      RECT  496800.0 1207200.0 507000.0 1221000.0 ;
      RECT  496800.0 1234800.0 507000.0 1221000.0 ;
      RECT  496800.0 1234800.0 507000.0 1248600.0 ;
      RECT  496800.0 1262400.0 507000.0 1248600.0 ;
      RECT  496800.0 1262400.0 507000.0 1276200.0 ;
      RECT  496800.0 1290000.0 507000.0 1276200.0 ;
      RECT  496800.0 1290000.0 507000.0 1303800.0 ;
      RECT  496800.0 1317600.0 507000.0 1303800.0 ;
      RECT  496800.0 1317600.0 507000.0 1331400.0 ;
      RECT  496800.0 1345200.0 507000.0 1331400.0 ;
      RECT  496800.0 1345200.0 507000.0 1359000.0 ;
      RECT  496800.0 1372800.0 507000.0 1359000.0 ;
      RECT  496800.0 1372800.0 507000.0 1386600.0 ;
      RECT  496800.0 1400400.0 507000.0 1386600.0 ;
      RECT  496800.0 1400400.0 507000.0 1414200.0 ;
      RECT  496800.0 1428000.0 507000.0 1414200.0 ;
      RECT  496800.0 1428000.0 507000.0 1441800.0 ;
      RECT  496800.0 1455600.0 507000.0 1441800.0 ;
      RECT  496800.0 1455600.0 507000.0 1469400.0 ;
      RECT  496800.0 1483200.0 507000.0 1469400.0 ;
      RECT  496800.0 1483200.0 507000.0 1497000.0 ;
      RECT  496800.0 1510800.0 507000.0 1497000.0 ;
      RECT  496800.0 1510800.0 507000.0 1524600.0 ;
      RECT  496800.0 1538400.0 507000.0 1524600.0 ;
      RECT  496800.0 1538400.0 507000.0 1552200.0 ;
      RECT  496800.0 1566000.0 507000.0 1552200.0 ;
      RECT  496800.0 1566000.0 507000.0 1579800.0 ;
      RECT  496800.0 1593600.0 507000.0 1579800.0 ;
      RECT  496800.0 1593600.0 507000.0 1607400.0 ;
      RECT  496800.0 1621200.0 507000.0 1607400.0 ;
      RECT  496800.0 1621200.0 507000.0 1635000.0 ;
      RECT  496800.0 1648800.0 507000.0 1635000.0 ;
      RECT  496800.0 1648800.0 507000.0 1662600.0 ;
      RECT  496800.0 1676400.0 507000.0 1662600.0 ;
      RECT  496800.0 1676400.0 507000.0 1690200.0 ;
      RECT  496800.0 1704000.0 507000.0 1690200.0 ;
      RECT  496800.0 1704000.0 507000.0 1717800.0 ;
      RECT  496800.0 1731600.0 507000.0 1717800.0 ;
      RECT  496800.0 1731600.0 507000.0 1745400.0 ;
      RECT  496800.0 1759200.0 507000.0 1745400.0 ;
      RECT  496800.0 1759200.0 507000.0 1773000.0 ;
      RECT  496800.0 1786800.0 507000.0 1773000.0 ;
      RECT  496800.0 1786800.0 507000.0 1800600.0 ;
      RECT  496800.0 1814400.0 507000.0 1800600.0 ;
      RECT  496800.0 1814400.0 507000.0 1828200.0 ;
      RECT  496800.0 1842000.0 507000.0 1828200.0 ;
      RECT  496800.0 1842000.0 507000.0 1855800.0 ;
      RECT  496800.0 1869600.0 507000.0 1855800.0 ;
      RECT  496800.0 1869600.0 507000.0 1883400.0 ;
      RECT  496800.0 1897200.0 507000.0 1883400.0 ;
      RECT  496800.0 1897200.0 507000.0 1911000.0 ;
      RECT  496800.0 1924800.0 507000.0 1911000.0 ;
      RECT  496800.0 1924800.0 507000.0 1938600.0 ;
      RECT  496800.0 1952400.0 507000.0 1938600.0 ;
      RECT  496800.0 1952400.0 507000.0 1966200.0 ;
      RECT  496800.0 1980000.0 507000.0 1966200.0 ;
      RECT  496800.0 1980000.0 507000.0 1993800.0 ;
      RECT  496800.0 2007600.0 507000.0 1993800.0 ;
      RECT  496800.0 2007600.0 507000.0 2021400.0 ;
      RECT  496800.0 2035200.0 507000.0 2021400.0 ;
      RECT  496800.0 2035200.0 507000.0 2049000.0 ;
      RECT  496800.0 2062800.0 507000.0 2049000.0 ;
      RECT  496800.0 2062800.0 507000.0 2076600.0 ;
      RECT  496800.0 2090400.0 507000.0 2076600.0 ;
      RECT  496800.0 2090400.0 507000.0 2104200.0 ;
      RECT  496800.0 2118000.0 507000.0 2104200.0 ;
      RECT  496800.0 2118000.0 507000.0 2131800.0 ;
      RECT  496800.0 2145600.0 507000.0 2131800.0 ;
      RECT  507000.0 379200.0 517200.0 393000.0 ;
      RECT  507000.0 406800.0 517200.0 393000.0 ;
      RECT  507000.0 406800.0 517200.0 420600.0 ;
      RECT  507000.0 434400.0 517200.0 420600.0 ;
      RECT  507000.0 434400.0 517200.0 448200.0 ;
      RECT  507000.0 462000.0 517200.0 448200.0 ;
      RECT  507000.0 462000.0 517200.0 475800.0 ;
      RECT  507000.0 489600.0 517200.0 475800.0 ;
      RECT  507000.0 489600.0 517200.0 503400.0 ;
      RECT  507000.0 517200.0 517200.0 503400.0 ;
      RECT  507000.0 517200.0 517200.0 531000.0 ;
      RECT  507000.0 544800.0 517200.0 531000.0 ;
      RECT  507000.0 544800.0 517200.0 558600.0 ;
      RECT  507000.0 572400.0 517200.0 558600.0 ;
      RECT  507000.0 572400.0 517200.0 586200.0 ;
      RECT  507000.0 600000.0 517200.0 586200.0 ;
      RECT  507000.0 600000.0 517200.0 613800.0 ;
      RECT  507000.0 627600.0 517200.0 613800.0 ;
      RECT  507000.0 627600.0 517200.0 641400.0 ;
      RECT  507000.0 655200.0 517200.0 641400.0 ;
      RECT  507000.0 655200.0 517200.0 669000.0 ;
      RECT  507000.0 682800.0 517200.0 669000.0 ;
      RECT  507000.0 682800.0 517200.0 696600.0 ;
      RECT  507000.0 710400.0 517200.0 696600.0 ;
      RECT  507000.0 710400.0 517200.0 724200.0 ;
      RECT  507000.0 738000.0 517200.0 724200.0 ;
      RECT  507000.0 738000.0 517200.0 751800.0 ;
      RECT  507000.0 765600.0 517200.0 751800.0 ;
      RECT  507000.0 765600.0 517200.0 779400.0 ;
      RECT  507000.0 793200.0 517200.0 779400.0 ;
      RECT  507000.0 793200.0 517200.0 807000.0 ;
      RECT  507000.0 820800.0 517200.0 807000.0 ;
      RECT  507000.0 820800.0 517200.0 834600.0 ;
      RECT  507000.0 848400.0 517200.0 834600.0 ;
      RECT  507000.0 848400.0 517200.0 862200.0 ;
      RECT  507000.0 876000.0 517200.0 862200.0 ;
      RECT  507000.0 876000.0 517200.0 889800.0 ;
      RECT  507000.0 903600.0 517200.0 889800.0 ;
      RECT  507000.0 903600.0 517200.0 917400.0 ;
      RECT  507000.0 931200.0 517200.0 917400.0 ;
      RECT  507000.0 931200.0 517200.0 945000.0 ;
      RECT  507000.0 958800.0 517200.0 945000.0 ;
      RECT  507000.0 958800.0 517200.0 972600.0 ;
      RECT  507000.0 986400.0 517200.0 972600.0 ;
      RECT  507000.0 986400.0 517200.0 1000200.0 ;
      RECT  507000.0 1014000.0 517200.0 1000200.0 ;
      RECT  507000.0 1014000.0 517200.0 1027800.0 ;
      RECT  507000.0 1041600.0 517200.0 1027800.0 ;
      RECT  507000.0 1041600.0 517200.0 1055400.0 ;
      RECT  507000.0 1069200.0 517200.0 1055400.0 ;
      RECT  507000.0 1069200.0 517200.0 1083000.0 ;
      RECT  507000.0 1096800.0 517200.0 1083000.0 ;
      RECT  507000.0 1096800.0 517200.0 1110600.0 ;
      RECT  507000.0 1124400.0 517200.0 1110600.0 ;
      RECT  507000.0 1124400.0 517200.0 1138200.0 ;
      RECT  507000.0 1152000.0 517200.0 1138200.0 ;
      RECT  507000.0 1152000.0 517200.0 1165800.0 ;
      RECT  507000.0 1179600.0 517200.0 1165800.0 ;
      RECT  507000.0 1179600.0 517200.0 1193400.0 ;
      RECT  507000.0 1207200.0 517200.0 1193400.0 ;
      RECT  507000.0 1207200.0 517200.0 1221000.0 ;
      RECT  507000.0 1234800.0 517200.0 1221000.0 ;
      RECT  507000.0 1234800.0 517200.0 1248600.0 ;
      RECT  507000.0 1262400.0 517200.0 1248600.0 ;
      RECT  507000.0 1262400.0 517200.0 1276200.0 ;
      RECT  507000.0 1290000.0 517200.0 1276200.0 ;
      RECT  507000.0 1290000.0 517200.0 1303800.0 ;
      RECT  507000.0 1317600.0 517200.0 1303800.0 ;
      RECT  507000.0 1317600.0 517200.0 1331400.0 ;
      RECT  507000.0 1345200.0 517200.0 1331400.0 ;
      RECT  507000.0 1345200.0 517200.0 1359000.0 ;
      RECT  507000.0 1372800.0 517200.0 1359000.0 ;
      RECT  507000.0 1372800.0 517200.0 1386600.0 ;
      RECT  507000.0 1400400.0 517200.0 1386600.0 ;
      RECT  507000.0 1400400.0 517200.0 1414200.0 ;
      RECT  507000.0 1428000.0 517200.0 1414200.0 ;
      RECT  507000.0 1428000.0 517200.0 1441800.0 ;
      RECT  507000.0 1455600.0 517200.0 1441800.0 ;
      RECT  507000.0 1455600.0 517200.0 1469400.0 ;
      RECT  507000.0 1483200.0 517200.0 1469400.0 ;
      RECT  507000.0 1483200.0 517200.0 1497000.0 ;
      RECT  507000.0 1510800.0 517200.0 1497000.0 ;
      RECT  507000.0 1510800.0 517200.0 1524600.0 ;
      RECT  507000.0 1538400.0 517200.0 1524600.0 ;
      RECT  507000.0 1538400.0 517200.0 1552200.0 ;
      RECT  507000.0 1566000.0 517200.0 1552200.0 ;
      RECT  507000.0 1566000.0 517200.0 1579800.0 ;
      RECT  507000.0 1593600.0 517200.0 1579800.0 ;
      RECT  507000.0 1593600.0 517200.0 1607400.0 ;
      RECT  507000.0 1621200.0 517200.0 1607400.0 ;
      RECT  507000.0 1621200.0 517200.0 1635000.0 ;
      RECT  507000.0 1648800.0 517200.0 1635000.0 ;
      RECT  507000.0 1648800.0 517200.0 1662600.0 ;
      RECT  507000.0 1676400.0 517200.0 1662600.0 ;
      RECT  507000.0 1676400.0 517200.0 1690200.0 ;
      RECT  507000.0 1704000.0 517200.0 1690200.0 ;
      RECT  507000.0 1704000.0 517200.0 1717800.0 ;
      RECT  507000.0 1731600.0 517200.0 1717800.0 ;
      RECT  507000.0 1731600.0 517200.0 1745400.0 ;
      RECT  507000.0 1759200.0 517200.0 1745400.0 ;
      RECT  507000.0 1759200.0 517200.0 1773000.0 ;
      RECT  507000.0 1786800.0 517200.0 1773000.0 ;
      RECT  507000.0 1786800.0 517200.0 1800600.0 ;
      RECT  507000.0 1814400.0 517200.0 1800600.0 ;
      RECT  507000.0 1814400.0 517200.0 1828200.0 ;
      RECT  507000.0 1842000.0 517200.0 1828200.0 ;
      RECT  507000.0 1842000.0 517200.0 1855800.0 ;
      RECT  507000.0 1869600.0 517200.0 1855800.0 ;
      RECT  507000.0 1869600.0 517200.0 1883400.0 ;
      RECT  507000.0 1897200.0 517200.0 1883400.0 ;
      RECT  507000.0 1897200.0 517200.0 1911000.0 ;
      RECT  507000.0 1924800.0 517200.0 1911000.0 ;
      RECT  507000.0 1924800.0 517200.0 1938600.0 ;
      RECT  507000.0 1952400.0 517200.0 1938600.0 ;
      RECT  507000.0 1952400.0 517200.0 1966200.0 ;
      RECT  507000.0 1980000.0 517200.0 1966200.0 ;
      RECT  507000.0 1980000.0 517200.0 1993800.0 ;
      RECT  507000.0 2007600.0 517200.0 1993800.0 ;
      RECT  507000.0 2007600.0 517200.0 2021400.0 ;
      RECT  507000.0 2035200.0 517200.0 2021400.0 ;
      RECT  507000.0 2035200.0 517200.0 2049000.0 ;
      RECT  507000.0 2062800.0 517200.0 2049000.0 ;
      RECT  507000.0 2062800.0 517200.0 2076600.0 ;
      RECT  507000.0 2090400.0 517200.0 2076600.0 ;
      RECT  507000.0 2090400.0 517200.0 2104200.0 ;
      RECT  507000.0 2118000.0 517200.0 2104200.0 ;
      RECT  507000.0 2118000.0 517200.0 2131800.0 ;
      RECT  507000.0 2145600.0 517200.0 2131800.0 ;
      RECT  517200.0 379200.0 527400.0 393000.0 ;
      RECT  517200.0 406800.0 527400.0 393000.0 ;
      RECT  517200.0 406800.0 527400.0 420600.0 ;
      RECT  517200.0 434400.0 527400.0 420600.0 ;
      RECT  517200.0 434400.0 527400.0 448200.0 ;
      RECT  517200.0 462000.0 527400.0 448200.0 ;
      RECT  517200.0 462000.0 527400.0 475800.0 ;
      RECT  517200.0 489600.0 527400.0 475800.0 ;
      RECT  517200.0 489600.0 527400.0 503400.0 ;
      RECT  517200.0 517200.0 527400.0 503400.0 ;
      RECT  517200.0 517200.0 527400.0 531000.0 ;
      RECT  517200.0 544800.0 527400.0 531000.0 ;
      RECT  517200.0 544800.0 527400.0 558600.0 ;
      RECT  517200.0 572400.0 527400.0 558600.0 ;
      RECT  517200.0 572400.0 527400.0 586200.0 ;
      RECT  517200.0 600000.0 527400.0 586200.0 ;
      RECT  517200.0 600000.0 527400.0 613800.0 ;
      RECT  517200.0 627600.0 527400.0 613800.0 ;
      RECT  517200.0 627600.0 527400.0 641400.0 ;
      RECT  517200.0 655200.0 527400.0 641400.0 ;
      RECT  517200.0 655200.0 527400.0 669000.0 ;
      RECT  517200.0 682800.0 527400.0 669000.0 ;
      RECT  517200.0 682800.0 527400.0 696600.0 ;
      RECT  517200.0 710400.0 527400.0 696600.0 ;
      RECT  517200.0 710400.0 527400.0 724200.0 ;
      RECT  517200.0 738000.0 527400.0 724200.0 ;
      RECT  517200.0 738000.0 527400.0 751800.0 ;
      RECT  517200.0 765600.0 527400.0 751800.0 ;
      RECT  517200.0 765600.0 527400.0 779400.0 ;
      RECT  517200.0 793200.0 527400.0 779400.0 ;
      RECT  517200.0 793200.0 527400.0 807000.0 ;
      RECT  517200.0 820800.0 527400.0 807000.0 ;
      RECT  517200.0 820800.0 527400.0 834600.0 ;
      RECT  517200.0 848400.0 527400.0 834600.0 ;
      RECT  517200.0 848400.0 527400.0 862200.0 ;
      RECT  517200.0 876000.0 527400.0 862200.0 ;
      RECT  517200.0 876000.0 527400.0 889800.0 ;
      RECT  517200.0 903600.0 527400.0 889800.0 ;
      RECT  517200.0 903600.0 527400.0 917400.0 ;
      RECT  517200.0 931200.0 527400.0 917400.0 ;
      RECT  517200.0 931200.0 527400.0 945000.0 ;
      RECT  517200.0 958800.0 527400.0 945000.0 ;
      RECT  517200.0 958800.0 527400.0 972600.0 ;
      RECT  517200.0 986400.0 527400.0 972600.0 ;
      RECT  517200.0 986400.0 527400.0 1000200.0 ;
      RECT  517200.0 1014000.0 527400.0 1000200.0 ;
      RECT  517200.0 1014000.0 527400.0 1027800.0 ;
      RECT  517200.0 1041600.0 527400.0 1027800.0 ;
      RECT  517200.0 1041600.0 527400.0 1055400.0 ;
      RECT  517200.0 1069200.0 527400.0 1055400.0 ;
      RECT  517200.0 1069200.0 527400.0 1083000.0 ;
      RECT  517200.0 1096800.0 527400.0 1083000.0 ;
      RECT  517200.0 1096800.0 527400.0 1110600.0 ;
      RECT  517200.0 1124400.0 527400.0 1110600.0 ;
      RECT  517200.0 1124400.0 527400.0 1138200.0 ;
      RECT  517200.0 1152000.0 527400.0 1138200.0 ;
      RECT  517200.0 1152000.0 527400.0 1165800.0 ;
      RECT  517200.0 1179600.0 527400.0 1165800.0 ;
      RECT  517200.0 1179600.0 527400.0 1193400.0 ;
      RECT  517200.0 1207200.0 527400.0 1193400.0 ;
      RECT  517200.0 1207200.0 527400.0 1221000.0 ;
      RECT  517200.0 1234800.0 527400.0 1221000.0 ;
      RECT  517200.0 1234800.0 527400.0 1248600.0 ;
      RECT  517200.0 1262400.0 527400.0 1248600.0 ;
      RECT  517200.0 1262400.0 527400.0 1276200.0 ;
      RECT  517200.0 1290000.0 527400.0 1276200.0 ;
      RECT  517200.0 1290000.0 527400.0 1303800.0 ;
      RECT  517200.0 1317600.0 527400.0 1303800.0 ;
      RECT  517200.0 1317600.0 527400.0 1331400.0 ;
      RECT  517200.0 1345200.0 527400.0 1331400.0 ;
      RECT  517200.0 1345200.0 527400.0 1359000.0 ;
      RECT  517200.0 1372800.0 527400.0 1359000.0 ;
      RECT  517200.0 1372800.0 527400.0 1386600.0 ;
      RECT  517200.0 1400400.0 527400.0 1386600.0 ;
      RECT  517200.0 1400400.0 527400.0 1414200.0 ;
      RECT  517200.0 1428000.0 527400.0 1414200.0 ;
      RECT  517200.0 1428000.0 527400.0 1441800.0 ;
      RECT  517200.0 1455600.0 527400.0 1441800.0 ;
      RECT  517200.0 1455600.0 527400.0 1469400.0 ;
      RECT  517200.0 1483200.0 527400.0 1469400.0 ;
      RECT  517200.0 1483200.0 527400.0 1497000.0 ;
      RECT  517200.0 1510800.0 527400.0 1497000.0 ;
      RECT  517200.0 1510800.0 527400.0 1524600.0 ;
      RECT  517200.0 1538400.0 527400.0 1524600.0 ;
      RECT  517200.0 1538400.0 527400.0 1552200.0 ;
      RECT  517200.0 1566000.0 527400.0 1552200.0 ;
      RECT  517200.0 1566000.0 527400.0 1579800.0 ;
      RECT  517200.0 1593600.0 527400.0 1579800.0 ;
      RECT  517200.0 1593600.0 527400.0 1607400.0 ;
      RECT  517200.0 1621200.0 527400.0 1607400.0 ;
      RECT  517200.0 1621200.0 527400.0 1635000.0 ;
      RECT  517200.0 1648800.0 527400.0 1635000.0 ;
      RECT  517200.0 1648800.0 527400.0 1662600.0 ;
      RECT  517200.0 1676400.0 527400.0 1662600.0 ;
      RECT  517200.0 1676400.0 527400.0 1690200.0 ;
      RECT  517200.0 1704000.0 527400.0 1690200.0 ;
      RECT  517200.0 1704000.0 527400.0 1717800.0 ;
      RECT  517200.0 1731600.0 527400.0 1717800.0 ;
      RECT  517200.0 1731600.0 527400.0 1745400.0 ;
      RECT  517200.0 1759200.0 527400.0 1745400.0 ;
      RECT  517200.0 1759200.0 527400.0 1773000.0 ;
      RECT  517200.0 1786800.0 527400.0 1773000.0 ;
      RECT  517200.0 1786800.0 527400.0 1800600.0 ;
      RECT  517200.0 1814400.0 527400.0 1800600.0 ;
      RECT  517200.0 1814400.0 527400.0 1828200.0 ;
      RECT  517200.0 1842000.0 527400.0 1828200.0 ;
      RECT  517200.0 1842000.0 527400.0 1855800.0 ;
      RECT  517200.0 1869600.0 527400.0 1855800.0 ;
      RECT  517200.0 1869600.0 527400.0 1883400.0 ;
      RECT  517200.0 1897200.0 527400.0 1883400.0 ;
      RECT  517200.0 1897200.0 527400.0 1911000.0 ;
      RECT  517200.0 1924800.0 527400.0 1911000.0 ;
      RECT  517200.0 1924800.0 527400.0 1938600.0 ;
      RECT  517200.0 1952400.0 527400.0 1938600.0 ;
      RECT  517200.0 1952400.0 527400.0 1966200.0 ;
      RECT  517200.0 1980000.0 527400.0 1966200.0 ;
      RECT  517200.0 1980000.0 527400.0 1993800.0 ;
      RECT  517200.0 2007600.0 527400.0 1993800.0 ;
      RECT  517200.0 2007600.0 527400.0 2021400.0 ;
      RECT  517200.0 2035200.0 527400.0 2021400.0 ;
      RECT  517200.0 2035200.0 527400.0 2049000.0 ;
      RECT  517200.0 2062800.0 527400.0 2049000.0 ;
      RECT  517200.0 2062800.0 527400.0 2076600.0 ;
      RECT  517200.0 2090400.0 527400.0 2076600.0 ;
      RECT  517200.0 2090400.0 527400.0 2104200.0 ;
      RECT  517200.0 2118000.0 527400.0 2104200.0 ;
      RECT  517200.0 2118000.0 527400.0 2131800.0 ;
      RECT  517200.0 2145600.0 527400.0 2131800.0 ;
      RECT  527400.0 379200.0 537600.0 393000.0 ;
      RECT  527400.0 406800.0 537600.0 393000.0 ;
      RECT  527400.0 406800.0 537600.0 420600.0 ;
      RECT  527400.0 434400.0 537600.0 420600.0 ;
      RECT  527400.0 434400.0 537600.0 448200.0 ;
      RECT  527400.0 462000.0 537600.0 448200.0 ;
      RECT  527400.0 462000.0 537600.0 475800.0 ;
      RECT  527400.0 489600.0 537600.0 475800.0 ;
      RECT  527400.0 489600.0 537600.0 503400.0 ;
      RECT  527400.0 517200.0 537600.0 503400.0 ;
      RECT  527400.0 517200.0 537600.0 531000.0 ;
      RECT  527400.0 544800.0 537600.0 531000.0 ;
      RECT  527400.0 544800.0 537600.0 558600.0 ;
      RECT  527400.0 572400.0 537600.0 558600.0 ;
      RECT  527400.0 572400.0 537600.0 586200.0 ;
      RECT  527400.0 600000.0 537600.0 586200.0 ;
      RECT  527400.0 600000.0 537600.0 613800.0 ;
      RECT  527400.0 627600.0 537600.0 613800.0 ;
      RECT  527400.0 627600.0 537600.0 641400.0 ;
      RECT  527400.0 655200.0 537600.0 641400.0 ;
      RECT  527400.0 655200.0 537600.0 669000.0 ;
      RECT  527400.0 682800.0 537600.0 669000.0 ;
      RECT  527400.0 682800.0 537600.0 696600.0 ;
      RECT  527400.0 710400.0 537600.0 696600.0 ;
      RECT  527400.0 710400.0 537600.0 724200.0 ;
      RECT  527400.0 738000.0 537600.0 724200.0 ;
      RECT  527400.0 738000.0 537600.0 751800.0 ;
      RECT  527400.0 765600.0 537600.0 751800.0 ;
      RECT  527400.0 765600.0 537600.0 779400.0 ;
      RECT  527400.0 793200.0 537600.0 779400.0 ;
      RECT  527400.0 793200.0 537600.0 807000.0 ;
      RECT  527400.0 820800.0 537600.0 807000.0 ;
      RECT  527400.0 820800.0 537600.0 834600.0 ;
      RECT  527400.0 848400.0 537600.0 834600.0 ;
      RECT  527400.0 848400.0 537600.0 862200.0 ;
      RECT  527400.0 876000.0 537600.0 862200.0 ;
      RECT  527400.0 876000.0 537600.0 889800.0 ;
      RECT  527400.0 903600.0 537600.0 889800.0 ;
      RECT  527400.0 903600.0 537600.0 917400.0 ;
      RECT  527400.0 931200.0 537600.0 917400.0 ;
      RECT  527400.0 931200.0 537600.0 945000.0 ;
      RECT  527400.0 958800.0 537600.0 945000.0 ;
      RECT  527400.0 958800.0 537600.0 972600.0 ;
      RECT  527400.0 986400.0 537600.0 972600.0 ;
      RECT  527400.0 986400.0 537600.0 1000200.0 ;
      RECT  527400.0 1014000.0 537600.0 1000200.0 ;
      RECT  527400.0 1014000.0 537600.0 1027800.0 ;
      RECT  527400.0 1041600.0 537600.0 1027800.0 ;
      RECT  527400.0 1041600.0 537600.0 1055400.0 ;
      RECT  527400.0 1069200.0 537600.0 1055400.0 ;
      RECT  527400.0 1069200.0 537600.0 1083000.0 ;
      RECT  527400.0 1096800.0 537600.0 1083000.0 ;
      RECT  527400.0 1096800.0 537600.0 1110600.0 ;
      RECT  527400.0 1124400.0 537600.0 1110600.0 ;
      RECT  527400.0 1124400.0 537600.0 1138200.0 ;
      RECT  527400.0 1152000.0 537600.0 1138200.0 ;
      RECT  527400.0 1152000.0 537600.0 1165800.0 ;
      RECT  527400.0 1179600.0 537600.0 1165800.0 ;
      RECT  527400.0 1179600.0 537600.0 1193400.0 ;
      RECT  527400.0 1207200.0 537600.0 1193400.0 ;
      RECT  527400.0 1207200.0 537600.0 1221000.0 ;
      RECT  527400.0 1234800.0 537600.0 1221000.0 ;
      RECT  527400.0 1234800.0 537600.0 1248600.0 ;
      RECT  527400.0 1262400.0 537600.0 1248600.0 ;
      RECT  527400.0 1262400.0 537600.0 1276200.0 ;
      RECT  527400.0 1290000.0 537600.0 1276200.0 ;
      RECT  527400.0 1290000.0 537600.0 1303800.0 ;
      RECT  527400.0 1317600.0 537600.0 1303800.0 ;
      RECT  527400.0 1317600.0 537600.0 1331400.0 ;
      RECT  527400.0 1345200.0 537600.0 1331400.0 ;
      RECT  527400.0 1345200.0 537600.0 1359000.0 ;
      RECT  527400.0 1372800.0 537600.0 1359000.0 ;
      RECT  527400.0 1372800.0 537600.0 1386600.0 ;
      RECT  527400.0 1400400.0 537600.0 1386600.0 ;
      RECT  527400.0 1400400.0 537600.0 1414200.0 ;
      RECT  527400.0 1428000.0 537600.0 1414200.0 ;
      RECT  527400.0 1428000.0 537600.0 1441800.0 ;
      RECT  527400.0 1455600.0 537600.0 1441800.0 ;
      RECT  527400.0 1455600.0 537600.0 1469400.0 ;
      RECT  527400.0 1483200.0 537600.0 1469400.0 ;
      RECT  527400.0 1483200.0 537600.0 1497000.0 ;
      RECT  527400.0 1510800.0 537600.0 1497000.0 ;
      RECT  527400.0 1510800.0 537600.0 1524600.0 ;
      RECT  527400.0 1538400.0 537600.0 1524600.0 ;
      RECT  527400.0 1538400.0 537600.0 1552200.0 ;
      RECT  527400.0 1566000.0 537600.0 1552200.0 ;
      RECT  527400.0 1566000.0 537600.0 1579800.0 ;
      RECT  527400.0 1593600.0 537600.0 1579800.0 ;
      RECT  527400.0 1593600.0 537600.0 1607400.0 ;
      RECT  527400.0 1621200.0 537600.0 1607400.0 ;
      RECT  527400.0 1621200.0 537600.0 1635000.0 ;
      RECT  527400.0 1648800.0 537600.0 1635000.0 ;
      RECT  527400.0 1648800.0 537600.0 1662600.0 ;
      RECT  527400.0 1676400.0 537600.0 1662600.0 ;
      RECT  527400.0 1676400.0 537600.0 1690200.0 ;
      RECT  527400.0 1704000.0 537600.0 1690200.0 ;
      RECT  527400.0 1704000.0 537600.0 1717800.0 ;
      RECT  527400.0 1731600.0 537600.0 1717800.0 ;
      RECT  527400.0 1731600.0 537600.0 1745400.0 ;
      RECT  527400.0 1759200.0 537600.0 1745400.0 ;
      RECT  527400.0 1759200.0 537600.0 1773000.0 ;
      RECT  527400.0 1786800.0 537600.0 1773000.0 ;
      RECT  527400.0 1786800.0 537600.0 1800600.0 ;
      RECT  527400.0 1814400.0 537600.0 1800600.0 ;
      RECT  527400.0 1814400.0 537600.0 1828200.0 ;
      RECT  527400.0 1842000.0 537600.0 1828200.0 ;
      RECT  527400.0 1842000.0 537600.0 1855800.0 ;
      RECT  527400.0 1869600.0 537600.0 1855800.0 ;
      RECT  527400.0 1869600.0 537600.0 1883400.0 ;
      RECT  527400.0 1897200.0 537600.0 1883400.0 ;
      RECT  527400.0 1897200.0 537600.0 1911000.0 ;
      RECT  527400.0 1924800.0 537600.0 1911000.0 ;
      RECT  527400.0 1924800.0 537600.0 1938600.0 ;
      RECT  527400.0 1952400.0 537600.0 1938600.0 ;
      RECT  527400.0 1952400.0 537600.0 1966200.0 ;
      RECT  527400.0 1980000.0 537600.0 1966200.0 ;
      RECT  527400.0 1980000.0 537600.0 1993800.0 ;
      RECT  527400.0 2007600.0 537600.0 1993800.0 ;
      RECT  527400.0 2007600.0 537600.0 2021400.0 ;
      RECT  527400.0 2035200.0 537600.0 2021400.0 ;
      RECT  527400.0 2035200.0 537600.0 2049000.0 ;
      RECT  527400.0 2062800.0 537600.0 2049000.0 ;
      RECT  527400.0 2062800.0 537600.0 2076600.0 ;
      RECT  527400.0 2090400.0 537600.0 2076600.0 ;
      RECT  527400.0 2090400.0 537600.0 2104200.0 ;
      RECT  527400.0 2118000.0 537600.0 2104200.0 ;
      RECT  527400.0 2118000.0 537600.0 2131800.0 ;
      RECT  527400.0 2145600.0 537600.0 2131800.0 ;
      RECT  537600.0 379200.0 547800.0 393000.0 ;
      RECT  537600.0 406800.0 547800.0 393000.0 ;
      RECT  537600.0 406800.0 547800.0 420600.0 ;
      RECT  537600.0 434400.0 547800.0 420600.0 ;
      RECT  537600.0 434400.0 547800.0 448200.0 ;
      RECT  537600.0 462000.0 547800.0 448200.0 ;
      RECT  537600.0 462000.0 547800.0 475800.0 ;
      RECT  537600.0 489600.0 547800.0 475800.0 ;
      RECT  537600.0 489600.0 547800.0 503400.0 ;
      RECT  537600.0 517200.0 547800.0 503400.0 ;
      RECT  537600.0 517200.0 547800.0 531000.0 ;
      RECT  537600.0 544800.0 547800.0 531000.0 ;
      RECT  537600.0 544800.0 547800.0 558600.0 ;
      RECT  537600.0 572400.0 547800.0 558600.0 ;
      RECT  537600.0 572400.0 547800.0 586200.0 ;
      RECT  537600.0 600000.0 547800.0 586200.0 ;
      RECT  537600.0 600000.0 547800.0 613800.0 ;
      RECT  537600.0 627600.0 547800.0 613800.0 ;
      RECT  537600.0 627600.0 547800.0 641400.0 ;
      RECT  537600.0 655200.0 547800.0 641400.0 ;
      RECT  537600.0 655200.0 547800.0 669000.0 ;
      RECT  537600.0 682800.0 547800.0 669000.0 ;
      RECT  537600.0 682800.0 547800.0 696600.0 ;
      RECT  537600.0 710400.0 547800.0 696600.0 ;
      RECT  537600.0 710400.0 547800.0 724200.0 ;
      RECT  537600.0 738000.0 547800.0 724200.0 ;
      RECT  537600.0 738000.0 547800.0 751800.0 ;
      RECT  537600.0 765600.0 547800.0 751800.0 ;
      RECT  537600.0 765600.0 547800.0 779400.0 ;
      RECT  537600.0 793200.0 547800.0 779400.0 ;
      RECT  537600.0 793200.0 547800.0 807000.0 ;
      RECT  537600.0 820800.0 547800.0 807000.0 ;
      RECT  537600.0 820800.0 547800.0 834600.0 ;
      RECT  537600.0 848400.0 547800.0 834600.0 ;
      RECT  537600.0 848400.0 547800.0 862200.0 ;
      RECT  537600.0 876000.0 547800.0 862200.0 ;
      RECT  537600.0 876000.0 547800.0 889800.0 ;
      RECT  537600.0 903600.0 547800.0 889800.0 ;
      RECT  537600.0 903600.0 547800.0 917400.0 ;
      RECT  537600.0 931200.0 547800.0 917400.0 ;
      RECT  537600.0 931200.0 547800.0 945000.0 ;
      RECT  537600.0 958800.0 547800.0 945000.0 ;
      RECT  537600.0 958800.0 547800.0 972600.0 ;
      RECT  537600.0 986400.0 547800.0 972600.0 ;
      RECT  537600.0 986400.0 547800.0 1000200.0 ;
      RECT  537600.0 1014000.0 547800.0 1000200.0 ;
      RECT  537600.0 1014000.0 547800.0 1027800.0 ;
      RECT  537600.0 1041600.0 547800.0 1027800.0 ;
      RECT  537600.0 1041600.0 547800.0 1055400.0 ;
      RECT  537600.0 1069200.0 547800.0 1055400.0 ;
      RECT  537600.0 1069200.0 547800.0 1083000.0 ;
      RECT  537600.0 1096800.0 547800.0 1083000.0 ;
      RECT  537600.0 1096800.0 547800.0 1110600.0 ;
      RECT  537600.0 1124400.0 547800.0 1110600.0 ;
      RECT  537600.0 1124400.0 547800.0 1138200.0 ;
      RECT  537600.0 1152000.0 547800.0 1138200.0 ;
      RECT  537600.0 1152000.0 547800.0 1165800.0 ;
      RECT  537600.0 1179600.0 547800.0 1165800.0 ;
      RECT  537600.0 1179600.0 547800.0 1193400.0 ;
      RECT  537600.0 1207200.0 547800.0 1193400.0 ;
      RECT  537600.0 1207200.0 547800.0 1221000.0 ;
      RECT  537600.0 1234800.0 547800.0 1221000.0 ;
      RECT  537600.0 1234800.0 547800.0 1248600.0 ;
      RECT  537600.0 1262400.0 547800.0 1248600.0 ;
      RECT  537600.0 1262400.0 547800.0 1276200.0 ;
      RECT  537600.0 1290000.0 547800.0 1276200.0 ;
      RECT  537600.0 1290000.0 547800.0 1303800.0 ;
      RECT  537600.0 1317600.0 547800.0 1303800.0 ;
      RECT  537600.0 1317600.0 547800.0 1331400.0 ;
      RECT  537600.0 1345200.0 547800.0 1331400.0 ;
      RECT  537600.0 1345200.0 547800.0 1359000.0 ;
      RECT  537600.0 1372800.0 547800.0 1359000.0 ;
      RECT  537600.0 1372800.0 547800.0 1386600.0 ;
      RECT  537600.0 1400400.0 547800.0 1386600.0 ;
      RECT  537600.0 1400400.0 547800.0 1414200.0 ;
      RECT  537600.0 1428000.0 547800.0 1414200.0 ;
      RECT  537600.0 1428000.0 547800.0 1441800.0 ;
      RECT  537600.0 1455600.0 547800.0 1441800.0 ;
      RECT  537600.0 1455600.0 547800.0 1469400.0 ;
      RECT  537600.0 1483200.0 547800.0 1469400.0 ;
      RECT  537600.0 1483200.0 547800.0 1497000.0 ;
      RECT  537600.0 1510800.0 547800.0 1497000.0 ;
      RECT  537600.0 1510800.0 547800.0 1524600.0 ;
      RECT  537600.0 1538400.0 547800.0 1524600.0 ;
      RECT  537600.0 1538400.0 547800.0 1552200.0 ;
      RECT  537600.0 1566000.0 547800.0 1552200.0 ;
      RECT  537600.0 1566000.0 547800.0 1579800.0 ;
      RECT  537600.0 1593600.0 547800.0 1579800.0 ;
      RECT  537600.0 1593600.0 547800.0 1607400.0 ;
      RECT  537600.0 1621200.0 547800.0 1607400.0 ;
      RECT  537600.0 1621200.0 547800.0 1635000.0 ;
      RECT  537600.0 1648800.0 547800.0 1635000.0 ;
      RECT  537600.0 1648800.0 547800.0 1662600.0 ;
      RECT  537600.0 1676400.0 547800.0 1662600.0 ;
      RECT  537600.0 1676400.0 547800.0 1690200.0 ;
      RECT  537600.0 1704000.0 547800.0 1690200.0 ;
      RECT  537600.0 1704000.0 547800.0 1717800.0 ;
      RECT  537600.0 1731600.0 547800.0 1717800.0 ;
      RECT  537600.0 1731600.0 547800.0 1745400.0 ;
      RECT  537600.0 1759200.0 547800.0 1745400.0 ;
      RECT  537600.0 1759200.0 547800.0 1773000.0 ;
      RECT  537600.0 1786800.0 547800.0 1773000.0 ;
      RECT  537600.0 1786800.0 547800.0 1800600.0 ;
      RECT  537600.0 1814400.0 547800.0 1800600.0 ;
      RECT  537600.0 1814400.0 547800.0 1828200.0 ;
      RECT  537600.0 1842000.0 547800.0 1828200.0 ;
      RECT  537600.0 1842000.0 547800.0 1855800.0 ;
      RECT  537600.0 1869600.0 547800.0 1855800.0 ;
      RECT  537600.0 1869600.0 547800.0 1883400.0 ;
      RECT  537600.0 1897200.0 547800.0 1883400.0 ;
      RECT  537600.0 1897200.0 547800.0 1911000.0 ;
      RECT  537600.0 1924800.0 547800.0 1911000.0 ;
      RECT  537600.0 1924800.0 547800.0 1938600.0 ;
      RECT  537600.0 1952400.0 547800.0 1938600.0 ;
      RECT  537600.0 1952400.0 547800.0 1966200.0 ;
      RECT  537600.0 1980000.0 547800.0 1966200.0 ;
      RECT  537600.0 1980000.0 547800.0 1993800.0 ;
      RECT  537600.0 2007600.0 547800.0 1993800.0 ;
      RECT  537600.0 2007600.0 547800.0 2021400.0 ;
      RECT  537600.0 2035200.0 547800.0 2021400.0 ;
      RECT  537600.0 2035200.0 547800.0 2049000.0 ;
      RECT  537600.0 2062800.0 547800.0 2049000.0 ;
      RECT  537600.0 2062800.0 547800.0 2076600.0 ;
      RECT  537600.0 2090400.0 547800.0 2076600.0 ;
      RECT  537600.0 2090400.0 547800.0 2104200.0 ;
      RECT  537600.0 2118000.0 547800.0 2104200.0 ;
      RECT  537600.0 2118000.0 547800.0 2131800.0 ;
      RECT  537600.0 2145600.0 547800.0 2131800.0 ;
      RECT  547800.0 379200.0 558000.0 393000.0 ;
      RECT  547800.0 406800.0 558000.0 393000.0 ;
      RECT  547800.0 406800.0 558000.0 420600.0 ;
      RECT  547800.0 434400.0 558000.0 420600.0 ;
      RECT  547800.0 434400.0 558000.0 448200.0 ;
      RECT  547800.0 462000.0 558000.0 448200.0 ;
      RECT  547800.0 462000.0 558000.0 475800.0 ;
      RECT  547800.0 489600.0 558000.0 475800.0 ;
      RECT  547800.0 489600.0 558000.0 503400.0 ;
      RECT  547800.0 517200.0 558000.0 503400.0 ;
      RECT  547800.0 517200.0 558000.0 531000.0 ;
      RECT  547800.0 544800.0 558000.0 531000.0 ;
      RECT  547800.0 544800.0 558000.0 558600.0 ;
      RECT  547800.0 572400.0 558000.0 558600.0 ;
      RECT  547800.0 572400.0 558000.0 586200.0 ;
      RECT  547800.0 600000.0 558000.0 586200.0 ;
      RECT  547800.0 600000.0 558000.0 613800.0 ;
      RECT  547800.0 627600.0 558000.0 613800.0 ;
      RECT  547800.0 627600.0 558000.0 641400.0 ;
      RECT  547800.0 655200.0 558000.0 641400.0 ;
      RECT  547800.0 655200.0 558000.0 669000.0 ;
      RECT  547800.0 682800.0 558000.0 669000.0 ;
      RECT  547800.0 682800.0 558000.0 696600.0 ;
      RECT  547800.0 710400.0 558000.0 696600.0 ;
      RECT  547800.0 710400.0 558000.0 724200.0 ;
      RECT  547800.0 738000.0 558000.0 724200.0 ;
      RECT  547800.0 738000.0 558000.0 751800.0 ;
      RECT  547800.0 765600.0 558000.0 751800.0 ;
      RECT  547800.0 765600.0 558000.0 779400.0 ;
      RECT  547800.0 793200.0 558000.0 779400.0 ;
      RECT  547800.0 793200.0 558000.0 807000.0 ;
      RECT  547800.0 820800.0 558000.0 807000.0 ;
      RECT  547800.0 820800.0 558000.0 834600.0 ;
      RECT  547800.0 848400.0 558000.0 834600.0 ;
      RECT  547800.0 848400.0 558000.0 862200.0 ;
      RECT  547800.0 876000.0 558000.0 862200.0 ;
      RECT  547800.0 876000.0 558000.0 889800.0 ;
      RECT  547800.0 903600.0 558000.0 889800.0 ;
      RECT  547800.0 903600.0 558000.0 917400.0 ;
      RECT  547800.0 931200.0 558000.0 917400.0 ;
      RECT  547800.0 931200.0 558000.0 945000.0 ;
      RECT  547800.0 958800.0 558000.0 945000.0 ;
      RECT  547800.0 958800.0 558000.0 972600.0 ;
      RECT  547800.0 986400.0 558000.0 972600.0 ;
      RECT  547800.0 986400.0 558000.0 1000200.0 ;
      RECT  547800.0 1014000.0 558000.0 1000200.0 ;
      RECT  547800.0 1014000.0 558000.0 1027800.0 ;
      RECT  547800.0 1041600.0 558000.0 1027800.0 ;
      RECT  547800.0 1041600.0 558000.0 1055400.0 ;
      RECT  547800.0 1069200.0 558000.0 1055400.0 ;
      RECT  547800.0 1069200.0 558000.0 1083000.0 ;
      RECT  547800.0 1096800.0 558000.0 1083000.0 ;
      RECT  547800.0 1096800.0 558000.0 1110600.0 ;
      RECT  547800.0 1124400.0 558000.0 1110600.0 ;
      RECT  547800.0 1124400.0 558000.0 1138200.0 ;
      RECT  547800.0 1152000.0 558000.0 1138200.0 ;
      RECT  547800.0 1152000.0 558000.0 1165800.0 ;
      RECT  547800.0 1179600.0 558000.0 1165800.0 ;
      RECT  547800.0 1179600.0 558000.0 1193400.0 ;
      RECT  547800.0 1207200.0 558000.0 1193400.0 ;
      RECT  547800.0 1207200.0 558000.0 1221000.0 ;
      RECT  547800.0 1234800.0 558000.0 1221000.0 ;
      RECT  547800.0 1234800.0 558000.0 1248600.0 ;
      RECT  547800.0 1262400.0 558000.0 1248600.0 ;
      RECT  547800.0 1262400.0 558000.0 1276200.0 ;
      RECT  547800.0 1290000.0 558000.0 1276200.0 ;
      RECT  547800.0 1290000.0 558000.0 1303800.0 ;
      RECT  547800.0 1317600.0 558000.0 1303800.0 ;
      RECT  547800.0 1317600.0 558000.0 1331400.0 ;
      RECT  547800.0 1345200.0 558000.0 1331400.0 ;
      RECT  547800.0 1345200.0 558000.0 1359000.0 ;
      RECT  547800.0 1372800.0 558000.0 1359000.0 ;
      RECT  547800.0 1372800.0 558000.0 1386600.0 ;
      RECT  547800.0 1400400.0 558000.0 1386600.0 ;
      RECT  547800.0 1400400.0 558000.0 1414200.0 ;
      RECT  547800.0 1428000.0 558000.0 1414200.0 ;
      RECT  547800.0 1428000.0 558000.0 1441800.0 ;
      RECT  547800.0 1455600.0 558000.0 1441800.0 ;
      RECT  547800.0 1455600.0 558000.0 1469400.0 ;
      RECT  547800.0 1483200.0 558000.0 1469400.0 ;
      RECT  547800.0 1483200.0 558000.0 1497000.0 ;
      RECT  547800.0 1510800.0 558000.0 1497000.0 ;
      RECT  547800.0 1510800.0 558000.0 1524600.0 ;
      RECT  547800.0 1538400.0 558000.0 1524600.0 ;
      RECT  547800.0 1538400.0 558000.0 1552200.0 ;
      RECT  547800.0 1566000.0 558000.0 1552200.0 ;
      RECT  547800.0 1566000.0 558000.0 1579800.0 ;
      RECT  547800.0 1593600.0 558000.0 1579800.0 ;
      RECT  547800.0 1593600.0 558000.0 1607400.0 ;
      RECT  547800.0 1621200.0 558000.0 1607400.0 ;
      RECT  547800.0 1621200.0 558000.0 1635000.0 ;
      RECT  547800.0 1648800.0 558000.0 1635000.0 ;
      RECT  547800.0 1648800.0 558000.0 1662600.0 ;
      RECT  547800.0 1676400.0 558000.0 1662600.0 ;
      RECT  547800.0 1676400.0 558000.0 1690200.0 ;
      RECT  547800.0 1704000.0 558000.0 1690200.0 ;
      RECT  547800.0 1704000.0 558000.0 1717800.0 ;
      RECT  547800.0 1731600.0 558000.0 1717800.0 ;
      RECT  547800.0 1731600.0 558000.0 1745400.0 ;
      RECT  547800.0 1759200.0 558000.0 1745400.0 ;
      RECT  547800.0 1759200.0 558000.0 1773000.0 ;
      RECT  547800.0 1786800.0 558000.0 1773000.0 ;
      RECT  547800.0 1786800.0 558000.0 1800600.0 ;
      RECT  547800.0 1814400.0 558000.0 1800600.0 ;
      RECT  547800.0 1814400.0 558000.0 1828200.0 ;
      RECT  547800.0 1842000.0 558000.0 1828200.0 ;
      RECT  547800.0 1842000.0 558000.0 1855800.0 ;
      RECT  547800.0 1869600.0 558000.0 1855800.0 ;
      RECT  547800.0 1869600.0 558000.0 1883400.0 ;
      RECT  547800.0 1897200.0 558000.0 1883400.0 ;
      RECT  547800.0 1897200.0 558000.0 1911000.0 ;
      RECT  547800.0 1924800.0 558000.0 1911000.0 ;
      RECT  547800.0 1924800.0 558000.0 1938600.0 ;
      RECT  547800.0 1952400.0 558000.0 1938600.0 ;
      RECT  547800.0 1952400.0 558000.0 1966200.0 ;
      RECT  547800.0 1980000.0 558000.0 1966200.0 ;
      RECT  547800.0 1980000.0 558000.0 1993800.0 ;
      RECT  547800.0 2007600.0 558000.0 1993800.0 ;
      RECT  547800.0 2007600.0 558000.0 2021400.0 ;
      RECT  547800.0 2035200.0 558000.0 2021400.0 ;
      RECT  547800.0 2035200.0 558000.0 2049000.0 ;
      RECT  547800.0 2062800.0 558000.0 2049000.0 ;
      RECT  547800.0 2062800.0 558000.0 2076600.0 ;
      RECT  547800.0 2090400.0 558000.0 2076600.0 ;
      RECT  547800.0 2090400.0 558000.0 2104200.0 ;
      RECT  547800.0 2118000.0 558000.0 2104200.0 ;
      RECT  547800.0 2118000.0 558000.0 2131800.0 ;
      RECT  547800.0 2145600.0 558000.0 2131800.0 ;
      RECT  558000.0 379200.0 568200.0 393000.0 ;
      RECT  558000.0 406800.0 568200.0 393000.0 ;
      RECT  558000.0 406800.0 568200.0 420600.0 ;
      RECT  558000.0 434400.0 568200.0 420600.0 ;
      RECT  558000.0 434400.0 568200.0 448200.0 ;
      RECT  558000.0 462000.0 568200.0 448200.0 ;
      RECT  558000.0 462000.0 568200.0 475800.0 ;
      RECT  558000.0 489600.0 568200.0 475800.0 ;
      RECT  558000.0 489600.0 568200.0 503400.0 ;
      RECT  558000.0 517200.0 568200.0 503400.0 ;
      RECT  558000.0 517200.0 568200.0 531000.0 ;
      RECT  558000.0 544800.0 568200.0 531000.0 ;
      RECT  558000.0 544800.0 568200.0 558600.0 ;
      RECT  558000.0 572400.0 568200.0 558600.0 ;
      RECT  558000.0 572400.0 568200.0 586200.0 ;
      RECT  558000.0 600000.0 568200.0 586200.0 ;
      RECT  558000.0 600000.0 568200.0 613800.0 ;
      RECT  558000.0 627600.0 568200.0 613800.0 ;
      RECT  558000.0 627600.0 568200.0 641400.0 ;
      RECT  558000.0 655200.0 568200.0 641400.0 ;
      RECT  558000.0 655200.0 568200.0 669000.0 ;
      RECT  558000.0 682800.0 568200.0 669000.0 ;
      RECT  558000.0 682800.0 568200.0 696600.0 ;
      RECT  558000.0 710400.0 568200.0 696600.0 ;
      RECT  558000.0 710400.0 568200.0 724200.0 ;
      RECT  558000.0 738000.0 568200.0 724200.0 ;
      RECT  558000.0 738000.0 568200.0 751800.0 ;
      RECT  558000.0 765600.0 568200.0 751800.0 ;
      RECT  558000.0 765600.0 568200.0 779400.0 ;
      RECT  558000.0 793200.0 568200.0 779400.0 ;
      RECT  558000.0 793200.0 568200.0 807000.0 ;
      RECT  558000.0 820800.0 568200.0 807000.0 ;
      RECT  558000.0 820800.0 568200.0 834600.0 ;
      RECT  558000.0 848400.0 568200.0 834600.0 ;
      RECT  558000.0 848400.0 568200.0 862200.0 ;
      RECT  558000.0 876000.0 568200.0 862200.0 ;
      RECT  558000.0 876000.0 568200.0 889800.0 ;
      RECT  558000.0 903600.0 568200.0 889800.0 ;
      RECT  558000.0 903600.0 568200.0 917400.0 ;
      RECT  558000.0 931200.0 568200.0 917400.0 ;
      RECT  558000.0 931200.0 568200.0 945000.0 ;
      RECT  558000.0 958800.0 568200.0 945000.0 ;
      RECT  558000.0 958800.0 568200.0 972600.0 ;
      RECT  558000.0 986400.0 568200.0 972600.0 ;
      RECT  558000.0 986400.0 568200.0 1000200.0 ;
      RECT  558000.0 1014000.0 568200.0 1000200.0 ;
      RECT  558000.0 1014000.0 568200.0 1027800.0 ;
      RECT  558000.0 1041600.0 568200.0 1027800.0 ;
      RECT  558000.0 1041600.0 568200.0 1055400.0 ;
      RECT  558000.0 1069200.0 568200.0 1055400.0 ;
      RECT  558000.0 1069200.0 568200.0 1083000.0 ;
      RECT  558000.0 1096800.0 568200.0 1083000.0 ;
      RECT  558000.0 1096800.0 568200.0 1110600.0 ;
      RECT  558000.0 1124400.0 568200.0 1110600.0 ;
      RECT  558000.0 1124400.0 568200.0 1138200.0 ;
      RECT  558000.0 1152000.0 568200.0 1138200.0 ;
      RECT  558000.0 1152000.0 568200.0 1165800.0 ;
      RECT  558000.0 1179600.0 568200.0 1165800.0 ;
      RECT  558000.0 1179600.0 568200.0 1193400.0 ;
      RECT  558000.0 1207200.0 568200.0 1193400.0 ;
      RECT  558000.0 1207200.0 568200.0 1221000.0 ;
      RECT  558000.0 1234800.0 568200.0 1221000.0 ;
      RECT  558000.0 1234800.0 568200.0 1248600.0 ;
      RECT  558000.0 1262400.0 568200.0 1248600.0 ;
      RECT  558000.0 1262400.0 568200.0 1276200.0 ;
      RECT  558000.0 1290000.0 568200.0 1276200.0 ;
      RECT  558000.0 1290000.0 568200.0 1303800.0 ;
      RECT  558000.0 1317600.0 568200.0 1303800.0 ;
      RECT  558000.0 1317600.0 568200.0 1331400.0 ;
      RECT  558000.0 1345200.0 568200.0 1331400.0 ;
      RECT  558000.0 1345200.0 568200.0 1359000.0 ;
      RECT  558000.0 1372800.0 568200.0 1359000.0 ;
      RECT  558000.0 1372800.0 568200.0 1386600.0 ;
      RECT  558000.0 1400400.0 568200.0 1386600.0 ;
      RECT  558000.0 1400400.0 568200.0 1414200.0 ;
      RECT  558000.0 1428000.0 568200.0 1414200.0 ;
      RECT  558000.0 1428000.0 568200.0 1441800.0 ;
      RECT  558000.0 1455600.0 568200.0 1441800.0 ;
      RECT  558000.0 1455600.0 568200.0 1469400.0 ;
      RECT  558000.0 1483200.0 568200.0 1469400.0 ;
      RECT  558000.0 1483200.0 568200.0 1497000.0 ;
      RECT  558000.0 1510800.0 568200.0 1497000.0 ;
      RECT  558000.0 1510800.0 568200.0 1524600.0 ;
      RECT  558000.0 1538400.0 568200.0 1524600.0 ;
      RECT  558000.0 1538400.0 568200.0 1552200.0 ;
      RECT  558000.0 1566000.0 568200.0 1552200.0 ;
      RECT  558000.0 1566000.0 568200.0 1579800.0 ;
      RECT  558000.0 1593600.0 568200.0 1579800.0 ;
      RECT  558000.0 1593600.0 568200.0 1607400.0 ;
      RECT  558000.0 1621200.0 568200.0 1607400.0 ;
      RECT  558000.0 1621200.0 568200.0 1635000.0 ;
      RECT  558000.0 1648800.0 568200.0 1635000.0 ;
      RECT  558000.0 1648800.0 568200.0 1662600.0 ;
      RECT  558000.0 1676400.0 568200.0 1662600.0 ;
      RECT  558000.0 1676400.0 568200.0 1690200.0 ;
      RECT  558000.0 1704000.0 568200.0 1690200.0 ;
      RECT  558000.0 1704000.0 568200.0 1717800.0 ;
      RECT  558000.0 1731600.0 568200.0 1717800.0 ;
      RECT  558000.0 1731600.0 568200.0 1745400.0 ;
      RECT  558000.0 1759200.0 568200.0 1745400.0 ;
      RECT  558000.0 1759200.0 568200.0 1773000.0 ;
      RECT  558000.0 1786800.0 568200.0 1773000.0 ;
      RECT  558000.0 1786800.0 568200.0 1800600.0 ;
      RECT  558000.0 1814400.0 568200.0 1800600.0 ;
      RECT  558000.0 1814400.0 568200.0 1828200.0 ;
      RECT  558000.0 1842000.0 568200.0 1828200.0 ;
      RECT  558000.0 1842000.0 568200.0 1855800.0 ;
      RECT  558000.0 1869600.0 568200.0 1855800.0 ;
      RECT  558000.0 1869600.0 568200.0 1883400.0 ;
      RECT  558000.0 1897200.0 568200.0 1883400.0 ;
      RECT  558000.0 1897200.0 568200.0 1911000.0 ;
      RECT  558000.0 1924800.0 568200.0 1911000.0 ;
      RECT  558000.0 1924800.0 568200.0 1938600.0 ;
      RECT  558000.0 1952400.0 568200.0 1938600.0 ;
      RECT  558000.0 1952400.0 568200.0 1966200.0 ;
      RECT  558000.0 1980000.0 568200.0 1966200.0 ;
      RECT  558000.0 1980000.0 568200.0 1993800.0 ;
      RECT  558000.0 2007600.0 568200.0 1993800.0 ;
      RECT  558000.0 2007600.0 568200.0 2021400.0 ;
      RECT  558000.0 2035200.0 568200.0 2021400.0 ;
      RECT  558000.0 2035200.0 568200.0 2049000.0 ;
      RECT  558000.0 2062800.0 568200.0 2049000.0 ;
      RECT  558000.0 2062800.0 568200.0 2076600.0 ;
      RECT  558000.0 2090400.0 568200.0 2076600.0 ;
      RECT  558000.0 2090400.0 568200.0 2104200.0 ;
      RECT  558000.0 2118000.0 568200.0 2104200.0 ;
      RECT  558000.0 2118000.0 568200.0 2131800.0 ;
      RECT  558000.0 2145600.0 568200.0 2131800.0 ;
      RECT  568200.0 379200.0 578400.0 393000.0 ;
      RECT  568200.0 406800.0 578400.0 393000.0 ;
      RECT  568200.0 406800.0 578400.0 420600.0 ;
      RECT  568200.0 434400.0 578400.0 420600.0 ;
      RECT  568200.0 434400.0 578400.0 448200.0 ;
      RECT  568200.0 462000.0 578400.0 448200.0 ;
      RECT  568200.0 462000.0 578400.0 475800.0 ;
      RECT  568200.0 489600.0 578400.0 475800.0 ;
      RECT  568200.0 489600.0 578400.0 503400.0 ;
      RECT  568200.0 517200.0 578400.0 503400.0 ;
      RECT  568200.0 517200.0 578400.0 531000.0 ;
      RECT  568200.0 544800.0 578400.0 531000.0 ;
      RECT  568200.0 544800.0 578400.0 558600.0 ;
      RECT  568200.0 572400.0 578400.0 558600.0 ;
      RECT  568200.0 572400.0 578400.0 586200.0 ;
      RECT  568200.0 600000.0 578400.0 586200.0 ;
      RECT  568200.0 600000.0 578400.0 613800.0 ;
      RECT  568200.0 627600.0 578400.0 613800.0 ;
      RECT  568200.0 627600.0 578400.0 641400.0 ;
      RECT  568200.0 655200.0 578400.0 641400.0 ;
      RECT  568200.0 655200.0 578400.0 669000.0 ;
      RECT  568200.0 682800.0 578400.0 669000.0 ;
      RECT  568200.0 682800.0 578400.0 696600.0 ;
      RECT  568200.0 710400.0 578400.0 696600.0 ;
      RECT  568200.0 710400.0 578400.0 724200.0 ;
      RECT  568200.0 738000.0 578400.0 724200.0 ;
      RECT  568200.0 738000.0 578400.0 751800.0 ;
      RECT  568200.0 765600.0 578400.0 751800.0 ;
      RECT  568200.0 765600.0 578400.0 779400.0 ;
      RECT  568200.0 793200.0 578400.0 779400.0 ;
      RECT  568200.0 793200.0 578400.0 807000.0 ;
      RECT  568200.0 820800.0 578400.0 807000.0 ;
      RECT  568200.0 820800.0 578400.0 834600.0 ;
      RECT  568200.0 848400.0 578400.0 834600.0 ;
      RECT  568200.0 848400.0 578400.0 862200.0 ;
      RECT  568200.0 876000.0 578400.0 862200.0 ;
      RECT  568200.0 876000.0 578400.0 889800.0 ;
      RECT  568200.0 903600.0 578400.0 889800.0 ;
      RECT  568200.0 903600.0 578400.0 917400.0 ;
      RECT  568200.0 931200.0 578400.0 917400.0 ;
      RECT  568200.0 931200.0 578400.0 945000.0 ;
      RECT  568200.0 958800.0 578400.0 945000.0 ;
      RECT  568200.0 958800.0 578400.0 972600.0 ;
      RECT  568200.0 986400.0 578400.0 972600.0 ;
      RECT  568200.0 986400.0 578400.0 1000200.0 ;
      RECT  568200.0 1014000.0 578400.0 1000200.0 ;
      RECT  568200.0 1014000.0 578400.0 1027800.0 ;
      RECT  568200.0 1041600.0 578400.0 1027800.0 ;
      RECT  568200.0 1041600.0 578400.0 1055400.0 ;
      RECT  568200.0 1069200.0 578400.0 1055400.0 ;
      RECT  568200.0 1069200.0 578400.0 1083000.0 ;
      RECT  568200.0 1096800.0 578400.0 1083000.0 ;
      RECT  568200.0 1096800.0 578400.0 1110600.0 ;
      RECT  568200.0 1124400.0 578400.0 1110600.0 ;
      RECT  568200.0 1124400.0 578400.0 1138200.0 ;
      RECT  568200.0 1152000.0 578400.0 1138200.0 ;
      RECT  568200.0 1152000.0 578400.0 1165800.0 ;
      RECT  568200.0 1179600.0 578400.0 1165800.0 ;
      RECT  568200.0 1179600.0 578400.0 1193400.0 ;
      RECT  568200.0 1207200.0 578400.0 1193400.0 ;
      RECT  568200.0 1207200.0 578400.0 1221000.0 ;
      RECT  568200.0 1234800.0 578400.0 1221000.0 ;
      RECT  568200.0 1234800.0 578400.0 1248600.0 ;
      RECT  568200.0 1262400.0 578400.0 1248600.0 ;
      RECT  568200.0 1262400.0 578400.0 1276200.0 ;
      RECT  568200.0 1290000.0 578400.0 1276200.0 ;
      RECT  568200.0 1290000.0 578400.0 1303800.0 ;
      RECT  568200.0 1317600.0 578400.0 1303800.0 ;
      RECT  568200.0 1317600.0 578400.0 1331400.0 ;
      RECT  568200.0 1345200.0 578400.0 1331400.0 ;
      RECT  568200.0 1345200.0 578400.0 1359000.0 ;
      RECT  568200.0 1372800.0 578400.0 1359000.0 ;
      RECT  568200.0 1372800.0 578400.0 1386600.0 ;
      RECT  568200.0 1400400.0 578400.0 1386600.0 ;
      RECT  568200.0 1400400.0 578400.0 1414200.0 ;
      RECT  568200.0 1428000.0 578400.0 1414200.0 ;
      RECT  568200.0 1428000.0 578400.0 1441800.0 ;
      RECT  568200.0 1455600.0 578400.0 1441800.0 ;
      RECT  568200.0 1455600.0 578400.0 1469400.0 ;
      RECT  568200.0 1483200.0 578400.0 1469400.0 ;
      RECT  568200.0 1483200.0 578400.0 1497000.0 ;
      RECT  568200.0 1510800.0 578400.0 1497000.0 ;
      RECT  568200.0 1510800.0 578400.0 1524600.0 ;
      RECT  568200.0 1538400.0 578400.0 1524600.0 ;
      RECT  568200.0 1538400.0 578400.0 1552200.0 ;
      RECT  568200.0 1566000.0 578400.0 1552200.0 ;
      RECT  568200.0 1566000.0 578400.0 1579800.0 ;
      RECT  568200.0 1593600.0 578400.0 1579800.0 ;
      RECT  568200.0 1593600.0 578400.0 1607400.0 ;
      RECT  568200.0 1621200.0 578400.0 1607400.0 ;
      RECT  568200.0 1621200.0 578400.0 1635000.0 ;
      RECT  568200.0 1648800.0 578400.0 1635000.0 ;
      RECT  568200.0 1648800.0 578400.0 1662600.0 ;
      RECT  568200.0 1676400.0 578400.0 1662600.0 ;
      RECT  568200.0 1676400.0 578400.0 1690200.0 ;
      RECT  568200.0 1704000.0 578400.0 1690200.0 ;
      RECT  568200.0 1704000.0 578400.0 1717800.0 ;
      RECT  568200.0 1731600.0 578400.0 1717800.0 ;
      RECT  568200.0 1731600.0 578400.0 1745400.0 ;
      RECT  568200.0 1759200.0 578400.0 1745400.0 ;
      RECT  568200.0 1759200.0 578400.0 1773000.0 ;
      RECT  568200.0 1786800.0 578400.0 1773000.0 ;
      RECT  568200.0 1786800.0 578400.0 1800600.0 ;
      RECT  568200.0 1814400.0 578400.0 1800600.0 ;
      RECT  568200.0 1814400.0 578400.0 1828200.0 ;
      RECT  568200.0 1842000.0 578400.0 1828200.0 ;
      RECT  568200.0 1842000.0 578400.0 1855800.0 ;
      RECT  568200.0 1869600.0 578400.0 1855800.0 ;
      RECT  568200.0 1869600.0 578400.0 1883400.0 ;
      RECT  568200.0 1897200.0 578400.0 1883400.0 ;
      RECT  568200.0 1897200.0 578400.0 1911000.0 ;
      RECT  568200.0 1924800.0 578400.0 1911000.0 ;
      RECT  568200.0 1924800.0 578400.0 1938600.0 ;
      RECT  568200.0 1952400.0 578400.0 1938600.0 ;
      RECT  568200.0 1952400.0 578400.0 1966200.0 ;
      RECT  568200.0 1980000.0 578400.0 1966200.0 ;
      RECT  568200.0 1980000.0 578400.0 1993800.0 ;
      RECT  568200.0 2007600.0 578400.0 1993800.0 ;
      RECT  568200.0 2007600.0 578400.0 2021400.0 ;
      RECT  568200.0 2035200.0 578400.0 2021400.0 ;
      RECT  568200.0 2035200.0 578400.0 2049000.0 ;
      RECT  568200.0 2062800.0 578400.0 2049000.0 ;
      RECT  568200.0 2062800.0 578400.0 2076600.0 ;
      RECT  568200.0 2090400.0 578400.0 2076600.0 ;
      RECT  568200.0 2090400.0 578400.0 2104200.0 ;
      RECT  568200.0 2118000.0 578400.0 2104200.0 ;
      RECT  568200.0 2118000.0 578400.0 2131800.0 ;
      RECT  568200.0 2145600.0 578400.0 2131800.0 ;
      RECT  578400.0 379200.0 588600.0 393000.0 ;
      RECT  578400.0 406800.0 588600.0 393000.0 ;
      RECT  578400.0 406800.0 588600.0 420600.0 ;
      RECT  578400.0 434400.0 588600.0 420600.0 ;
      RECT  578400.0 434400.0 588600.0 448200.0 ;
      RECT  578400.0 462000.0 588600.0 448200.0 ;
      RECT  578400.0 462000.0 588600.0 475800.0 ;
      RECT  578400.0 489600.0 588600.0 475800.0 ;
      RECT  578400.0 489600.0 588600.0 503400.0 ;
      RECT  578400.0 517200.0 588600.0 503400.0 ;
      RECT  578400.0 517200.0 588600.0 531000.0 ;
      RECT  578400.0 544800.0 588600.0 531000.0 ;
      RECT  578400.0 544800.0 588600.0 558600.0 ;
      RECT  578400.0 572400.0 588600.0 558600.0 ;
      RECT  578400.0 572400.0 588600.0 586200.0 ;
      RECT  578400.0 600000.0 588600.0 586200.0 ;
      RECT  578400.0 600000.0 588600.0 613800.0 ;
      RECT  578400.0 627600.0 588600.0 613800.0 ;
      RECT  578400.0 627600.0 588600.0 641400.0 ;
      RECT  578400.0 655200.0 588600.0 641400.0 ;
      RECT  578400.0 655200.0 588600.0 669000.0 ;
      RECT  578400.0 682800.0 588600.0 669000.0 ;
      RECT  578400.0 682800.0 588600.0 696600.0 ;
      RECT  578400.0 710400.0 588600.0 696600.0 ;
      RECT  578400.0 710400.0 588600.0 724200.0 ;
      RECT  578400.0 738000.0 588600.0 724200.0 ;
      RECT  578400.0 738000.0 588600.0 751800.0 ;
      RECT  578400.0 765600.0 588600.0 751800.0 ;
      RECT  578400.0 765600.0 588600.0 779400.0 ;
      RECT  578400.0 793200.0 588600.0 779400.0 ;
      RECT  578400.0 793200.0 588600.0 807000.0 ;
      RECT  578400.0 820800.0 588600.0 807000.0 ;
      RECT  578400.0 820800.0 588600.0 834600.0 ;
      RECT  578400.0 848400.0 588600.0 834600.0 ;
      RECT  578400.0 848400.0 588600.0 862200.0 ;
      RECT  578400.0 876000.0 588600.0 862200.0 ;
      RECT  578400.0 876000.0 588600.0 889800.0 ;
      RECT  578400.0 903600.0 588600.0 889800.0 ;
      RECT  578400.0 903600.0 588600.0 917400.0 ;
      RECT  578400.0 931200.0 588600.0 917400.0 ;
      RECT  578400.0 931200.0 588600.0 945000.0 ;
      RECT  578400.0 958800.0 588600.0 945000.0 ;
      RECT  578400.0 958800.0 588600.0 972600.0 ;
      RECT  578400.0 986400.0 588600.0 972600.0 ;
      RECT  578400.0 986400.0 588600.0 1000200.0 ;
      RECT  578400.0 1014000.0 588600.0 1000200.0 ;
      RECT  578400.0 1014000.0 588600.0 1027800.0 ;
      RECT  578400.0 1041600.0 588600.0 1027800.0 ;
      RECT  578400.0 1041600.0 588600.0 1055400.0 ;
      RECT  578400.0 1069200.0 588600.0 1055400.0 ;
      RECT  578400.0 1069200.0 588600.0 1083000.0 ;
      RECT  578400.0 1096800.0 588600.0 1083000.0 ;
      RECT  578400.0 1096800.0 588600.0 1110600.0 ;
      RECT  578400.0 1124400.0 588600.0 1110600.0 ;
      RECT  578400.0 1124400.0 588600.0 1138200.0 ;
      RECT  578400.0 1152000.0 588600.0 1138200.0 ;
      RECT  578400.0 1152000.0 588600.0 1165800.0 ;
      RECT  578400.0 1179600.0 588600.0 1165800.0 ;
      RECT  578400.0 1179600.0 588600.0 1193400.0 ;
      RECT  578400.0 1207200.0 588600.0 1193400.0 ;
      RECT  578400.0 1207200.0 588600.0 1221000.0 ;
      RECT  578400.0 1234800.0 588600.0 1221000.0 ;
      RECT  578400.0 1234800.0 588600.0 1248600.0 ;
      RECT  578400.0 1262400.0 588600.0 1248600.0 ;
      RECT  578400.0 1262400.0 588600.0 1276200.0 ;
      RECT  578400.0 1290000.0 588600.0 1276200.0 ;
      RECT  578400.0 1290000.0 588600.0 1303800.0 ;
      RECT  578400.0 1317600.0 588600.0 1303800.0 ;
      RECT  578400.0 1317600.0 588600.0 1331400.0 ;
      RECT  578400.0 1345200.0 588600.0 1331400.0 ;
      RECT  578400.0 1345200.0 588600.0 1359000.0 ;
      RECT  578400.0 1372800.0 588600.0 1359000.0 ;
      RECT  578400.0 1372800.0 588600.0 1386600.0 ;
      RECT  578400.0 1400400.0 588600.0 1386600.0 ;
      RECT  578400.0 1400400.0 588600.0 1414200.0 ;
      RECT  578400.0 1428000.0 588600.0 1414200.0 ;
      RECT  578400.0 1428000.0 588600.0 1441800.0 ;
      RECT  578400.0 1455600.0 588600.0 1441800.0 ;
      RECT  578400.0 1455600.0 588600.0 1469400.0 ;
      RECT  578400.0 1483200.0 588600.0 1469400.0 ;
      RECT  578400.0 1483200.0 588600.0 1497000.0 ;
      RECT  578400.0 1510800.0 588600.0 1497000.0 ;
      RECT  578400.0 1510800.0 588600.0 1524600.0 ;
      RECT  578400.0 1538400.0 588600.0 1524600.0 ;
      RECT  578400.0 1538400.0 588600.0 1552200.0 ;
      RECT  578400.0 1566000.0 588600.0 1552200.0 ;
      RECT  578400.0 1566000.0 588600.0 1579800.0 ;
      RECT  578400.0 1593600.0 588600.0 1579800.0 ;
      RECT  578400.0 1593600.0 588600.0 1607400.0 ;
      RECT  578400.0 1621200.0 588600.0 1607400.0 ;
      RECT  578400.0 1621200.0 588600.0 1635000.0 ;
      RECT  578400.0 1648800.0 588600.0 1635000.0 ;
      RECT  578400.0 1648800.0 588600.0 1662600.0 ;
      RECT  578400.0 1676400.0 588600.0 1662600.0 ;
      RECT  578400.0 1676400.0 588600.0 1690200.0 ;
      RECT  578400.0 1704000.0 588600.0 1690200.0 ;
      RECT  578400.0 1704000.0 588600.0 1717800.0 ;
      RECT  578400.0 1731600.0 588600.0 1717800.0 ;
      RECT  578400.0 1731600.0 588600.0 1745400.0 ;
      RECT  578400.0 1759200.0 588600.0 1745400.0 ;
      RECT  578400.0 1759200.0 588600.0 1773000.0 ;
      RECT  578400.0 1786800.0 588600.0 1773000.0 ;
      RECT  578400.0 1786800.0 588600.0 1800600.0 ;
      RECT  578400.0 1814400.0 588600.0 1800600.0 ;
      RECT  578400.0 1814400.0 588600.0 1828200.0 ;
      RECT  578400.0 1842000.0 588600.0 1828200.0 ;
      RECT  578400.0 1842000.0 588600.0 1855800.0 ;
      RECT  578400.0 1869600.0 588600.0 1855800.0 ;
      RECT  578400.0 1869600.0 588600.0 1883400.0 ;
      RECT  578400.0 1897200.0 588600.0 1883400.0 ;
      RECT  578400.0 1897200.0 588600.0 1911000.0 ;
      RECT  578400.0 1924800.0 588600.0 1911000.0 ;
      RECT  578400.0 1924800.0 588600.0 1938600.0 ;
      RECT  578400.0 1952400.0 588600.0 1938600.0 ;
      RECT  578400.0 1952400.0 588600.0 1966200.0 ;
      RECT  578400.0 1980000.0 588600.0 1966200.0 ;
      RECT  578400.0 1980000.0 588600.0 1993800.0 ;
      RECT  578400.0 2007600.0 588600.0 1993800.0 ;
      RECT  578400.0 2007600.0 588600.0 2021400.0 ;
      RECT  578400.0 2035200.0 588600.0 2021400.0 ;
      RECT  578400.0 2035200.0 588600.0 2049000.0 ;
      RECT  578400.0 2062800.0 588600.0 2049000.0 ;
      RECT  578400.0 2062800.0 588600.0 2076600.0 ;
      RECT  578400.0 2090400.0 588600.0 2076600.0 ;
      RECT  578400.0 2090400.0 588600.0 2104200.0 ;
      RECT  578400.0 2118000.0 588600.0 2104200.0 ;
      RECT  578400.0 2118000.0 588600.0 2131800.0 ;
      RECT  578400.0 2145600.0 588600.0 2131800.0 ;
      RECT  588600.0 379200.0 598800.0 393000.0 ;
      RECT  588600.0 406800.0 598800.0 393000.0 ;
      RECT  588600.0 406800.0 598800.0 420600.0 ;
      RECT  588600.0 434400.0 598800.0 420600.0 ;
      RECT  588600.0 434400.0 598800.0 448200.0 ;
      RECT  588600.0 462000.0 598800.0 448200.0 ;
      RECT  588600.0 462000.0 598800.0 475800.0 ;
      RECT  588600.0 489600.0 598800.0 475800.0 ;
      RECT  588600.0 489600.0 598800.0 503400.0 ;
      RECT  588600.0 517200.0 598800.0 503400.0 ;
      RECT  588600.0 517200.0 598800.0 531000.0 ;
      RECT  588600.0 544800.0 598800.0 531000.0 ;
      RECT  588600.0 544800.0 598800.0 558600.0 ;
      RECT  588600.0 572400.0 598800.0 558600.0 ;
      RECT  588600.0 572400.0 598800.0 586200.0 ;
      RECT  588600.0 600000.0 598800.0 586200.0 ;
      RECT  588600.0 600000.0 598800.0 613800.0 ;
      RECT  588600.0 627600.0 598800.0 613800.0 ;
      RECT  588600.0 627600.0 598800.0 641400.0 ;
      RECT  588600.0 655200.0 598800.0 641400.0 ;
      RECT  588600.0 655200.0 598800.0 669000.0 ;
      RECT  588600.0 682800.0 598800.0 669000.0 ;
      RECT  588600.0 682800.0 598800.0 696600.0 ;
      RECT  588600.0 710400.0 598800.0 696600.0 ;
      RECT  588600.0 710400.0 598800.0 724200.0 ;
      RECT  588600.0 738000.0 598800.0 724200.0 ;
      RECT  588600.0 738000.0 598800.0 751800.0 ;
      RECT  588600.0 765600.0 598800.0 751800.0 ;
      RECT  588600.0 765600.0 598800.0 779400.0 ;
      RECT  588600.0 793200.0 598800.0 779400.0 ;
      RECT  588600.0 793200.0 598800.0 807000.0 ;
      RECT  588600.0 820800.0 598800.0 807000.0 ;
      RECT  588600.0 820800.0 598800.0 834600.0 ;
      RECT  588600.0 848400.0 598800.0 834600.0 ;
      RECT  588600.0 848400.0 598800.0 862200.0 ;
      RECT  588600.0 876000.0 598800.0 862200.0 ;
      RECT  588600.0 876000.0 598800.0 889800.0 ;
      RECT  588600.0 903600.0 598800.0 889800.0 ;
      RECT  588600.0 903600.0 598800.0 917400.0 ;
      RECT  588600.0 931200.0 598800.0 917400.0 ;
      RECT  588600.0 931200.0 598800.0 945000.0 ;
      RECT  588600.0 958800.0 598800.0 945000.0 ;
      RECT  588600.0 958800.0 598800.0 972600.0 ;
      RECT  588600.0 986400.0 598800.0 972600.0 ;
      RECT  588600.0 986400.0 598800.0 1000200.0 ;
      RECT  588600.0 1014000.0 598800.0 1000200.0 ;
      RECT  588600.0 1014000.0 598800.0 1027800.0 ;
      RECT  588600.0 1041600.0 598800.0 1027800.0 ;
      RECT  588600.0 1041600.0 598800.0 1055400.0 ;
      RECT  588600.0 1069200.0 598800.0 1055400.0 ;
      RECT  588600.0 1069200.0 598800.0 1083000.0 ;
      RECT  588600.0 1096800.0 598800.0 1083000.0 ;
      RECT  588600.0 1096800.0 598800.0 1110600.0 ;
      RECT  588600.0 1124400.0 598800.0 1110600.0 ;
      RECT  588600.0 1124400.0 598800.0 1138200.0 ;
      RECT  588600.0 1152000.0 598800.0 1138200.0 ;
      RECT  588600.0 1152000.0 598800.0 1165800.0 ;
      RECT  588600.0 1179600.0 598800.0 1165800.0 ;
      RECT  588600.0 1179600.0 598800.0 1193400.0 ;
      RECT  588600.0 1207200.0 598800.0 1193400.0 ;
      RECT  588600.0 1207200.0 598800.0 1221000.0 ;
      RECT  588600.0 1234800.0 598800.0 1221000.0 ;
      RECT  588600.0 1234800.0 598800.0 1248600.0 ;
      RECT  588600.0 1262400.0 598800.0 1248600.0 ;
      RECT  588600.0 1262400.0 598800.0 1276200.0 ;
      RECT  588600.0 1290000.0 598800.0 1276200.0 ;
      RECT  588600.0 1290000.0 598800.0 1303800.0 ;
      RECT  588600.0 1317600.0 598800.0 1303800.0 ;
      RECT  588600.0 1317600.0 598800.0 1331400.0 ;
      RECT  588600.0 1345200.0 598800.0 1331400.0 ;
      RECT  588600.0 1345200.0 598800.0 1359000.0 ;
      RECT  588600.0 1372800.0 598800.0 1359000.0 ;
      RECT  588600.0 1372800.0 598800.0 1386600.0 ;
      RECT  588600.0 1400400.0 598800.0 1386600.0 ;
      RECT  588600.0 1400400.0 598800.0 1414200.0 ;
      RECT  588600.0 1428000.0 598800.0 1414200.0 ;
      RECT  588600.0 1428000.0 598800.0 1441800.0 ;
      RECT  588600.0 1455600.0 598800.0 1441800.0 ;
      RECT  588600.0 1455600.0 598800.0 1469400.0 ;
      RECT  588600.0 1483200.0 598800.0 1469400.0 ;
      RECT  588600.0 1483200.0 598800.0 1497000.0 ;
      RECT  588600.0 1510800.0 598800.0 1497000.0 ;
      RECT  588600.0 1510800.0 598800.0 1524600.0 ;
      RECT  588600.0 1538400.0 598800.0 1524600.0 ;
      RECT  588600.0 1538400.0 598800.0 1552200.0 ;
      RECT  588600.0 1566000.0 598800.0 1552200.0 ;
      RECT  588600.0 1566000.0 598800.0 1579800.0 ;
      RECT  588600.0 1593600.0 598800.0 1579800.0 ;
      RECT  588600.0 1593600.0 598800.0 1607400.0 ;
      RECT  588600.0 1621200.0 598800.0 1607400.0 ;
      RECT  588600.0 1621200.0 598800.0 1635000.0 ;
      RECT  588600.0 1648800.0 598800.0 1635000.0 ;
      RECT  588600.0 1648800.0 598800.0 1662600.0 ;
      RECT  588600.0 1676400.0 598800.0 1662600.0 ;
      RECT  588600.0 1676400.0 598800.0 1690200.0 ;
      RECT  588600.0 1704000.0 598800.0 1690200.0 ;
      RECT  588600.0 1704000.0 598800.0 1717800.0 ;
      RECT  588600.0 1731600.0 598800.0 1717800.0 ;
      RECT  588600.0 1731600.0 598800.0 1745400.0 ;
      RECT  588600.0 1759200.0 598800.0 1745400.0 ;
      RECT  588600.0 1759200.0 598800.0 1773000.0 ;
      RECT  588600.0 1786800.0 598800.0 1773000.0 ;
      RECT  588600.0 1786800.0 598800.0 1800600.0 ;
      RECT  588600.0 1814400.0 598800.0 1800600.0 ;
      RECT  588600.0 1814400.0 598800.0 1828200.0 ;
      RECT  588600.0 1842000.0 598800.0 1828200.0 ;
      RECT  588600.0 1842000.0 598800.0 1855800.0 ;
      RECT  588600.0 1869600.0 598800.0 1855800.0 ;
      RECT  588600.0 1869600.0 598800.0 1883400.0 ;
      RECT  588600.0 1897200.0 598800.0 1883400.0 ;
      RECT  588600.0 1897200.0 598800.0 1911000.0 ;
      RECT  588600.0 1924800.0 598800.0 1911000.0 ;
      RECT  588600.0 1924800.0 598800.0 1938600.0 ;
      RECT  588600.0 1952400.0 598800.0 1938600.0 ;
      RECT  588600.0 1952400.0 598800.0 1966200.0 ;
      RECT  588600.0 1980000.0 598800.0 1966200.0 ;
      RECT  588600.0 1980000.0 598800.0 1993800.0 ;
      RECT  588600.0 2007600.0 598800.0 1993800.0 ;
      RECT  588600.0 2007600.0 598800.0 2021400.0 ;
      RECT  588600.0 2035200.0 598800.0 2021400.0 ;
      RECT  588600.0 2035200.0 598800.0 2049000.0 ;
      RECT  588600.0 2062800.0 598800.0 2049000.0 ;
      RECT  588600.0 2062800.0 598800.0 2076600.0 ;
      RECT  588600.0 2090400.0 598800.0 2076600.0 ;
      RECT  588600.0 2090400.0 598800.0 2104200.0 ;
      RECT  588600.0 2118000.0 598800.0 2104200.0 ;
      RECT  588600.0 2118000.0 598800.0 2131800.0 ;
      RECT  588600.0 2145600.0 598800.0 2131800.0 ;
      RECT  598800.0 379200.0 609000.0 393000.0 ;
      RECT  598800.0 406800.0 609000.0 393000.0 ;
      RECT  598800.0 406800.0 609000.0 420600.0 ;
      RECT  598800.0 434400.0 609000.0 420600.0 ;
      RECT  598800.0 434400.0 609000.0 448200.0 ;
      RECT  598800.0 462000.0 609000.0 448200.0 ;
      RECT  598800.0 462000.0 609000.0 475800.0 ;
      RECT  598800.0 489600.0 609000.0 475800.0 ;
      RECT  598800.0 489600.0 609000.0 503400.0 ;
      RECT  598800.0 517200.0 609000.0 503400.0 ;
      RECT  598800.0 517200.0 609000.0 531000.0 ;
      RECT  598800.0 544800.0 609000.0 531000.0 ;
      RECT  598800.0 544800.0 609000.0 558600.0 ;
      RECT  598800.0 572400.0 609000.0 558600.0 ;
      RECT  598800.0 572400.0 609000.0 586200.0 ;
      RECT  598800.0 600000.0 609000.0 586200.0 ;
      RECT  598800.0 600000.0 609000.0 613800.0 ;
      RECT  598800.0 627600.0 609000.0 613800.0 ;
      RECT  598800.0 627600.0 609000.0 641400.0 ;
      RECT  598800.0 655200.0 609000.0 641400.0 ;
      RECT  598800.0 655200.0 609000.0 669000.0 ;
      RECT  598800.0 682800.0 609000.0 669000.0 ;
      RECT  598800.0 682800.0 609000.0 696600.0 ;
      RECT  598800.0 710400.0 609000.0 696600.0 ;
      RECT  598800.0 710400.0 609000.0 724200.0 ;
      RECT  598800.0 738000.0 609000.0 724200.0 ;
      RECT  598800.0 738000.0 609000.0 751800.0 ;
      RECT  598800.0 765600.0 609000.0 751800.0 ;
      RECT  598800.0 765600.0 609000.0 779400.0 ;
      RECT  598800.0 793200.0 609000.0 779400.0 ;
      RECT  598800.0 793200.0 609000.0 807000.0 ;
      RECT  598800.0 820800.0 609000.0 807000.0 ;
      RECT  598800.0 820800.0 609000.0 834600.0 ;
      RECT  598800.0 848400.0 609000.0 834600.0 ;
      RECT  598800.0 848400.0 609000.0 862200.0 ;
      RECT  598800.0 876000.0 609000.0 862200.0 ;
      RECT  598800.0 876000.0 609000.0 889800.0 ;
      RECT  598800.0 903600.0 609000.0 889800.0 ;
      RECT  598800.0 903600.0 609000.0 917400.0 ;
      RECT  598800.0 931200.0 609000.0 917400.0 ;
      RECT  598800.0 931200.0 609000.0 945000.0 ;
      RECT  598800.0 958800.0 609000.0 945000.0 ;
      RECT  598800.0 958800.0 609000.0 972600.0 ;
      RECT  598800.0 986400.0 609000.0 972600.0 ;
      RECT  598800.0 986400.0 609000.0 1000200.0 ;
      RECT  598800.0 1014000.0 609000.0 1000200.0 ;
      RECT  598800.0 1014000.0 609000.0 1027800.0 ;
      RECT  598800.0 1041600.0 609000.0 1027800.0 ;
      RECT  598800.0 1041600.0 609000.0 1055400.0 ;
      RECT  598800.0 1069200.0 609000.0 1055400.0 ;
      RECT  598800.0 1069200.0 609000.0 1083000.0 ;
      RECT  598800.0 1096800.0 609000.0 1083000.0 ;
      RECT  598800.0 1096800.0 609000.0 1110600.0 ;
      RECT  598800.0 1124400.0 609000.0 1110600.0 ;
      RECT  598800.0 1124400.0 609000.0 1138200.0 ;
      RECT  598800.0 1152000.0 609000.0 1138200.0 ;
      RECT  598800.0 1152000.0 609000.0 1165800.0 ;
      RECT  598800.0 1179600.0 609000.0 1165800.0 ;
      RECT  598800.0 1179600.0 609000.0 1193400.0 ;
      RECT  598800.0 1207200.0 609000.0 1193400.0 ;
      RECT  598800.0 1207200.0 609000.0 1221000.0 ;
      RECT  598800.0 1234800.0 609000.0 1221000.0 ;
      RECT  598800.0 1234800.0 609000.0 1248600.0 ;
      RECT  598800.0 1262400.0 609000.0 1248600.0 ;
      RECT  598800.0 1262400.0 609000.0 1276200.0 ;
      RECT  598800.0 1290000.0 609000.0 1276200.0 ;
      RECT  598800.0 1290000.0 609000.0 1303800.0 ;
      RECT  598800.0 1317600.0 609000.0 1303800.0 ;
      RECT  598800.0 1317600.0 609000.0 1331400.0 ;
      RECT  598800.0 1345200.0 609000.0 1331400.0 ;
      RECT  598800.0 1345200.0 609000.0 1359000.0 ;
      RECT  598800.0 1372800.0 609000.0 1359000.0 ;
      RECT  598800.0 1372800.0 609000.0 1386600.0 ;
      RECT  598800.0 1400400.0 609000.0 1386600.0 ;
      RECT  598800.0 1400400.0 609000.0 1414200.0 ;
      RECT  598800.0 1428000.0 609000.0 1414200.0 ;
      RECT  598800.0 1428000.0 609000.0 1441800.0 ;
      RECT  598800.0 1455600.0 609000.0 1441800.0 ;
      RECT  598800.0 1455600.0 609000.0 1469400.0 ;
      RECT  598800.0 1483200.0 609000.0 1469400.0 ;
      RECT  598800.0 1483200.0 609000.0 1497000.0 ;
      RECT  598800.0 1510800.0 609000.0 1497000.0 ;
      RECT  598800.0 1510800.0 609000.0 1524600.0 ;
      RECT  598800.0 1538400.0 609000.0 1524600.0 ;
      RECT  598800.0 1538400.0 609000.0 1552200.0 ;
      RECT  598800.0 1566000.0 609000.0 1552200.0 ;
      RECT  598800.0 1566000.0 609000.0 1579800.0 ;
      RECT  598800.0 1593600.0 609000.0 1579800.0 ;
      RECT  598800.0 1593600.0 609000.0 1607400.0 ;
      RECT  598800.0 1621200.0 609000.0 1607400.0 ;
      RECT  598800.0 1621200.0 609000.0 1635000.0 ;
      RECT  598800.0 1648800.0 609000.0 1635000.0 ;
      RECT  598800.0 1648800.0 609000.0 1662600.0 ;
      RECT  598800.0 1676400.0 609000.0 1662600.0 ;
      RECT  598800.0 1676400.0 609000.0 1690200.0 ;
      RECT  598800.0 1704000.0 609000.0 1690200.0 ;
      RECT  598800.0 1704000.0 609000.0 1717800.0 ;
      RECT  598800.0 1731600.0 609000.0 1717800.0 ;
      RECT  598800.0 1731600.0 609000.0 1745400.0 ;
      RECT  598800.0 1759200.0 609000.0 1745400.0 ;
      RECT  598800.0 1759200.0 609000.0 1773000.0 ;
      RECT  598800.0 1786800.0 609000.0 1773000.0 ;
      RECT  598800.0 1786800.0 609000.0 1800600.0 ;
      RECT  598800.0 1814400.0 609000.0 1800600.0 ;
      RECT  598800.0 1814400.0 609000.0 1828200.0 ;
      RECT  598800.0 1842000.0 609000.0 1828200.0 ;
      RECT  598800.0 1842000.0 609000.0 1855800.0 ;
      RECT  598800.0 1869600.0 609000.0 1855800.0 ;
      RECT  598800.0 1869600.0 609000.0 1883400.0 ;
      RECT  598800.0 1897200.0 609000.0 1883400.0 ;
      RECT  598800.0 1897200.0 609000.0 1911000.0 ;
      RECT  598800.0 1924800.0 609000.0 1911000.0 ;
      RECT  598800.0 1924800.0 609000.0 1938600.0 ;
      RECT  598800.0 1952400.0 609000.0 1938600.0 ;
      RECT  598800.0 1952400.0 609000.0 1966200.0 ;
      RECT  598800.0 1980000.0 609000.0 1966200.0 ;
      RECT  598800.0 1980000.0 609000.0 1993800.0 ;
      RECT  598800.0 2007600.0 609000.0 1993800.0 ;
      RECT  598800.0 2007600.0 609000.0 2021400.0 ;
      RECT  598800.0 2035200.0 609000.0 2021400.0 ;
      RECT  598800.0 2035200.0 609000.0 2049000.0 ;
      RECT  598800.0 2062800.0 609000.0 2049000.0 ;
      RECT  598800.0 2062800.0 609000.0 2076600.0 ;
      RECT  598800.0 2090400.0 609000.0 2076600.0 ;
      RECT  598800.0 2090400.0 609000.0 2104200.0 ;
      RECT  598800.0 2118000.0 609000.0 2104200.0 ;
      RECT  598800.0 2118000.0 609000.0 2131800.0 ;
      RECT  598800.0 2145600.0 609000.0 2131800.0 ;
      RECT  609000.0 379200.0 619200.0 393000.0 ;
      RECT  609000.0 406800.0 619200.0 393000.0 ;
      RECT  609000.0 406800.0 619200.0 420600.0 ;
      RECT  609000.0 434400.0 619200.0 420600.0 ;
      RECT  609000.0 434400.0 619200.0 448200.0 ;
      RECT  609000.0 462000.0 619200.0 448200.0 ;
      RECT  609000.0 462000.0 619200.0 475800.0 ;
      RECT  609000.0 489600.0 619200.0 475800.0 ;
      RECT  609000.0 489600.0 619200.0 503400.0 ;
      RECT  609000.0 517200.0 619200.0 503400.0 ;
      RECT  609000.0 517200.0 619200.0 531000.0 ;
      RECT  609000.0 544800.0 619200.0 531000.0 ;
      RECT  609000.0 544800.0 619200.0 558600.0 ;
      RECT  609000.0 572400.0 619200.0 558600.0 ;
      RECT  609000.0 572400.0 619200.0 586200.0 ;
      RECT  609000.0 600000.0 619200.0 586200.0 ;
      RECT  609000.0 600000.0 619200.0 613800.0 ;
      RECT  609000.0 627600.0 619200.0 613800.0 ;
      RECT  609000.0 627600.0 619200.0 641400.0 ;
      RECT  609000.0 655200.0 619200.0 641400.0 ;
      RECT  609000.0 655200.0 619200.0 669000.0 ;
      RECT  609000.0 682800.0 619200.0 669000.0 ;
      RECT  609000.0 682800.0 619200.0 696600.0 ;
      RECT  609000.0 710400.0 619200.0 696600.0 ;
      RECT  609000.0 710400.0 619200.0 724200.0 ;
      RECT  609000.0 738000.0 619200.0 724200.0 ;
      RECT  609000.0 738000.0 619200.0 751800.0 ;
      RECT  609000.0 765600.0 619200.0 751800.0 ;
      RECT  609000.0 765600.0 619200.0 779400.0 ;
      RECT  609000.0 793200.0 619200.0 779400.0 ;
      RECT  609000.0 793200.0 619200.0 807000.0 ;
      RECT  609000.0 820800.0 619200.0 807000.0 ;
      RECT  609000.0 820800.0 619200.0 834600.0 ;
      RECT  609000.0 848400.0 619200.0 834600.0 ;
      RECT  609000.0 848400.0 619200.0 862200.0 ;
      RECT  609000.0 876000.0 619200.0 862200.0 ;
      RECT  609000.0 876000.0 619200.0 889800.0 ;
      RECT  609000.0 903600.0 619200.0 889800.0 ;
      RECT  609000.0 903600.0 619200.0 917400.0 ;
      RECT  609000.0 931200.0 619200.0 917400.0 ;
      RECT  609000.0 931200.0 619200.0 945000.0 ;
      RECT  609000.0 958800.0 619200.0 945000.0 ;
      RECT  609000.0 958800.0 619200.0 972600.0 ;
      RECT  609000.0 986400.0 619200.0 972600.0 ;
      RECT  609000.0 986400.0 619200.0 1000200.0 ;
      RECT  609000.0 1014000.0 619200.0 1000200.0 ;
      RECT  609000.0 1014000.0 619200.0 1027800.0 ;
      RECT  609000.0 1041600.0 619200.0 1027800.0 ;
      RECT  609000.0 1041600.0 619200.0 1055400.0 ;
      RECT  609000.0 1069200.0 619200.0 1055400.0 ;
      RECT  609000.0 1069200.0 619200.0 1083000.0 ;
      RECT  609000.0 1096800.0 619200.0 1083000.0 ;
      RECT  609000.0 1096800.0 619200.0 1110600.0 ;
      RECT  609000.0 1124400.0 619200.0 1110600.0 ;
      RECT  609000.0 1124400.0 619200.0 1138200.0 ;
      RECT  609000.0 1152000.0 619200.0 1138200.0 ;
      RECT  609000.0 1152000.0 619200.0 1165800.0 ;
      RECT  609000.0 1179600.0 619200.0 1165800.0 ;
      RECT  609000.0 1179600.0 619200.0 1193400.0 ;
      RECT  609000.0 1207200.0 619200.0 1193400.0 ;
      RECT  609000.0 1207200.0 619200.0 1221000.0 ;
      RECT  609000.0 1234800.0 619200.0 1221000.0 ;
      RECT  609000.0 1234800.0 619200.0 1248600.0 ;
      RECT  609000.0 1262400.0 619200.0 1248600.0 ;
      RECT  609000.0 1262400.0 619200.0 1276200.0 ;
      RECT  609000.0 1290000.0 619200.0 1276200.0 ;
      RECT  609000.0 1290000.0 619200.0 1303800.0 ;
      RECT  609000.0 1317600.0 619200.0 1303800.0 ;
      RECT  609000.0 1317600.0 619200.0 1331400.0 ;
      RECT  609000.0 1345200.0 619200.0 1331400.0 ;
      RECT  609000.0 1345200.0 619200.0 1359000.0 ;
      RECT  609000.0 1372800.0 619200.0 1359000.0 ;
      RECT  609000.0 1372800.0 619200.0 1386600.0 ;
      RECT  609000.0 1400400.0 619200.0 1386600.0 ;
      RECT  609000.0 1400400.0 619200.0 1414200.0 ;
      RECT  609000.0 1428000.0 619200.0 1414200.0 ;
      RECT  609000.0 1428000.0 619200.0 1441800.0 ;
      RECT  609000.0 1455600.0 619200.0 1441800.0 ;
      RECT  609000.0 1455600.0 619200.0 1469400.0 ;
      RECT  609000.0 1483200.0 619200.0 1469400.0 ;
      RECT  609000.0 1483200.0 619200.0 1497000.0 ;
      RECT  609000.0 1510800.0 619200.0 1497000.0 ;
      RECT  609000.0 1510800.0 619200.0 1524600.0 ;
      RECT  609000.0 1538400.0 619200.0 1524600.0 ;
      RECT  609000.0 1538400.0 619200.0 1552200.0 ;
      RECT  609000.0 1566000.0 619200.0 1552200.0 ;
      RECT  609000.0 1566000.0 619200.0 1579800.0 ;
      RECT  609000.0 1593600.0 619200.0 1579800.0 ;
      RECT  609000.0 1593600.0 619200.0 1607400.0 ;
      RECT  609000.0 1621200.0 619200.0 1607400.0 ;
      RECT  609000.0 1621200.0 619200.0 1635000.0 ;
      RECT  609000.0 1648800.0 619200.0 1635000.0 ;
      RECT  609000.0 1648800.0 619200.0 1662600.0 ;
      RECT  609000.0 1676400.0 619200.0 1662600.0 ;
      RECT  609000.0 1676400.0 619200.0 1690200.0 ;
      RECT  609000.0 1704000.0 619200.0 1690200.0 ;
      RECT  609000.0 1704000.0 619200.0 1717800.0 ;
      RECT  609000.0 1731600.0 619200.0 1717800.0 ;
      RECT  609000.0 1731600.0 619200.0 1745400.0 ;
      RECT  609000.0 1759200.0 619200.0 1745400.0 ;
      RECT  609000.0 1759200.0 619200.0 1773000.0 ;
      RECT  609000.0 1786800.0 619200.0 1773000.0 ;
      RECT  609000.0 1786800.0 619200.0 1800600.0 ;
      RECT  609000.0 1814400.0 619200.0 1800600.0 ;
      RECT  609000.0 1814400.0 619200.0 1828200.0 ;
      RECT  609000.0 1842000.0 619200.0 1828200.0 ;
      RECT  609000.0 1842000.0 619200.0 1855800.0 ;
      RECT  609000.0 1869600.0 619200.0 1855800.0 ;
      RECT  609000.0 1869600.0 619200.0 1883400.0 ;
      RECT  609000.0 1897200.0 619200.0 1883400.0 ;
      RECT  609000.0 1897200.0 619200.0 1911000.0 ;
      RECT  609000.0 1924800.0 619200.0 1911000.0 ;
      RECT  609000.0 1924800.0 619200.0 1938600.0 ;
      RECT  609000.0 1952400.0 619200.0 1938600.0 ;
      RECT  609000.0 1952400.0 619200.0 1966200.0 ;
      RECT  609000.0 1980000.0 619200.0 1966200.0 ;
      RECT  609000.0 1980000.0 619200.0 1993800.0 ;
      RECT  609000.0 2007600.0 619200.0 1993800.0 ;
      RECT  609000.0 2007600.0 619200.0 2021400.0 ;
      RECT  609000.0 2035200.0 619200.0 2021400.0 ;
      RECT  609000.0 2035200.0 619200.0 2049000.0 ;
      RECT  609000.0 2062800.0 619200.0 2049000.0 ;
      RECT  609000.0 2062800.0 619200.0 2076600.0 ;
      RECT  609000.0 2090400.0 619200.0 2076600.0 ;
      RECT  609000.0 2090400.0 619200.0 2104200.0 ;
      RECT  609000.0 2118000.0 619200.0 2104200.0 ;
      RECT  609000.0 2118000.0 619200.0 2131800.0 ;
      RECT  609000.0 2145600.0 619200.0 2131800.0 ;
      RECT  619200.0 379200.0 629400.0 393000.0 ;
      RECT  619200.0 406800.0 629400.0 393000.0 ;
      RECT  619200.0 406800.0 629400.0 420600.0 ;
      RECT  619200.0 434400.0 629400.0 420600.0 ;
      RECT  619200.0 434400.0 629400.0 448200.0 ;
      RECT  619200.0 462000.0 629400.0 448200.0 ;
      RECT  619200.0 462000.0 629400.0 475800.0 ;
      RECT  619200.0 489600.0 629400.0 475800.0 ;
      RECT  619200.0 489600.0 629400.0 503400.0 ;
      RECT  619200.0 517200.0 629400.0 503400.0 ;
      RECT  619200.0 517200.0 629400.0 531000.0 ;
      RECT  619200.0 544800.0 629400.0 531000.0 ;
      RECT  619200.0 544800.0 629400.0 558600.0 ;
      RECT  619200.0 572400.0 629400.0 558600.0 ;
      RECT  619200.0 572400.0 629400.0 586200.0 ;
      RECT  619200.0 600000.0 629400.0 586200.0 ;
      RECT  619200.0 600000.0 629400.0 613800.0 ;
      RECT  619200.0 627600.0 629400.0 613800.0 ;
      RECT  619200.0 627600.0 629400.0 641400.0 ;
      RECT  619200.0 655200.0 629400.0 641400.0 ;
      RECT  619200.0 655200.0 629400.0 669000.0 ;
      RECT  619200.0 682800.0 629400.0 669000.0 ;
      RECT  619200.0 682800.0 629400.0 696600.0 ;
      RECT  619200.0 710400.0 629400.0 696600.0 ;
      RECT  619200.0 710400.0 629400.0 724200.0 ;
      RECT  619200.0 738000.0 629400.0 724200.0 ;
      RECT  619200.0 738000.0 629400.0 751800.0 ;
      RECT  619200.0 765600.0 629400.0 751800.0 ;
      RECT  619200.0 765600.0 629400.0 779400.0 ;
      RECT  619200.0 793200.0 629400.0 779400.0 ;
      RECT  619200.0 793200.0 629400.0 807000.0 ;
      RECT  619200.0 820800.0 629400.0 807000.0 ;
      RECT  619200.0 820800.0 629400.0 834600.0 ;
      RECT  619200.0 848400.0 629400.0 834600.0 ;
      RECT  619200.0 848400.0 629400.0 862200.0 ;
      RECT  619200.0 876000.0 629400.0 862200.0 ;
      RECT  619200.0 876000.0 629400.0 889800.0 ;
      RECT  619200.0 903600.0 629400.0 889800.0 ;
      RECT  619200.0 903600.0 629400.0 917400.0 ;
      RECT  619200.0 931200.0 629400.0 917400.0 ;
      RECT  619200.0 931200.0 629400.0 945000.0 ;
      RECT  619200.0 958800.0 629400.0 945000.0 ;
      RECT  619200.0 958800.0 629400.0 972600.0 ;
      RECT  619200.0 986400.0 629400.0 972600.0 ;
      RECT  619200.0 986400.0 629400.0 1000200.0 ;
      RECT  619200.0 1014000.0 629400.0 1000200.0 ;
      RECT  619200.0 1014000.0 629400.0 1027800.0 ;
      RECT  619200.0 1041600.0 629400.0 1027800.0 ;
      RECT  619200.0 1041600.0 629400.0 1055400.0 ;
      RECT  619200.0 1069200.0 629400.0 1055400.0 ;
      RECT  619200.0 1069200.0 629400.0 1083000.0 ;
      RECT  619200.0 1096800.0 629400.0 1083000.0 ;
      RECT  619200.0 1096800.0 629400.0 1110600.0 ;
      RECT  619200.0 1124400.0 629400.0 1110600.0 ;
      RECT  619200.0 1124400.0 629400.0 1138200.0 ;
      RECT  619200.0 1152000.0 629400.0 1138200.0 ;
      RECT  619200.0 1152000.0 629400.0 1165800.0 ;
      RECT  619200.0 1179600.0 629400.0 1165800.0 ;
      RECT  619200.0 1179600.0 629400.0 1193400.0 ;
      RECT  619200.0 1207200.0 629400.0 1193400.0 ;
      RECT  619200.0 1207200.0 629400.0 1221000.0 ;
      RECT  619200.0 1234800.0 629400.0 1221000.0 ;
      RECT  619200.0 1234800.0 629400.0 1248600.0 ;
      RECT  619200.0 1262400.0 629400.0 1248600.0 ;
      RECT  619200.0 1262400.0 629400.0 1276200.0 ;
      RECT  619200.0 1290000.0 629400.0 1276200.0 ;
      RECT  619200.0 1290000.0 629400.0 1303800.0 ;
      RECT  619200.0 1317600.0 629400.0 1303800.0 ;
      RECT  619200.0 1317600.0 629400.0 1331400.0 ;
      RECT  619200.0 1345200.0 629400.0 1331400.0 ;
      RECT  619200.0 1345200.0 629400.0 1359000.0 ;
      RECT  619200.0 1372800.0 629400.0 1359000.0 ;
      RECT  619200.0 1372800.0 629400.0 1386600.0 ;
      RECT  619200.0 1400400.0 629400.0 1386600.0 ;
      RECT  619200.0 1400400.0 629400.0 1414200.0 ;
      RECT  619200.0 1428000.0 629400.0 1414200.0 ;
      RECT  619200.0 1428000.0 629400.0 1441800.0 ;
      RECT  619200.0 1455600.0 629400.0 1441800.0 ;
      RECT  619200.0 1455600.0 629400.0 1469400.0 ;
      RECT  619200.0 1483200.0 629400.0 1469400.0 ;
      RECT  619200.0 1483200.0 629400.0 1497000.0 ;
      RECT  619200.0 1510800.0 629400.0 1497000.0 ;
      RECT  619200.0 1510800.0 629400.0 1524600.0 ;
      RECT  619200.0 1538400.0 629400.0 1524600.0 ;
      RECT  619200.0 1538400.0 629400.0 1552200.0 ;
      RECT  619200.0 1566000.0 629400.0 1552200.0 ;
      RECT  619200.0 1566000.0 629400.0 1579800.0 ;
      RECT  619200.0 1593600.0 629400.0 1579800.0 ;
      RECT  619200.0 1593600.0 629400.0 1607400.0 ;
      RECT  619200.0 1621200.0 629400.0 1607400.0 ;
      RECT  619200.0 1621200.0 629400.0 1635000.0 ;
      RECT  619200.0 1648800.0 629400.0 1635000.0 ;
      RECT  619200.0 1648800.0 629400.0 1662600.0 ;
      RECT  619200.0 1676400.0 629400.0 1662600.0 ;
      RECT  619200.0 1676400.0 629400.0 1690200.0 ;
      RECT  619200.0 1704000.0 629400.0 1690200.0 ;
      RECT  619200.0 1704000.0 629400.0 1717800.0 ;
      RECT  619200.0 1731600.0 629400.0 1717800.0 ;
      RECT  619200.0 1731600.0 629400.0 1745400.0 ;
      RECT  619200.0 1759200.0 629400.0 1745400.0 ;
      RECT  619200.0 1759200.0 629400.0 1773000.0 ;
      RECT  619200.0 1786800.0 629400.0 1773000.0 ;
      RECT  619200.0 1786800.0 629400.0 1800600.0 ;
      RECT  619200.0 1814400.0 629400.0 1800600.0 ;
      RECT  619200.0 1814400.0 629400.0 1828200.0 ;
      RECT  619200.0 1842000.0 629400.0 1828200.0 ;
      RECT  619200.0 1842000.0 629400.0 1855800.0 ;
      RECT  619200.0 1869600.0 629400.0 1855800.0 ;
      RECT  619200.0 1869600.0 629400.0 1883400.0 ;
      RECT  619200.0 1897200.0 629400.0 1883400.0 ;
      RECT  619200.0 1897200.0 629400.0 1911000.0 ;
      RECT  619200.0 1924800.0 629400.0 1911000.0 ;
      RECT  619200.0 1924800.0 629400.0 1938600.0 ;
      RECT  619200.0 1952400.0 629400.0 1938600.0 ;
      RECT  619200.0 1952400.0 629400.0 1966200.0 ;
      RECT  619200.0 1980000.0 629400.0 1966200.0 ;
      RECT  619200.0 1980000.0 629400.0 1993800.0 ;
      RECT  619200.0 2007600.0 629400.0 1993800.0 ;
      RECT  619200.0 2007600.0 629400.0 2021400.0 ;
      RECT  619200.0 2035200.0 629400.0 2021400.0 ;
      RECT  619200.0 2035200.0 629400.0 2049000.0 ;
      RECT  619200.0 2062800.0 629400.0 2049000.0 ;
      RECT  619200.0 2062800.0 629400.0 2076600.0 ;
      RECT  619200.0 2090400.0 629400.0 2076600.0 ;
      RECT  619200.0 2090400.0 629400.0 2104200.0 ;
      RECT  619200.0 2118000.0 629400.0 2104200.0 ;
      RECT  619200.0 2118000.0 629400.0 2131800.0 ;
      RECT  619200.0 2145600.0 629400.0 2131800.0 ;
      RECT  629400.0 379200.0 639600.0 393000.0 ;
      RECT  629400.0 406800.0 639600.0 393000.0 ;
      RECT  629400.0 406800.0 639600.0 420600.0 ;
      RECT  629400.0 434400.0 639600.0 420600.0 ;
      RECT  629400.0 434400.0 639600.0 448200.0 ;
      RECT  629400.0 462000.0 639600.0 448200.0 ;
      RECT  629400.0 462000.0 639600.0 475800.0 ;
      RECT  629400.0 489600.0 639600.0 475800.0 ;
      RECT  629400.0 489600.0 639600.0 503400.0 ;
      RECT  629400.0 517200.0 639600.0 503400.0 ;
      RECT  629400.0 517200.0 639600.0 531000.0 ;
      RECT  629400.0 544800.0 639600.0 531000.0 ;
      RECT  629400.0 544800.0 639600.0 558600.0 ;
      RECT  629400.0 572400.0 639600.0 558600.0 ;
      RECT  629400.0 572400.0 639600.0 586200.0 ;
      RECT  629400.0 600000.0 639600.0 586200.0 ;
      RECT  629400.0 600000.0 639600.0 613800.0 ;
      RECT  629400.0 627600.0 639600.0 613800.0 ;
      RECT  629400.0 627600.0 639600.0 641400.0 ;
      RECT  629400.0 655200.0 639600.0 641400.0 ;
      RECT  629400.0 655200.0 639600.0 669000.0 ;
      RECT  629400.0 682800.0 639600.0 669000.0 ;
      RECT  629400.0 682800.0 639600.0 696600.0 ;
      RECT  629400.0 710400.0 639600.0 696600.0 ;
      RECT  629400.0 710400.0 639600.0 724200.0 ;
      RECT  629400.0 738000.0 639600.0 724200.0 ;
      RECT  629400.0 738000.0 639600.0 751800.0 ;
      RECT  629400.0 765600.0 639600.0 751800.0 ;
      RECT  629400.0 765600.0 639600.0 779400.0 ;
      RECT  629400.0 793200.0 639600.0 779400.0 ;
      RECT  629400.0 793200.0 639600.0 807000.0 ;
      RECT  629400.0 820800.0 639600.0 807000.0 ;
      RECT  629400.0 820800.0 639600.0 834600.0 ;
      RECT  629400.0 848400.0 639600.0 834600.0 ;
      RECT  629400.0 848400.0 639600.0 862200.0 ;
      RECT  629400.0 876000.0 639600.0 862200.0 ;
      RECT  629400.0 876000.0 639600.0 889800.0 ;
      RECT  629400.0 903600.0 639600.0 889800.0 ;
      RECT  629400.0 903600.0 639600.0 917400.0 ;
      RECT  629400.0 931200.0 639600.0 917400.0 ;
      RECT  629400.0 931200.0 639600.0 945000.0 ;
      RECT  629400.0 958800.0 639600.0 945000.0 ;
      RECT  629400.0 958800.0 639600.0 972600.0 ;
      RECT  629400.0 986400.0 639600.0 972600.0 ;
      RECT  629400.0 986400.0 639600.0 1000200.0 ;
      RECT  629400.0 1014000.0 639600.0 1000200.0 ;
      RECT  629400.0 1014000.0 639600.0 1027800.0 ;
      RECT  629400.0 1041600.0 639600.0 1027800.0 ;
      RECT  629400.0 1041600.0 639600.0 1055400.0 ;
      RECT  629400.0 1069200.0 639600.0 1055400.0 ;
      RECT  629400.0 1069200.0 639600.0 1083000.0 ;
      RECT  629400.0 1096800.0 639600.0 1083000.0 ;
      RECT  629400.0 1096800.0 639600.0 1110600.0 ;
      RECT  629400.0 1124400.0 639600.0 1110600.0 ;
      RECT  629400.0 1124400.0 639600.0 1138200.0 ;
      RECT  629400.0 1152000.0 639600.0 1138200.0 ;
      RECT  629400.0 1152000.0 639600.0 1165800.0 ;
      RECT  629400.0 1179600.0 639600.0 1165800.0 ;
      RECT  629400.0 1179600.0 639600.0 1193400.0 ;
      RECT  629400.0 1207200.0 639600.0 1193400.0 ;
      RECT  629400.0 1207200.0 639600.0 1221000.0 ;
      RECT  629400.0 1234800.0 639600.0 1221000.0 ;
      RECT  629400.0 1234800.0 639600.0 1248600.0 ;
      RECT  629400.0 1262400.0 639600.0 1248600.0 ;
      RECT  629400.0 1262400.0 639600.0 1276200.0 ;
      RECT  629400.0 1290000.0 639600.0 1276200.0 ;
      RECT  629400.0 1290000.0 639600.0 1303800.0 ;
      RECT  629400.0 1317600.0 639600.0 1303800.0 ;
      RECT  629400.0 1317600.0 639600.0 1331400.0 ;
      RECT  629400.0 1345200.0 639600.0 1331400.0 ;
      RECT  629400.0 1345200.0 639600.0 1359000.0 ;
      RECT  629400.0 1372800.0 639600.0 1359000.0 ;
      RECT  629400.0 1372800.0 639600.0 1386600.0 ;
      RECT  629400.0 1400400.0 639600.0 1386600.0 ;
      RECT  629400.0 1400400.0 639600.0 1414200.0 ;
      RECT  629400.0 1428000.0 639600.0 1414200.0 ;
      RECT  629400.0 1428000.0 639600.0 1441800.0 ;
      RECT  629400.0 1455600.0 639600.0 1441800.0 ;
      RECT  629400.0 1455600.0 639600.0 1469400.0 ;
      RECT  629400.0 1483200.0 639600.0 1469400.0 ;
      RECT  629400.0 1483200.0 639600.0 1497000.0 ;
      RECT  629400.0 1510800.0 639600.0 1497000.0 ;
      RECT  629400.0 1510800.0 639600.0 1524600.0 ;
      RECT  629400.0 1538400.0 639600.0 1524600.0 ;
      RECT  629400.0 1538400.0 639600.0 1552200.0 ;
      RECT  629400.0 1566000.0 639600.0 1552200.0 ;
      RECT  629400.0 1566000.0 639600.0 1579800.0 ;
      RECT  629400.0 1593600.0 639600.0 1579800.0 ;
      RECT  629400.0 1593600.0 639600.0 1607400.0 ;
      RECT  629400.0 1621200.0 639600.0 1607400.0 ;
      RECT  629400.0 1621200.0 639600.0 1635000.0 ;
      RECT  629400.0 1648800.0 639600.0 1635000.0 ;
      RECT  629400.0 1648800.0 639600.0 1662600.0 ;
      RECT  629400.0 1676400.0 639600.0 1662600.0 ;
      RECT  629400.0 1676400.0 639600.0 1690200.0 ;
      RECT  629400.0 1704000.0 639600.0 1690200.0 ;
      RECT  629400.0 1704000.0 639600.0 1717800.0 ;
      RECT  629400.0 1731600.0 639600.0 1717800.0 ;
      RECT  629400.0 1731600.0 639600.0 1745400.0 ;
      RECT  629400.0 1759200.0 639600.0 1745400.0 ;
      RECT  629400.0 1759200.0 639600.0 1773000.0 ;
      RECT  629400.0 1786800.0 639600.0 1773000.0 ;
      RECT  629400.0 1786800.0 639600.0 1800600.0 ;
      RECT  629400.0 1814400.0 639600.0 1800600.0 ;
      RECT  629400.0 1814400.0 639600.0 1828200.0 ;
      RECT  629400.0 1842000.0 639600.0 1828200.0 ;
      RECT  629400.0 1842000.0 639600.0 1855800.0 ;
      RECT  629400.0 1869600.0 639600.0 1855800.0 ;
      RECT  629400.0 1869600.0 639600.0 1883400.0 ;
      RECT  629400.0 1897200.0 639600.0 1883400.0 ;
      RECT  629400.0 1897200.0 639600.0 1911000.0 ;
      RECT  629400.0 1924800.0 639600.0 1911000.0 ;
      RECT  629400.0 1924800.0 639600.0 1938600.0 ;
      RECT  629400.0 1952400.0 639600.0 1938600.0 ;
      RECT  629400.0 1952400.0 639600.0 1966200.0 ;
      RECT  629400.0 1980000.0 639600.0 1966200.0 ;
      RECT  629400.0 1980000.0 639600.0 1993800.0 ;
      RECT  629400.0 2007600.0 639600.0 1993800.0 ;
      RECT  629400.0 2007600.0 639600.0 2021400.0 ;
      RECT  629400.0 2035200.0 639600.0 2021400.0 ;
      RECT  629400.0 2035200.0 639600.0 2049000.0 ;
      RECT  629400.0 2062800.0 639600.0 2049000.0 ;
      RECT  629400.0 2062800.0 639600.0 2076600.0 ;
      RECT  629400.0 2090400.0 639600.0 2076600.0 ;
      RECT  629400.0 2090400.0 639600.0 2104200.0 ;
      RECT  629400.0 2118000.0 639600.0 2104200.0 ;
      RECT  629400.0 2118000.0 639600.0 2131800.0 ;
      RECT  629400.0 2145600.0 639600.0 2131800.0 ;
      RECT  639600.0 379200.0 649800.0 393000.0 ;
      RECT  639600.0 406800.0 649800.0 393000.0 ;
      RECT  639600.0 406800.0 649800.0 420600.0 ;
      RECT  639600.0 434400.0 649800.0 420600.0 ;
      RECT  639600.0 434400.0 649800.0 448200.0 ;
      RECT  639600.0 462000.0 649800.0 448200.0 ;
      RECT  639600.0 462000.0 649800.0 475800.0 ;
      RECT  639600.0 489600.0 649800.0 475800.0 ;
      RECT  639600.0 489600.0 649800.0 503400.0 ;
      RECT  639600.0 517200.0 649800.0 503400.0 ;
      RECT  639600.0 517200.0 649800.0 531000.0 ;
      RECT  639600.0 544800.0 649800.0 531000.0 ;
      RECT  639600.0 544800.0 649800.0 558600.0 ;
      RECT  639600.0 572400.0 649800.0 558600.0 ;
      RECT  639600.0 572400.0 649800.0 586200.0 ;
      RECT  639600.0 600000.0 649800.0 586200.0 ;
      RECT  639600.0 600000.0 649800.0 613800.0 ;
      RECT  639600.0 627600.0 649800.0 613800.0 ;
      RECT  639600.0 627600.0 649800.0 641400.0 ;
      RECT  639600.0 655200.0 649800.0 641400.0 ;
      RECT  639600.0 655200.0 649800.0 669000.0 ;
      RECT  639600.0 682800.0 649800.0 669000.0 ;
      RECT  639600.0 682800.0 649800.0 696600.0 ;
      RECT  639600.0 710400.0 649800.0 696600.0 ;
      RECT  639600.0 710400.0 649800.0 724200.0 ;
      RECT  639600.0 738000.0 649800.0 724200.0 ;
      RECT  639600.0 738000.0 649800.0 751800.0 ;
      RECT  639600.0 765600.0 649800.0 751800.0 ;
      RECT  639600.0 765600.0 649800.0 779400.0 ;
      RECT  639600.0 793200.0 649800.0 779400.0 ;
      RECT  639600.0 793200.0 649800.0 807000.0 ;
      RECT  639600.0 820800.0 649800.0 807000.0 ;
      RECT  639600.0 820800.0 649800.0 834600.0 ;
      RECT  639600.0 848400.0 649800.0 834600.0 ;
      RECT  639600.0 848400.0 649800.0 862200.0 ;
      RECT  639600.0 876000.0 649800.0 862200.0 ;
      RECT  639600.0 876000.0 649800.0 889800.0 ;
      RECT  639600.0 903600.0 649800.0 889800.0 ;
      RECT  639600.0 903600.0 649800.0 917400.0 ;
      RECT  639600.0 931200.0 649800.0 917400.0 ;
      RECT  639600.0 931200.0 649800.0 945000.0 ;
      RECT  639600.0 958800.0 649800.0 945000.0 ;
      RECT  639600.0 958800.0 649800.0 972600.0 ;
      RECT  639600.0 986400.0 649800.0 972600.0 ;
      RECT  639600.0 986400.0 649800.0 1000200.0 ;
      RECT  639600.0 1014000.0 649800.0 1000200.0 ;
      RECT  639600.0 1014000.0 649800.0 1027800.0 ;
      RECT  639600.0 1041600.0 649800.0 1027800.0 ;
      RECT  639600.0 1041600.0 649800.0 1055400.0 ;
      RECT  639600.0 1069200.0 649800.0 1055400.0 ;
      RECT  639600.0 1069200.0 649800.0 1083000.0 ;
      RECT  639600.0 1096800.0 649800.0 1083000.0 ;
      RECT  639600.0 1096800.0 649800.0 1110600.0 ;
      RECT  639600.0 1124400.0 649800.0 1110600.0 ;
      RECT  639600.0 1124400.0 649800.0 1138200.0 ;
      RECT  639600.0 1152000.0 649800.0 1138200.0 ;
      RECT  639600.0 1152000.0 649800.0 1165800.0 ;
      RECT  639600.0 1179600.0 649800.0 1165800.0 ;
      RECT  639600.0 1179600.0 649800.0 1193400.0 ;
      RECT  639600.0 1207200.0 649800.0 1193400.0 ;
      RECT  639600.0 1207200.0 649800.0 1221000.0 ;
      RECT  639600.0 1234800.0 649800.0 1221000.0 ;
      RECT  639600.0 1234800.0 649800.0 1248600.0 ;
      RECT  639600.0 1262400.0 649800.0 1248600.0 ;
      RECT  639600.0 1262400.0 649800.0 1276200.0 ;
      RECT  639600.0 1290000.0 649800.0 1276200.0 ;
      RECT  639600.0 1290000.0 649800.0 1303800.0 ;
      RECT  639600.0 1317600.0 649800.0 1303800.0 ;
      RECT  639600.0 1317600.0 649800.0 1331400.0 ;
      RECT  639600.0 1345200.0 649800.0 1331400.0 ;
      RECT  639600.0 1345200.0 649800.0 1359000.0 ;
      RECT  639600.0 1372800.0 649800.0 1359000.0 ;
      RECT  639600.0 1372800.0 649800.0 1386600.0 ;
      RECT  639600.0 1400400.0 649800.0 1386600.0 ;
      RECT  639600.0 1400400.0 649800.0 1414200.0 ;
      RECT  639600.0 1428000.0 649800.0 1414200.0 ;
      RECT  639600.0 1428000.0 649800.0 1441800.0 ;
      RECT  639600.0 1455600.0 649800.0 1441800.0 ;
      RECT  639600.0 1455600.0 649800.0 1469400.0 ;
      RECT  639600.0 1483200.0 649800.0 1469400.0 ;
      RECT  639600.0 1483200.0 649800.0 1497000.0 ;
      RECT  639600.0 1510800.0 649800.0 1497000.0 ;
      RECT  639600.0 1510800.0 649800.0 1524600.0 ;
      RECT  639600.0 1538400.0 649800.0 1524600.0 ;
      RECT  639600.0 1538400.0 649800.0 1552200.0 ;
      RECT  639600.0 1566000.0 649800.0 1552200.0 ;
      RECT  639600.0 1566000.0 649800.0 1579800.0 ;
      RECT  639600.0 1593600.0 649800.0 1579800.0 ;
      RECT  639600.0 1593600.0 649800.0 1607400.0 ;
      RECT  639600.0 1621200.0 649800.0 1607400.0 ;
      RECT  639600.0 1621200.0 649800.0 1635000.0 ;
      RECT  639600.0 1648800.0 649800.0 1635000.0 ;
      RECT  639600.0 1648800.0 649800.0 1662600.0 ;
      RECT  639600.0 1676400.0 649800.0 1662600.0 ;
      RECT  639600.0 1676400.0 649800.0 1690200.0 ;
      RECT  639600.0 1704000.0 649800.0 1690200.0 ;
      RECT  639600.0 1704000.0 649800.0 1717800.0 ;
      RECT  639600.0 1731600.0 649800.0 1717800.0 ;
      RECT  639600.0 1731600.0 649800.0 1745400.0 ;
      RECT  639600.0 1759200.0 649800.0 1745400.0 ;
      RECT  639600.0 1759200.0 649800.0 1773000.0 ;
      RECT  639600.0 1786800.0 649800.0 1773000.0 ;
      RECT  639600.0 1786800.0 649800.0 1800600.0 ;
      RECT  639600.0 1814400.0 649800.0 1800600.0 ;
      RECT  639600.0 1814400.0 649800.0 1828200.0 ;
      RECT  639600.0 1842000.0 649800.0 1828200.0 ;
      RECT  639600.0 1842000.0 649800.0 1855800.0 ;
      RECT  639600.0 1869600.0 649800.0 1855800.0 ;
      RECT  639600.0 1869600.0 649800.0 1883400.0 ;
      RECT  639600.0 1897200.0 649800.0 1883400.0 ;
      RECT  639600.0 1897200.0 649800.0 1911000.0 ;
      RECT  639600.0 1924800.0 649800.0 1911000.0 ;
      RECT  639600.0 1924800.0 649800.0 1938600.0 ;
      RECT  639600.0 1952400.0 649800.0 1938600.0 ;
      RECT  639600.0 1952400.0 649800.0 1966200.0 ;
      RECT  639600.0 1980000.0 649800.0 1966200.0 ;
      RECT  639600.0 1980000.0 649800.0 1993800.0 ;
      RECT  639600.0 2007600.0 649800.0 1993800.0 ;
      RECT  639600.0 2007600.0 649800.0 2021400.0 ;
      RECT  639600.0 2035200.0 649800.0 2021400.0 ;
      RECT  639600.0 2035200.0 649800.0 2049000.0 ;
      RECT  639600.0 2062800.0 649800.0 2049000.0 ;
      RECT  639600.0 2062800.0 649800.0 2076600.0 ;
      RECT  639600.0 2090400.0 649800.0 2076600.0 ;
      RECT  639600.0 2090400.0 649800.0 2104200.0 ;
      RECT  639600.0 2118000.0 649800.0 2104200.0 ;
      RECT  639600.0 2118000.0 649800.0 2131800.0 ;
      RECT  639600.0 2145600.0 649800.0 2131800.0 ;
      RECT  649800.0 379200.0 660000.0 393000.0 ;
      RECT  649800.0 406800.0 660000.0 393000.0 ;
      RECT  649800.0 406800.0 660000.0 420600.0 ;
      RECT  649800.0 434400.0 660000.0 420600.0 ;
      RECT  649800.0 434400.0 660000.0 448200.0 ;
      RECT  649800.0 462000.0 660000.0 448200.0 ;
      RECT  649800.0 462000.0 660000.0 475800.0 ;
      RECT  649800.0 489600.0 660000.0 475800.0 ;
      RECT  649800.0 489600.0 660000.0 503400.0 ;
      RECT  649800.0 517200.0 660000.0 503400.0 ;
      RECT  649800.0 517200.0 660000.0 531000.0 ;
      RECT  649800.0 544800.0 660000.0 531000.0 ;
      RECT  649800.0 544800.0 660000.0 558600.0 ;
      RECT  649800.0 572400.0 660000.0 558600.0 ;
      RECT  649800.0 572400.0 660000.0 586200.0 ;
      RECT  649800.0 600000.0 660000.0 586200.0 ;
      RECT  649800.0 600000.0 660000.0 613800.0 ;
      RECT  649800.0 627600.0 660000.0 613800.0 ;
      RECT  649800.0 627600.0 660000.0 641400.0 ;
      RECT  649800.0 655200.0 660000.0 641400.0 ;
      RECT  649800.0 655200.0 660000.0 669000.0 ;
      RECT  649800.0 682800.0 660000.0 669000.0 ;
      RECT  649800.0 682800.0 660000.0 696600.0 ;
      RECT  649800.0 710400.0 660000.0 696600.0 ;
      RECT  649800.0 710400.0 660000.0 724200.0 ;
      RECT  649800.0 738000.0 660000.0 724200.0 ;
      RECT  649800.0 738000.0 660000.0 751800.0 ;
      RECT  649800.0 765600.0 660000.0 751800.0 ;
      RECT  649800.0 765600.0 660000.0 779400.0 ;
      RECT  649800.0 793200.0 660000.0 779400.0 ;
      RECT  649800.0 793200.0 660000.0 807000.0 ;
      RECT  649800.0 820800.0 660000.0 807000.0 ;
      RECT  649800.0 820800.0 660000.0 834600.0 ;
      RECT  649800.0 848400.0 660000.0 834600.0 ;
      RECT  649800.0 848400.0 660000.0 862200.0 ;
      RECT  649800.0 876000.0 660000.0 862200.0 ;
      RECT  649800.0 876000.0 660000.0 889800.0 ;
      RECT  649800.0 903600.0 660000.0 889800.0 ;
      RECT  649800.0 903600.0 660000.0 917400.0 ;
      RECT  649800.0 931200.0 660000.0 917400.0 ;
      RECT  649800.0 931200.0 660000.0 945000.0 ;
      RECT  649800.0 958800.0 660000.0 945000.0 ;
      RECT  649800.0 958800.0 660000.0 972600.0 ;
      RECT  649800.0 986400.0 660000.0 972600.0 ;
      RECT  649800.0 986400.0 660000.0 1000200.0 ;
      RECT  649800.0 1014000.0 660000.0 1000200.0 ;
      RECT  649800.0 1014000.0 660000.0 1027800.0 ;
      RECT  649800.0 1041600.0 660000.0 1027800.0 ;
      RECT  649800.0 1041600.0 660000.0 1055400.0 ;
      RECT  649800.0 1069200.0 660000.0 1055400.0 ;
      RECT  649800.0 1069200.0 660000.0 1083000.0 ;
      RECT  649800.0 1096800.0 660000.0 1083000.0 ;
      RECT  649800.0 1096800.0 660000.0 1110600.0 ;
      RECT  649800.0 1124400.0 660000.0 1110600.0 ;
      RECT  649800.0 1124400.0 660000.0 1138200.0 ;
      RECT  649800.0 1152000.0 660000.0 1138200.0 ;
      RECT  649800.0 1152000.0 660000.0 1165800.0 ;
      RECT  649800.0 1179600.0 660000.0 1165800.0 ;
      RECT  649800.0 1179600.0 660000.0 1193400.0 ;
      RECT  649800.0 1207200.0 660000.0 1193400.0 ;
      RECT  649800.0 1207200.0 660000.0 1221000.0 ;
      RECT  649800.0 1234800.0 660000.0 1221000.0 ;
      RECT  649800.0 1234800.0 660000.0 1248600.0 ;
      RECT  649800.0 1262400.0 660000.0 1248600.0 ;
      RECT  649800.0 1262400.0 660000.0 1276200.0 ;
      RECT  649800.0 1290000.0 660000.0 1276200.0 ;
      RECT  649800.0 1290000.0 660000.0 1303800.0 ;
      RECT  649800.0 1317600.0 660000.0 1303800.0 ;
      RECT  649800.0 1317600.0 660000.0 1331400.0 ;
      RECT  649800.0 1345200.0 660000.0 1331400.0 ;
      RECT  649800.0 1345200.0 660000.0 1359000.0 ;
      RECT  649800.0 1372800.0 660000.0 1359000.0 ;
      RECT  649800.0 1372800.0 660000.0 1386600.0 ;
      RECT  649800.0 1400400.0 660000.0 1386600.0 ;
      RECT  649800.0 1400400.0 660000.0 1414200.0 ;
      RECT  649800.0 1428000.0 660000.0 1414200.0 ;
      RECT  649800.0 1428000.0 660000.0 1441800.0 ;
      RECT  649800.0 1455600.0 660000.0 1441800.0 ;
      RECT  649800.0 1455600.0 660000.0 1469400.0 ;
      RECT  649800.0 1483200.0 660000.0 1469400.0 ;
      RECT  649800.0 1483200.0 660000.0 1497000.0 ;
      RECT  649800.0 1510800.0 660000.0 1497000.0 ;
      RECT  649800.0 1510800.0 660000.0 1524600.0 ;
      RECT  649800.0 1538400.0 660000.0 1524600.0 ;
      RECT  649800.0 1538400.0 660000.0 1552200.0 ;
      RECT  649800.0 1566000.0 660000.0 1552200.0 ;
      RECT  649800.0 1566000.0 660000.0 1579800.0 ;
      RECT  649800.0 1593600.0 660000.0 1579800.0 ;
      RECT  649800.0 1593600.0 660000.0 1607400.0 ;
      RECT  649800.0 1621200.0 660000.0 1607400.0 ;
      RECT  649800.0 1621200.0 660000.0 1635000.0 ;
      RECT  649800.0 1648800.0 660000.0 1635000.0 ;
      RECT  649800.0 1648800.0 660000.0 1662600.0 ;
      RECT  649800.0 1676400.0 660000.0 1662600.0 ;
      RECT  649800.0 1676400.0 660000.0 1690200.0 ;
      RECT  649800.0 1704000.0 660000.0 1690200.0 ;
      RECT  649800.0 1704000.0 660000.0 1717800.0 ;
      RECT  649800.0 1731600.0 660000.0 1717800.0 ;
      RECT  649800.0 1731600.0 660000.0 1745400.0 ;
      RECT  649800.0 1759200.0 660000.0 1745400.0 ;
      RECT  649800.0 1759200.0 660000.0 1773000.0 ;
      RECT  649800.0 1786800.0 660000.0 1773000.0 ;
      RECT  649800.0 1786800.0 660000.0 1800600.0 ;
      RECT  649800.0 1814400.0 660000.0 1800600.0 ;
      RECT  649800.0 1814400.0 660000.0 1828200.0 ;
      RECT  649800.0 1842000.0 660000.0 1828200.0 ;
      RECT  649800.0 1842000.0 660000.0 1855800.0 ;
      RECT  649800.0 1869600.0 660000.0 1855800.0 ;
      RECT  649800.0 1869600.0 660000.0 1883400.0 ;
      RECT  649800.0 1897200.0 660000.0 1883400.0 ;
      RECT  649800.0 1897200.0 660000.0 1911000.0 ;
      RECT  649800.0 1924800.0 660000.0 1911000.0 ;
      RECT  649800.0 1924800.0 660000.0 1938600.0 ;
      RECT  649800.0 1952400.0 660000.0 1938600.0 ;
      RECT  649800.0 1952400.0 660000.0 1966200.0 ;
      RECT  649800.0 1980000.0 660000.0 1966200.0 ;
      RECT  649800.0 1980000.0 660000.0 1993800.0 ;
      RECT  649800.0 2007600.0 660000.0 1993800.0 ;
      RECT  649800.0 2007600.0 660000.0 2021400.0 ;
      RECT  649800.0 2035200.0 660000.0 2021400.0 ;
      RECT  649800.0 2035200.0 660000.0 2049000.0 ;
      RECT  649800.0 2062800.0 660000.0 2049000.0 ;
      RECT  649800.0 2062800.0 660000.0 2076600.0 ;
      RECT  649800.0 2090400.0 660000.0 2076600.0 ;
      RECT  649800.0 2090400.0 660000.0 2104200.0 ;
      RECT  649800.0 2118000.0 660000.0 2104200.0 ;
      RECT  649800.0 2118000.0 660000.0 2131800.0 ;
      RECT  649800.0 2145600.0 660000.0 2131800.0 ;
      RECT  660000.0 379200.0 670200.0 393000.0 ;
      RECT  660000.0 406800.0 670200.0 393000.0 ;
      RECT  660000.0 406800.0 670200.0 420600.0 ;
      RECT  660000.0 434400.0 670200.0 420600.0 ;
      RECT  660000.0 434400.0 670200.0 448200.0 ;
      RECT  660000.0 462000.0 670200.0 448200.0 ;
      RECT  660000.0 462000.0 670200.0 475800.0 ;
      RECT  660000.0 489600.0 670200.0 475800.0 ;
      RECT  660000.0 489600.0 670200.0 503400.0 ;
      RECT  660000.0 517200.0 670200.0 503400.0 ;
      RECT  660000.0 517200.0 670200.0 531000.0 ;
      RECT  660000.0 544800.0 670200.0 531000.0 ;
      RECT  660000.0 544800.0 670200.0 558600.0 ;
      RECT  660000.0 572400.0 670200.0 558600.0 ;
      RECT  660000.0 572400.0 670200.0 586200.0 ;
      RECT  660000.0 600000.0 670200.0 586200.0 ;
      RECT  660000.0 600000.0 670200.0 613800.0 ;
      RECT  660000.0 627600.0 670200.0 613800.0 ;
      RECT  660000.0 627600.0 670200.0 641400.0 ;
      RECT  660000.0 655200.0 670200.0 641400.0 ;
      RECT  660000.0 655200.0 670200.0 669000.0 ;
      RECT  660000.0 682800.0 670200.0 669000.0 ;
      RECT  660000.0 682800.0 670200.0 696600.0 ;
      RECT  660000.0 710400.0 670200.0 696600.0 ;
      RECT  660000.0 710400.0 670200.0 724200.0 ;
      RECT  660000.0 738000.0 670200.0 724200.0 ;
      RECT  660000.0 738000.0 670200.0 751800.0 ;
      RECT  660000.0 765600.0 670200.0 751800.0 ;
      RECT  660000.0 765600.0 670200.0 779400.0 ;
      RECT  660000.0 793200.0 670200.0 779400.0 ;
      RECT  660000.0 793200.0 670200.0 807000.0 ;
      RECT  660000.0 820800.0 670200.0 807000.0 ;
      RECT  660000.0 820800.0 670200.0 834600.0 ;
      RECT  660000.0 848400.0 670200.0 834600.0 ;
      RECT  660000.0 848400.0 670200.0 862200.0 ;
      RECT  660000.0 876000.0 670200.0 862200.0 ;
      RECT  660000.0 876000.0 670200.0 889800.0 ;
      RECT  660000.0 903600.0 670200.0 889800.0 ;
      RECT  660000.0 903600.0 670200.0 917400.0 ;
      RECT  660000.0 931200.0 670200.0 917400.0 ;
      RECT  660000.0 931200.0 670200.0 945000.0 ;
      RECT  660000.0 958800.0 670200.0 945000.0 ;
      RECT  660000.0 958800.0 670200.0 972600.0 ;
      RECT  660000.0 986400.0 670200.0 972600.0 ;
      RECT  660000.0 986400.0 670200.0 1000200.0 ;
      RECT  660000.0 1014000.0 670200.0 1000200.0 ;
      RECT  660000.0 1014000.0 670200.0 1027800.0 ;
      RECT  660000.0 1041600.0 670200.0 1027800.0 ;
      RECT  660000.0 1041600.0 670200.0 1055400.0 ;
      RECT  660000.0 1069200.0 670200.0 1055400.0 ;
      RECT  660000.0 1069200.0 670200.0 1083000.0 ;
      RECT  660000.0 1096800.0 670200.0 1083000.0 ;
      RECT  660000.0 1096800.0 670200.0 1110600.0 ;
      RECT  660000.0 1124400.0 670200.0 1110600.0 ;
      RECT  660000.0 1124400.0 670200.0 1138200.0 ;
      RECT  660000.0 1152000.0 670200.0 1138200.0 ;
      RECT  660000.0 1152000.0 670200.0 1165800.0 ;
      RECT  660000.0 1179600.0 670200.0 1165800.0 ;
      RECT  660000.0 1179600.0 670200.0 1193400.0 ;
      RECT  660000.0 1207200.0 670200.0 1193400.0 ;
      RECT  660000.0 1207200.0 670200.0 1221000.0 ;
      RECT  660000.0 1234800.0 670200.0 1221000.0 ;
      RECT  660000.0 1234800.0 670200.0 1248600.0 ;
      RECT  660000.0 1262400.0 670200.0 1248600.0 ;
      RECT  660000.0 1262400.0 670200.0 1276200.0 ;
      RECT  660000.0 1290000.0 670200.0 1276200.0 ;
      RECT  660000.0 1290000.0 670200.0 1303800.0 ;
      RECT  660000.0 1317600.0 670200.0 1303800.0 ;
      RECT  660000.0 1317600.0 670200.0 1331400.0 ;
      RECT  660000.0 1345200.0 670200.0 1331400.0 ;
      RECT  660000.0 1345200.0 670200.0 1359000.0 ;
      RECT  660000.0 1372800.0 670200.0 1359000.0 ;
      RECT  660000.0 1372800.0 670200.0 1386600.0 ;
      RECT  660000.0 1400400.0 670200.0 1386600.0 ;
      RECT  660000.0 1400400.0 670200.0 1414200.0 ;
      RECT  660000.0 1428000.0 670200.0 1414200.0 ;
      RECT  660000.0 1428000.0 670200.0 1441800.0 ;
      RECT  660000.0 1455600.0 670200.0 1441800.0 ;
      RECT  660000.0 1455600.0 670200.0 1469400.0 ;
      RECT  660000.0 1483200.0 670200.0 1469400.0 ;
      RECT  660000.0 1483200.0 670200.0 1497000.0 ;
      RECT  660000.0 1510800.0 670200.0 1497000.0 ;
      RECT  660000.0 1510800.0 670200.0 1524600.0 ;
      RECT  660000.0 1538400.0 670200.0 1524600.0 ;
      RECT  660000.0 1538400.0 670200.0 1552200.0 ;
      RECT  660000.0 1566000.0 670200.0 1552200.0 ;
      RECT  660000.0 1566000.0 670200.0 1579800.0 ;
      RECT  660000.0 1593600.0 670200.0 1579800.0 ;
      RECT  660000.0 1593600.0 670200.0 1607400.0 ;
      RECT  660000.0 1621200.0 670200.0 1607400.0 ;
      RECT  660000.0 1621200.0 670200.0 1635000.0 ;
      RECT  660000.0 1648800.0 670200.0 1635000.0 ;
      RECT  660000.0 1648800.0 670200.0 1662600.0 ;
      RECT  660000.0 1676400.0 670200.0 1662600.0 ;
      RECT  660000.0 1676400.0 670200.0 1690200.0 ;
      RECT  660000.0 1704000.0 670200.0 1690200.0 ;
      RECT  660000.0 1704000.0 670200.0 1717800.0 ;
      RECT  660000.0 1731600.0 670200.0 1717800.0 ;
      RECT  660000.0 1731600.0 670200.0 1745400.0 ;
      RECT  660000.0 1759200.0 670200.0 1745400.0 ;
      RECT  660000.0 1759200.0 670200.0 1773000.0 ;
      RECT  660000.0 1786800.0 670200.0 1773000.0 ;
      RECT  660000.0 1786800.0 670200.0 1800600.0 ;
      RECT  660000.0 1814400.0 670200.0 1800600.0 ;
      RECT  660000.0 1814400.0 670200.0 1828200.0 ;
      RECT  660000.0 1842000.0 670200.0 1828200.0 ;
      RECT  660000.0 1842000.0 670200.0 1855800.0 ;
      RECT  660000.0 1869600.0 670200.0 1855800.0 ;
      RECT  660000.0 1869600.0 670200.0 1883400.0 ;
      RECT  660000.0 1897200.0 670200.0 1883400.0 ;
      RECT  660000.0 1897200.0 670200.0 1911000.0 ;
      RECT  660000.0 1924800.0 670200.0 1911000.0 ;
      RECT  660000.0 1924800.0 670200.0 1938600.0 ;
      RECT  660000.0 1952400.0 670200.0 1938600.0 ;
      RECT  660000.0 1952400.0 670200.0 1966200.0 ;
      RECT  660000.0 1980000.0 670200.0 1966200.0 ;
      RECT  660000.0 1980000.0 670200.0 1993800.0 ;
      RECT  660000.0 2007600.0 670200.0 1993800.0 ;
      RECT  660000.0 2007600.0 670200.0 2021400.0 ;
      RECT  660000.0 2035200.0 670200.0 2021400.0 ;
      RECT  660000.0 2035200.0 670200.0 2049000.0 ;
      RECT  660000.0 2062800.0 670200.0 2049000.0 ;
      RECT  660000.0 2062800.0 670200.0 2076600.0 ;
      RECT  660000.0 2090400.0 670200.0 2076600.0 ;
      RECT  660000.0 2090400.0 670200.0 2104200.0 ;
      RECT  660000.0 2118000.0 670200.0 2104200.0 ;
      RECT  660000.0 2118000.0 670200.0 2131800.0 ;
      RECT  660000.0 2145600.0 670200.0 2131800.0 ;
      RECT  670200.0 379200.0 680400.0 393000.0 ;
      RECT  670200.0 406800.0 680400.0 393000.0 ;
      RECT  670200.0 406800.0 680400.0 420600.0 ;
      RECT  670200.0 434400.0 680400.0 420600.0 ;
      RECT  670200.0 434400.0 680400.0 448200.0 ;
      RECT  670200.0 462000.0 680400.0 448200.0 ;
      RECT  670200.0 462000.0 680400.0 475800.0 ;
      RECT  670200.0 489600.0 680400.0 475800.0 ;
      RECT  670200.0 489600.0 680400.0 503400.0 ;
      RECT  670200.0 517200.0 680400.0 503400.0 ;
      RECT  670200.0 517200.0 680400.0 531000.0 ;
      RECT  670200.0 544800.0 680400.0 531000.0 ;
      RECT  670200.0 544800.0 680400.0 558600.0 ;
      RECT  670200.0 572400.0 680400.0 558600.0 ;
      RECT  670200.0 572400.0 680400.0 586200.0 ;
      RECT  670200.0 600000.0 680400.0 586200.0 ;
      RECT  670200.0 600000.0 680400.0 613800.0 ;
      RECT  670200.0 627600.0 680400.0 613800.0 ;
      RECT  670200.0 627600.0 680400.0 641400.0 ;
      RECT  670200.0 655200.0 680400.0 641400.0 ;
      RECT  670200.0 655200.0 680400.0 669000.0 ;
      RECT  670200.0 682800.0 680400.0 669000.0 ;
      RECT  670200.0 682800.0 680400.0 696600.0 ;
      RECT  670200.0 710400.0 680400.0 696600.0 ;
      RECT  670200.0 710400.0 680400.0 724200.0 ;
      RECT  670200.0 738000.0 680400.0 724200.0 ;
      RECT  670200.0 738000.0 680400.0 751800.0 ;
      RECT  670200.0 765600.0 680400.0 751800.0 ;
      RECT  670200.0 765600.0 680400.0 779400.0 ;
      RECT  670200.0 793200.0 680400.0 779400.0 ;
      RECT  670200.0 793200.0 680400.0 807000.0 ;
      RECT  670200.0 820800.0 680400.0 807000.0 ;
      RECT  670200.0 820800.0 680400.0 834600.0 ;
      RECT  670200.0 848400.0 680400.0 834600.0 ;
      RECT  670200.0 848400.0 680400.0 862200.0 ;
      RECT  670200.0 876000.0 680400.0 862200.0 ;
      RECT  670200.0 876000.0 680400.0 889800.0 ;
      RECT  670200.0 903600.0 680400.0 889800.0 ;
      RECT  670200.0 903600.0 680400.0 917400.0 ;
      RECT  670200.0 931200.0 680400.0 917400.0 ;
      RECT  670200.0 931200.0 680400.0 945000.0 ;
      RECT  670200.0 958800.0 680400.0 945000.0 ;
      RECT  670200.0 958800.0 680400.0 972600.0 ;
      RECT  670200.0 986400.0 680400.0 972600.0 ;
      RECT  670200.0 986400.0 680400.0 1000200.0 ;
      RECT  670200.0 1014000.0 680400.0 1000200.0 ;
      RECT  670200.0 1014000.0 680400.0 1027800.0 ;
      RECT  670200.0 1041600.0 680400.0 1027800.0 ;
      RECT  670200.0 1041600.0 680400.0 1055400.0 ;
      RECT  670200.0 1069200.0 680400.0 1055400.0 ;
      RECT  670200.0 1069200.0 680400.0 1083000.0 ;
      RECT  670200.0 1096800.0 680400.0 1083000.0 ;
      RECT  670200.0 1096800.0 680400.0 1110600.0 ;
      RECT  670200.0 1124400.0 680400.0 1110600.0 ;
      RECT  670200.0 1124400.0 680400.0 1138200.0 ;
      RECT  670200.0 1152000.0 680400.0 1138200.0 ;
      RECT  670200.0 1152000.0 680400.0 1165800.0 ;
      RECT  670200.0 1179600.0 680400.0 1165800.0 ;
      RECT  670200.0 1179600.0 680400.0 1193400.0 ;
      RECT  670200.0 1207200.0 680400.0 1193400.0 ;
      RECT  670200.0 1207200.0 680400.0 1221000.0 ;
      RECT  670200.0 1234800.0 680400.0 1221000.0 ;
      RECT  670200.0 1234800.0 680400.0 1248600.0 ;
      RECT  670200.0 1262400.0 680400.0 1248600.0 ;
      RECT  670200.0 1262400.0 680400.0 1276200.0 ;
      RECT  670200.0 1290000.0 680400.0 1276200.0 ;
      RECT  670200.0 1290000.0 680400.0 1303800.0 ;
      RECT  670200.0 1317600.0 680400.0 1303800.0 ;
      RECT  670200.0 1317600.0 680400.0 1331400.0 ;
      RECT  670200.0 1345200.0 680400.0 1331400.0 ;
      RECT  670200.0 1345200.0 680400.0 1359000.0 ;
      RECT  670200.0 1372800.0 680400.0 1359000.0 ;
      RECT  670200.0 1372800.0 680400.0 1386600.0 ;
      RECT  670200.0 1400400.0 680400.0 1386600.0 ;
      RECT  670200.0 1400400.0 680400.0 1414200.0 ;
      RECT  670200.0 1428000.0 680400.0 1414200.0 ;
      RECT  670200.0 1428000.0 680400.0 1441800.0 ;
      RECT  670200.0 1455600.0 680400.0 1441800.0 ;
      RECT  670200.0 1455600.0 680400.0 1469400.0 ;
      RECT  670200.0 1483200.0 680400.0 1469400.0 ;
      RECT  670200.0 1483200.0 680400.0 1497000.0 ;
      RECT  670200.0 1510800.0 680400.0 1497000.0 ;
      RECT  670200.0 1510800.0 680400.0 1524600.0 ;
      RECT  670200.0 1538400.0 680400.0 1524600.0 ;
      RECT  670200.0 1538400.0 680400.0 1552200.0 ;
      RECT  670200.0 1566000.0 680400.0 1552200.0 ;
      RECT  670200.0 1566000.0 680400.0 1579800.0 ;
      RECT  670200.0 1593600.0 680400.0 1579800.0 ;
      RECT  670200.0 1593600.0 680400.0 1607400.0 ;
      RECT  670200.0 1621200.0 680400.0 1607400.0 ;
      RECT  670200.0 1621200.0 680400.0 1635000.0 ;
      RECT  670200.0 1648800.0 680400.0 1635000.0 ;
      RECT  670200.0 1648800.0 680400.0 1662600.0 ;
      RECT  670200.0 1676400.0 680400.0 1662600.0 ;
      RECT  670200.0 1676400.0 680400.0 1690200.0 ;
      RECT  670200.0 1704000.0 680400.0 1690200.0 ;
      RECT  670200.0 1704000.0 680400.0 1717800.0 ;
      RECT  670200.0 1731600.0 680400.0 1717800.0 ;
      RECT  670200.0 1731600.0 680400.0 1745400.0 ;
      RECT  670200.0 1759200.0 680400.0 1745400.0 ;
      RECT  670200.0 1759200.0 680400.0 1773000.0 ;
      RECT  670200.0 1786800.0 680400.0 1773000.0 ;
      RECT  670200.0 1786800.0 680400.0 1800600.0 ;
      RECT  670200.0 1814400.0 680400.0 1800600.0 ;
      RECT  670200.0 1814400.0 680400.0 1828200.0 ;
      RECT  670200.0 1842000.0 680400.0 1828200.0 ;
      RECT  670200.0 1842000.0 680400.0 1855800.0 ;
      RECT  670200.0 1869600.0 680400.0 1855800.0 ;
      RECT  670200.0 1869600.0 680400.0 1883400.0 ;
      RECT  670200.0 1897200.0 680400.0 1883400.0 ;
      RECT  670200.0 1897200.0 680400.0 1911000.0 ;
      RECT  670200.0 1924800.0 680400.0 1911000.0 ;
      RECT  670200.0 1924800.0 680400.0 1938600.0 ;
      RECT  670200.0 1952400.0 680400.0 1938600.0 ;
      RECT  670200.0 1952400.0 680400.0 1966200.0 ;
      RECT  670200.0 1980000.0 680400.0 1966200.0 ;
      RECT  670200.0 1980000.0 680400.0 1993800.0 ;
      RECT  670200.0 2007600.0 680400.0 1993800.0 ;
      RECT  670200.0 2007600.0 680400.0 2021400.0 ;
      RECT  670200.0 2035200.0 680400.0 2021400.0 ;
      RECT  670200.0 2035200.0 680400.0 2049000.0 ;
      RECT  670200.0 2062800.0 680400.0 2049000.0 ;
      RECT  670200.0 2062800.0 680400.0 2076600.0 ;
      RECT  670200.0 2090400.0 680400.0 2076600.0 ;
      RECT  670200.0 2090400.0 680400.0 2104200.0 ;
      RECT  670200.0 2118000.0 680400.0 2104200.0 ;
      RECT  670200.0 2118000.0 680400.0 2131800.0 ;
      RECT  670200.0 2145600.0 680400.0 2131800.0 ;
      RECT  680400.0 379200.0 690600.0 393000.0 ;
      RECT  680400.0 406800.0 690600.0 393000.0 ;
      RECT  680400.0 406800.0 690600.0 420600.0 ;
      RECT  680400.0 434400.0 690600.0 420600.0 ;
      RECT  680400.0 434400.0 690600.0 448200.0 ;
      RECT  680400.0 462000.0 690600.0 448200.0 ;
      RECT  680400.0 462000.0 690600.0 475800.0 ;
      RECT  680400.0 489600.0 690600.0 475800.0 ;
      RECT  680400.0 489600.0 690600.0 503400.0 ;
      RECT  680400.0 517200.0 690600.0 503400.0 ;
      RECT  680400.0 517200.0 690600.0 531000.0 ;
      RECT  680400.0 544800.0 690600.0 531000.0 ;
      RECT  680400.0 544800.0 690600.0 558600.0 ;
      RECT  680400.0 572400.0 690600.0 558600.0 ;
      RECT  680400.0 572400.0 690600.0 586200.0 ;
      RECT  680400.0 600000.0 690600.0 586200.0 ;
      RECT  680400.0 600000.0 690600.0 613800.0 ;
      RECT  680400.0 627600.0 690600.0 613800.0 ;
      RECT  680400.0 627600.0 690600.0 641400.0 ;
      RECT  680400.0 655200.0 690600.0 641400.0 ;
      RECT  680400.0 655200.0 690600.0 669000.0 ;
      RECT  680400.0 682800.0 690600.0 669000.0 ;
      RECT  680400.0 682800.0 690600.0 696600.0 ;
      RECT  680400.0 710400.0 690600.0 696600.0 ;
      RECT  680400.0 710400.0 690600.0 724200.0 ;
      RECT  680400.0 738000.0 690600.0 724200.0 ;
      RECT  680400.0 738000.0 690600.0 751800.0 ;
      RECT  680400.0 765600.0 690600.0 751800.0 ;
      RECT  680400.0 765600.0 690600.0 779400.0 ;
      RECT  680400.0 793200.0 690600.0 779400.0 ;
      RECT  680400.0 793200.0 690600.0 807000.0 ;
      RECT  680400.0 820800.0 690600.0 807000.0 ;
      RECT  680400.0 820800.0 690600.0 834600.0 ;
      RECT  680400.0 848400.0 690600.0 834600.0 ;
      RECT  680400.0 848400.0 690600.0 862200.0 ;
      RECT  680400.0 876000.0 690600.0 862200.0 ;
      RECT  680400.0 876000.0 690600.0 889800.0 ;
      RECT  680400.0 903600.0 690600.0 889800.0 ;
      RECT  680400.0 903600.0 690600.0 917400.0 ;
      RECT  680400.0 931200.0 690600.0 917400.0 ;
      RECT  680400.0 931200.0 690600.0 945000.0 ;
      RECT  680400.0 958800.0 690600.0 945000.0 ;
      RECT  680400.0 958800.0 690600.0 972600.0 ;
      RECT  680400.0 986400.0 690600.0 972600.0 ;
      RECT  680400.0 986400.0 690600.0 1000200.0 ;
      RECT  680400.0 1014000.0 690600.0 1000200.0 ;
      RECT  680400.0 1014000.0 690600.0 1027800.0 ;
      RECT  680400.0 1041600.0 690600.0 1027800.0 ;
      RECT  680400.0 1041600.0 690600.0 1055400.0 ;
      RECT  680400.0 1069200.0 690600.0 1055400.0 ;
      RECT  680400.0 1069200.0 690600.0 1083000.0 ;
      RECT  680400.0 1096800.0 690600.0 1083000.0 ;
      RECT  680400.0 1096800.0 690600.0 1110600.0 ;
      RECT  680400.0 1124400.0 690600.0 1110600.0 ;
      RECT  680400.0 1124400.0 690600.0 1138200.0 ;
      RECT  680400.0 1152000.0 690600.0 1138200.0 ;
      RECT  680400.0 1152000.0 690600.0 1165800.0 ;
      RECT  680400.0 1179600.0 690600.0 1165800.0 ;
      RECT  680400.0 1179600.0 690600.0 1193400.0 ;
      RECT  680400.0 1207200.0 690600.0 1193400.0 ;
      RECT  680400.0 1207200.0 690600.0 1221000.0 ;
      RECT  680400.0 1234800.0 690600.0 1221000.0 ;
      RECT  680400.0 1234800.0 690600.0 1248600.0 ;
      RECT  680400.0 1262400.0 690600.0 1248600.0 ;
      RECT  680400.0 1262400.0 690600.0 1276200.0 ;
      RECT  680400.0 1290000.0 690600.0 1276200.0 ;
      RECT  680400.0 1290000.0 690600.0 1303800.0 ;
      RECT  680400.0 1317600.0 690600.0 1303800.0 ;
      RECT  680400.0 1317600.0 690600.0 1331400.0 ;
      RECT  680400.0 1345200.0 690600.0 1331400.0 ;
      RECT  680400.0 1345200.0 690600.0 1359000.0 ;
      RECT  680400.0 1372800.0 690600.0 1359000.0 ;
      RECT  680400.0 1372800.0 690600.0 1386600.0 ;
      RECT  680400.0 1400400.0 690600.0 1386600.0 ;
      RECT  680400.0 1400400.0 690600.0 1414200.0 ;
      RECT  680400.0 1428000.0 690600.0 1414200.0 ;
      RECT  680400.0 1428000.0 690600.0 1441800.0 ;
      RECT  680400.0 1455600.0 690600.0 1441800.0 ;
      RECT  680400.0 1455600.0 690600.0 1469400.0 ;
      RECT  680400.0 1483200.0 690600.0 1469400.0 ;
      RECT  680400.0 1483200.0 690600.0 1497000.0 ;
      RECT  680400.0 1510800.0 690600.0 1497000.0 ;
      RECT  680400.0 1510800.0 690600.0 1524600.0 ;
      RECT  680400.0 1538400.0 690600.0 1524600.0 ;
      RECT  680400.0 1538400.0 690600.0 1552200.0 ;
      RECT  680400.0 1566000.0 690600.0 1552200.0 ;
      RECT  680400.0 1566000.0 690600.0 1579800.0 ;
      RECT  680400.0 1593600.0 690600.0 1579800.0 ;
      RECT  680400.0 1593600.0 690600.0 1607400.0 ;
      RECT  680400.0 1621200.0 690600.0 1607400.0 ;
      RECT  680400.0 1621200.0 690600.0 1635000.0 ;
      RECT  680400.0 1648800.0 690600.0 1635000.0 ;
      RECT  680400.0 1648800.0 690600.0 1662600.0 ;
      RECT  680400.0 1676400.0 690600.0 1662600.0 ;
      RECT  680400.0 1676400.0 690600.0 1690200.0 ;
      RECT  680400.0 1704000.0 690600.0 1690200.0 ;
      RECT  680400.0 1704000.0 690600.0 1717800.0 ;
      RECT  680400.0 1731600.0 690600.0 1717800.0 ;
      RECT  680400.0 1731600.0 690600.0 1745400.0 ;
      RECT  680400.0 1759200.0 690600.0 1745400.0 ;
      RECT  680400.0 1759200.0 690600.0 1773000.0 ;
      RECT  680400.0 1786800.0 690600.0 1773000.0 ;
      RECT  680400.0 1786800.0 690600.0 1800600.0 ;
      RECT  680400.0 1814400.0 690600.0 1800600.0 ;
      RECT  680400.0 1814400.0 690600.0 1828200.0 ;
      RECT  680400.0 1842000.0 690600.0 1828200.0 ;
      RECT  680400.0 1842000.0 690600.0 1855800.0 ;
      RECT  680400.0 1869600.0 690600.0 1855800.0 ;
      RECT  680400.0 1869600.0 690600.0 1883400.0 ;
      RECT  680400.0 1897200.0 690600.0 1883400.0 ;
      RECT  680400.0 1897200.0 690600.0 1911000.0 ;
      RECT  680400.0 1924800.0 690600.0 1911000.0 ;
      RECT  680400.0 1924800.0 690600.0 1938600.0 ;
      RECT  680400.0 1952400.0 690600.0 1938600.0 ;
      RECT  680400.0 1952400.0 690600.0 1966200.0 ;
      RECT  680400.0 1980000.0 690600.0 1966200.0 ;
      RECT  680400.0 1980000.0 690600.0 1993800.0 ;
      RECT  680400.0 2007600.0 690600.0 1993800.0 ;
      RECT  680400.0 2007600.0 690600.0 2021400.0 ;
      RECT  680400.0 2035200.0 690600.0 2021400.0 ;
      RECT  680400.0 2035200.0 690600.0 2049000.0 ;
      RECT  680400.0 2062800.0 690600.0 2049000.0 ;
      RECT  680400.0 2062800.0 690600.0 2076600.0 ;
      RECT  680400.0 2090400.0 690600.0 2076600.0 ;
      RECT  680400.0 2090400.0 690600.0 2104200.0 ;
      RECT  680400.0 2118000.0 690600.0 2104200.0 ;
      RECT  680400.0 2118000.0 690600.0 2131800.0 ;
      RECT  680400.0 2145600.0 690600.0 2131800.0 ;
      RECT  690600.0 379200.0 700800.0 393000.0 ;
      RECT  690600.0 406800.0 700800.0 393000.0 ;
      RECT  690600.0 406800.0 700800.0 420600.0 ;
      RECT  690600.0 434400.0 700800.0 420600.0 ;
      RECT  690600.0 434400.0 700800.0 448200.0 ;
      RECT  690600.0 462000.0 700800.0 448200.0 ;
      RECT  690600.0 462000.0 700800.0 475800.0 ;
      RECT  690600.0 489600.0 700800.0 475800.0 ;
      RECT  690600.0 489600.0 700800.0 503400.0 ;
      RECT  690600.0 517200.0 700800.0 503400.0 ;
      RECT  690600.0 517200.0 700800.0 531000.0 ;
      RECT  690600.0 544800.0 700800.0 531000.0 ;
      RECT  690600.0 544800.0 700800.0 558600.0 ;
      RECT  690600.0 572400.0 700800.0 558600.0 ;
      RECT  690600.0 572400.0 700800.0 586200.0 ;
      RECT  690600.0 600000.0 700800.0 586200.0 ;
      RECT  690600.0 600000.0 700800.0 613800.0 ;
      RECT  690600.0 627600.0 700800.0 613800.0 ;
      RECT  690600.0 627600.0 700800.0 641400.0 ;
      RECT  690600.0 655200.0 700800.0 641400.0 ;
      RECT  690600.0 655200.0 700800.0 669000.0 ;
      RECT  690600.0 682800.0 700800.0 669000.0 ;
      RECT  690600.0 682800.0 700800.0 696600.0 ;
      RECT  690600.0 710400.0 700800.0 696600.0 ;
      RECT  690600.0 710400.0 700800.0 724200.0 ;
      RECT  690600.0 738000.0 700800.0 724200.0 ;
      RECT  690600.0 738000.0 700800.0 751800.0 ;
      RECT  690600.0 765600.0 700800.0 751800.0 ;
      RECT  690600.0 765600.0 700800.0 779400.0 ;
      RECT  690600.0 793200.0 700800.0 779400.0 ;
      RECT  690600.0 793200.0 700800.0 807000.0 ;
      RECT  690600.0 820800.0 700800.0 807000.0 ;
      RECT  690600.0 820800.0 700800.0 834600.0 ;
      RECT  690600.0 848400.0 700800.0 834600.0 ;
      RECT  690600.0 848400.0 700800.0 862200.0 ;
      RECT  690600.0 876000.0 700800.0 862200.0 ;
      RECT  690600.0 876000.0 700800.0 889800.0 ;
      RECT  690600.0 903600.0 700800.0 889800.0 ;
      RECT  690600.0 903600.0 700800.0 917400.0 ;
      RECT  690600.0 931200.0 700800.0 917400.0 ;
      RECT  690600.0 931200.0 700800.0 945000.0 ;
      RECT  690600.0 958800.0 700800.0 945000.0 ;
      RECT  690600.0 958800.0 700800.0 972600.0 ;
      RECT  690600.0 986400.0 700800.0 972600.0 ;
      RECT  690600.0 986400.0 700800.0 1000200.0 ;
      RECT  690600.0 1014000.0 700800.0 1000200.0 ;
      RECT  690600.0 1014000.0 700800.0 1027800.0 ;
      RECT  690600.0 1041600.0 700800.0 1027800.0 ;
      RECT  690600.0 1041600.0 700800.0 1055400.0 ;
      RECT  690600.0 1069200.0 700800.0 1055400.0 ;
      RECT  690600.0 1069200.0 700800.0 1083000.0 ;
      RECT  690600.0 1096800.0 700800.0 1083000.0 ;
      RECT  690600.0 1096800.0 700800.0 1110600.0 ;
      RECT  690600.0 1124400.0 700800.0 1110600.0 ;
      RECT  690600.0 1124400.0 700800.0 1138200.0 ;
      RECT  690600.0 1152000.0 700800.0 1138200.0 ;
      RECT  690600.0 1152000.0 700800.0 1165800.0 ;
      RECT  690600.0 1179600.0 700800.0 1165800.0 ;
      RECT  690600.0 1179600.0 700800.0 1193400.0 ;
      RECT  690600.0 1207200.0 700800.0 1193400.0 ;
      RECT  690600.0 1207200.0 700800.0 1221000.0 ;
      RECT  690600.0 1234800.0 700800.0 1221000.0 ;
      RECT  690600.0 1234800.0 700800.0 1248600.0 ;
      RECT  690600.0 1262400.0 700800.0 1248600.0 ;
      RECT  690600.0 1262400.0 700800.0 1276200.0 ;
      RECT  690600.0 1290000.0 700800.0 1276200.0 ;
      RECT  690600.0 1290000.0 700800.0 1303800.0 ;
      RECT  690600.0 1317600.0 700800.0 1303800.0 ;
      RECT  690600.0 1317600.0 700800.0 1331400.0 ;
      RECT  690600.0 1345200.0 700800.0 1331400.0 ;
      RECT  690600.0 1345200.0 700800.0 1359000.0 ;
      RECT  690600.0 1372800.0 700800.0 1359000.0 ;
      RECT  690600.0 1372800.0 700800.0 1386600.0 ;
      RECT  690600.0 1400400.0 700800.0 1386600.0 ;
      RECT  690600.0 1400400.0 700800.0 1414200.0 ;
      RECT  690600.0 1428000.0 700800.0 1414200.0 ;
      RECT  690600.0 1428000.0 700800.0 1441800.0 ;
      RECT  690600.0 1455600.0 700800.0 1441800.0 ;
      RECT  690600.0 1455600.0 700800.0 1469400.0 ;
      RECT  690600.0 1483200.0 700800.0 1469400.0 ;
      RECT  690600.0 1483200.0 700800.0 1497000.0 ;
      RECT  690600.0 1510800.0 700800.0 1497000.0 ;
      RECT  690600.0 1510800.0 700800.0 1524600.0 ;
      RECT  690600.0 1538400.0 700800.0 1524600.0 ;
      RECT  690600.0 1538400.0 700800.0 1552200.0 ;
      RECT  690600.0 1566000.0 700800.0 1552200.0 ;
      RECT  690600.0 1566000.0 700800.0 1579800.0 ;
      RECT  690600.0 1593600.0 700800.0 1579800.0 ;
      RECT  690600.0 1593600.0 700800.0 1607400.0 ;
      RECT  690600.0 1621200.0 700800.0 1607400.0 ;
      RECT  690600.0 1621200.0 700800.0 1635000.0 ;
      RECT  690600.0 1648800.0 700800.0 1635000.0 ;
      RECT  690600.0 1648800.0 700800.0 1662600.0 ;
      RECT  690600.0 1676400.0 700800.0 1662600.0 ;
      RECT  690600.0 1676400.0 700800.0 1690200.0 ;
      RECT  690600.0 1704000.0 700800.0 1690200.0 ;
      RECT  690600.0 1704000.0 700800.0 1717800.0 ;
      RECT  690600.0 1731600.0 700800.0 1717800.0 ;
      RECT  690600.0 1731600.0 700800.0 1745400.0 ;
      RECT  690600.0 1759200.0 700800.0 1745400.0 ;
      RECT  690600.0 1759200.0 700800.0 1773000.0 ;
      RECT  690600.0 1786800.0 700800.0 1773000.0 ;
      RECT  690600.0 1786800.0 700800.0 1800600.0 ;
      RECT  690600.0 1814400.0 700800.0 1800600.0 ;
      RECT  690600.0 1814400.0 700800.0 1828200.0 ;
      RECT  690600.0 1842000.0 700800.0 1828200.0 ;
      RECT  690600.0 1842000.0 700800.0 1855800.0 ;
      RECT  690600.0 1869600.0 700800.0 1855800.0 ;
      RECT  690600.0 1869600.0 700800.0 1883400.0 ;
      RECT  690600.0 1897200.0 700800.0 1883400.0 ;
      RECT  690600.0 1897200.0 700800.0 1911000.0 ;
      RECT  690600.0 1924800.0 700800.0 1911000.0 ;
      RECT  690600.0 1924800.0 700800.0 1938600.0 ;
      RECT  690600.0 1952400.0 700800.0 1938600.0 ;
      RECT  690600.0 1952400.0 700800.0 1966200.0 ;
      RECT  690600.0 1980000.0 700800.0 1966200.0 ;
      RECT  690600.0 1980000.0 700800.0 1993800.0 ;
      RECT  690600.0 2007600.0 700800.0 1993800.0 ;
      RECT  690600.0 2007600.0 700800.0 2021400.0 ;
      RECT  690600.0 2035200.0 700800.0 2021400.0 ;
      RECT  690600.0 2035200.0 700800.0 2049000.0 ;
      RECT  690600.0 2062800.0 700800.0 2049000.0 ;
      RECT  690600.0 2062800.0 700800.0 2076600.0 ;
      RECT  690600.0 2090400.0 700800.0 2076600.0 ;
      RECT  690600.0 2090400.0 700800.0 2104200.0 ;
      RECT  690600.0 2118000.0 700800.0 2104200.0 ;
      RECT  690600.0 2118000.0 700800.0 2131800.0 ;
      RECT  690600.0 2145600.0 700800.0 2131800.0 ;
      RECT  700800.0 379200.0 711000.0 393000.0 ;
      RECT  700800.0 406800.0 711000.0 393000.0 ;
      RECT  700800.0 406800.0 711000.0 420600.0 ;
      RECT  700800.0 434400.0 711000.0 420600.0 ;
      RECT  700800.0 434400.0 711000.0 448200.0 ;
      RECT  700800.0 462000.0 711000.0 448200.0 ;
      RECT  700800.0 462000.0 711000.0 475800.0 ;
      RECT  700800.0 489600.0 711000.0 475800.0 ;
      RECT  700800.0 489600.0 711000.0 503400.0 ;
      RECT  700800.0 517200.0 711000.0 503400.0 ;
      RECT  700800.0 517200.0 711000.0 531000.0 ;
      RECT  700800.0 544800.0 711000.0 531000.0 ;
      RECT  700800.0 544800.0 711000.0 558600.0 ;
      RECT  700800.0 572400.0 711000.0 558600.0 ;
      RECT  700800.0 572400.0 711000.0 586200.0 ;
      RECT  700800.0 600000.0 711000.0 586200.0 ;
      RECT  700800.0 600000.0 711000.0 613800.0 ;
      RECT  700800.0 627600.0 711000.0 613800.0 ;
      RECT  700800.0 627600.0 711000.0 641400.0 ;
      RECT  700800.0 655200.0 711000.0 641400.0 ;
      RECT  700800.0 655200.0 711000.0 669000.0 ;
      RECT  700800.0 682800.0 711000.0 669000.0 ;
      RECT  700800.0 682800.0 711000.0 696600.0 ;
      RECT  700800.0 710400.0 711000.0 696600.0 ;
      RECT  700800.0 710400.0 711000.0 724200.0 ;
      RECT  700800.0 738000.0 711000.0 724200.0 ;
      RECT  700800.0 738000.0 711000.0 751800.0 ;
      RECT  700800.0 765600.0 711000.0 751800.0 ;
      RECT  700800.0 765600.0 711000.0 779400.0 ;
      RECT  700800.0 793200.0 711000.0 779400.0 ;
      RECT  700800.0 793200.0 711000.0 807000.0 ;
      RECT  700800.0 820800.0 711000.0 807000.0 ;
      RECT  700800.0 820800.0 711000.0 834600.0 ;
      RECT  700800.0 848400.0 711000.0 834600.0 ;
      RECT  700800.0 848400.0 711000.0 862200.0 ;
      RECT  700800.0 876000.0 711000.0 862200.0 ;
      RECT  700800.0 876000.0 711000.0 889800.0 ;
      RECT  700800.0 903600.0 711000.0 889800.0 ;
      RECT  700800.0 903600.0 711000.0 917400.0 ;
      RECT  700800.0 931200.0 711000.0 917400.0 ;
      RECT  700800.0 931200.0 711000.0 945000.0 ;
      RECT  700800.0 958800.0 711000.0 945000.0 ;
      RECT  700800.0 958800.0 711000.0 972600.0 ;
      RECT  700800.0 986400.0 711000.0 972600.0 ;
      RECT  700800.0 986400.0 711000.0 1000200.0 ;
      RECT  700800.0 1014000.0 711000.0 1000200.0 ;
      RECT  700800.0 1014000.0 711000.0 1027800.0 ;
      RECT  700800.0 1041600.0 711000.0 1027800.0 ;
      RECT  700800.0 1041600.0 711000.0 1055400.0 ;
      RECT  700800.0 1069200.0 711000.0 1055400.0 ;
      RECT  700800.0 1069200.0 711000.0 1083000.0 ;
      RECT  700800.0 1096800.0 711000.0 1083000.0 ;
      RECT  700800.0 1096800.0 711000.0 1110600.0 ;
      RECT  700800.0 1124400.0 711000.0 1110600.0 ;
      RECT  700800.0 1124400.0 711000.0 1138200.0 ;
      RECT  700800.0 1152000.0 711000.0 1138200.0 ;
      RECT  700800.0 1152000.0 711000.0 1165800.0 ;
      RECT  700800.0 1179600.0 711000.0 1165800.0 ;
      RECT  700800.0 1179600.0 711000.0 1193400.0 ;
      RECT  700800.0 1207200.0 711000.0 1193400.0 ;
      RECT  700800.0 1207200.0 711000.0 1221000.0 ;
      RECT  700800.0 1234800.0 711000.0 1221000.0 ;
      RECT  700800.0 1234800.0 711000.0 1248600.0 ;
      RECT  700800.0 1262400.0 711000.0 1248600.0 ;
      RECT  700800.0 1262400.0 711000.0 1276200.0 ;
      RECT  700800.0 1290000.0 711000.0 1276200.0 ;
      RECT  700800.0 1290000.0 711000.0 1303800.0 ;
      RECT  700800.0 1317600.0 711000.0 1303800.0 ;
      RECT  700800.0 1317600.0 711000.0 1331400.0 ;
      RECT  700800.0 1345200.0 711000.0 1331400.0 ;
      RECT  700800.0 1345200.0 711000.0 1359000.0 ;
      RECT  700800.0 1372800.0 711000.0 1359000.0 ;
      RECT  700800.0 1372800.0 711000.0 1386600.0 ;
      RECT  700800.0 1400400.0 711000.0 1386600.0 ;
      RECT  700800.0 1400400.0 711000.0 1414200.0 ;
      RECT  700800.0 1428000.0 711000.0 1414200.0 ;
      RECT  700800.0 1428000.0 711000.0 1441800.0 ;
      RECT  700800.0 1455600.0 711000.0 1441800.0 ;
      RECT  700800.0 1455600.0 711000.0 1469400.0 ;
      RECT  700800.0 1483200.0 711000.0 1469400.0 ;
      RECT  700800.0 1483200.0 711000.0 1497000.0 ;
      RECT  700800.0 1510800.0 711000.0 1497000.0 ;
      RECT  700800.0 1510800.0 711000.0 1524600.0 ;
      RECT  700800.0 1538400.0 711000.0 1524600.0 ;
      RECT  700800.0 1538400.0 711000.0 1552200.0 ;
      RECT  700800.0 1566000.0 711000.0 1552200.0 ;
      RECT  700800.0 1566000.0 711000.0 1579800.0 ;
      RECT  700800.0 1593600.0 711000.0 1579800.0 ;
      RECT  700800.0 1593600.0 711000.0 1607400.0 ;
      RECT  700800.0 1621200.0 711000.0 1607400.0 ;
      RECT  700800.0 1621200.0 711000.0 1635000.0 ;
      RECT  700800.0 1648800.0 711000.0 1635000.0 ;
      RECT  700800.0 1648800.0 711000.0 1662600.0 ;
      RECT  700800.0 1676400.0 711000.0 1662600.0 ;
      RECT  700800.0 1676400.0 711000.0 1690200.0 ;
      RECT  700800.0 1704000.0 711000.0 1690200.0 ;
      RECT  700800.0 1704000.0 711000.0 1717800.0 ;
      RECT  700800.0 1731600.0 711000.0 1717800.0 ;
      RECT  700800.0 1731600.0 711000.0 1745400.0 ;
      RECT  700800.0 1759200.0 711000.0 1745400.0 ;
      RECT  700800.0 1759200.0 711000.0 1773000.0 ;
      RECT  700800.0 1786800.0 711000.0 1773000.0 ;
      RECT  700800.0 1786800.0 711000.0 1800600.0 ;
      RECT  700800.0 1814400.0 711000.0 1800600.0 ;
      RECT  700800.0 1814400.0 711000.0 1828200.0 ;
      RECT  700800.0 1842000.0 711000.0 1828200.0 ;
      RECT  700800.0 1842000.0 711000.0 1855800.0 ;
      RECT  700800.0 1869600.0 711000.0 1855800.0 ;
      RECT  700800.0 1869600.0 711000.0 1883400.0 ;
      RECT  700800.0 1897200.0 711000.0 1883400.0 ;
      RECT  700800.0 1897200.0 711000.0 1911000.0 ;
      RECT  700800.0 1924800.0 711000.0 1911000.0 ;
      RECT  700800.0 1924800.0 711000.0 1938600.0 ;
      RECT  700800.0 1952400.0 711000.0 1938600.0 ;
      RECT  700800.0 1952400.0 711000.0 1966200.0 ;
      RECT  700800.0 1980000.0 711000.0 1966200.0 ;
      RECT  700800.0 1980000.0 711000.0 1993800.0 ;
      RECT  700800.0 2007600.0 711000.0 1993800.0 ;
      RECT  700800.0 2007600.0 711000.0 2021400.0 ;
      RECT  700800.0 2035200.0 711000.0 2021400.0 ;
      RECT  700800.0 2035200.0 711000.0 2049000.0 ;
      RECT  700800.0 2062800.0 711000.0 2049000.0 ;
      RECT  700800.0 2062800.0 711000.0 2076600.0 ;
      RECT  700800.0 2090400.0 711000.0 2076600.0 ;
      RECT  700800.0 2090400.0 711000.0 2104200.0 ;
      RECT  700800.0 2118000.0 711000.0 2104200.0 ;
      RECT  700800.0 2118000.0 711000.0 2131800.0 ;
      RECT  700800.0 2145600.0 711000.0 2131800.0 ;
      RECT  711000.0 379200.0 721200.0 393000.0 ;
      RECT  711000.0 406800.0 721200.0 393000.0 ;
      RECT  711000.0 406800.0 721200.0 420600.0 ;
      RECT  711000.0 434400.0 721200.0 420600.0 ;
      RECT  711000.0 434400.0 721200.0 448200.0 ;
      RECT  711000.0 462000.0 721200.0 448200.0 ;
      RECT  711000.0 462000.0 721200.0 475800.0 ;
      RECT  711000.0 489600.0 721200.0 475800.0 ;
      RECT  711000.0 489600.0 721200.0 503400.0 ;
      RECT  711000.0 517200.0 721200.0 503400.0 ;
      RECT  711000.0 517200.0 721200.0 531000.0 ;
      RECT  711000.0 544800.0 721200.0 531000.0 ;
      RECT  711000.0 544800.0 721200.0 558600.0 ;
      RECT  711000.0 572400.0 721200.0 558600.0 ;
      RECT  711000.0 572400.0 721200.0 586200.0 ;
      RECT  711000.0 600000.0 721200.0 586200.0 ;
      RECT  711000.0 600000.0 721200.0 613800.0 ;
      RECT  711000.0 627600.0 721200.0 613800.0 ;
      RECT  711000.0 627600.0 721200.0 641400.0 ;
      RECT  711000.0 655200.0 721200.0 641400.0 ;
      RECT  711000.0 655200.0 721200.0 669000.0 ;
      RECT  711000.0 682800.0 721200.0 669000.0 ;
      RECT  711000.0 682800.0 721200.0 696600.0 ;
      RECT  711000.0 710400.0 721200.0 696600.0 ;
      RECT  711000.0 710400.0 721200.0 724200.0 ;
      RECT  711000.0 738000.0 721200.0 724200.0 ;
      RECT  711000.0 738000.0 721200.0 751800.0 ;
      RECT  711000.0 765600.0 721200.0 751800.0 ;
      RECT  711000.0 765600.0 721200.0 779400.0 ;
      RECT  711000.0 793200.0 721200.0 779400.0 ;
      RECT  711000.0 793200.0 721200.0 807000.0 ;
      RECT  711000.0 820800.0 721200.0 807000.0 ;
      RECT  711000.0 820800.0 721200.0 834600.0 ;
      RECT  711000.0 848400.0 721200.0 834600.0 ;
      RECT  711000.0 848400.0 721200.0 862200.0 ;
      RECT  711000.0 876000.0 721200.0 862200.0 ;
      RECT  711000.0 876000.0 721200.0 889800.0 ;
      RECT  711000.0 903600.0 721200.0 889800.0 ;
      RECT  711000.0 903600.0 721200.0 917400.0 ;
      RECT  711000.0 931200.0 721200.0 917400.0 ;
      RECT  711000.0 931200.0 721200.0 945000.0 ;
      RECT  711000.0 958800.0 721200.0 945000.0 ;
      RECT  711000.0 958800.0 721200.0 972600.0 ;
      RECT  711000.0 986400.0 721200.0 972600.0 ;
      RECT  711000.0 986400.0 721200.0 1000200.0 ;
      RECT  711000.0 1014000.0 721200.0 1000200.0 ;
      RECT  711000.0 1014000.0 721200.0 1027800.0 ;
      RECT  711000.0 1041600.0 721200.0 1027800.0 ;
      RECT  711000.0 1041600.0 721200.0 1055400.0 ;
      RECT  711000.0 1069200.0 721200.0 1055400.0 ;
      RECT  711000.0 1069200.0 721200.0 1083000.0 ;
      RECT  711000.0 1096800.0 721200.0 1083000.0 ;
      RECT  711000.0 1096800.0 721200.0 1110600.0 ;
      RECT  711000.0 1124400.0 721200.0 1110600.0 ;
      RECT  711000.0 1124400.0 721200.0 1138200.0 ;
      RECT  711000.0 1152000.0 721200.0 1138200.0 ;
      RECT  711000.0 1152000.0 721200.0 1165800.0 ;
      RECT  711000.0 1179600.0 721200.0 1165800.0 ;
      RECT  711000.0 1179600.0 721200.0 1193400.0 ;
      RECT  711000.0 1207200.0 721200.0 1193400.0 ;
      RECT  711000.0 1207200.0 721200.0 1221000.0 ;
      RECT  711000.0 1234800.0 721200.0 1221000.0 ;
      RECT  711000.0 1234800.0 721200.0 1248600.0 ;
      RECT  711000.0 1262400.0 721200.0 1248600.0 ;
      RECT  711000.0 1262400.0 721200.0 1276200.0 ;
      RECT  711000.0 1290000.0 721200.0 1276200.0 ;
      RECT  711000.0 1290000.0 721200.0 1303800.0 ;
      RECT  711000.0 1317600.0 721200.0 1303800.0 ;
      RECT  711000.0 1317600.0 721200.0 1331400.0 ;
      RECT  711000.0 1345200.0 721200.0 1331400.0 ;
      RECT  711000.0 1345200.0 721200.0 1359000.0 ;
      RECT  711000.0 1372800.0 721200.0 1359000.0 ;
      RECT  711000.0 1372800.0 721200.0 1386600.0 ;
      RECT  711000.0 1400400.0 721200.0 1386600.0 ;
      RECT  711000.0 1400400.0 721200.0 1414200.0 ;
      RECT  711000.0 1428000.0 721200.0 1414200.0 ;
      RECT  711000.0 1428000.0 721200.0 1441800.0 ;
      RECT  711000.0 1455600.0 721200.0 1441800.0 ;
      RECT  711000.0 1455600.0 721200.0 1469400.0 ;
      RECT  711000.0 1483200.0 721200.0 1469400.0 ;
      RECT  711000.0 1483200.0 721200.0 1497000.0 ;
      RECT  711000.0 1510800.0 721200.0 1497000.0 ;
      RECT  711000.0 1510800.0 721200.0 1524600.0 ;
      RECT  711000.0 1538400.0 721200.0 1524600.0 ;
      RECT  711000.0 1538400.0 721200.0 1552200.0 ;
      RECT  711000.0 1566000.0 721200.0 1552200.0 ;
      RECT  711000.0 1566000.0 721200.0 1579800.0 ;
      RECT  711000.0 1593600.0 721200.0 1579800.0 ;
      RECT  711000.0 1593600.0 721200.0 1607400.0 ;
      RECT  711000.0 1621200.0 721200.0 1607400.0 ;
      RECT  711000.0 1621200.0 721200.0 1635000.0 ;
      RECT  711000.0 1648800.0 721200.0 1635000.0 ;
      RECT  711000.0 1648800.0 721200.0 1662600.0 ;
      RECT  711000.0 1676400.0 721200.0 1662600.0 ;
      RECT  711000.0 1676400.0 721200.0 1690200.0 ;
      RECT  711000.0 1704000.0 721200.0 1690200.0 ;
      RECT  711000.0 1704000.0 721200.0 1717800.0 ;
      RECT  711000.0 1731600.0 721200.0 1717800.0 ;
      RECT  711000.0 1731600.0 721200.0 1745400.0 ;
      RECT  711000.0 1759200.0 721200.0 1745400.0 ;
      RECT  711000.0 1759200.0 721200.0 1773000.0 ;
      RECT  711000.0 1786800.0 721200.0 1773000.0 ;
      RECT  711000.0 1786800.0 721200.0 1800600.0 ;
      RECT  711000.0 1814400.0 721200.0 1800600.0 ;
      RECT  711000.0 1814400.0 721200.0 1828200.0 ;
      RECT  711000.0 1842000.0 721200.0 1828200.0 ;
      RECT  711000.0 1842000.0 721200.0 1855800.0 ;
      RECT  711000.0 1869600.0 721200.0 1855800.0 ;
      RECT  711000.0 1869600.0 721200.0 1883400.0 ;
      RECT  711000.0 1897200.0 721200.0 1883400.0 ;
      RECT  711000.0 1897200.0 721200.0 1911000.0 ;
      RECT  711000.0 1924800.0 721200.0 1911000.0 ;
      RECT  711000.0 1924800.0 721200.0 1938600.0 ;
      RECT  711000.0 1952400.0 721200.0 1938600.0 ;
      RECT  711000.0 1952400.0 721200.0 1966200.0 ;
      RECT  711000.0 1980000.0 721200.0 1966200.0 ;
      RECT  711000.0 1980000.0 721200.0 1993800.0 ;
      RECT  711000.0 2007600.0 721200.0 1993800.0 ;
      RECT  711000.0 2007600.0 721200.0 2021400.0 ;
      RECT  711000.0 2035200.0 721200.0 2021400.0 ;
      RECT  711000.0 2035200.0 721200.0 2049000.0 ;
      RECT  711000.0 2062800.0 721200.0 2049000.0 ;
      RECT  711000.0 2062800.0 721200.0 2076600.0 ;
      RECT  711000.0 2090400.0 721200.0 2076600.0 ;
      RECT  711000.0 2090400.0 721200.0 2104200.0 ;
      RECT  711000.0 2118000.0 721200.0 2104200.0 ;
      RECT  711000.0 2118000.0 721200.0 2131800.0 ;
      RECT  711000.0 2145600.0 721200.0 2131800.0 ;
      RECT  721200.0 379200.0 731400.0 393000.0 ;
      RECT  721200.0 406800.0 731400.0 393000.0 ;
      RECT  721200.0 406800.0 731400.0 420600.0 ;
      RECT  721200.0 434400.0 731400.0 420600.0 ;
      RECT  721200.0 434400.0 731400.0 448200.0 ;
      RECT  721200.0 462000.0 731400.0 448200.0 ;
      RECT  721200.0 462000.0 731400.0 475800.0 ;
      RECT  721200.0 489600.0 731400.0 475800.0 ;
      RECT  721200.0 489600.0 731400.0 503400.0 ;
      RECT  721200.0 517200.0 731400.0 503400.0 ;
      RECT  721200.0 517200.0 731400.0 531000.0 ;
      RECT  721200.0 544800.0 731400.0 531000.0 ;
      RECT  721200.0 544800.0 731400.0 558600.0 ;
      RECT  721200.0 572400.0 731400.0 558600.0 ;
      RECT  721200.0 572400.0 731400.0 586200.0 ;
      RECT  721200.0 600000.0 731400.0 586200.0 ;
      RECT  721200.0 600000.0 731400.0 613800.0 ;
      RECT  721200.0 627600.0 731400.0 613800.0 ;
      RECT  721200.0 627600.0 731400.0 641400.0 ;
      RECT  721200.0 655200.0 731400.0 641400.0 ;
      RECT  721200.0 655200.0 731400.0 669000.0 ;
      RECT  721200.0 682800.0 731400.0 669000.0 ;
      RECT  721200.0 682800.0 731400.0 696600.0 ;
      RECT  721200.0 710400.0 731400.0 696600.0 ;
      RECT  721200.0 710400.0 731400.0 724200.0 ;
      RECT  721200.0 738000.0 731400.0 724200.0 ;
      RECT  721200.0 738000.0 731400.0 751800.0 ;
      RECT  721200.0 765600.0 731400.0 751800.0 ;
      RECT  721200.0 765600.0 731400.0 779400.0 ;
      RECT  721200.0 793200.0 731400.0 779400.0 ;
      RECT  721200.0 793200.0 731400.0 807000.0 ;
      RECT  721200.0 820800.0 731400.0 807000.0 ;
      RECT  721200.0 820800.0 731400.0 834600.0 ;
      RECT  721200.0 848400.0 731400.0 834600.0 ;
      RECT  721200.0 848400.0 731400.0 862200.0 ;
      RECT  721200.0 876000.0 731400.0 862200.0 ;
      RECT  721200.0 876000.0 731400.0 889800.0 ;
      RECT  721200.0 903600.0 731400.0 889800.0 ;
      RECT  721200.0 903600.0 731400.0 917400.0 ;
      RECT  721200.0 931200.0 731400.0 917400.0 ;
      RECT  721200.0 931200.0 731400.0 945000.0 ;
      RECT  721200.0 958800.0 731400.0 945000.0 ;
      RECT  721200.0 958800.0 731400.0 972600.0 ;
      RECT  721200.0 986400.0 731400.0 972600.0 ;
      RECT  721200.0 986400.0 731400.0 1000200.0 ;
      RECT  721200.0 1014000.0 731400.0 1000200.0 ;
      RECT  721200.0 1014000.0 731400.0 1027800.0 ;
      RECT  721200.0 1041600.0 731400.0 1027800.0 ;
      RECT  721200.0 1041600.0 731400.0 1055400.0 ;
      RECT  721200.0 1069200.0 731400.0 1055400.0 ;
      RECT  721200.0 1069200.0 731400.0 1083000.0 ;
      RECT  721200.0 1096800.0 731400.0 1083000.0 ;
      RECT  721200.0 1096800.0 731400.0 1110600.0 ;
      RECT  721200.0 1124400.0 731400.0 1110600.0 ;
      RECT  721200.0 1124400.0 731400.0 1138200.0 ;
      RECT  721200.0 1152000.0 731400.0 1138200.0 ;
      RECT  721200.0 1152000.0 731400.0 1165800.0 ;
      RECT  721200.0 1179600.0 731400.0 1165800.0 ;
      RECT  721200.0 1179600.0 731400.0 1193400.0 ;
      RECT  721200.0 1207200.0 731400.0 1193400.0 ;
      RECT  721200.0 1207200.0 731400.0 1221000.0 ;
      RECT  721200.0 1234800.0 731400.0 1221000.0 ;
      RECT  721200.0 1234800.0 731400.0 1248600.0 ;
      RECT  721200.0 1262400.0 731400.0 1248600.0 ;
      RECT  721200.0 1262400.0 731400.0 1276200.0 ;
      RECT  721200.0 1290000.0 731400.0 1276200.0 ;
      RECT  721200.0 1290000.0 731400.0 1303800.0 ;
      RECT  721200.0 1317600.0 731400.0 1303800.0 ;
      RECT  721200.0 1317600.0 731400.0 1331400.0 ;
      RECT  721200.0 1345200.0 731400.0 1331400.0 ;
      RECT  721200.0 1345200.0 731400.0 1359000.0 ;
      RECT  721200.0 1372800.0 731400.0 1359000.0 ;
      RECT  721200.0 1372800.0 731400.0 1386600.0 ;
      RECT  721200.0 1400400.0 731400.0 1386600.0 ;
      RECT  721200.0 1400400.0 731400.0 1414200.0 ;
      RECT  721200.0 1428000.0 731400.0 1414200.0 ;
      RECT  721200.0 1428000.0 731400.0 1441800.0 ;
      RECT  721200.0 1455600.0 731400.0 1441800.0 ;
      RECT  721200.0 1455600.0 731400.0 1469400.0 ;
      RECT  721200.0 1483200.0 731400.0 1469400.0 ;
      RECT  721200.0 1483200.0 731400.0 1497000.0 ;
      RECT  721200.0 1510800.0 731400.0 1497000.0 ;
      RECT  721200.0 1510800.0 731400.0 1524600.0 ;
      RECT  721200.0 1538400.0 731400.0 1524600.0 ;
      RECT  721200.0 1538400.0 731400.0 1552200.0 ;
      RECT  721200.0 1566000.0 731400.0 1552200.0 ;
      RECT  721200.0 1566000.0 731400.0 1579800.0 ;
      RECT  721200.0 1593600.0 731400.0 1579800.0 ;
      RECT  721200.0 1593600.0 731400.0 1607400.0 ;
      RECT  721200.0 1621200.0 731400.0 1607400.0 ;
      RECT  721200.0 1621200.0 731400.0 1635000.0 ;
      RECT  721200.0 1648800.0 731400.0 1635000.0 ;
      RECT  721200.0 1648800.0 731400.0 1662600.0 ;
      RECT  721200.0 1676400.0 731400.0 1662600.0 ;
      RECT  721200.0 1676400.0 731400.0 1690200.0 ;
      RECT  721200.0 1704000.0 731400.0 1690200.0 ;
      RECT  721200.0 1704000.0 731400.0 1717800.0 ;
      RECT  721200.0 1731600.0 731400.0 1717800.0 ;
      RECT  721200.0 1731600.0 731400.0 1745400.0 ;
      RECT  721200.0 1759200.0 731400.0 1745400.0 ;
      RECT  721200.0 1759200.0 731400.0 1773000.0 ;
      RECT  721200.0 1786800.0 731400.0 1773000.0 ;
      RECT  721200.0 1786800.0 731400.0 1800600.0 ;
      RECT  721200.0 1814400.0 731400.0 1800600.0 ;
      RECT  721200.0 1814400.0 731400.0 1828200.0 ;
      RECT  721200.0 1842000.0 731400.0 1828200.0 ;
      RECT  721200.0 1842000.0 731400.0 1855800.0 ;
      RECT  721200.0 1869600.0 731400.0 1855800.0 ;
      RECT  721200.0 1869600.0 731400.0 1883400.0 ;
      RECT  721200.0 1897200.0 731400.0 1883400.0 ;
      RECT  721200.0 1897200.0 731400.0 1911000.0 ;
      RECT  721200.0 1924800.0 731400.0 1911000.0 ;
      RECT  721200.0 1924800.0 731400.0 1938600.0 ;
      RECT  721200.0 1952400.0 731400.0 1938600.0 ;
      RECT  721200.0 1952400.0 731400.0 1966200.0 ;
      RECT  721200.0 1980000.0 731400.0 1966200.0 ;
      RECT  721200.0 1980000.0 731400.0 1993800.0 ;
      RECT  721200.0 2007600.0 731400.0 1993800.0 ;
      RECT  721200.0 2007600.0 731400.0 2021400.0 ;
      RECT  721200.0 2035200.0 731400.0 2021400.0 ;
      RECT  721200.0 2035200.0 731400.0 2049000.0 ;
      RECT  721200.0 2062800.0 731400.0 2049000.0 ;
      RECT  721200.0 2062800.0 731400.0 2076600.0 ;
      RECT  721200.0 2090400.0 731400.0 2076600.0 ;
      RECT  721200.0 2090400.0 731400.0 2104200.0 ;
      RECT  721200.0 2118000.0 731400.0 2104200.0 ;
      RECT  721200.0 2118000.0 731400.0 2131800.0 ;
      RECT  721200.0 2145600.0 731400.0 2131800.0 ;
      RECT  731400.0 379200.0 741600.0 393000.0 ;
      RECT  731400.0 406800.0 741600.0 393000.0 ;
      RECT  731400.0 406800.0 741600.0 420600.0 ;
      RECT  731400.0 434400.0 741600.0 420600.0 ;
      RECT  731400.0 434400.0 741600.0 448200.0 ;
      RECT  731400.0 462000.0 741600.0 448200.0 ;
      RECT  731400.0 462000.0 741600.0 475800.0 ;
      RECT  731400.0 489600.0 741600.0 475800.0 ;
      RECT  731400.0 489600.0 741600.0 503400.0 ;
      RECT  731400.0 517200.0 741600.0 503400.0 ;
      RECT  731400.0 517200.0 741600.0 531000.0 ;
      RECT  731400.0 544800.0 741600.0 531000.0 ;
      RECT  731400.0 544800.0 741600.0 558600.0 ;
      RECT  731400.0 572400.0 741600.0 558600.0 ;
      RECT  731400.0 572400.0 741600.0 586200.0 ;
      RECT  731400.0 600000.0 741600.0 586200.0 ;
      RECT  731400.0 600000.0 741600.0 613800.0 ;
      RECT  731400.0 627600.0 741600.0 613800.0 ;
      RECT  731400.0 627600.0 741600.0 641400.0 ;
      RECT  731400.0 655200.0 741600.0 641400.0 ;
      RECT  731400.0 655200.0 741600.0 669000.0 ;
      RECT  731400.0 682800.0 741600.0 669000.0 ;
      RECT  731400.0 682800.0 741600.0 696600.0 ;
      RECT  731400.0 710400.0 741600.0 696600.0 ;
      RECT  731400.0 710400.0 741600.0 724200.0 ;
      RECT  731400.0 738000.0 741600.0 724200.0 ;
      RECT  731400.0 738000.0 741600.0 751800.0 ;
      RECT  731400.0 765600.0 741600.0 751800.0 ;
      RECT  731400.0 765600.0 741600.0 779400.0 ;
      RECT  731400.0 793200.0 741600.0 779400.0 ;
      RECT  731400.0 793200.0 741600.0 807000.0 ;
      RECT  731400.0 820800.0 741600.0 807000.0 ;
      RECT  731400.0 820800.0 741600.0 834600.0 ;
      RECT  731400.0 848400.0 741600.0 834600.0 ;
      RECT  731400.0 848400.0 741600.0 862200.0 ;
      RECT  731400.0 876000.0 741600.0 862200.0 ;
      RECT  731400.0 876000.0 741600.0 889800.0 ;
      RECT  731400.0 903600.0 741600.0 889800.0 ;
      RECT  731400.0 903600.0 741600.0 917400.0 ;
      RECT  731400.0 931200.0 741600.0 917400.0 ;
      RECT  731400.0 931200.0 741600.0 945000.0 ;
      RECT  731400.0 958800.0 741600.0 945000.0 ;
      RECT  731400.0 958800.0 741600.0 972600.0 ;
      RECT  731400.0 986400.0 741600.0 972600.0 ;
      RECT  731400.0 986400.0 741600.0 1000200.0 ;
      RECT  731400.0 1014000.0 741600.0 1000200.0 ;
      RECT  731400.0 1014000.0 741600.0 1027800.0 ;
      RECT  731400.0 1041600.0 741600.0 1027800.0 ;
      RECT  731400.0 1041600.0 741600.0 1055400.0 ;
      RECT  731400.0 1069200.0 741600.0 1055400.0 ;
      RECT  731400.0 1069200.0 741600.0 1083000.0 ;
      RECT  731400.0 1096800.0 741600.0 1083000.0 ;
      RECT  731400.0 1096800.0 741600.0 1110600.0 ;
      RECT  731400.0 1124400.0 741600.0 1110600.0 ;
      RECT  731400.0 1124400.0 741600.0 1138200.0 ;
      RECT  731400.0 1152000.0 741600.0 1138200.0 ;
      RECT  731400.0 1152000.0 741600.0 1165800.0 ;
      RECT  731400.0 1179600.0 741600.0 1165800.0 ;
      RECT  731400.0 1179600.0 741600.0 1193400.0 ;
      RECT  731400.0 1207200.0 741600.0 1193400.0 ;
      RECT  731400.0 1207200.0 741600.0 1221000.0 ;
      RECT  731400.0 1234800.0 741600.0 1221000.0 ;
      RECT  731400.0 1234800.0 741600.0 1248600.0 ;
      RECT  731400.0 1262400.0 741600.0 1248600.0 ;
      RECT  731400.0 1262400.0 741600.0 1276200.0 ;
      RECT  731400.0 1290000.0 741600.0 1276200.0 ;
      RECT  731400.0 1290000.0 741600.0 1303800.0 ;
      RECT  731400.0 1317600.0 741600.0 1303800.0 ;
      RECT  731400.0 1317600.0 741600.0 1331400.0 ;
      RECT  731400.0 1345200.0 741600.0 1331400.0 ;
      RECT  731400.0 1345200.0 741600.0 1359000.0 ;
      RECT  731400.0 1372800.0 741600.0 1359000.0 ;
      RECT  731400.0 1372800.0 741600.0 1386600.0 ;
      RECT  731400.0 1400400.0 741600.0 1386600.0 ;
      RECT  731400.0 1400400.0 741600.0 1414200.0 ;
      RECT  731400.0 1428000.0 741600.0 1414200.0 ;
      RECT  731400.0 1428000.0 741600.0 1441800.0 ;
      RECT  731400.0 1455600.0 741600.0 1441800.0 ;
      RECT  731400.0 1455600.0 741600.0 1469400.0 ;
      RECT  731400.0 1483200.0 741600.0 1469400.0 ;
      RECT  731400.0 1483200.0 741600.0 1497000.0 ;
      RECT  731400.0 1510800.0 741600.0 1497000.0 ;
      RECT  731400.0 1510800.0 741600.0 1524600.0 ;
      RECT  731400.0 1538400.0 741600.0 1524600.0 ;
      RECT  731400.0 1538400.0 741600.0 1552200.0 ;
      RECT  731400.0 1566000.0 741600.0 1552200.0 ;
      RECT  731400.0 1566000.0 741600.0 1579800.0 ;
      RECT  731400.0 1593600.0 741600.0 1579800.0 ;
      RECT  731400.0 1593600.0 741600.0 1607400.0 ;
      RECT  731400.0 1621200.0 741600.0 1607400.0 ;
      RECT  731400.0 1621200.0 741600.0 1635000.0 ;
      RECT  731400.0 1648800.0 741600.0 1635000.0 ;
      RECT  731400.0 1648800.0 741600.0 1662600.0 ;
      RECT  731400.0 1676400.0 741600.0 1662600.0 ;
      RECT  731400.0 1676400.0 741600.0 1690200.0 ;
      RECT  731400.0 1704000.0 741600.0 1690200.0 ;
      RECT  731400.0 1704000.0 741600.0 1717800.0 ;
      RECT  731400.0 1731600.0 741600.0 1717800.0 ;
      RECT  731400.0 1731600.0 741600.0 1745400.0 ;
      RECT  731400.0 1759200.0 741600.0 1745400.0 ;
      RECT  731400.0 1759200.0 741600.0 1773000.0 ;
      RECT  731400.0 1786800.0 741600.0 1773000.0 ;
      RECT  731400.0 1786800.0 741600.0 1800600.0 ;
      RECT  731400.0 1814400.0 741600.0 1800600.0 ;
      RECT  731400.0 1814400.0 741600.0 1828200.0 ;
      RECT  731400.0 1842000.0 741600.0 1828200.0 ;
      RECT  731400.0 1842000.0 741600.0 1855800.0 ;
      RECT  731400.0 1869600.0 741600.0 1855800.0 ;
      RECT  731400.0 1869600.0 741600.0 1883400.0 ;
      RECT  731400.0 1897200.0 741600.0 1883400.0 ;
      RECT  731400.0 1897200.0 741600.0 1911000.0 ;
      RECT  731400.0 1924800.0 741600.0 1911000.0 ;
      RECT  731400.0 1924800.0 741600.0 1938600.0 ;
      RECT  731400.0 1952400.0 741600.0 1938600.0 ;
      RECT  731400.0 1952400.0 741600.0 1966200.0 ;
      RECT  731400.0 1980000.0 741600.0 1966200.0 ;
      RECT  731400.0 1980000.0 741600.0 1993800.0 ;
      RECT  731400.0 2007600.0 741600.0 1993800.0 ;
      RECT  731400.0 2007600.0 741600.0 2021400.0 ;
      RECT  731400.0 2035200.0 741600.0 2021400.0 ;
      RECT  731400.0 2035200.0 741600.0 2049000.0 ;
      RECT  731400.0 2062800.0 741600.0 2049000.0 ;
      RECT  731400.0 2062800.0 741600.0 2076600.0 ;
      RECT  731400.0 2090400.0 741600.0 2076600.0 ;
      RECT  731400.0 2090400.0 741600.0 2104200.0 ;
      RECT  731400.0 2118000.0 741600.0 2104200.0 ;
      RECT  731400.0 2118000.0 741600.0 2131800.0 ;
      RECT  731400.0 2145600.0 741600.0 2131800.0 ;
      RECT  741600.0 379200.0 751800.0 393000.0 ;
      RECT  741600.0 406800.0 751800.0 393000.0 ;
      RECT  741600.0 406800.0 751800.0 420600.0 ;
      RECT  741600.0 434400.0 751800.0 420600.0 ;
      RECT  741600.0 434400.0 751800.0 448200.0 ;
      RECT  741600.0 462000.0 751800.0 448200.0 ;
      RECT  741600.0 462000.0 751800.0 475800.0 ;
      RECT  741600.0 489600.0 751800.0 475800.0 ;
      RECT  741600.0 489600.0 751800.0 503400.0 ;
      RECT  741600.0 517200.0 751800.0 503400.0 ;
      RECT  741600.0 517200.0 751800.0 531000.0 ;
      RECT  741600.0 544800.0 751800.0 531000.0 ;
      RECT  741600.0 544800.0 751800.0 558600.0 ;
      RECT  741600.0 572400.0 751800.0 558600.0 ;
      RECT  741600.0 572400.0 751800.0 586200.0 ;
      RECT  741600.0 600000.0 751800.0 586200.0 ;
      RECT  741600.0 600000.0 751800.0 613800.0 ;
      RECT  741600.0 627600.0 751800.0 613800.0 ;
      RECT  741600.0 627600.0 751800.0 641400.0 ;
      RECT  741600.0 655200.0 751800.0 641400.0 ;
      RECT  741600.0 655200.0 751800.0 669000.0 ;
      RECT  741600.0 682800.0 751800.0 669000.0 ;
      RECT  741600.0 682800.0 751800.0 696600.0 ;
      RECT  741600.0 710400.0 751800.0 696600.0 ;
      RECT  741600.0 710400.0 751800.0 724200.0 ;
      RECT  741600.0 738000.0 751800.0 724200.0 ;
      RECT  741600.0 738000.0 751800.0 751800.0 ;
      RECT  741600.0 765600.0 751800.0 751800.0 ;
      RECT  741600.0 765600.0 751800.0 779400.0 ;
      RECT  741600.0 793200.0 751800.0 779400.0 ;
      RECT  741600.0 793200.0 751800.0 807000.0 ;
      RECT  741600.0 820800.0 751800.0 807000.0 ;
      RECT  741600.0 820800.0 751800.0 834600.0 ;
      RECT  741600.0 848400.0 751800.0 834600.0 ;
      RECT  741600.0 848400.0 751800.0 862200.0 ;
      RECT  741600.0 876000.0 751800.0 862200.0 ;
      RECT  741600.0 876000.0 751800.0 889800.0 ;
      RECT  741600.0 903600.0 751800.0 889800.0 ;
      RECT  741600.0 903600.0 751800.0 917400.0 ;
      RECT  741600.0 931200.0 751800.0 917400.0 ;
      RECT  741600.0 931200.0 751800.0 945000.0 ;
      RECT  741600.0 958800.0 751800.0 945000.0 ;
      RECT  741600.0 958800.0 751800.0 972600.0 ;
      RECT  741600.0 986400.0 751800.0 972600.0 ;
      RECT  741600.0 986400.0 751800.0 1000200.0 ;
      RECT  741600.0 1014000.0 751800.0 1000200.0 ;
      RECT  741600.0 1014000.0 751800.0 1027800.0 ;
      RECT  741600.0 1041600.0 751800.0 1027800.0 ;
      RECT  741600.0 1041600.0 751800.0 1055400.0 ;
      RECT  741600.0 1069200.0 751800.0 1055400.0 ;
      RECT  741600.0 1069200.0 751800.0 1083000.0 ;
      RECT  741600.0 1096800.0 751800.0 1083000.0 ;
      RECT  741600.0 1096800.0 751800.0 1110600.0 ;
      RECT  741600.0 1124400.0 751800.0 1110600.0 ;
      RECT  741600.0 1124400.0 751800.0 1138200.0 ;
      RECT  741600.0 1152000.0 751800.0 1138200.0 ;
      RECT  741600.0 1152000.0 751800.0 1165800.0 ;
      RECT  741600.0 1179600.0 751800.0 1165800.0 ;
      RECT  741600.0 1179600.0 751800.0 1193400.0 ;
      RECT  741600.0 1207200.0 751800.0 1193400.0 ;
      RECT  741600.0 1207200.0 751800.0 1221000.0 ;
      RECT  741600.0 1234800.0 751800.0 1221000.0 ;
      RECT  741600.0 1234800.0 751800.0 1248600.0 ;
      RECT  741600.0 1262400.0 751800.0 1248600.0 ;
      RECT  741600.0 1262400.0 751800.0 1276200.0 ;
      RECT  741600.0 1290000.0 751800.0 1276200.0 ;
      RECT  741600.0 1290000.0 751800.0 1303800.0 ;
      RECT  741600.0 1317600.0 751800.0 1303800.0 ;
      RECT  741600.0 1317600.0 751800.0 1331400.0 ;
      RECT  741600.0 1345200.0 751800.0 1331400.0 ;
      RECT  741600.0 1345200.0 751800.0 1359000.0 ;
      RECT  741600.0 1372800.0 751800.0 1359000.0 ;
      RECT  741600.0 1372800.0 751800.0 1386600.0 ;
      RECT  741600.0 1400400.0 751800.0 1386600.0 ;
      RECT  741600.0 1400400.0 751800.0 1414200.0 ;
      RECT  741600.0 1428000.0 751800.0 1414200.0 ;
      RECT  741600.0 1428000.0 751800.0 1441800.0 ;
      RECT  741600.0 1455600.0 751800.0 1441800.0 ;
      RECT  741600.0 1455600.0 751800.0 1469400.0 ;
      RECT  741600.0 1483200.0 751800.0 1469400.0 ;
      RECT  741600.0 1483200.0 751800.0 1497000.0 ;
      RECT  741600.0 1510800.0 751800.0 1497000.0 ;
      RECT  741600.0 1510800.0 751800.0 1524600.0 ;
      RECT  741600.0 1538400.0 751800.0 1524600.0 ;
      RECT  741600.0 1538400.0 751800.0 1552200.0 ;
      RECT  741600.0 1566000.0 751800.0 1552200.0 ;
      RECT  741600.0 1566000.0 751800.0 1579800.0 ;
      RECT  741600.0 1593600.0 751800.0 1579800.0 ;
      RECT  741600.0 1593600.0 751800.0 1607400.0 ;
      RECT  741600.0 1621200.0 751800.0 1607400.0 ;
      RECT  741600.0 1621200.0 751800.0 1635000.0 ;
      RECT  741600.0 1648800.0 751800.0 1635000.0 ;
      RECT  741600.0 1648800.0 751800.0 1662600.0 ;
      RECT  741600.0 1676400.0 751800.0 1662600.0 ;
      RECT  741600.0 1676400.0 751800.0 1690200.0 ;
      RECT  741600.0 1704000.0 751800.0 1690200.0 ;
      RECT  741600.0 1704000.0 751800.0 1717800.0 ;
      RECT  741600.0 1731600.0 751800.0 1717800.0 ;
      RECT  741600.0 1731600.0 751800.0 1745400.0 ;
      RECT  741600.0 1759200.0 751800.0 1745400.0 ;
      RECT  741600.0 1759200.0 751800.0 1773000.0 ;
      RECT  741600.0 1786800.0 751800.0 1773000.0 ;
      RECT  741600.0 1786800.0 751800.0 1800600.0 ;
      RECT  741600.0 1814400.0 751800.0 1800600.0 ;
      RECT  741600.0 1814400.0 751800.0 1828200.0 ;
      RECT  741600.0 1842000.0 751800.0 1828200.0 ;
      RECT  741600.0 1842000.0 751800.0 1855800.0 ;
      RECT  741600.0 1869600.0 751800.0 1855800.0 ;
      RECT  741600.0 1869600.0 751800.0 1883400.0 ;
      RECT  741600.0 1897200.0 751800.0 1883400.0 ;
      RECT  741600.0 1897200.0 751800.0 1911000.0 ;
      RECT  741600.0 1924800.0 751800.0 1911000.0 ;
      RECT  741600.0 1924800.0 751800.0 1938600.0 ;
      RECT  741600.0 1952400.0 751800.0 1938600.0 ;
      RECT  741600.0 1952400.0 751800.0 1966200.0 ;
      RECT  741600.0 1980000.0 751800.0 1966200.0 ;
      RECT  741600.0 1980000.0 751800.0 1993800.0 ;
      RECT  741600.0 2007600.0 751800.0 1993800.0 ;
      RECT  741600.0 2007600.0 751800.0 2021400.0 ;
      RECT  741600.0 2035200.0 751800.0 2021400.0 ;
      RECT  741600.0 2035200.0 751800.0 2049000.0 ;
      RECT  741600.0 2062800.0 751800.0 2049000.0 ;
      RECT  741600.0 2062800.0 751800.0 2076600.0 ;
      RECT  741600.0 2090400.0 751800.0 2076600.0 ;
      RECT  741600.0 2090400.0 751800.0 2104200.0 ;
      RECT  741600.0 2118000.0 751800.0 2104200.0 ;
      RECT  741600.0 2118000.0 751800.0 2131800.0 ;
      RECT  741600.0 2145600.0 751800.0 2131800.0 ;
      RECT  751800.0 379200.0 762000.0 393000.0 ;
      RECT  751800.0 406800.0 762000.0 393000.0 ;
      RECT  751800.0 406800.0 762000.0 420600.0 ;
      RECT  751800.0 434400.0 762000.0 420600.0 ;
      RECT  751800.0 434400.0 762000.0 448200.0 ;
      RECT  751800.0 462000.0 762000.0 448200.0 ;
      RECT  751800.0 462000.0 762000.0 475800.0 ;
      RECT  751800.0 489600.0 762000.0 475800.0 ;
      RECT  751800.0 489600.0 762000.0 503400.0 ;
      RECT  751800.0 517200.0 762000.0 503400.0 ;
      RECT  751800.0 517200.0 762000.0 531000.0 ;
      RECT  751800.0 544800.0 762000.0 531000.0 ;
      RECT  751800.0 544800.0 762000.0 558600.0 ;
      RECT  751800.0 572400.0 762000.0 558600.0 ;
      RECT  751800.0 572400.0 762000.0 586200.0 ;
      RECT  751800.0 600000.0 762000.0 586200.0 ;
      RECT  751800.0 600000.0 762000.0 613800.0 ;
      RECT  751800.0 627600.0 762000.0 613800.0 ;
      RECT  751800.0 627600.0 762000.0 641400.0 ;
      RECT  751800.0 655200.0 762000.0 641400.0 ;
      RECT  751800.0 655200.0 762000.0 669000.0 ;
      RECT  751800.0 682800.0 762000.0 669000.0 ;
      RECT  751800.0 682800.0 762000.0 696600.0 ;
      RECT  751800.0 710400.0 762000.0 696600.0 ;
      RECT  751800.0 710400.0 762000.0 724200.0 ;
      RECT  751800.0 738000.0 762000.0 724200.0 ;
      RECT  751800.0 738000.0 762000.0 751800.0 ;
      RECT  751800.0 765600.0 762000.0 751800.0 ;
      RECT  751800.0 765600.0 762000.0 779400.0 ;
      RECT  751800.0 793200.0 762000.0 779400.0 ;
      RECT  751800.0 793200.0 762000.0 807000.0 ;
      RECT  751800.0 820800.0 762000.0 807000.0 ;
      RECT  751800.0 820800.0 762000.0 834600.0 ;
      RECT  751800.0 848400.0 762000.0 834600.0 ;
      RECT  751800.0 848400.0 762000.0 862200.0 ;
      RECT  751800.0 876000.0 762000.0 862200.0 ;
      RECT  751800.0 876000.0 762000.0 889800.0 ;
      RECT  751800.0 903600.0 762000.0 889800.0 ;
      RECT  751800.0 903600.0 762000.0 917400.0 ;
      RECT  751800.0 931200.0 762000.0 917400.0 ;
      RECT  751800.0 931200.0 762000.0 945000.0 ;
      RECT  751800.0 958800.0 762000.0 945000.0 ;
      RECT  751800.0 958800.0 762000.0 972600.0 ;
      RECT  751800.0 986400.0 762000.0 972600.0 ;
      RECT  751800.0 986400.0 762000.0 1000200.0 ;
      RECT  751800.0 1014000.0 762000.0 1000200.0 ;
      RECT  751800.0 1014000.0 762000.0 1027800.0 ;
      RECT  751800.0 1041600.0 762000.0 1027800.0 ;
      RECT  751800.0 1041600.0 762000.0 1055400.0 ;
      RECT  751800.0 1069200.0 762000.0 1055400.0 ;
      RECT  751800.0 1069200.0 762000.0 1083000.0 ;
      RECT  751800.0 1096800.0 762000.0 1083000.0 ;
      RECT  751800.0 1096800.0 762000.0 1110600.0 ;
      RECT  751800.0 1124400.0 762000.0 1110600.0 ;
      RECT  751800.0 1124400.0 762000.0 1138200.0 ;
      RECT  751800.0 1152000.0 762000.0 1138200.0 ;
      RECT  751800.0 1152000.0 762000.0 1165800.0 ;
      RECT  751800.0 1179600.0 762000.0 1165800.0 ;
      RECT  751800.0 1179600.0 762000.0 1193400.0 ;
      RECT  751800.0 1207200.0 762000.0 1193400.0 ;
      RECT  751800.0 1207200.0 762000.0 1221000.0 ;
      RECT  751800.0 1234800.0 762000.0 1221000.0 ;
      RECT  751800.0 1234800.0 762000.0 1248600.0 ;
      RECT  751800.0 1262400.0 762000.0 1248600.0 ;
      RECT  751800.0 1262400.0 762000.0 1276200.0 ;
      RECT  751800.0 1290000.0 762000.0 1276200.0 ;
      RECT  751800.0 1290000.0 762000.0 1303800.0 ;
      RECT  751800.0 1317600.0 762000.0 1303800.0 ;
      RECT  751800.0 1317600.0 762000.0 1331400.0 ;
      RECT  751800.0 1345200.0 762000.0 1331400.0 ;
      RECT  751800.0 1345200.0 762000.0 1359000.0 ;
      RECT  751800.0 1372800.0 762000.0 1359000.0 ;
      RECT  751800.0 1372800.0 762000.0 1386600.0 ;
      RECT  751800.0 1400400.0 762000.0 1386600.0 ;
      RECT  751800.0 1400400.0 762000.0 1414200.0 ;
      RECT  751800.0 1428000.0 762000.0 1414200.0 ;
      RECT  751800.0 1428000.0 762000.0 1441800.0 ;
      RECT  751800.0 1455600.0 762000.0 1441800.0 ;
      RECT  751800.0 1455600.0 762000.0 1469400.0 ;
      RECT  751800.0 1483200.0 762000.0 1469400.0 ;
      RECT  751800.0 1483200.0 762000.0 1497000.0 ;
      RECT  751800.0 1510800.0 762000.0 1497000.0 ;
      RECT  751800.0 1510800.0 762000.0 1524600.0 ;
      RECT  751800.0 1538400.0 762000.0 1524600.0 ;
      RECT  751800.0 1538400.0 762000.0 1552200.0 ;
      RECT  751800.0 1566000.0 762000.0 1552200.0 ;
      RECT  751800.0 1566000.0 762000.0 1579800.0 ;
      RECT  751800.0 1593600.0 762000.0 1579800.0 ;
      RECT  751800.0 1593600.0 762000.0 1607400.0 ;
      RECT  751800.0 1621200.0 762000.0 1607400.0 ;
      RECT  751800.0 1621200.0 762000.0 1635000.0 ;
      RECT  751800.0 1648800.0 762000.0 1635000.0 ;
      RECT  751800.0 1648800.0 762000.0 1662600.0 ;
      RECT  751800.0 1676400.0 762000.0 1662600.0 ;
      RECT  751800.0 1676400.0 762000.0 1690200.0 ;
      RECT  751800.0 1704000.0 762000.0 1690200.0 ;
      RECT  751800.0 1704000.0 762000.0 1717800.0 ;
      RECT  751800.0 1731600.0 762000.0 1717800.0 ;
      RECT  751800.0 1731600.0 762000.0 1745400.0 ;
      RECT  751800.0 1759200.0 762000.0 1745400.0 ;
      RECT  751800.0 1759200.0 762000.0 1773000.0 ;
      RECT  751800.0 1786800.0 762000.0 1773000.0 ;
      RECT  751800.0 1786800.0 762000.0 1800600.0 ;
      RECT  751800.0 1814400.0 762000.0 1800600.0 ;
      RECT  751800.0 1814400.0 762000.0 1828200.0 ;
      RECT  751800.0 1842000.0 762000.0 1828200.0 ;
      RECT  751800.0 1842000.0 762000.0 1855800.0 ;
      RECT  751800.0 1869600.0 762000.0 1855800.0 ;
      RECT  751800.0 1869600.0 762000.0 1883400.0 ;
      RECT  751800.0 1897200.0 762000.0 1883400.0 ;
      RECT  751800.0 1897200.0 762000.0 1911000.0 ;
      RECT  751800.0 1924800.0 762000.0 1911000.0 ;
      RECT  751800.0 1924800.0 762000.0 1938600.0 ;
      RECT  751800.0 1952400.0 762000.0 1938600.0 ;
      RECT  751800.0 1952400.0 762000.0 1966200.0 ;
      RECT  751800.0 1980000.0 762000.0 1966200.0 ;
      RECT  751800.0 1980000.0 762000.0 1993800.0 ;
      RECT  751800.0 2007600.0 762000.0 1993800.0 ;
      RECT  751800.0 2007600.0 762000.0 2021400.0 ;
      RECT  751800.0 2035200.0 762000.0 2021400.0 ;
      RECT  751800.0 2035200.0 762000.0 2049000.0 ;
      RECT  751800.0 2062800.0 762000.0 2049000.0 ;
      RECT  751800.0 2062800.0 762000.0 2076600.0 ;
      RECT  751800.0 2090400.0 762000.0 2076600.0 ;
      RECT  751800.0 2090400.0 762000.0 2104200.0 ;
      RECT  751800.0 2118000.0 762000.0 2104200.0 ;
      RECT  751800.0 2118000.0 762000.0 2131800.0 ;
      RECT  751800.0 2145600.0 762000.0 2131800.0 ;
      RECT  762000.0 379200.0 772200.0 393000.0 ;
      RECT  762000.0 406800.0 772200.0 393000.0 ;
      RECT  762000.0 406800.0 772200.0 420600.0 ;
      RECT  762000.0 434400.0 772200.0 420600.0 ;
      RECT  762000.0 434400.0 772200.0 448200.0 ;
      RECT  762000.0 462000.0 772200.0 448200.0 ;
      RECT  762000.0 462000.0 772200.0 475800.0 ;
      RECT  762000.0 489600.0 772200.0 475800.0 ;
      RECT  762000.0 489600.0 772200.0 503400.0 ;
      RECT  762000.0 517200.0 772200.0 503400.0 ;
      RECT  762000.0 517200.0 772200.0 531000.0 ;
      RECT  762000.0 544800.0 772200.0 531000.0 ;
      RECT  762000.0 544800.0 772200.0 558600.0 ;
      RECT  762000.0 572400.0 772200.0 558600.0 ;
      RECT  762000.0 572400.0 772200.0 586200.0 ;
      RECT  762000.0 600000.0 772200.0 586200.0 ;
      RECT  762000.0 600000.0 772200.0 613800.0 ;
      RECT  762000.0 627600.0 772200.0 613800.0 ;
      RECT  762000.0 627600.0 772200.0 641400.0 ;
      RECT  762000.0 655200.0 772200.0 641400.0 ;
      RECT  762000.0 655200.0 772200.0 669000.0 ;
      RECT  762000.0 682800.0 772200.0 669000.0 ;
      RECT  762000.0 682800.0 772200.0 696600.0 ;
      RECT  762000.0 710400.0 772200.0 696600.0 ;
      RECT  762000.0 710400.0 772200.0 724200.0 ;
      RECT  762000.0 738000.0 772200.0 724200.0 ;
      RECT  762000.0 738000.0 772200.0 751800.0 ;
      RECT  762000.0 765600.0 772200.0 751800.0 ;
      RECT  762000.0 765600.0 772200.0 779400.0 ;
      RECT  762000.0 793200.0 772200.0 779400.0 ;
      RECT  762000.0 793200.0 772200.0 807000.0 ;
      RECT  762000.0 820800.0 772200.0 807000.0 ;
      RECT  762000.0 820800.0 772200.0 834600.0 ;
      RECT  762000.0 848400.0 772200.0 834600.0 ;
      RECT  762000.0 848400.0 772200.0 862200.0 ;
      RECT  762000.0 876000.0 772200.0 862200.0 ;
      RECT  762000.0 876000.0 772200.0 889800.0 ;
      RECT  762000.0 903600.0 772200.0 889800.0 ;
      RECT  762000.0 903600.0 772200.0 917400.0 ;
      RECT  762000.0 931200.0 772200.0 917400.0 ;
      RECT  762000.0 931200.0 772200.0 945000.0 ;
      RECT  762000.0 958800.0 772200.0 945000.0 ;
      RECT  762000.0 958800.0 772200.0 972600.0 ;
      RECT  762000.0 986400.0 772200.0 972600.0 ;
      RECT  762000.0 986400.0 772200.0 1000200.0 ;
      RECT  762000.0 1014000.0 772200.0 1000200.0 ;
      RECT  762000.0 1014000.0 772200.0 1027800.0 ;
      RECT  762000.0 1041600.0 772200.0 1027800.0 ;
      RECT  762000.0 1041600.0 772200.0 1055400.0 ;
      RECT  762000.0 1069200.0 772200.0 1055400.0 ;
      RECT  762000.0 1069200.0 772200.0 1083000.0 ;
      RECT  762000.0 1096800.0 772200.0 1083000.0 ;
      RECT  762000.0 1096800.0 772200.0 1110600.0 ;
      RECT  762000.0 1124400.0 772200.0 1110600.0 ;
      RECT  762000.0 1124400.0 772200.0 1138200.0 ;
      RECT  762000.0 1152000.0 772200.0 1138200.0 ;
      RECT  762000.0 1152000.0 772200.0 1165800.0 ;
      RECT  762000.0 1179600.0 772200.0 1165800.0 ;
      RECT  762000.0 1179600.0 772200.0 1193400.0 ;
      RECT  762000.0 1207200.0 772200.0 1193400.0 ;
      RECT  762000.0 1207200.0 772200.0 1221000.0 ;
      RECT  762000.0 1234800.0 772200.0 1221000.0 ;
      RECT  762000.0 1234800.0 772200.0 1248600.0 ;
      RECT  762000.0 1262400.0 772200.0 1248600.0 ;
      RECT  762000.0 1262400.0 772200.0 1276200.0 ;
      RECT  762000.0 1290000.0 772200.0 1276200.0 ;
      RECT  762000.0 1290000.0 772200.0 1303800.0 ;
      RECT  762000.0 1317600.0 772200.0 1303800.0 ;
      RECT  762000.0 1317600.0 772200.0 1331400.0 ;
      RECT  762000.0 1345200.0 772200.0 1331400.0 ;
      RECT  762000.0 1345200.0 772200.0 1359000.0 ;
      RECT  762000.0 1372800.0 772200.0 1359000.0 ;
      RECT  762000.0 1372800.0 772200.0 1386600.0 ;
      RECT  762000.0 1400400.0 772200.0 1386600.0 ;
      RECT  762000.0 1400400.0 772200.0 1414200.0 ;
      RECT  762000.0 1428000.0 772200.0 1414200.0 ;
      RECT  762000.0 1428000.0 772200.0 1441800.0 ;
      RECT  762000.0 1455600.0 772200.0 1441800.0 ;
      RECT  762000.0 1455600.0 772200.0 1469400.0 ;
      RECT  762000.0 1483200.0 772200.0 1469400.0 ;
      RECT  762000.0 1483200.0 772200.0 1497000.0 ;
      RECT  762000.0 1510800.0 772200.0 1497000.0 ;
      RECT  762000.0 1510800.0 772200.0 1524600.0 ;
      RECT  762000.0 1538400.0 772200.0 1524600.0 ;
      RECT  762000.0 1538400.0 772200.0 1552200.0 ;
      RECT  762000.0 1566000.0 772200.0 1552200.0 ;
      RECT  762000.0 1566000.0 772200.0 1579800.0 ;
      RECT  762000.0 1593600.0 772200.0 1579800.0 ;
      RECT  762000.0 1593600.0 772200.0 1607400.0 ;
      RECT  762000.0 1621200.0 772200.0 1607400.0 ;
      RECT  762000.0 1621200.0 772200.0 1635000.0 ;
      RECT  762000.0 1648800.0 772200.0 1635000.0 ;
      RECT  762000.0 1648800.0 772200.0 1662600.0 ;
      RECT  762000.0 1676400.0 772200.0 1662600.0 ;
      RECT  762000.0 1676400.0 772200.0 1690200.0 ;
      RECT  762000.0 1704000.0 772200.0 1690200.0 ;
      RECT  762000.0 1704000.0 772200.0 1717800.0 ;
      RECT  762000.0 1731600.0 772200.0 1717800.0 ;
      RECT  762000.0 1731600.0 772200.0 1745400.0 ;
      RECT  762000.0 1759200.0 772200.0 1745400.0 ;
      RECT  762000.0 1759200.0 772200.0 1773000.0 ;
      RECT  762000.0 1786800.0 772200.0 1773000.0 ;
      RECT  762000.0 1786800.0 772200.0 1800600.0 ;
      RECT  762000.0 1814400.0 772200.0 1800600.0 ;
      RECT  762000.0 1814400.0 772200.0 1828200.0 ;
      RECT  762000.0 1842000.0 772200.0 1828200.0 ;
      RECT  762000.0 1842000.0 772200.0 1855800.0 ;
      RECT  762000.0 1869600.0 772200.0 1855800.0 ;
      RECT  762000.0 1869600.0 772200.0 1883400.0 ;
      RECT  762000.0 1897200.0 772200.0 1883400.0 ;
      RECT  762000.0 1897200.0 772200.0 1911000.0 ;
      RECT  762000.0 1924800.0 772200.0 1911000.0 ;
      RECT  762000.0 1924800.0 772200.0 1938600.0 ;
      RECT  762000.0 1952400.0 772200.0 1938600.0 ;
      RECT  762000.0 1952400.0 772200.0 1966200.0 ;
      RECT  762000.0 1980000.0 772200.0 1966200.0 ;
      RECT  762000.0 1980000.0 772200.0 1993800.0 ;
      RECT  762000.0 2007600.0 772200.0 1993800.0 ;
      RECT  762000.0 2007600.0 772200.0 2021400.0 ;
      RECT  762000.0 2035200.0 772200.0 2021400.0 ;
      RECT  762000.0 2035200.0 772200.0 2049000.0 ;
      RECT  762000.0 2062800.0 772200.0 2049000.0 ;
      RECT  762000.0 2062800.0 772200.0 2076600.0 ;
      RECT  762000.0 2090400.0 772200.0 2076600.0 ;
      RECT  762000.0 2090400.0 772200.0 2104200.0 ;
      RECT  762000.0 2118000.0 772200.0 2104200.0 ;
      RECT  762000.0 2118000.0 772200.0 2131800.0 ;
      RECT  762000.0 2145600.0 772200.0 2131800.0 ;
      RECT  772200.0 379200.0 782400.0 393000.0 ;
      RECT  772200.0 406800.0 782400.0 393000.0 ;
      RECT  772200.0 406800.0 782400.0 420600.0 ;
      RECT  772200.0 434400.0 782400.0 420600.0 ;
      RECT  772200.0 434400.0 782400.0 448200.0 ;
      RECT  772200.0 462000.0 782400.0 448200.0 ;
      RECT  772200.0 462000.0 782400.0 475800.0 ;
      RECT  772200.0 489600.0 782400.0 475800.0 ;
      RECT  772200.0 489600.0 782400.0 503400.0 ;
      RECT  772200.0 517200.0 782400.0 503400.0 ;
      RECT  772200.0 517200.0 782400.0 531000.0 ;
      RECT  772200.0 544800.0 782400.0 531000.0 ;
      RECT  772200.0 544800.0 782400.0 558600.0 ;
      RECT  772200.0 572400.0 782400.0 558600.0 ;
      RECT  772200.0 572400.0 782400.0 586200.0 ;
      RECT  772200.0 600000.0 782400.0 586200.0 ;
      RECT  772200.0 600000.0 782400.0 613800.0 ;
      RECT  772200.0 627600.0 782400.0 613800.0 ;
      RECT  772200.0 627600.0 782400.0 641400.0 ;
      RECT  772200.0 655200.0 782400.0 641400.0 ;
      RECT  772200.0 655200.0 782400.0 669000.0 ;
      RECT  772200.0 682800.0 782400.0 669000.0 ;
      RECT  772200.0 682800.0 782400.0 696600.0 ;
      RECT  772200.0 710400.0 782400.0 696600.0 ;
      RECT  772200.0 710400.0 782400.0 724200.0 ;
      RECT  772200.0 738000.0 782400.0 724200.0 ;
      RECT  772200.0 738000.0 782400.0 751800.0 ;
      RECT  772200.0 765600.0 782400.0 751800.0 ;
      RECT  772200.0 765600.0 782400.0 779400.0 ;
      RECT  772200.0 793200.0 782400.0 779400.0 ;
      RECT  772200.0 793200.0 782400.0 807000.0 ;
      RECT  772200.0 820800.0 782400.0 807000.0 ;
      RECT  772200.0 820800.0 782400.0 834600.0 ;
      RECT  772200.0 848400.0 782400.0 834600.0 ;
      RECT  772200.0 848400.0 782400.0 862200.0 ;
      RECT  772200.0 876000.0 782400.0 862200.0 ;
      RECT  772200.0 876000.0 782400.0 889800.0 ;
      RECT  772200.0 903600.0 782400.0 889800.0 ;
      RECT  772200.0 903600.0 782400.0 917400.0 ;
      RECT  772200.0 931200.0 782400.0 917400.0 ;
      RECT  772200.0 931200.0 782400.0 945000.0 ;
      RECT  772200.0 958800.0 782400.0 945000.0 ;
      RECT  772200.0 958800.0 782400.0 972600.0 ;
      RECT  772200.0 986400.0 782400.0 972600.0 ;
      RECT  772200.0 986400.0 782400.0 1000200.0 ;
      RECT  772200.0 1014000.0 782400.0 1000200.0 ;
      RECT  772200.0 1014000.0 782400.0 1027800.0 ;
      RECT  772200.0 1041600.0 782400.0 1027800.0 ;
      RECT  772200.0 1041600.0 782400.0 1055400.0 ;
      RECT  772200.0 1069200.0 782400.0 1055400.0 ;
      RECT  772200.0 1069200.0 782400.0 1083000.0 ;
      RECT  772200.0 1096800.0 782400.0 1083000.0 ;
      RECT  772200.0 1096800.0 782400.0 1110600.0 ;
      RECT  772200.0 1124400.0 782400.0 1110600.0 ;
      RECT  772200.0 1124400.0 782400.0 1138200.0 ;
      RECT  772200.0 1152000.0 782400.0 1138200.0 ;
      RECT  772200.0 1152000.0 782400.0 1165800.0 ;
      RECT  772200.0 1179600.0 782400.0 1165800.0 ;
      RECT  772200.0 1179600.0 782400.0 1193400.0 ;
      RECT  772200.0 1207200.0 782400.0 1193400.0 ;
      RECT  772200.0 1207200.0 782400.0 1221000.0 ;
      RECT  772200.0 1234800.0 782400.0 1221000.0 ;
      RECT  772200.0 1234800.0 782400.0 1248600.0 ;
      RECT  772200.0 1262400.0 782400.0 1248600.0 ;
      RECT  772200.0 1262400.0 782400.0 1276200.0 ;
      RECT  772200.0 1290000.0 782400.0 1276200.0 ;
      RECT  772200.0 1290000.0 782400.0 1303800.0 ;
      RECT  772200.0 1317600.0 782400.0 1303800.0 ;
      RECT  772200.0 1317600.0 782400.0 1331400.0 ;
      RECT  772200.0 1345200.0 782400.0 1331400.0 ;
      RECT  772200.0 1345200.0 782400.0 1359000.0 ;
      RECT  772200.0 1372800.0 782400.0 1359000.0 ;
      RECT  772200.0 1372800.0 782400.0 1386600.0 ;
      RECT  772200.0 1400400.0 782400.0 1386600.0 ;
      RECT  772200.0 1400400.0 782400.0 1414200.0 ;
      RECT  772200.0 1428000.0 782400.0 1414200.0 ;
      RECT  772200.0 1428000.0 782400.0 1441800.0 ;
      RECT  772200.0 1455600.0 782400.0 1441800.0 ;
      RECT  772200.0 1455600.0 782400.0 1469400.0 ;
      RECT  772200.0 1483200.0 782400.0 1469400.0 ;
      RECT  772200.0 1483200.0 782400.0 1497000.0 ;
      RECT  772200.0 1510800.0 782400.0 1497000.0 ;
      RECT  772200.0 1510800.0 782400.0 1524600.0 ;
      RECT  772200.0 1538400.0 782400.0 1524600.0 ;
      RECT  772200.0 1538400.0 782400.0 1552200.0 ;
      RECT  772200.0 1566000.0 782400.0 1552200.0 ;
      RECT  772200.0 1566000.0 782400.0 1579800.0 ;
      RECT  772200.0 1593600.0 782400.0 1579800.0 ;
      RECT  772200.0 1593600.0 782400.0 1607400.0 ;
      RECT  772200.0 1621200.0 782400.0 1607400.0 ;
      RECT  772200.0 1621200.0 782400.0 1635000.0 ;
      RECT  772200.0 1648800.0 782400.0 1635000.0 ;
      RECT  772200.0 1648800.0 782400.0 1662600.0 ;
      RECT  772200.0 1676400.0 782400.0 1662600.0 ;
      RECT  772200.0 1676400.0 782400.0 1690200.0 ;
      RECT  772200.0 1704000.0 782400.0 1690200.0 ;
      RECT  772200.0 1704000.0 782400.0 1717800.0 ;
      RECT  772200.0 1731600.0 782400.0 1717800.0 ;
      RECT  772200.0 1731600.0 782400.0 1745400.0 ;
      RECT  772200.0 1759200.0 782400.0 1745400.0 ;
      RECT  772200.0 1759200.0 782400.0 1773000.0 ;
      RECT  772200.0 1786800.0 782400.0 1773000.0 ;
      RECT  772200.0 1786800.0 782400.0 1800600.0 ;
      RECT  772200.0 1814400.0 782400.0 1800600.0 ;
      RECT  772200.0 1814400.0 782400.0 1828200.0 ;
      RECT  772200.0 1842000.0 782400.0 1828200.0 ;
      RECT  772200.0 1842000.0 782400.0 1855800.0 ;
      RECT  772200.0 1869600.0 782400.0 1855800.0 ;
      RECT  772200.0 1869600.0 782400.0 1883400.0 ;
      RECT  772200.0 1897200.0 782400.0 1883400.0 ;
      RECT  772200.0 1897200.0 782400.0 1911000.0 ;
      RECT  772200.0 1924800.0 782400.0 1911000.0 ;
      RECT  772200.0 1924800.0 782400.0 1938600.0 ;
      RECT  772200.0 1952400.0 782400.0 1938600.0 ;
      RECT  772200.0 1952400.0 782400.0 1966200.0 ;
      RECT  772200.0 1980000.0 782400.0 1966200.0 ;
      RECT  772200.0 1980000.0 782400.0 1993800.0 ;
      RECT  772200.0 2007600.0 782400.0 1993800.0 ;
      RECT  772200.0 2007600.0 782400.0 2021400.0 ;
      RECT  772200.0 2035200.0 782400.0 2021400.0 ;
      RECT  772200.0 2035200.0 782400.0 2049000.0 ;
      RECT  772200.0 2062800.0 782400.0 2049000.0 ;
      RECT  772200.0 2062800.0 782400.0 2076600.0 ;
      RECT  772200.0 2090400.0 782400.0 2076600.0 ;
      RECT  772200.0 2090400.0 782400.0 2104200.0 ;
      RECT  772200.0 2118000.0 782400.0 2104200.0 ;
      RECT  772200.0 2118000.0 782400.0 2131800.0 ;
      RECT  772200.0 2145600.0 782400.0 2131800.0 ;
      RECT  782400.0 379200.0 792600.0 393000.0 ;
      RECT  782400.0 406800.0 792600.0 393000.0 ;
      RECT  782400.0 406800.0 792600.0 420600.0 ;
      RECT  782400.0 434400.0 792600.0 420600.0 ;
      RECT  782400.0 434400.0 792600.0 448200.0 ;
      RECT  782400.0 462000.0 792600.0 448200.0 ;
      RECT  782400.0 462000.0 792600.0 475800.0 ;
      RECT  782400.0 489600.0 792600.0 475800.0 ;
      RECT  782400.0 489600.0 792600.0 503400.0 ;
      RECT  782400.0 517200.0 792600.0 503400.0 ;
      RECT  782400.0 517200.0 792600.0 531000.0 ;
      RECT  782400.0 544800.0 792600.0 531000.0 ;
      RECT  782400.0 544800.0 792600.0 558600.0 ;
      RECT  782400.0 572400.0 792600.0 558600.0 ;
      RECT  782400.0 572400.0 792600.0 586200.0 ;
      RECT  782400.0 600000.0 792600.0 586200.0 ;
      RECT  782400.0 600000.0 792600.0 613800.0 ;
      RECT  782400.0 627600.0 792600.0 613800.0 ;
      RECT  782400.0 627600.0 792600.0 641400.0 ;
      RECT  782400.0 655200.0 792600.0 641400.0 ;
      RECT  782400.0 655200.0 792600.0 669000.0 ;
      RECT  782400.0 682800.0 792600.0 669000.0 ;
      RECT  782400.0 682800.0 792600.0 696600.0 ;
      RECT  782400.0 710400.0 792600.0 696600.0 ;
      RECT  782400.0 710400.0 792600.0 724200.0 ;
      RECT  782400.0 738000.0 792600.0 724200.0 ;
      RECT  782400.0 738000.0 792600.0 751800.0 ;
      RECT  782400.0 765600.0 792600.0 751800.0 ;
      RECT  782400.0 765600.0 792600.0 779400.0 ;
      RECT  782400.0 793200.0 792600.0 779400.0 ;
      RECT  782400.0 793200.0 792600.0 807000.0 ;
      RECT  782400.0 820800.0 792600.0 807000.0 ;
      RECT  782400.0 820800.0 792600.0 834600.0 ;
      RECT  782400.0 848400.0 792600.0 834600.0 ;
      RECT  782400.0 848400.0 792600.0 862200.0 ;
      RECT  782400.0 876000.0 792600.0 862200.0 ;
      RECT  782400.0 876000.0 792600.0 889800.0 ;
      RECT  782400.0 903600.0 792600.0 889800.0 ;
      RECT  782400.0 903600.0 792600.0 917400.0 ;
      RECT  782400.0 931200.0 792600.0 917400.0 ;
      RECT  782400.0 931200.0 792600.0 945000.0 ;
      RECT  782400.0 958800.0 792600.0 945000.0 ;
      RECT  782400.0 958800.0 792600.0 972600.0 ;
      RECT  782400.0 986400.0 792600.0 972600.0 ;
      RECT  782400.0 986400.0 792600.0 1000200.0 ;
      RECT  782400.0 1014000.0 792600.0 1000200.0 ;
      RECT  782400.0 1014000.0 792600.0 1027800.0 ;
      RECT  782400.0 1041600.0 792600.0 1027800.0 ;
      RECT  782400.0 1041600.0 792600.0 1055400.0 ;
      RECT  782400.0 1069200.0 792600.0 1055400.0 ;
      RECT  782400.0 1069200.0 792600.0 1083000.0 ;
      RECT  782400.0 1096800.0 792600.0 1083000.0 ;
      RECT  782400.0 1096800.0 792600.0 1110600.0 ;
      RECT  782400.0 1124400.0 792600.0 1110600.0 ;
      RECT  782400.0 1124400.0 792600.0 1138200.0 ;
      RECT  782400.0 1152000.0 792600.0 1138200.0 ;
      RECT  782400.0 1152000.0 792600.0 1165800.0 ;
      RECT  782400.0 1179600.0 792600.0 1165800.0 ;
      RECT  782400.0 1179600.0 792600.0 1193400.0 ;
      RECT  782400.0 1207200.0 792600.0 1193400.0 ;
      RECT  782400.0 1207200.0 792600.0 1221000.0 ;
      RECT  782400.0 1234800.0 792600.0 1221000.0 ;
      RECT  782400.0 1234800.0 792600.0 1248600.0 ;
      RECT  782400.0 1262400.0 792600.0 1248600.0 ;
      RECT  782400.0 1262400.0 792600.0 1276200.0 ;
      RECT  782400.0 1290000.0 792600.0 1276200.0 ;
      RECT  782400.0 1290000.0 792600.0 1303800.0 ;
      RECT  782400.0 1317600.0 792600.0 1303800.0 ;
      RECT  782400.0 1317600.0 792600.0 1331400.0 ;
      RECT  782400.0 1345200.0 792600.0 1331400.0 ;
      RECT  782400.0 1345200.0 792600.0 1359000.0 ;
      RECT  782400.0 1372800.0 792600.0 1359000.0 ;
      RECT  782400.0 1372800.0 792600.0 1386600.0 ;
      RECT  782400.0 1400400.0 792600.0 1386600.0 ;
      RECT  782400.0 1400400.0 792600.0 1414200.0 ;
      RECT  782400.0 1428000.0 792600.0 1414200.0 ;
      RECT  782400.0 1428000.0 792600.0 1441800.0 ;
      RECT  782400.0 1455600.0 792600.0 1441800.0 ;
      RECT  782400.0 1455600.0 792600.0 1469400.0 ;
      RECT  782400.0 1483200.0 792600.0 1469400.0 ;
      RECT  782400.0 1483200.0 792600.0 1497000.0 ;
      RECT  782400.0 1510800.0 792600.0 1497000.0 ;
      RECT  782400.0 1510800.0 792600.0 1524600.0 ;
      RECT  782400.0 1538400.0 792600.0 1524600.0 ;
      RECT  782400.0 1538400.0 792600.0 1552200.0 ;
      RECT  782400.0 1566000.0 792600.0 1552200.0 ;
      RECT  782400.0 1566000.0 792600.0 1579800.0 ;
      RECT  782400.0 1593600.0 792600.0 1579800.0 ;
      RECT  782400.0 1593600.0 792600.0 1607400.0 ;
      RECT  782400.0 1621200.0 792600.0 1607400.0 ;
      RECT  782400.0 1621200.0 792600.0 1635000.0 ;
      RECT  782400.0 1648800.0 792600.0 1635000.0 ;
      RECT  782400.0 1648800.0 792600.0 1662600.0 ;
      RECT  782400.0 1676400.0 792600.0 1662600.0 ;
      RECT  782400.0 1676400.0 792600.0 1690200.0 ;
      RECT  782400.0 1704000.0 792600.0 1690200.0 ;
      RECT  782400.0 1704000.0 792600.0 1717800.0 ;
      RECT  782400.0 1731600.0 792600.0 1717800.0 ;
      RECT  782400.0 1731600.0 792600.0 1745400.0 ;
      RECT  782400.0 1759200.0 792600.0 1745400.0 ;
      RECT  782400.0 1759200.0 792600.0 1773000.0 ;
      RECT  782400.0 1786800.0 792600.0 1773000.0 ;
      RECT  782400.0 1786800.0 792600.0 1800600.0 ;
      RECT  782400.0 1814400.0 792600.0 1800600.0 ;
      RECT  782400.0 1814400.0 792600.0 1828200.0 ;
      RECT  782400.0 1842000.0 792600.0 1828200.0 ;
      RECT  782400.0 1842000.0 792600.0 1855800.0 ;
      RECT  782400.0 1869600.0 792600.0 1855800.0 ;
      RECT  782400.0 1869600.0 792600.0 1883400.0 ;
      RECT  782400.0 1897200.0 792600.0 1883400.0 ;
      RECT  782400.0 1897200.0 792600.0 1911000.0 ;
      RECT  782400.0 1924800.0 792600.0 1911000.0 ;
      RECT  782400.0 1924800.0 792600.0 1938600.0 ;
      RECT  782400.0 1952400.0 792600.0 1938600.0 ;
      RECT  782400.0 1952400.0 792600.0 1966200.0 ;
      RECT  782400.0 1980000.0 792600.0 1966200.0 ;
      RECT  782400.0 1980000.0 792600.0 1993800.0 ;
      RECT  782400.0 2007600.0 792600.0 1993800.0 ;
      RECT  782400.0 2007600.0 792600.0 2021400.0 ;
      RECT  782400.0 2035200.0 792600.0 2021400.0 ;
      RECT  782400.0 2035200.0 792600.0 2049000.0 ;
      RECT  782400.0 2062800.0 792600.0 2049000.0 ;
      RECT  782400.0 2062800.0 792600.0 2076600.0 ;
      RECT  782400.0 2090400.0 792600.0 2076600.0 ;
      RECT  782400.0 2090400.0 792600.0 2104200.0 ;
      RECT  782400.0 2118000.0 792600.0 2104200.0 ;
      RECT  782400.0 2118000.0 792600.0 2131800.0 ;
      RECT  782400.0 2145600.0 792600.0 2131800.0 ;
      RECT  792600.0 379200.0 802800.0 393000.0 ;
      RECT  792600.0 406800.0 802800.0 393000.0 ;
      RECT  792600.0 406800.0 802800.0 420600.0 ;
      RECT  792600.0 434400.0 802800.0 420600.0 ;
      RECT  792600.0 434400.0 802800.0 448200.0 ;
      RECT  792600.0 462000.0 802800.0 448200.0 ;
      RECT  792600.0 462000.0 802800.0 475800.0 ;
      RECT  792600.0 489600.0 802800.0 475800.0 ;
      RECT  792600.0 489600.0 802800.0 503400.0 ;
      RECT  792600.0 517200.0 802800.0 503400.0 ;
      RECT  792600.0 517200.0 802800.0 531000.0 ;
      RECT  792600.0 544800.0 802800.0 531000.0 ;
      RECT  792600.0 544800.0 802800.0 558600.0 ;
      RECT  792600.0 572400.0 802800.0 558600.0 ;
      RECT  792600.0 572400.0 802800.0 586200.0 ;
      RECT  792600.0 600000.0 802800.0 586200.0 ;
      RECT  792600.0 600000.0 802800.0 613800.0 ;
      RECT  792600.0 627600.0 802800.0 613800.0 ;
      RECT  792600.0 627600.0 802800.0 641400.0 ;
      RECT  792600.0 655200.0 802800.0 641400.0 ;
      RECT  792600.0 655200.0 802800.0 669000.0 ;
      RECT  792600.0 682800.0 802800.0 669000.0 ;
      RECT  792600.0 682800.0 802800.0 696600.0 ;
      RECT  792600.0 710400.0 802800.0 696600.0 ;
      RECT  792600.0 710400.0 802800.0 724200.0 ;
      RECT  792600.0 738000.0 802800.0 724200.0 ;
      RECT  792600.0 738000.0 802800.0 751800.0 ;
      RECT  792600.0 765600.0 802800.0 751800.0 ;
      RECT  792600.0 765600.0 802800.0 779400.0 ;
      RECT  792600.0 793200.0 802800.0 779400.0 ;
      RECT  792600.0 793200.0 802800.0 807000.0 ;
      RECT  792600.0 820800.0 802800.0 807000.0 ;
      RECT  792600.0 820800.0 802800.0 834600.0 ;
      RECT  792600.0 848400.0 802800.0 834600.0 ;
      RECT  792600.0 848400.0 802800.0 862200.0 ;
      RECT  792600.0 876000.0 802800.0 862200.0 ;
      RECT  792600.0 876000.0 802800.0 889800.0 ;
      RECT  792600.0 903600.0 802800.0 889800.0 ;
      RECT  792600.0 903600.0 802800.0 917400.0 ;
      RECT  792600.0 931200.0 802800.0 917400.0 ;
      RECT  792600.0 931200.0 802800.0 945000.0 ;
      RECT  792600.0 958800.0 802800.0 945000.0 ;
      RECT  792600.0 958800.0 802800.0 972600.0 ;
      RECT  792600.0 986400.0 802800.0 972600.0 ;
      RECT  792600.0 986400.0 802800.0 1000200.0 ;
      RECT  792600.0 1014000.0 802800.0 1000200.0 ;
      RECT  792600.0 1014000.0 802800.0 1027800.0 ;
      RECT  792600.0 1041600.0 802800.0 1027800.0 ;
      RECT  792600.0 1041600.0 802800.0 1055400.0 ;
      RECT  792600.0 1069200.0 802800.0 1055400.0 ;
      RECT  792600.0 1069200.0 802800.0 1083000.0 ;
      RECT  792600.0 1096800.0 802800.0 1083000.0 ;
      RECT  792600.0 1096800.0 802800.0 1110600.0 ;
      RECT  792600.0 1124400.0 802800.0 1110600.0 ;
      RECT  792600.0 1124400.0 802800.0 1138200.0 ;
      RECT  792600.0 1152000.0 802800.0 1138200.0 ;
      RECT  792600.0 1152000.0 802800.0 1165800.0 ;
      RECT  792600.0 1179600.0 802800.0 1165800.0 ;
      RECT  792600.0 1179600.0 802800.0 1193400.0 ;
      RECT  792600.0 1207200.0 802800.0 1193400.0 ;
      RECT  792600.0 1207200.0 802800.0 1221000.0 ;
      RECT  792600.0 1234800.0 802800.0 1221000.0 ;
      RECT  792600.0 1234800.0 802800.0 1248600.0 ;
      RECT  792600.0 1262400.0 802800.0 1248600.0 ;
      RECT  792600.0 1262400.0 802800.0 1276200.0 ;
      RECT  792600.0 1290000.0 802800.0 1276200.0 ;
      RECT  792600.0 1290000.0 802800.0 1303800.0 ;
      RECT  792600.0 1317600.0 802800.0 1303800.0 ;
      RECT  792600.0 1317600.0 802800.0 1331400.0 ;
      RECT  792600.0 1345200.0 802800.0 1331400.0 ;
      RECT  792600.0 1345200.0 802800.0 1359000.0 ;
      RECT  792600.0 1372800.0 802800.0 1359000.0 ;
      RECT  792600.0 1372800.0 802800.0 1386600.0 ;
      RECT  792600.0 1400400.0 802800.0 1386600.0 ;
      RECT  792600.0 1400400.0 802800.0 1414200.0 ;
      RECT  792600.0 1428000.0 802800.0 1414200.0 ;
      RECT  792600.0 1428000.0 802800.0 1441800.0 ;
      RECT  792600.0 1455600.0 802800.0 1441800.0 ;
      RECT  792600.0 1455600.0 802800.0 1469400.0 ;
      RECT  792600.0 1483200.0 802800.0 1469400.0 ;
      RECT  792600.0 1483200.0 802800.0 1497000.0 ;
      RECT  792600.0 1510800.0 802800.0 1497000.0 ;
      RECT  792600.0 1510800.0 802800.0 1524600.0 ;
      RECT  792600.0 1538400.0 802800.0 1524600.0 ;
      RECT  792600.0 1538400.0 802800.0 1552200.0 ;
      RECT  792600.0 1566000.0 802800.0 1552200.0 ;
      RECT  792600.0 1566000.0 802800.0 1579800.0 ;
      RECT  792600.0 1593600.0 802800.0 1579800.0 ;
      RECT  792600.0 1593600.0 802800.0 1607400.0 ;
      RECT  792600.0 1621200.0 802800.0 1607400.0 ;
      RECT  792600.0 1621200.0 802800.0 1635000.0 ;
      RECT  792600.0 1648800.0 802800.0 1635000.0 ;
      RECT  792600.0 1648800.0 802800.0 1662600.0 ;
      RECT  792600.0 1676400.0 802800.0 1662600.0 ;
      RECT  792600.0 1676400.0 802800.0 1690200.0 ;
      RECT  792600.0 1704000.0 802800.0 1690200.0 ;
      RECT  792600.0 1704000.0 802800.0 1717800.0 ;
      RECT  792600.0 1731600.0 802800.0 1717800.0 ;
      RECT  792600.0 1731600.0 802800.0 1745400.0 ;
      RECT  792600.0 1759200.0 802800.0 1745400.0 ;
      RECT  792600.0 1759200.0 802800.0 1773000.0 ;
      RECT  792600.0 1786800.0 802800.0 1773000.0 ;
      RECT  792600.0 1786800.0 802800.0 1800600.0 ;
      RECT  792600.0 1814400.0 802800.0 1800600.0 ;
      RECT  792600.0 1814400.0 802800.0 1828200.0 ;
      RECT  792600.0 1842000.0 802800.0 1828200.0 ;
      RECT  792600.0 1842000.0 802800.0 1855800.0 ;
      RECT  792600.0 1869600.0 802800.0 1855800.0 ;
      RECT  792600.0 1869600.0 802800.0 1883400.0 ;
      RECT  792600.0 1897200.0 802800.0 1883400.0 ;
      RECT  792600.0 1897200.0 802800.0 1911000.0 ;
      RECT  792600.0 1924800.0 802800.0 1911000.0 ;
      RECT  792600.0 1924800.0 802800.0 1938600.0 ;
      RECT  792600.0 1952400.0 802800.0 1938600.0 ;
      RECT  792600.0 1952400.0 802800.0 1966200.0 ;
      RECT  792600.0 1980000.0 802800.0 1966200.0 ;
      RECT  792600.0 1980000.0 802800.0 1993800.0 ;
      RECT  792600.0 2007600.0 802800.0 1993800.0 ;
      RECT  792600.0 2007600.0 802800.0 2021400.0 ;
      RECT  792600.0 2035200.0 802800.0 2021400.0 ;
      RECT  792600.0 2035200.0 802800.0 2049000.0 ;
      RECT  792600.0 2062800.0 802800.0 2049000.0 ;
      RECT  792600.0 2062800.0 802800.0 2076600.0 ;
      RECT  792600.0 2090400.0 802800.0 2076600.0 ;
      RECT  792600.0 2090400.0 802800.0 2104200.0 ;
      RECT  792600.0 2118000.0 802800.0 2104200.0 ;
      RECT  792600.0 2118000.0 802800.0 2131800.0 ;
      RECT  792600.0 2145600.0 802800.0 2131800.0 ;
      RECT  802800.0 379200.0 813000.0 393000.0 ;
      RECT  802800.0 406800.0 813000.0 393000.0 ;
      RECT  802800.0 406800.0 813000.0 420600.0 ;
      RECT  802800.0 434400.0 813000.0 420600.0 ;
      RECT  802800.0 434400.0 813000.0 448200.0 ;
      RECT  802800.0 462000.0 813000.0 448200.0 ;
      RECT  802800.0 462000.0 813000.0 475800.0 ;
      RECT  802800.0 489600.0 813000.0 475800.0 ;
      RECT  802800.0 489600.0 813000.0 503400.0 ;
      RECT  802800.0 517200.0 813000.0 503400.0 ;
      RECT  802800.0 517200.0 813000.0 531000.0 ;
      RECT  802800.0 544800.0 813000.0 531000.0 ;
      RECT  802800.0 544800.0 813000.0 558600.0 ;
      RECT  802800.0 572400.0 813000.0 558600.0 ;
      RECT  802800.0 572400.0 813000.0 586200.0 ;
      RECT  802800.0 600000.0 813000.0 586200.0 ;
      RECT  802800.0 600000.0 813000.0 613800.0 ;
      RECT  802800.0 627600.0 813000.0 613800.0 ;
      RECT  802800.0 627600.0 813000.0 641400.0 ;
      RECT  802800.0 655200.0 813000.0 641400.0 ;
      RECT  802800.0 655200.0 813000.0 669000.0 ;
      RECT  802800.0 682800.0 813000.0 669000.0 ;
      RECT  802800.0 682800.0 813000.0 696600.0 ;
      RECT  802800.0 710400.0 813000.0 696600.0 ;
      RECT  802800.0 710400.0 813000.0 724200.0 ;
      RECT  802800.0 738000.0 813000.0 724200.0 ;
      RECT  802800.0 738000.0 813000.0 751800.0 ;
      RECT  802800.0 765600.0 813000.0 751800.0 ;
      RECT  802800.0 765600.0 813000.0 779400.0 ;
      RECT  802800.0 793200.0 813000.0 779400.0 ;
      RECT  802800.0 793200.0 813000.0 807000.0 ;
      RECT  802800.0 820800.0 813000.0 807000.0 ;
      RECT  802800.0 820800.0 813000.0 834600.0 ;
      RECT  802800.0 848400.0 813000.0 834600.0 ;
      RECT  802800.0 848400.0 813000.0 862200.0 ;
      RECT  802800.0 876000.0 813000.0 862200.0 ;
      RECT  802800.0 876000.0 813000.0 889800.0 ;
      RECT  802800.0 903600.0 813000.0 889800.0 ;
      RECT  802800.0 903600.0 813000.0 917400.0 ;
      RECT  802800.0 931200.0 813000.0 917400.0 ;
      RECT  802800.0 931200.0 813000.0 945000.0 ;
      RECT  802800.0 958800.0 813000.0 945000.0 ;
      RECT  802800.0 958800.0 813000.0 972600.0 ;
      RECT  802800.0 986400.0 813000.0 972600.0 ;
      RECT  802800.0 986400.0 813000.0 1000200.0 ;
      RECT  802800.0 1014000.0 813000.0 1000200.0 ;
      RECT  802800.0 1014000.0 813000.0 1027800.0 ;
      RECT  802800.0 1041600.0 813000.0 1027800.0 ;
      RECT  802800.0 1041600.0 813000.0 1055400.0 ;
      RECT  802800.0 1069200.0 813000.0 1055400.0 ;
      RECT  802800.0 1069200.0 813000.0 1083000.0 ;
      RECT  802800.0 1096800.0 813000.0 1083000.0 ;
      RECT  802800.0 1096800.0 813000.0 1110600.0 ;
      RECT  802800.0 1124400.0 813000.0 1110600.0 ;
      RECT  802800.0 1124400.0 813000.0 1138200.0 ;
      RECT  802800.0 1152000.0 813000.0 1138200.0 ;
      RECT  802800.0 1152000.0 813000.0 1165800.0 ;
      RECT  802800.0 1179600.0 813000.0 1165800.0 ;
      RECT  802800.0 1179600.0 813000.0 1193400.0 ;
      RECT  802800.0 1207200.0 813000.0 1193400.0 ;
      RECT  802800.0 1207200.0 813000.0 1221000.0 ;
      RECT  802800.0 1234800.0 813000.0 1221000.0 ;
      RECT  802800.0 1234800.0 813000.0 1248600.0 ;
      RECT  802800.0 1262400.0 813000.0 1248600.0 ;
      RECT  802800.0 1262400.0 813000.0 1276200.0 ;
      RECT  802800.0 1290000.0 813000.0 1276200.0 ;
      RECT  802800.0 1290000.0 813000.0 1303800.0 ;
      RECT  802800.0 1317600.0 813000.0 1303800.0 ;
      RECT  802800.0 1317600.0 813000.0 1331400.0 ;
      RECT  802800.0 1345200.0 813000.0 1331400.0 ;
      RECT  802800.0 1345200.0 813000.0 1359000.0 ;
      RECT  802800.0 1372800.0 813000.0 1359000.0 ;
      RECT  802800.0 1372800.0 813000.0 1386600.0 ;
      RECT  802800.0 1400400.0 813000.0 1386600.0 ;
      RECT  802800.0 1400400.0 813000.0 1414200.0 ;
      RECT  802800.0 1428000.0 813000.0 1414200.0 ;
      RECT  802800.0 1428000.0 813000.0 1441800.0 ;
      RECT  802800.0 1455600.0 813000.0 1441800.0 ;
      RECT  802800.0 1455600.0 813000.0 1469400.0 ;
      RECT  802800.0 1483200.0 813000.0 1469400.0 ;
      RECT  802800.0 1483200.0 813000.0 1497000.0 ;
      RECT  802800.0 1510800.0 813000.0 1497000.0 ;
      RECT  802800.0 1510800.0 813000.0 1524600.0 ;
      RECT  802800.0 1538400.0 813000.0 1524600.0 ;
      RECT  802800.0 1538400.0 813000.0 1552200.0 ;
      RECT  802800.0 1566000.0 813000.0 1552200.0 ;
      RECT  802800.0 1566000.0 813000.0 1579800.0 ;
      RECT  802800.0 1593600.0 813000.0 1579800.0 ;
      RECT  802800.0 1593600.0 813000.0 1607400.0 ;
      RECT  802800.0 1621200.0 813000.0 1607400.0 ;
      RECT  802800.0 1621200.0 813000.0 1635000.0 ;
      RECT  802800.0 1648800.0 813000.0 1635000.0 ;
      RECT  802800.0 1648800.0 813000.0 1662600.0 ;
      RECT  802800.0 1676400.0 813000.0 1662600.0 ;
      RECT  802800.0 1676400.0 813000.0 1690200.0 ;
      RECT  802800.0 1704000.0 813000.0 1690200.0 ;
      RECT  802800.0 1704000.0 813000.0 1717800.0 ;
      RECT  802800.0 1731600.0 813000.0 1717800.0 ;
      RECT  802800.0 1731600.0 813000.0 1745400.0 ;
      RECT  802800.0 1759200.0 813000.0 1745400.0 ;
      RECT  802800.0 1759200.0 813000.0 1773000.0 ;
      RECT  802800.0 1786800.0 813000.0 1773000.0 ;
      RECT  802800.0 1786800.0 813000.0 1800600.0 ;
      RECT  802800.0 1814400.0 813000.0 1800600.0 ;
      RECT  802800.0 1814400.0 813000.0 1828200.0 ;
      RECT  802800.0 1842000.0 813000.0 1828200.0 ;
      RECT  802800.0 1842000.0 813000.0 1855800.0 ;
      RECT  802800.0 1869600.0 813000.0 1855800.0 ;
      RECT  802800.0 1869600.0 813000.0 1883400.0 ;
      RECT  802800.0 1897200.0 813000.0 1883400.0 ;
      RECT  802800.0 1897200.0 813000.0 1911000.0 ;
      RECT  802800.0 1924800.0 813000.0 1911000.0 ;
      RECT  802800.0 1924800.0 813000.0 1938600.0 ;
      RECT  802800.0 1952400.0 813000.0 1938600.0 ;
      RECT  802800.0 1952400.0 813000.0 1966200.0 ;
      RECT  802800.0 1980000.0 813000.0 1966200.0 ;
      RECT  802800.0 1980000.0 813000.0 1993800.0 ;
      RECT  802800.0 2007600.0 813000.0 1993800.0 ;
      RECT  802800.0 2007600.0 813000.0 2021400.0 ;
      RECT  802800.0 2035200.0 813000.0 2021400.0 ;
      RECT  802800.0 2035200.0 813000.0 2049000.0 ;
      RECT  802800.0 2062800.0 813000.0 2049000.0 ;
      RECT  802800.0 2062800.0 813000.0 2076600.0 ;
      RECT  802800.0 2090400.0 813000.0 2076600.0 ;
      RECT  802800.0 2090400.0 813000.0 2104200.0 ;
      RECT  802800.0 2118000.0 813000.0 2104200.0 ;
      RECT  802800.0 2118000.0 813000.0 2131800.0 ;
      RECT  802800.0 2145600.0 813000.0 2131800.0 ;
      RECT  813000.0 379200.0 823200.0 393000.0 ;
      RECT  813000.0 406800.0 823200.0 393000.0 ;
      RECT  813000.0 406800.0 823200.0 420600.0 ;
      RECT  813000.0 434400.0 823200.0 420600.0 ;
      RECT  813000.0 434400.0 823200.0 448200.0 ;
      RECT  813000.0 462000.0 823200.0 448200.0 ;
      RECT  813000.0 462000.0 823200.0 475800.0 ;
      RECT  813000.0 489600.0 823200.0 475800.0 ;
      RECT  813000.0 489600.0 823200.0 503400.0 ;
      RECT  813000.0 517200.0 823200.0 503400.0 ;
      RECT  813000.0 517200.0 823200.0 531000.0 ;
      RECT  813000.0 544800.0 823200.0 531000.0 ;
      RECT  813000.0 544800.0 823200.0 558600.0 ;
      RECT  813000.0 572400.0 823200.0 558600.0 ;
      RECT  813000.0 572400.0 823200.0 586200.0 ;
      RECT  813000.0 600000.0 823200.0 586200.0 ;
      RECT  813000.0 600000.0 823200.0 613800.0 ;
      RECT  813000.0 627600.0 823200.0 613800.0 ;
      RECT  813000.0 627600.0 823200.0 641400.0 ;
      RECT  813000.0 655200.0 823200.0 641400.0 ;
      RECT  813000.0 655200.0 823200.0 669000.0 ;
      RECT  813000.0 682800.0 823200.0 669000.0 ;
      RECT  813000.0 682800.0 823200.0 696600.0 ;
      RECT  813000.0 710400.0 823200.0 696600.0 ;
      RECT  813000.0 710400.0 823200.0 724200.0 ;
      RECT  813000.0 738000.0 823200.0 724200.0 ;
      RECT  813000.0 738000.0 823200.0 751800.0 ;
      RECT  813000.0 765600.0 823200.0 751800.0 ;
      RECT  813000.0 765600.0 823200.0 779400.0 ;
      RECT  813000.0 793200.0 823200.0 779400.0 ;
      RECT  813000.0 793200.0 823200.0 807000.0 ;
      RECT  813000.0 820800.0 823200.0 807000.0 ;
      RECT  813000.0 820800.0 823200.0 834600.0 ;
      RECT  813000.0 848400.0 823200.0 834600.0 ;
      RECT  813000.0 848400.0 823200.0 862200.0 ;
      RECT  813000.0 876000.0 823200.0 862200.0 ;
      RECT  813000.0 876000.0 823200.0 889800.0 ;
      RECT  813000.0 903600.0 823200.0 889800.0 ;
      RECT  813000.0 903600.0 823200.0 917400.0 ;
      RECT  813000.0 931200.0 823200.0 917400.0 ;
      RECT  813000.0 931200.0 823200.0 945000.0 ;
      RECT  813000.0 958800.0 823200.0 945000.0 ;
      RECT  813000.0 958800.0 823200.0 972600.0 ;
      RECT  813000.0 986400.0 823200.0 972600.0 ;
      RECT  813000.0 986400.0 823200.0 1000200.0 ;
      RECT  813000.0 1014000.0 823200.0 1000200.0 ;
      RECT  813000.0 1014000.0 823200.0 1027800.0 ;
      RECT  813000.0 1041600.0 823200.0 1027800.0 ;
      RECT  813000.0 1041600.0 823200.0 1055400.0 ;
      RECT  813000.0 1069200.0 823200.0 1055400.0 ;
      RECT  813000.0 1069200.0 823200.0 1083000.0 ;
      RECT  813000.0 1096800.0 823200.0 1083000.0 ;
      RECT  813000.0 1096800.0 823200.0 1110600.0 ;
      RECT  813000.0 1124400.0 823200.0 1110600.0 ;
      RECT  813000.0 1124400.0 823200.0 1138200.0 ;
      RECT  813000.0 1152000.0 823200.0 1138200.0 ;
      RECT  813000.0 1152000.0 823200.0 1165800.0 ;
      RECT  813000.0 1179600.0 823200.0 1165800.0 ;
      RECT  813000.0 1179600.0 823200.0 1193400.0 ;
      RECT  813000.0 1207200.0 823200.0 1193400.0 ;
      RECT  813000.0 1207200.0 823200.0 1221000.0 ;
      RECT  813000.0 1234800.0 823200.0 1221000.0 ;
      RECT  813000.0 1234800.0 823200.0 1248600.0 ;
      RECT  813000.0 1262400.0 823200.0 1248600.0 ;
      RECT  813000.0 1262400.0 823200.0 1276200.0 ;
      RECT  813000.0 1290000.0 823200.0 1276200.0 ;
      RECT  813000.0 1290000.0 823200.0 1303800.0 ;
      RECT  813000.0 1317600.0 823200.0 1303800.0 ;
      RECT  813000.0 1317600.0 823200.0 1331400.0 ;
      RECT  813000.0 1345200.0 823200.0 1331400.0 ;
      RECT  813000.0 1345200.0 823200.0 1359000.0 ;
      RECT  813000.0 1372800.0 823200.0 1359000.0 ;
      RECT  813000.0 1372800.0 823200.0 1386600.0 ;
      RECT  813000.0 1400400.0 823200.0 1386600.0 ;
      RECT  813000.0 1400400.0 823200.0 1414200.0 ;
      RECT  813000.0 1428000.0 823200.0 1414200.0 ;
      RECT  813000.0 1428000.0 823200.0 1441800.0 ;
      RECT  813000.0 1455600.0 823200.0 1441800.0 ;
      RECT  813000.0 1455600.0 823200.0 1469400.0 ;
      RECT  813000.0 1483200.0 823200.0 1469400.0 ;
      RECT  813000.0 1483200.0 823200.0 1497000.0 ;
      RECT  813000.0 1510800.0 823200.0 1497000.0 ;
      RECT  813000.0 1510800.0 823200.0 1524600.0 ;
      RECT  813000.0 1538400.0 823200.0 1524600.0 ;
      RECT  813000.0 1538400.0 823200.0 1552200.0 ;
      RECT  813000.0 1566000.0 823200.0 1552200.0 ;
      RECT  813000.0 1566000.0 823200.0 1579800.0 ;
      RECT  813000.0 1593600.0 823200.0 1579800.0 ;
      RECT  813000.0 1593600.0 823200.0 1607400.0 ;
      RECT  813000.0 1621200.0 823200.0 1607400.0 ;
      RECT  813000.0 1621200.0 823200.0 1635000.0 ;
      RECT  813000.0 1648800.0 823200.0 1635000.0 ;
      RECT  813000.0 1648800.0 823200.0 1662600.0 ;
      RECT  813000.0 1676400.0 823200.0 1662600.0 ;
      RECT  813000.0 1676400.0 823200.0 1690200.0 ;
      RECT  813000.0 1704000.0 823200.0 1690200.0 ;
      RECT  813000.0 1704000.0 823200.0 1717800.0 ;
      RECT  813000.0 1731600.0 823200.0 1717800.0 ;
      RECT  813000.0 1731600.0 823200.0 1745400.0 ;
      RECT  813000.0 1759200.0 823200.0 1745400.0 ;
      RECT  813000.0 1759200.0 823200.0 1773000.0 ;
      RECT  813000.0 1786800.0 823200.0 1773000.0 ;
      RECT  813000.0 1786800.0 823200.0 1800600.0 ;
      RECT  813000.0 1814400.0 823200.0 1800600.0 ;
      RECT  813000.0 1814400.0 823200.0 1828200.0 ;
      RECT  813000.0 1842000.0 823200.0 1828200.0 ;
      RECT  813000.0 1842000.0 823200.0 1855800.0 ;
      RECT  813000.0 1869600.0 823200.0 1855800.0 ;
      RECT  813000.0 1869600.0 823200.0 1883400.0 ;
      RECT  813000.0 1897200.0 823200.0 1883400.0 ;
      RECT  813000.0 1897200.0 823200.0 1911000.0 ;
      RECT  813000.0 1924800.0 823200.0 1911000.0 ;
      RECT  813000.0 1924800.0 823200.0 1938600.0 ;
      RECT  813000.0 1952400.0 823200.0 1938600.0 ;
      RECT  813000.0 1952400.0 823200.0 1966200.0 ;
      RECT  813000.0 1980000.0 823200.0 1966200.0 ;
      RECT  813000.0 1980000.0 823200.0 1993800.0 ;
      RECT  813000.0 2007600.0 823200.0 1993800.0 ;
      RECT  813000.0 2007600.0 823200.0 2021400.0 ;
      RECT  813000.0 2035200.0 823200.0 2021400.0 ;
      RECT  813000.0 2035200.0 823200.0 2049000.0 ;
      RECT  813000.0 2062800.0 823200.0 2049000.0 ;
      RECT  813000.0 2062800.0 823200.0 2076600.0 ;
      RECT  813000.0 2090400.0 823200.0 2076600.0 ;
      RECT  813000.0 2090400.0 823200.0 2104200.0 ;
      RECT  813000.0 2118000.0 823200.0 2104200.0 ;
      RECT  813000.0 2118000.0 823200.0 2131800.0 ;
      RECT  813000.0 2145600.0 823200.0 2131800.0 ;
      RECT  823200.0 379200.0 833400.0 393000.0 ;
      RECT  823200.0 406800.0 833400.0 393000.0 ;
      RECT  823200.0 406800.0 833400.0 420600.0 ;
      RECT  823200.0 434400.0 833400.0 420600.0 ;
      RECT  823200.0 434400.0 833400.0 448200.0 ;
      RECT  823200.0 462000.0 833400.0 448200.0 ;
      RECT  823200.0 462000.0 833400.0 475800.0 ;
      RECT  823200.0 489600.0 833400.0 475800.0 ;
      RECT  823200.0 489600.0 833400.0 503400.0 ;
      RECT  823200.0 517200.0 833400.0 503400.0 ;
      RECT  823200.0 517200.0 833400.0 531000.0 ;
      RECT  823200.0 544800.0 833400.0 531000.0 ;
      RECT  823200.0 544800.0 833400.0 558600.0 ;
      RECT  823200.0 572400.0 833400.0 558600.0 ;
      RECT  823200.0 572400.0 833400.0 586200.0 ;
      RECT  823200.0 600000.0 833400.0 586200.0 ;
      RECT  823200.0 600000.0 833400.0 613800.0 ;
      RECT  823200.0 627600.0 833400.0 613800.0 ;
      RECT  823200.0 627600.0 833400.0 641400.0 ;
      RECT  823200.0 655200.0 833400.0 641400.0 ;
      RECT  823200.0 655200.0 833400.0 669000.0 ;
      RECT  823200.0 682800.0 833400.0 669000.0 ;
      RECT  823200.0 682800.0 833400.0 696600.0 ;
      RECT  823200.0 710400.0 833400.0 696600.0 ;
      RECT  823200.0 710400.0 833400.0 724200.0 ;
      RECT  823200.0 738000.0 833400.0 724200.0 ;
      RECT  823200.0 738000.0 833400.0 751800.0 ;
      RECT  823200.0 765600.0 833400.0 751800.0 ;
      RECT  823200.0 765600.0 833400.0 779400.0 ;
      RECT  823200.0 793200.0 833400.0 779400.0 ;
      RECT  823200.0 793200.0 833400.0 807000.0 ;
      RECT  823200.0 820800.0 833400.0 807000.0 ;
      RECT  823200.0 820800.0 833400.0 834600.0 ;
      RECT  823200.0 848400.0 833400.0 834600.0 ;
      RECT  823200.0 848400.0 833400.0 862200.0 ;
      RECT  823200.0 876000.0 833400.0 862200.0 ;
      RECT  823200.0 876000.0 833400.0 889800.0 ;
      RECT  823200.0 903600.0 833400.0 889800.0 ;
      RECT  823200.0 903600.0 833400.0 917400.0 ;
      RECT  823200.0 931200.0 833400.0 917400.0 ;
      RECT  823200.0 931200.0 833400.0 945000.0 ;
      RECT  823200.0 958800.0 833400.0 945000.0 ;
      RECT  823200.0 958800.0 833400.0 972600.0 ;
      RECT  823200.0 986400.0 833400.0 972600.0 ;
      RECT  823200.0 986400.0 833400.0 1000200.0 ;
      RECT  823200.0 1014000.0 833400.0 1000200.0 ;
      RECT  823200.0 1014000.0 833400.0 1027800.0 ;
      RECT  823200.0 1041600.0 833400.0 1027800.0 ;
      RECT  823200.0 1041600.0 833400.0 1055400.0 ;
      RECT  823200.0 1069200.0 833400.0 1055400.0 ;
      RECT  823200.0 1069200.0 833400.0 1083000.0 ;
      RECT  823200.0 1096800.0 833400.0 1083000.0 ;
      RECT  823200.0 1096800.0 833400.0 1110600.0 ;
      RECT  823200.0 1124400.0 833400.0 1110600.0 ;
      RECT  823200.0 1124400.0 833400.0 1138200.0 ;
      RECT  823200.0 1152000.0 833400.0 1138200.0 ;
      RECT  823200.0 1152000.0 833400.0 1165800.0 ;
      RECT  823200.0 1179600.0 833400.0 1165800.0 ;
      RECT  823200.0 1179600.0 833400.0 1193400.0 ;
      RECT  823200.0 1207200.0 833400.0 1193400.0 ;
      RECT  823200.0 1207200.0 833400.0 1221000.0 ;
      RECT  823200.0 1234800.0 833400.0 1221000.0 ;
      RECT  823200.0 1234800.0 833400.0 1248600.0 ;
      RECT  823200.0 1262400.0 833400.0 1248600.0 ;
      RECT  823200.0 1262400.0 833400.0 1276200.0 ;
      RECT  823200.0 1290000.0 833400.0 1276200.0 ;
      RECT  823200.0 1290000.0 833400.0 1303800.0 ;
      RECT  823200.0 1317600.0 833400.0 1303800.0 ;
      RECT  823200.0 1317600.0 833400.0 1331400.0 ;
      RECT  823200.0 1345200.0 833400.0 1331400.0 ;
      RECT  823200.0 1345200.0 833400.0 1359000.0 ;
      RECT  823200.0 1372800.0 833400.0 1359000.0 ;
      RECT  823200.0 1372800.0 833400.0 1386600.0 ;
      RECT  823200.0 1400400.0 833400.0 1386600.0 ;
      RECT  823200.0 1400400.0 833400.0 1414200.0 ;
      RECT  823200.0 1428000.0 833400.0 1414200.0 ;
      RECT  823200.0 1428000.0 833400.0 1441800.0 ;
      RECT  823200.0 1455600.0 833400.0 1441800.0 ;
      RECT  823200.0 1455600.0 833400.0 1469400.0 ;
      RECT  823200.0 1483200.0 833400.0 1469400.0 ;
      RECT  823200.0 1483200.0 833400.0 1497000.0 ;
      RECT  823200.0 1510800.0 833400.0 1497000.0 ;
      RECT  823200.0 1510800.0 833400.0 1524600.0 ;
      RECT  823200.0 1538400.0 833400.0 1524600.0 ;
      RECT  823200.0 1538400.0 833400.0 1552200.0 ;
      RECT  823200.0 1566000.0 833400.0 1552200.0 ;
      RECT  823200.0 1566000.0 833400.0 1579800.0 ;
      RECT  823200.0 1593600.0 833400.0 1579800.0 ;
      RECT  823200.0 1593600.0 833400.0 1607400.0 ;
      RECT  823200.0 1621200.0 833400.0 1607400.0 ;
      RECT  823200.0 1621200.0 833400.0 1635000.0 ;
      RECT  823200.0 1648800.0 833400.0 1635000.0 ;
      RECT  823200.0 1648800.0 833400.0 1662600.0 ;
      RECT  823200.0 1676400.0 833400.0 1662600.0 ;
      RECT  823200.0 1676400.0 833400.0 1690200.0 ;
      RECT  823200.0 1704000.0 833400.0 1690200.0 ;
      RECT  823200.0 1704000.0 833400.0 1717800.0 ;
      RECT  823200.0 1731600.0 833400.0 1717800.0 ;
      RECT  823200.0 1731600.0 833400.0 1745400.0 ;
      RECT  823200.0 1759200.0 833400.0 1745400.0 ;
      RECT  823200.0 1759200.0 833400.0 1773000.0 ;
      RECT  823200.0 1786800.0 833400.0 1773000.0 ;
      RECT  823200.0 1786800.0 833400.0 1800600.0 ;
      RECT  823200.0 1814400.0 833400.0 1800600.0 ;
      RECT  823200.0 1814400.0 833400.0 1828200.0 ;
      RECT  823200.0 1842000.0 833400.0 1828200.0 ;
      RECT  823200.0 1842000.0 833400.0 1855800.0 ;
      RECT  823200.0 1869600.0 833400.0 1855800.0 ;
      RECT  823200.0 1869600.0 833400.0 1883400.0 ;
      RECT  823200.0 1897200.0 833400.0 1883400.0 ;
      RECT  823200.0 1897200.0 833400.0 1911000.0 ;
      RECT  823200.0 1924800.0 833400.0 1911000.0 ;
      RECT  823200.0 1924800.0 833400.0 1938600.0 ;
      RECT  823200.0 1952400.0 833400.0 1938600.0 ;
      RECT  823200.0 1952400.0 833400.0 1966200.0 ;
      RECT  823200.0 1980000.0 833400.0 1966200.0 ;
      RECT  823200.0 1980000.0 833400.0 1993800.0 ;
      RECT  823200.0 2007600.0 833400.0 1993800.0 ;
      RECT  823200.0 2007600.0 833400.0 2021400.0 ;
      RECT  823200.0 2035200.0 833400.0 2021400.0 ;
      RECT  823200.0 2035200.0 833400.0 2049000.0 ;
      RECT  823200.0 2062800.0 833400.0 2049000.0 ;
      RECT  823200.0 2062800.0 833400.0 2076600.0 ;
      RECT  823200.0 2090400.0 833400.0 2076600.0 ;
      RECT  823200.0 2090400.0 833400.0 2104200.0 ;
      RECT  823200.0 2118000.0 833400.0 2104200.0 ;
      RECT  823200.0 2118000.0 833400.0 2131800.0 ;
      RECT  823200.0 2145600.0 833400.0 2131800.0 ;
      RECT  833400.0 379200.0 843600.0 393000.0 ;
      RECT  833400.0 406800.0 843600.0 393000.0 ;
      RECT  833400.0 406800.0 843600.0 420600.0 ;
      RECT  833400.0 434400.0 843600.0 420600.0 ;
      RECT  833400.0 434400.0 843600.0 448200.0 ;
      RECT  833400.0 462000.0 843600.0 448200.0 ;
      RECT  833400.0 462000.0 843600.0 475800.0 ;
      RECT  833400.0 489600.0 843600.0 475800.0 ;
      RECT  833400.0 489600.0 843600.0 503400.0 ;
      RECT  833400.0 517200.0 843600.0 503400.0 ;
      RECT  833400.0 517200.0 843600.0 531000.0 ;
      RECT  833400.0 544800.0 843600.0 531000.0 ;
      RECT  833400.0 544800.0 843600.0 558600.0 ;
      RECT  833400.0 572400.0 843600.0 558600.0 ;
      RECT  833400.0 572400.0 843600.0 586200.0 ;
      RECT  833400.0 600000.0 843600.0 586200.0 ;
      RECT  833400.0 600000.0 843600.0 613800.0 ;
      RECT  833400.0 627600.0 843600.0 613800.0 ;
      RECT  833400.0 627600.0 843600.0 641400.0 ;
      RECT  833400.0 655200.0 843600.0 641400.0 ;
      RECT  833400.0 655200.0 843600.0 669000.0 ;
      RECT  833400.0 682800.0 843600.0 669000.0 ;
      RECT  833400.0 682800.0 843600.0 696600.0 ;
      RECT  833400.0 710400.0 843600.0 696600.0 ;
      RECT  833400.0 710400.0 843600.0 724200.0 ;
      RECT  833400.0 738000.0 843600.0 724200.0 ;
      RECT  833400.0 738000.0 843600.0 751800.0 ;
      RECT  833400.0 765600.0 843600.0 751800.0 ;
      RECT  833400.0 765600.0 843600.0 779400.0 ;
      RECT  833400.0 793200.0 843600.0 779400.0 ;
      RECT  833400.0 793200.0 843600.0 807000.0 ;
      RECT  833400.0 820800.0 843600.0 807000.0 ;
      RECT  833400.0 820800.0 843600.0 834600.0 ;
      RECT  833400.0 848400.0 843600.0 834600.0 ;
      RECT  833400.0 848400.0 843600.0 862200.0 ;
      RECT  833400.0 876000.0 843600.0 862200.0 ;
      RECT  833400.0 876000.0 843600.0 889800.0 ;
      RECT  833400.0 903600.0 843600.0 889800.0 ;
      RECT  833400.0 903600.0 843600.0 917400.0 ;
      RECT  833400.0 931200.0 843600.0 917400.0 ;
      RECT  833400.0 931200.0 843600.0 945000.0 ;
      RECT  833400.0 958800.0 843600.0 945000.0 ;
      RECT  833400.0 958800.0 843600.0 972600.0 ;
      RECT  833400.0 986400.0 843600.0 972600.0 ;
      RECT  833400.0 986400.0 843600.0 1000200.0 ;
      RECT  833400.0 1014000.0 843600.0 1000200.0 ;
      RECT  833400.0 1014000.0 843600.0 1027800.0 ;
      RECT  833400.0 1041600.0 843600.0 1027800.0 ;
      RECT  833400.0 1041600.0 843600.0 1055400.0 ;
      RECT  833400.0 1069200.0 843600.0 1055400.0 ;
      RECT  833400.0 1069200.0 843600.0 1083000.0 ;
      RECT  833400.0 1096800.0 843600.0 1083000.0 ;
      RECT  833400.0 1096800.0 843600.0 1110600.0 ;
      RECT  833400.0 1124400.0 843600.0 1110600.0 ;
      RECT  833400.0 1124400.0 843600.0 1138200.0 ;
      RECT  833400.0 1152000.0 843600.0 1138200.0 ;
      RECT  833400.0 1152000.0 843600.0 1165800.0 ;
      RECT  833400.0 1179600.0 843600.0 1165800.0 ;
      RECT  833400.0 1179600.0 843600.0 1193400.0 ;
      RECT  833400.0 1207200.0 843600.0 1193400.0 ;
      RECT  833400.0 1207200.0 843600.0 1221000.0 ;
      RECT  833400.0 1234800.0 843600.0 1221000.0 ;
      RECT  833400.0 1234800.0 843600.0 1248600.0 ;
      RECT  833400.0 1262400.0 843600.0 1248600.0 ;
      RECT  833400.0 1262400.0 843600.0 1276200.0 ;
      RECT  833400.0 1290000.0 843600.0 1276200.0 ;
      RECT  833400.0 1290000.0 843600.0 1303800.0 ;
      RECT  833400.0 1317600.0 843600.0 1303800.0 ;
      RECT  833400.0 1317600.0 843600.0 1331400.0 ;
      RECT  833400.0 1345200.0 843600.0 1331400.0 ;
      RECT  833400.0 1345200.0 843600.0 1359000.0 ;
      RECT  833400.0 1372800.0 843600.0 1359000.0 ;
      RECT  833400.0 1372800.0 843600.0 1386600.0 ;
      RECT  833400.0 1400400.0 843600.0 1386600.0 ;
      RECT  833400.0 1400400.0 843600.0 1414200.0 ;
      RECT  833400.0 1428000.0 843600.0 1414200.0 ;
      RECT  833400.0 1428000.0 843600.0 1441800.0 ;
      RECT  833400.0 1455600.0 843600.0 1441800.0 ;
      RECT  833400.0 1455600.0 843600.0 1469400.0 ;
      RECT  833400.0 1483200.0 843600.0 1469400.0 ;
      RECT  833400.0 1483200.0 843600.0 1497000.0 ;
      RECT  833400.0 1510800.0 843600.0 1497000.0 ;
      RECT  833400.0 1510800.0 843600.0 1524600.0 ;
      RECT  833400.0 1538400.0 843600.0 1524600.0 ;
      RECT  833400.0 1538400.0 843600.0 1552200.0 ;
      RECT  833400.0 1566000.0 843600.0 1552200.0 ;
      RECT  833400.0 1566000.0 843600.0 1579800.0 ;
      RECT  833400.0 1593600.0 843600.0 1579800.0 ;
      RECT  833400.0 1593600.0 843600.0 1607400.0 ;
      RECT  833400.0 1621200.0 843600.0 1607400.0 ;
      RECT  833400.0 1621200.0 843600.0 1635000.0 ;
      RECT  833400.0 1648800.0 843600.0 1635000.0 ;
      RECT  833400.0 1648800.0 843600.0 1662600.0 ;
      RECT  833400.0 1676400.0 843600.0 1662600.0 ;
      RECT  833400.0 1676400.0 843600.0 1690200.0 ;
      RECT  833400.0 1704000.0 843600.0 1690200.0 ;
      RECT  833400.0 1704000.0 843600.0 1717800.0 ;
      RECT  833400.0 1731600.0 843600.0 1717800.0 ;
      RECT  833400.0 1731600.0 843600.0 1745400.0 ;
      RECT  833400.0 1759200.0 843600.0 1745400.0 ;
      RECT  833400.0 1759200.0 843600.0 1773000.0 ;
      RECT  833400.0 1786800.0 843600.0 1773000.0 ;
      RECT  833400.0 1786800.0 843600.0 1800600.0 ;
      RECT  833400.0 1814400.0 843600.0 1800600.0 ;
      RECT  833400.0 1814400.0 843600.0 1828200.0 ;
      RECT  833400.0 1842000.0 843600.0 1828200.0 ;
      RECT  833400.0 1842000.0 843600.0 1855800.0 ;
      RECT  833400.0 1869600.0 843600.0 1855800.0 ;
      RECT  833400.0 1869600.0 843600.0 1883400.0 ;
      RECT  833400.0 1897200.0 843600.0 1883400.0 ;
      RECT  833400.0 1897200.0 843600.0 1911000.0 ;
      RECT  833400.0 1924800.0 843600.0 1911000.0 ;
      RECT  833400.0 1924800.0 843600.0 1938600.0 ;
      RECT  833400.0 1952400.0 843600.0 1938600.0 ;
      RECT  833400.0 1952400.0 843600.0 1966200.0 ;
      RECT  833400.0 1980000.0 843600.0 1966200.0 ;
      RECT  833400.0 1980000.0 843600.0 1993800.0 ;
      RECT  833400.0 2007600.0 843600.0 1993800.0 ;
      RECT  833400.0 2007600.0 843600.0 2021400.0 ;
      RECT  833400.0 2035200.0 843600.0 2021400.0 ;
      RECT  833400.0 2035200.0 843600.0 2049000.0 ;
      RECT  833400.0 2062800.0 843600.0 2049000.0 ;
      RECT  833400.0 2062800.0 843600.0 2076600.0 ;
      RECT  833400.0 2090400.0 843600.0 2076600.0 ;
      RECT  833400.0 2090400.0 843600.0 2104200.0 ;
      RECT  833400.0 2118000.0 843600.0 2104200.0 ;
      RECT  833400.0 2118000.0 843600.0 2131800.0 ;
      RECT  833400.0 2145600.0 843600.0 2131800.0 ;
      RECT  843600.0 379200.0 853800.0 393000.0 ;
      RECT  843600.0 406800.0 853800.0 393000.0 ;
      RECT  843600.0 406800.0 853800.0 420600.0 ;
      RECT  843600.0 434400.0 853800.0 420600.0 ;
      RECT  843600.0 434400.0 853800.0 448200.0 ;
      RECT  843600.0 462000.0 853800.0 448200.0 ;
      RECT  843600.0 462000.0 853800.0 475800.0 ;
      RECT  843600.0 489600.0 853800.0 475800.0 ;
      RECT  843600.0 489600.0 853800.0 503400.0 ;
      RECT  843600.0 517200.0 853800.0 503400.0 ;
      RECT  843600.0 517200.0 853800.0 531000.0 ;
      RECT  843600.0 544800.0 853800.0 531000.0 ;
      RECT  843600.0 544800.0 853800.0 558600.0 ;
      RECT  843600.0 572400.0 853800.0 558600.0 ;
      RECT  843600.0 572400.0 853800.0 586200.0 ;
      RECT  843600.0 600000.0 853800.0 586200.0 ;
      RECT  843600.0 600000.0 853800.0 613800.0 ;
      RECT  843600.0 627600.0 853800.0 613800.0 ;
      RECT  843600.0 627600.0 853800.0 641400.0 ;
      RECT  843600.0 655200.0 853800.0 641400.0 ;
      RECT  843600.0 655200.0 853800.0 669000.0 ;
      RECT  843600.0 682800.0 853800.0 669000.0 ;
      RECT  843600.0 682800.0 853800.0 696600.0 ;
      RECT  843600.0 710400.0 853800.0 696600.0 ;
      RECT  843600.0 710400.0 853800.0 724200.0 ;
      RECT  843600.0 738000.0 853800.0 724200.0 ;
      RECT  843600.0 738000.0 853800.0 751800.0 ;
      RECT  843600.0 765600.0 853800.0 751800.0 ;
      RECT  843600.0 765600.0 853800.0 779400.0 ;
      RECT  843600.0 793200.0 853800.0 779400.0 ;
      RECT  843600.0 793200.0 853800.0 807000.0 ;
      RECT  843600.0 820800.0 853800.0 807000.0 ;
      RECT  843600.0 820800.0 853800.0 834600.0 ;
      RECT  843600.0 848400.0 853800.0 834600.0 ;
      RECT  843600.0 848400.0 853800.0 862200.0 ;
      RECT  843600.0 876000.0 853800.0 862200.0 ;
      RECT  843600.0 876000.0 853800.0 889800.0 ;
      RECT  843600.0 903600.0 853800.0 889800.0 ;
      RECT  843600.0 903600.0 853800.0 917400.0 ;
      RECT  843600.0 931200.0 853800.0 917400.0 ;
      RECT  843600.0 931200.0 853800.0 945000.0 ;
      RECT  843600.0 958800.0 853800.0 945000.0 ;
      RECT  843600.0 958800.0 853800.0 972600.0 ;
      RECT  843600.0 986400.0 853800.0 972600.0 ;
      RECT  843600.0 986400.0 853800.0 1000200.0 ;
      RECT  843600.0 1014000.0 853800.0 1000200.0 ;
      RECT  843600.0 1014000.0 853800.0 1027800.0 ;
      RECT  843600.0 1041600.0 853800.0 1027800.0 ;
      RECT  843600.0 1041600.0 853800.0 1055400.0 ;
      RECT  843600.0 1069200.0 853800.0 1055400.0 ;
      RECT  843600.0 1069200.0 853800.0 1083000.0 ;
      RECT  843600.0 1096800.0 853800.0 1083000.0 ;
      RECT  843600.0 1096800.0 853800.0 1110600.0 ;
      RECT  843600.0 1124400.0 853800.0 1110600.0 ;
      RECT  843600.0 1124400.0 853800.0 1138200.0 ;
      RECT  843600.0 1152000.0 853800.0 1138200.0 ;
      RECT  843600.0 1152000.0 853800.0 1165800.0 ;
      RECT  843600.0 1179600.0 853800.0 1165800.0 ;
      RECT  843600.0 1179600.0 853800.0 1193400.0 ;
      RECT  843600.0 1207200.0 853800.0 1193400.0 ;
      RECT  843600.0 1207200.0 853800.0 1221000.0 ;
      RECT  843600.0 1234800.0 853800.0 1221000.0 ;
      RECT  843600.0 1234800.0 853800.0 1248600.0 ;
      RECT  843600.0 1262400.0 853800.0 1248600.0 ;
      RECT  843600.0 1262400.0 853800.0 1276200.0 ;
      RECT  843600.0 1290000.0 853800.0 1276200.0 ;
      RECT  843600.0 1290000.0 853800.0 1303800.0 ;
      RECT  843600.0 1317600.0 853800.0 1303800.0 ;
      RECT  843600.0 1317600.0 853800.0 1331400.0 ;
      RECT  843600.0 1345200.0 853800.0 1331400.0 ;
      RECT  843600.0 1345200.0 853800.0 1359000.0 ;
      RECT  843600.0 1372800.0 853800.0 1359000.0 ;
      RECT  843600.0 1372800.0 853800.0 1386600.0 ;
      RECT  843600.0 1400400.0 853800.0 1386600.0 ;
      RECT  843600.0 1400400.0 853800.0 1414200.0 ;
      RECT  843600.0 1428000.0 853800.0 1414200.0 ;
      RECT  843600.0 1428000.0 853800.0 1441800.0 ;
      RECT  843600.0 1455600.0 853800.0 1441800.0 ;
      RECT  843600.0 1455600.0 853800.0 1469400.0 ;
      RECT  843600.0 1483200.0 853800.0 1469400.0 ;
      RECT  843600.0 1483200.0 853800.0 1497000.0 ;
      RECT  843600.0 1510800.0 853800.0 1497000.0 ;
      RECT  843600.0 1510800.0 853800.0 1524600.0 ;
      RECT  843600.0 1538400.0 853800.0 1524600.0 ;
      RECT  843600.0 1538400.0 853800.0 1552200.0 ;
      RECT  843600.0 1566000.0 853800.0 1552200.0 ;
      RECT  843600.0 1566000.0 853800.0 1579800.0 ;
      RECT  843600.0 1593600.0 853800.0 1579800.0 ;
      RECT  843600.0 1593600.0 853800.0 1607400.0 ;
      RECT  843600.0 1621200.0 853800.0 1607400.0 ;
      RECT  843600.0 1621200.0 853800.0 1635000.0 ;
      RECT  843600.0 1648800.0 853800.0 1635000.0 ;
      RECT  843600.0 1648800.0 853800.0 1662600.0 ;
      RECT  843600.0 1676400.0 853800.0 1662600.0 ;
      RECT  843600.0 1676400.0 853800.0 1690200.0 ;
      RECT  843600.0 1704000.0 853800.0 1690200.0 ;
      RECT  843600.0 1704000.0 853800.0 1717800.0 ;
      RECT  843600.0 1731600.0 853800.0 1717800.0 ;
      RECT  843600.0 1731600.0 853800.0 1745400.0 ;
      RECT  843600.0 1759200.0 853800.0 1745400.0 ;
      RECT  843600.0 1759200.0 853800.0 1773000.0 ;
      RECT  843600.0 1786800.0 853800.0 1773000.0 ;
      RECT  843600.0 1786800.0 853800.0 1800600.0 ;
      RECT  843600.0 1814400.0 853800.0 1800600.0 ;
      RECT  843600.0 1814400.0 853800.0 1828200.0 ;
      RECT  843600.0 1842000.0 853800.0 1828200.0 ;
      RECT  843600.0 1842000.0 853800.0 1855800.0 ;
      RECT  843600.0 1869600.0 853800.0 1855800.0 ;
      RECT  843600.0 1869600.0 853800.0 1883400.0 ;
      RECT  843600.0 1897200.0 853800.0 1883400.0 ;
      RECT  843600.0 1897200.0 853800.0 1911000.0 ;
      RECT  843600.0 1924800.0 853800.0 1911000.0 ;
      RECT  843600.0 1924800.0 853800.0 1938600.0 ;
      RECT  843600.0 1952400.0 853800.0 1938600.0 ;
      RECT  843600.0 1952400.0 853800.0 1966200.0 ;
      RECT  843600.0 1980000.0 853800.0 1966200.0 ;
      RECT  843600.0 1980000.0 853800.0 1993800.0 ;
      RECT  843600.0 2007600.0 853800.0 1993800.0 ;
      RECT  843600.0 2007600.0 853800.0 2021400.0 ;
      RECT  843600.0 2035200.0 853800.0 2021400.0 ;
      RECT  843600.0 2035200.0 853800.0 2049000.0 ;
      RECT  843600.0 2062800.0 853800.0 2049000.0 ;
      RECT  843600.0 2062800.0 853800.0 2076600.0 ;
      RECT  843600.0 2090400.0 853800.0 2076600.0 ;
      RECT  843600.0 2090400.0 853800.0 2104200.0 ;
      RECT  843600.0 2118000.0 853800.0 2104200.0 ;
      RECT  843600.0 2118000.0 853800.0 2131800.0 ;
      RECT  843600.0 2145600.0 853800.0 2131800.0 ;
      RECT  853800.0 379200.0 864000.0 393000.0 ;
      RECT  853800.0 406800.0 864000.0 393000.0 ;
      RECT  853800.0 406800.0 864000.0 420600.0 ;
      RECT  853800.0 434400.0 864000.0 420600.0 ;
      RECT  853800.0 434400.0 864000.0 448200.0 ;
      RECT  853800.0 462000.0 864000.0 448200.0 ;
      RECT  853800.0 462000.0 864000.0 475800.0 ;
      RECT  853800.0 489600.0 864000.0 475800.0 ;
      RECT  853800.0 489600.0 864000.0 503400.0 ;
      RECT  853800.0 517200.0 864000.0 503400.0 ;
      RECT  853800.0 517200.0 864000.0 531000.0 ;
      RECT  853800.0 544800.0 864000.0 531000.0 ;
      RECT  853800.0 544800.0 864000.0 558600.0 ;
      RECT  853800.0 572400.0 864000.0 558600.0 ;
      RECT  853800.0 572400.0 864000.0 586200.0 ;
      RECT  853800.0 600000.0 864000.0 586200.0 ;
      RECT  853800.0 600000.0 864000.0 613800.0 ;
      RECT  853800.0 627600.0 864000.0 613800.0 ;
      RECT  853800.0 627600.0 864000.0 641400.0 ;
      RECT  853800.0 655200.0 864000.0 641400.0 ;
      RECT  853800.0 655200.0 864000.0 669000.0 ;
      RECT  853800.0 682800.0 864000.0 669000.0 ;
      RECT  853800.0 682800.0 864000.0 696600.0 ;
      RECT  853800.0 710400.0 864000.0 696600.0 ;
      RECT  853800.0 710400.0 864000.0 724200.0 ;
      RECT  853800.0 738000.0 864000.0 724200.0 ;
      RECT  853800.0 738000.0 864000.0 751800.0 ;
      RECT  853800.0 765600.0 864000.0 751800.0 ;
      RECT  853800.0 765600.0 864000.0 779400.0 ;
      RECT  853800.0 793200.0 864000.0 779400.0 ;
      RECT  853800.0 793200.0 864000.0 807000.0 ;
      RECT  853800.0 820800.0 864000.0 807000.0 ;
      RECT  853800.0 820800.0 864000.0 834600.0 ;
      RECT  853800.0 848400.0 864000.0 834600.0 ;
      RECT  853800.0 848400.0 864000.0 862200.0 ;
      RECT  853800.0 876000.0 864000.0 862200.0 ;
      RECT  853800.0 876000.0 864000.0 889800.0 ;
      RECT  853800.0 903600.0 864000.0 889800.0 ;
      RECT  853800.0 903600.0 864000.0 917400.0 ;
      RECT  853800.0 931200.0 864000.0 917400.0 ;
      RECT  853800.0 931200.0 864000.0 945000.0 ;
      RECT  853800.0 958800.0 864000.0 945000.0 ;
      RECT  853800.0 958800.0 864000.0 972600.0 ;
      RECT  853800.0 986400.0 864000.0 972600.0 ;
      RECT  853800.0 986400.0 864000.0 1000200.0 ;
      RECT  853800.0 1014000.0 864000.0 1000200.0 ;
      RECT  853800.0 1014000.0 864000.0 1027800.0 ;
      RECT  853800.0 1041600.0 864000.0 1027800.0 ;
      RECT  853800.0 1041600.0 864000.0 1055400.0 ;
      RECT  853800.0 1069200.0 864000.0 1055400.0 ;
      RECT  853800.0 1069200.0 864000.0 1083000.0 ;
      RECT  853800.0 1096800.0 864000.0 1083000.0 ;
      RECT  853800.0 1096800.0 864000.0 1110600.0 ;
      RECT  853800.0 1124400.0 864000.0 1110600.0 ;
      RECT  853800.0 1124400.0 864000.0 1138200.0 ;
      RECT  853800.0 1152000.0 864000.0 1138200.0 ;
      RECT  853800.0 1152000.0 864000.0 1165800.0 ;
      RECT  853800.0 1179600.0 864000.0 1165800.0 ;
      RECT  853800.0 1179600.0 864000.0 1193400.0 ;
      RECT  853800.0 1207200.0 864000.0 1193400.0 ;
      RECT  853800.0 1207200.0 864000.0 1221000.0 ;
      RECT  853800.0 1234800.0 864000.0 1221000.0 ;
      RECT  853800.0 1234800.0 864000.0 1248600.0 ;
      RECT  853800.0 1262400.0 864000.0 1248600.0 ;
      RECT  853800.0 1262400.0 864000.0 1276200.0 ;
      RECT  853800.0 1290000.0 864000.0 1276200.0 ;
      RECT  853800.0 1290000.0 864000.0 1303800.0 ;
      RECT  853800.0 1317600.0 864000.0 1303800.0 ;
      RECT  853800.0 1317600.0 864000.0 1331400.0 ;
      RECT  853800.0 1345200.0 864000.0 1331400.0 ;
      RECT  853800.0 1345200.0 864000.0 1359000.0 ;
      RECT  853800.0 1372800.0 864000.0 1359000.0 ;
      RECT  853800.0 1372800.0 864000.0 1386600.0 ;
      RECT  853800.0 1400400.0 864000.0 1386600.0 ;
      RECT  853800.0 1400400.0 864000.0 1414200.0 ;
      RECT  853800.0 1428000.0 864000.0 1414200.0 ;
      RECT  853800.0 1428000.0 864000.0 1441800.0 ;
      RECT  853800.0 1455600.0 864000.0 1441800.0 ;
      RECT  853800.0 1455600.0 864000.0 1469400.0 ;
      RECT  853800.0 1483200.0 864000.0 1469400.0 ;
      RECT  853800.0 1483200.0 864000.0 1497000.0 ;
      RECT  853800.0 1510800.0 864000.0 1497000.0 ;
      RECT  853800.0 1510800.0 864000.0 1524600.0 ;
      RECT  853800.0 1538400.0 864000.0 1524600.0 ;
      RECT  853800.0 1538400.0 864000.0 1552200.0 ;
      RECT  853800.0 1566000.0 864000.0 1552200.0 ;
      RECT  853800.0 1566000.0 864000.0 1579800.0 ;
      RECT  853800.0 1593600.0 864000.0 1579800.0 ;
      RECT  853800.0 1593600.0 864000.0 1607400.0 ;
      RECT  853800.0 1621200.0 864000.0 1607400.0 ;
      RECT  853800.0 1621200.0 864000.0 1635000.0 ;
      RECT  853800.0 1648800.0 864000.0 1635000.0 ;
      RECT  853800.0 1648800.0 864000.0 1662600.0 ;
      RECT  853800.0 1676400.0 864000.0 1662600.0 ;
      RECT  853800.0 1676400.0 864000.0 1690200.0 ;
      RECT  853800.0 1704000.0 864000.0 1690200.0 ;
      RECT  853800.0 1704000.0 864000.0 1717800.0 ;
      RECT  853800.0 1731600.0 864000.0 1717800.0 ;
      RECT  853800.0 1731600.0 864000.0 1745400.0 ;
      RECT  853800.0 1759200.0 864000.0 1745400.0 ;
      RECT  853800.0 1759200.0 864000.0 1773000.0 ;
      RECT  853800.0 1786800.0 864000.0 1773000.0 ;
      RECT  853800.0 1786800.0 864000.0 1800600.0 ;
      RECT  853800.0 1814400.0 864000.0 1800600.0 ;
      RECT  853800.0 1814400.0 864000.0 1828200.0 ;
      RECT  853800.0 1842000.0 864000.0 1828200.0 ;
      RECT  853800.0 1842000.0 864000.0 1855800.0 ;
      RECT  853800.0 1869600.0 864000.0 1855800.0 ;
      RECT  853800.0 1869600.0 864000.0 1883400.0 ;
      RECT  853800.0 1897200.0 864000.0 1883400.0 ;
      RECT  853800.0 1897200.0 864000.0 1911000.0 ;
      RECT  853800.0 1924800.0 864000.0 1911000.0 ;
      RECT  853800.0 1924800.0 864000.0 1938600.0 ;
      RECT  853800.0 1952400.0 864000.0 1938600.0 ;
      RECT  853800.0 1952400.0 864000.0 1966200.0 ;
      RECT  853800.0 1980000.0 864000.0 1966200.0 ;
      RECT  853800.0 1980000.0 864000.0 1993800.0 ;
      RECT  853800.0 2007600.0 864000.0 1993800.0 ;
      RECT  853800.0 2007600.0 864000.0 2021400.0 ;
      RECT  853800.0 2035200.0 864000.0 2021400.0 ;
      RECT  853800.0 2035200.0 864000.0 2049000.0 ;
      RECT  853800.0 2062800.0 864000.0 2049000.0 ;
      RECT  853800.0 2062800.0 864000.0 2076600.0 ;
      RECT  853800.0 2090400.0 864000.0 2076600.0 ;
      RECT  853800.0 2090400.0 864000.0 2104200.0 ;
      RECT  853800.0 2118000.0 864000.0 2104200.0 ;
      RECT  853800.0 2118000.0 864000.0 2131800.0 ;
      RECT  853800.0 2145600.0 864000.0 2131800.0 ;
      RECT  864000.0 379200.0 874200.0 393000.0 ;
      RECT  864000.0 406800.0 874200.0 393000.0 ;
      RECT  864000.0 406800.0 874200.0 420600.0 ;
      RECT  864000.0 434400.0 874200.0 420600.0 ;
      RECT  864000.0 434400.0 874200.0 448200.0 ;
      RECT  864000.0 462000.0 874200.0 448200.0 ;
      RECT  864000.0 462000.0 874200.0 475800.0 ;
      RECT  864000.0 489600.0 874200.0 475800.0 ;
      RECT  864000.0 489600.0 874200.0 503400.0 ;
      RECT  864000.0 517200.0 874200.0 503400.0 ;
      RECT  864000.0 517200.0 874200.0 531000.0 ;
      RECT  864000.0 544800.0 874200.0 531000.0 ;
      RECT  864000.0 544800.0 874200.0 558600.0 ;
      RECT  864000.0 572400.0 874200.0 558600.0 ;
      RECT  864000.0 572400.0 874200.0 586200.0 ;
      RECT  864000.0 600000.0 874200.0 586200.0 ;
      RECT  864000.0 600000.0 874200.0 613800.0 ;
      RECT  864000.0 627600.0 874200.0 613800.0 ;
      RECT  864000.0 627600.0 874200.0 641400.0 ;
      RECT  864000.0 655200.0 874200.0 641400.0 ;
      RECT  864000.0 655200.0 874200.0 669000.0 ;
      RECT  864000.0 682800.0 874200.0 669000.0 ;
      RECT  864000.0 682800.0 874200.0 696600.0 ;
      RECT  864000.0 710400.0 874200.0 696600.0 ;
      RECT  864000.0 710400.0 874200.0 724200.0 ;
      RECT  864000.0 738000.0 874200.0 724200.0 ;
      RECT  864000.0 738000.0 874200.0 751800.0 ;
      RECT  864000.0 765600.0 874200.0 751800.0 ;
      RECT  864000.0 765600.0 874200.0 779400.0 ;
      RECT  864000.0 793200.0 874200.0 779400.0 ;
      RECT  864000.0 793200.0 874200.0 807000.0 ;
      RECT  864000.0 820800.0 874200.0 807000.0 ;
      RECT  864000.0 820800.0 874200.0 834600.0 ;
      RECT  864000.0 848400.0 874200.0 834600.0 ;
      RECT  864000.0 848400.0 874200.0 862200.0 ;
      RECT  864000.0 876000.0 874200.0 862200.0 ;
      RECT  864000.0 876000.0 874200.0 889800.0 ;
      RECT  864000.0 903600.0 874200.0 889800.0 ;
      RECT  864000.0 903600.0 874200.0 917400.0 ;
      RECT  864000.0 931200.0 874200.0 917400.0 ;
      RECT  864000.0 931200.0 874200.0 945000.0 ;
      RECT  864000.0 958800.0 874200.0 945000.0 ;
      RECT  864000.0 958800.0 874200.0 972600.0 ;
      RECT  864000.0 986400.0 874200.0 972600.0 ;
      RECT  864000.0 986400.0 874200.0 1000200.0 ;
      RECT  864000.0 1014000.0 874200.0 1000200.0 ;
      RECT  864000.0 1014000.0 874200.0 1027800.0 ;
      RECT  864000.0 1041600.0 874200.0 1027800.0 ;
      RECT  864000.0 1041600.0 874200.0 1055400.0 ;
      RECT  864000.0 1069200.0 874200.0 1055400.0 ;
      RECT  864000.0 1069200.0 874200.0 1083000.0 ;
      RECT  864000.0 1096800.0 874200.0 1083000.0 ;
      RECT  864000.0 1096800.0 874200.0 1110600.0 ;
      RECT  864000.0 1124400.0 874200.0 1110600.0 ;
      RECT  864000.0 1124400.0 874200.0 1138200.0 ;
      RECT  864000.0 1152000.0 874200.0 1138200.0 ;
      RECT  864000.0 1152000.0 874200.0 1165800.0 ;
      RECT  864000.0 1179600.0 874200.0 1165800.0 ;
      RECT  864000.0 1179600.0 874200.0 1193400.0 ;
      RECT  864000.0 1207200.0 874200.0 1193400.0 ;
      RECT  864000.0 1207200.0 874200.0 1221000.0 ;
      RECT  864000.0 1234800.0 874200.0 1221000.0 ;
      RECT  864000.0 1234800.0 874200.0 1248600.0 ;
      RECT  864000.0 1262400.0 874200.0 1248600.0 ;
      RECT  864000.0 1262400.0 874200.0 1276200.0 ;
      RECT  864000.0 1290000.0 874200.0 1276200.0 ;
      RECT  864000.0 1290000.0 874200.0 1303800.0 ;
      RECT  864000.0 1317600.0 874200.0 1303800.0 ;
      RECT  864000.0 1317600.0 874200.0 1331400.0 ;
      RECT  864000.0 1345200.0 874200.0 1331400.0 ;
      RECT  864000.0 1345200.0 874200.0 1359000.0 ;
      RECT  864000.0 1372800.0 874200.0 1359000.0 ;
      RECT  864000.0 1372800.0 874200.0 1386600.0 ;
      RECT  864000.0 1400400.0 874200.0 1386600.0 ;
      RECT  864000.0 1400400.0 874200.0 1414200.0 ;
      RECT  864000.0 1428000.0 874200.0 1414200.0 ;
      RECT  864000.0 1428000.0 874200.0 1441800.0 ;
      RECT  864000.0 1455600.0 874200.0 1441800.0 ;
      RECT  864000.0 1455600.0 874200.0 1469400.0 ;
      RECT  864000.0 1483200.0 874200.0 1469400.0 ;
      RECT  864000.0 1483200.0 874200.0 1497000.0 ;
      RECT  864000.0 1510800.0 874200.0 1497000.0 ;
      RECT  864000.0 1510800.0 874200.0 1524600.0 ;
      RECT  864000.0 1538400.0 874200.0 1524600.0 ;
      RECT  864000.0 1538400.0 874200.0 1552200.0 ;
      RECT  864000.0 1566000.0 874200.0 1552200.0 ;
      RECT  864000.0 1566000.0 874200.0 1579800.0 ;
      RECT  864000.0 1593600.0 874200.0 1579800.0 ;
      RECT  864000.0 1593600.0 874200.0 1607400.0 ;
      RECT  864000.0 1621200.0 874200.0 1607400.0 ;
      RECT  864000.0 1621200.0 874200.0 1635000.0 ;
      RECT  864000.0 1648800.0 874200.0 1635000.0 ;
      RECT  864000.0 1648800.0 874200.0 1662600.0 ;
      RECT  864000.0 1676400.0 874200.0 1662600.0 ;
      RECT  864000.0 1676400.0 874200.0 1690200.0 ;
      RECT  864000.0 1704000.0 874200.0 1690200.0 ;
      RECT  864000.0 1704000.0 874200.0 1717800.0 ;
      RECT  864000.0 1731600.0 874200.0 1717800.0 ;
      RECT  864000.0 1731600.0 874200.0 1745400.0 ;
      RECT  864000.0 1759200.0 874200.0 1745400.0 ;
      RECT  864000.0 1759200.0 874200.0 1773000.0 ;
      RECT  864000.0 1786800.0 874200.0 1773000.0 ;
      RECT  864000.0 1786800.0 874200.0 1800600.0 ;
      RECT  864000.0 1814400.0 874200.0 1800600.0 ;
      RECT  864000.0 1814400.0 874200.0 1828200.0 ;
      RECT  864000.0 1842000.0 874200.0 1828200.0 ;
      RECT  864000.0 1842000.0 874200.0 1855800.0 ;
      RECT  864000.0 1869600.0 874200.0 1855800.0 ;
      RECT  864000.0 1869600.0 874200.0 1883400.0 ;
      RECT  864000.0 1897200.0 874200.0 1883400.0 ;
      RECT  864000.0 1897200.0 874200.0 1911000.0 ;
      RECT  864000.0 1924800.0 874200.0 1911000.0 ;
      RECT  864000.0 1924800.0 874200.0 1938600.0 ;
      RECT  864000.0 1952400.0 874200.0 1938600.0 ;
      RECT  864000.0 1952400.0 874200.0 1966200.0 ;
      RECT  864000.0 1980000.0 874200.0 1966200.0 ;
      RECT  864000.0 1980000.0 874200.0 1993800.0 ;
      RECT  864000.0 2007600.0 874200.0 1993800.0 ;
      RECT  864000.0 2007600.0 874200.0 2021400.0 ;
      RECT  864000.0 2035200.0 874200.0 2021400.0 ;
      RECT  864000.0 2035200.0 874200.0 2049000.0 ;
      RECT  864000.0 2062800.0 874200.0 2049000.0 ;
      RECT  864000.0 2062800.0 874200.0 2076600.0 ;
      RECT  864000.0 2090400.0 874200.0 2076600.0 ;
      RECT  864000.0 2090400.0 874200.0 2104200.0 ;
      RECT  864000.0 2118000.0 874200.0 2104200.0 ;
      RECT  864000.0 2118000.0 874200.0 2131800.0 ;
      RECT  864000.0 2145600.0 874200.0 2131800.0 ;
      RECT  874200.0 379200.0 884400.0 393000.0 ;
      RECT  874200.0 406800.0 884400.0 393000.0 ;
      RECT  874200.0 406800.0 884400.0 420600.0 ;
      RECT  874200.0 434400.0 884400.0 420600.0 ;
      RECT  874200.0 434400.0 884400.0 448200.0 ;
      RECT  874200.0 462000.0 884400.0 448200.0 ;
      RECT  874200.0 462000.0 884400.0 475800.0 ;
      RECT  874200.0 489600.0 884400.0 475800.0 ;
      RECT  874200.0 489600.0 884400.0 503400.0 ;
      RECT  874200.0 517200.0 884400.0 503400.0 ;
      RECT  874200.0 517200.0 884400.0 531000.0 ;
      RECT  874200.0 544800.0 884400.0 531000.0 ;
      RECT  874200.0 544800.0 884400.0 558600.0 ;
      RECT  874200.0 572400.0 884400.0 558600.0 ;
      RECT  874200.0 572400.0 884400.0 586200.0 ;
      RECT  874200.0 600000.0 884400.0 586200.0 ;
      RECT  874200.0 600000.0 884400.0 613800.0 ;
      RECT  874200.0 627600.0 884400.0 613800.0 ;
      RECT  874200.0 627600.0 884400.0 641400.0 ;
      RECT  874200.0 655200.0 884400.0 641400.0 ;
      RECT  874200.0 655200.0 884400.0 669000.0 ;
      RECT  874200.0 682800.0 884400.0 669000.0 ;
      RECT  874200.0 682800.0 884400.0 696600.0 ;
      RECT  874200.0 710400.0 884400.0 696600.0 ;
      RECT  874200.0 710400.0 884400.0 724200.0 ;
      RECT  874200.0 738000.0 884400.0 724200.0 ;
      RECT  874200.0 738000.0 884400.0 751800.0 ;
      RECT  874200.0 765600.0 884400.0 751800.0 ;
      RECT  874200.0 765600.0 884400.0 779400.0 ;
      RECT  874200.0 793200.0 884400.0 779400.0 ;
      RECT  874200.0 793200.0 884400.0 807000.0 ;
      RECT  874200.0 820800.0 884400.0 807000.0 ;
      RECT  874200.0 820800.0 884400.0 834600.0 ;
      RECT  874200.0 848400.0 884400.0 834600.0 ;
      RECT  874200.0 848400.0 884400.0 862200.0 ;
      RECT  874200.0 876000.0 884400.0 862200.0 ;
      RECT  874200.0 876000.0 884400.0 889800.0 ;
      RECT  874200.0 903600.0 884400.0 889800.0 ;
      RECT  874200.0 903600.0 884400.0 917400.0 ;
      RECT  874200.0 931200.0 884400.0 917400.0 ;
      RECT  874200.0 931200.0 884400.0 945000.0 ;
      RECT  874200.0 958800.0 884400.0 945000.0 ;
      RECT  874200.0 958800.0 884400.0 972600.0 ;
      RECT  874200.0 986400.0 884400.0 972600.0 ;
      RECT  874200.0 986400.0 884400.0 1000200.0 ;
      RECT  874200.0 1014000.0 884400.0 1000200.0 ;
      RECT  874200.0 1014000.0 884400.0 1027800.0 ;
      RECT  874200.0 1041600.0 884400.0 1027800.0 ;
      RECT  874200.0 1041600.0 884400.0 1055400.0 ;
      RECT  874200.0 1069200.0 884400.0 1055400.0 ;
      RECT  874200.0 1069200.0 884400.0 1083000.0 ;
      RECT  874200.0 1096800.0 884400.0 1083000.0 ;
      RECT  874200.0 1096800.0 884400.0 1110600.0 ;
      RECT  874200.0 1124400.0 884400.0 1110600.0 ;
      RECT  874200.0 1124400.0 884400.0 1138200.0 ;
      RECT  874200.0 1152000.0 884400.0 1138200.0 ;
      RECT  874200.0 1152000.0 884400.0 1165800.0 ;
      RECT  874200.0 1179600.0 884400.0 1165800.0 ;
      RECT  874200.0 1179600.0 884400.0 1193400.0 ;
      RECT  874200.0 1207200.0 884400.0 1193400.0 ;
      RECT  874200.0 1207200.0 884400.0 1221000.0 ;
      RECT  874200.0 1234800.0 884400.0 1221000.0 ;
      RECT  874200.0 1234800.0 884400.0 1248600.0 ;
      RECT  874200.0 1262400.0 884400.0 1248600.0 ;
      RECT  874200.0 1262400.0 884400.0 1276200.0 ;
      RECT  874200.0 1290000.0 884400.0 1276200.0 ;
      RECT  874200.0 1290000.0 884400.0 1303800.0 ;
      RECT  874200.0 1317600.0 884400.0 1303800.0 ;
      RECT  874200.0 1317600.0 884400.0 1331400.0 ;
      RECT  874200.0 1345200.0 884400.0 1331400.0 ;
      RECT  874200.0 1345200.0 884400.0 1359000.0 ;
      RECT  874200.0 1372800.0 884400.0 1359000.0 ;
      RECT  874200.0 1372800.0 884400.0 1386600.0 ;
      RECT  874200.0 1400400.0 884400.0 1386600.0 ;
      RECT  874200.0 1400400.0 884400.0 1414200.0 ;
      RECT  874200.0 1428000.0 884400.0 1414200.0 ;
      RECT  874200.0 1428000.0 884400.0 1441800.0 ;
      RECT  874200.0 1455600.0 884400.0 1441800.0 ;
      RECT  874200.0 1455600.0 884400.0 1469400.0 ;
      RECT  874200.0 1483200.0 884400.0 1469400.0 ;
      RECT  874200.0 1483200.0 884400.0 1497000.0 ;
      RECT  874200.0 1510800.0 884400.0 1497000.0 ;
      RECT  874200.0 1510800.0 884400.0 1524600.0 ;
      RECT  874200.0 1538400.0 884400.0 1524600.0 ;
      RECT  874200.0 1538400.0 884400.0 1552200.0 ;
      RECT  874200.0 1566000.0 884400.0 1552200.0 ;
      RECT  874200.0 1566000.0 884400.0 1579800.0 ;
      RECT  874200.0 1593600.0 884400.0 1579800.0 ;
      RECT  874200.0 1593600.0 884400.0 1607400.0 ;
      RECT  874200.0 1621200.0 884400.0 1607400.0 ;
      RECT  874200.0 1621200.0 884400.0 1635000.0 ;
      RECT  874200.0 1648800.0 884400.0 1635000.0 ;
      RECT  874200.0 1648800.0 884400.0 1662600.0 ;
      RECT  874200.0 1676400.0 884400.0 1662600.0 ;
      RECT  874200.0 1676400.0 884400.0 1690200.0 ;
      RECT  874200.0 1704000.0 884400.0 1690200.0 ;
      RECT  874200.0 1704000.0 884400.0 1717800.0 ;
      RECT  874200.0 1731600.0 884400.0 1717800.0 ;
      RECT  874200.0 1731600.0 884400.0 1745400.0 ;
      RECT  874200.0 1759200.0 884400.0 1745400.0 ;
      RECT  874200.0 1759200.0 884400.0 1773000.0 ;
      RECT  874200.0 1786800.0 884400.0 1773000.0 ;
      RECT  874200.0 1786800.0 884400.0 1800600.0 ;
      RECT  874200.0 1814400.0 884400.0 1800600.0 ;
      RECT  874200.0 1814400.0 884400.0 1828200.0 ;
      RECT  874200.0 1842000.0 884400.0 1828200.0 ;
      RECT  874200.0 1842000.0 884400.0 1855800.0 ;
      RECT  874200.0 1869600.0 884400.0 1855800.0 ;
      RECT  874200.0 1869600.0 884400.0 1883400.0 ;
      RECT  874200.0 1897200.0 884400.0 1883400.0 ;
      RECT  874200.0 1897200.0 884400.0 1911000.0 ;
      RECT  874200.0 1924800.0 884400.0 1911000.0 ;
      RECT  874200.0 1924800.0 884400.0 1938600.0 ;
      RECT  874200.0 1952400.0 884400.0 1938600.0 ;
      RECT  874200.0 1952400.0 884400.0 1966200.0 ;
      RECT  874200.0 1980000.0 884400.0 1966200.0 ;
      RECT  874200.0 1980000.0 884400.0 1993800.0 ;
      RECT  874200.0 2007600.0 884400.0 1993800.0 ;
      RECT  874200.0 2007600.0 884400.0 2021400.0 ;
      RECT  874200.0 2035200.0 884400.0 2021400.0 ;
      RECT  874200.0 2035200.0 884400.0 2049000.0 ;
      RECT  874200.0 2062800.0 884400.0 2049000.0 ;
      RECT  874200.0 2062800.0 884400.0 2076600.0 ;
      RECT  874200.0 2090400.0 884400.0 2076600.0 ;
      RECT  874200.0 2090400.0 884400.0 2104200.0 ;
      RECT  874200.0 2118000.0 884400.0 2104200.0 ;
      RECT  874200.0 2118000.0 884400.0 2131800.0 ;
      RECT  874200.0 2145600.0 884400.0 2131800.0 ;
      RECT  884400.0 379200.0 894600.0 393000.0 ;
      RECT  884400.0 406800.0 894600.0 393000.0 ;
      RECT  884400.0 406800.0 894600.0 420600.0 ;
      RECT  884400.0 434400.0 894600.0 420600.0 ;
      RECT  884400.0 434400.0 894600.0 448200.0 ;
      RECT  884400.0 462000.0 894600.0 448200.0 ;
      RECT  884400.0 462000.0 894600.0 475800.0 ;
      RECT  884400.0 489600.0 894600.0 475800.0 ;
      RECT  884400.0 489600.0 894600.0 503400.0 ;
      RECT  884400.0 517200.0 894600.0 503400.0 ;
      RECT  884400.0 517200.0 894600.0 531000.0 ;
      RECT  884400.0 544800.0 894600.0 531000.0 ;
      RECT  884400.0 544800.0 894600.0 558600.0 ;
      RECT  884400.0 572400.0 894600.0 558600.0 ;
      RECT  884400.0 572400.0 894600.0 586200.0 ;
      RECT  884400.0 600000.0 894600.0 586200.0 ;
      RECT  884400.0 600000.0 894600.0 613800.0 ;
      RECT  884400.0 627600.0 894600.0 613800.0 ;
      RECT  884400.0 627600.0 894600.0 641400.0 ;
      RECT  884400.0 655200.0 894600.0 641400.0 ;
      RECT  884400.0 655200.0 894600.0 669000.0 ;
      RECT  884400.0 682800.0 894600.0 669000.0 ;
      RECT  884400.0 682800.0 894600.0 696600.0 ;
      RECT  884400.0 710400.0 894600.0 696600.0 ;
      RECT  884400.0 710400.0 894600.0 724200.0 ;
      RECT  884400.0 738000.0 894600.0 724200.0 ;
      RECT  884400.0 738000.0 894600.0 751800.0 ;
      RECT  884400.0 765600.0 894600.0 751800.0 ;
      RECT  884400.0 765600.0 894600.0 779400.0 ;
      RECT  884400.0 793200.0 894600.0 779400.0 ;
      RECT  884400.0 793200.0 894600.0 807000.0 ;
      RECT  884400.0 820800.0 894600.0 807000.0 ;
      RECT  884400.0 820800.0 894600.0 834600.0 ;
      RECT  884400.0 848400.0 894600.0 834600.0 ;
      RECT  884400.0 848400.0 894600.0 862200.0 ;
      RECT  884400.0 876000.0 894600.0 862200.0 ;
      RECT  884400.0 876000.0 894600.0 889800.0 ;
      RECT  884400.0 903600.0 894600.0 889800.0 ;
      RECT  884400.0 903600.0 894600.0 917400.0 ;
      RECT  884400.0 931200.0 894600.0 917400.0 ;
      RECT  884400.0 931200.0 894600.0 945000.0 ;
      RECT  884400.0 958800.0 894600.0 945000.0 ;
      RECT  884400.0 958800.0 894600.0 972600.0 ;
      RECT  884400.0 986400.0 894600.0 972600.0 ;
      RECT  884400.0 986400.0 894600.0 1000200.0 ;
      RECT  884400.0 1014000.0 894600.0 1000200.0 ;
      RECT  884400.0 1014000.0 894600.0 1027800.0 ;
      RECT  884400.0 1041600.0 894600.0 1027800.0 ;
      RECT  884400.0 1041600.0 894600.0 1055400.0 ;
      RECT  884400.0 1069200.0 894600.0 1055400.0 ;
      RECT  884400.0 1069200.0 894600.0 1083000.0 ;
      RECT  884400.0 1096800.0 894600.0 1083000.0 ;
      RECT  884400.0 1096800.0 894600.0 1110600.0 ;
      RECT  884400.0 1124400.0 894600.0 1110600.0 ;
      RECT  884400.0 1124400.0 894600.0 1138200.0 ;
      RECT  884400.0 1152000.0 894600.0 1138200.0 ;
      RECT  884400.0 1152000.0 894600.0 1165800.0 ;
      RECT  884400.0 1179600.0 894600.0 1165800.0 ;
      RECT  884400.0 1179600.0 894600.0 1193400.0 ;
      RECT  884400.0 1207200.0 894600.0 1193400.0 ;
      RECT  884400.0 1207200.0 894600.0 1221000.0 ;
      RECT  884400.0 1234800.0 894600.0 1221000.0 ;
      RECT  884400.0 1234800.0 894600.0 1248600.0 ;
      RECT  884400.0 1262400.0 894600.0 1248600.0 ;
      RECT  884400.0 1262400.0 894600.0 1276200.0 ;
      RECT  884400.0 1290000.0 894600.0 1276200.0 ;
      RECT  884400.0 1290000.0 894600.0 1303800.0 ;
      RECT  884400.0 1317600.0 894600.0 1303800.0 ;
      RECT  884400.0 1317600.0 894600.0 1331400.0 ;
      RECT  884400.0 1345200.0 894600.0 1331400.0 ;
      RECT  884400.0 1345200.0 894600.0 1359000.0 ;
      RECT  884400.0 1372800.0 894600.0 1359000.0 ;
      RECT  884400.0 1372800.0 894600.0 1386600.0 ;
      RECT  884400.0 1400400.0 894600.0 1386600.0 ;
      RECT  884400.0 1400400.0 894600.0 1414200.0 ;
      RECT  884400.0 1428000.0 894600.0 1414200.0 ;
      RECT  884400.0 1428000.0 894600.0 1441800.0 ;
      RECT  884400.0 1455600.0 894600.0 1441800.0 ;
      RECT  884400.0 1455600.0 894600.0 1469400.0 ;
      RECT  884400.0 1483200.0 894600.0 1469400.0 ;
      RECT  884400.0 1483200.0 894600.0 1497000.0 ;
      RECT  884400.0 1510800.0 894600.0 1497000.0 ;
      RECT  884400.0 1510800.0 894600.0 1524600.0 ;
      RECT  884400.0 1538400.0 894600.0 1524600.0 ;
      RECT  884400.0 1538400.0 894600.0 1552200.0 ;
      RECT  884400.0 1566000.0 894600.0 1552200.0 ;
      RECT  884400.0 1566000.0 894600.0 1579800.0 ;
      RECT  884400.0 1593600.0 894600.0 1579800.0 ;
      RECT  884400.0 1593600.0 894600.0 1607400.0 ;
      RECT  884400.0 1621200.0 894600.0 1607400.0 ;
      RECT  884400.0 1621200.0 894600.0 1635000.0 ;
      RECT  884400.0 1648800.0 894600.0 1635000.0 ;
      RECT  884400.0 1648800.0 894600.0 1662600.0 ;
      RECT  884400.0 1676400.0 894600.0 1662600.0 ;
      RECT  884400.0 1676400.0 894600.0 1690200.0 ;
      RECT  884400.0 1704000.0 894600.0 1690200.0 ;
      RECT  884400.0 1704000.0 894600.0 1717800.0 ;
      RECT  884400.0 1731600.0 894600.0 1717800.0 ;
      RECT  884400.0 1731600.0 894600.0 1745400.0 ;
      RECT  884400.0 1759200.0 894600.0 1745400.0 ;
      RECT  884400.0 1759200.0 894600.0 1773000.0 ;
      RECT  884400.0 1786800.0 894600.0 1773000.0 ;
      RECT  884400.0 1786800.0 894600.0 1800600.0 ;
      RECT  884400.0 1814400.0 894600.0 1800600.0 ;
      RECT  884400.0 1814400.0 894600.0 1828200.0 ;
      RECT  884400.0 1842000.0 894600.0 1828200.0 ;
      RECT  884400.0 1842000.0 894600.0 1855800.0 ;
      RECT  884400.0 1869600.0 894600.0 1855800.0 ;
      RECT  884400.0 1869600.0 894600.0 1883400.0 ;
      RECT  884400.0 1897200.0 894600.0 1883400.0 ;
      RECT  884400.0 1897200.0 894600.0 1911000.0 ;
      RECT  884400.0 1924800.0 894600.0 1911000.0 ;
      RECT  884400.0 1924800.0 894600.0 1938600.0 ;
      RECT  884400.0 1952400.0 894600.0 1938600.0 ;
      RECT  884400.0 1952400.0 894600.0 1966200.0 ;
      RECT  884400.0 1980000.0 894600.0 1966200.0 ;
      RECT  884400.0 1980000.0 894600.0 1993800.0 ;
      RECT  884400.0 2007600.0 894600.0 1993800.0 ;
      RECT  884400.0 2007600.0 894600.0 2021400.0 ;
      RECT  884400.0 2035200.0 894600.0 2021400.0 ;
      RECT  884400.0 2035200.0 894600.0 2049000.0 ;
      RECT  884400.0 2062800.0 894600.0 2049000.0 ;
      RECT  884400.0 2062800.0 894600.0 2076600.0 ;
      RECT  884400.0 2090400.0 894600.0 2076600.0 ;
      RECT  884400.0 2090400.0 894600.0 2104200.0 ;
      RECT  884400.0 2118000.0 894600.0 2104200.0 ;
      RECT  884400.0 2118000.0 894600.0 2131800.0 ;
      RECT  884400.0 2145600.0 894600.0 2131800.0 ;
      RECT  894600.0 379200.0 904800.0 393000.0 ;
      RECT  894600.0 406800.0 904800.0 393000.0 ;
      RECT  894600.0 406800.0 904800.0 420600.0 ;
      RECT  894600.0 434400.0 904800.0 420600.0 ;
      RECT  894600.0 434400.0 904800.0 448200.0 ;
      RECT  894600.0 462000.0 904800.0 448200.0 ;
      RECT  894600.0 462000.0 904800.0 475800.0 ;
      RECT  894600.0 489600.0 904800.0 475800.0 ;
      RECT  894600.0 489600.0 904800.0 503400.0 ;
      RECT  894600.0 517200.0 904800.0 503400.0 ;
      RECT  894600.0 517200.0 904800.0 531000.0 ;
      RECT  894600.0 544800.0 904800.0 531000.0 ;
      RECT  894600.0 544800.0 904800.0 558600.0 ;
      RECT  894600.0 572400.0 904800.0 558600.0 ;
      RECT  894600.0 572400.0 904800.0 586200.0 ;
      RECT  894600.0 600000.0 904800.0 586200.0 ;
      RECT  894600.0 600000.0 904800.0 613800.0 ;
      RECT  894600.0 627600.0 904800.0 613800.0 ;
      RECT  894600.0 627600.0 904800.0 641400.0 ;
      RECT  894600.0 655200.0 904800.0 641400.0 ;
      RECT  894600.0 655200.0 904800.0 669000.0 ;
      RECT  894600.0 682800.0 904800.0 669000.0 ;
      RECT  894600.0 682800.0 904800.0 696600.0 ;
      RECT  894600.0 710400.0 904800.0 696600.0 ;
      RECT  894600.0 710400.0 904800.0 724200.0 ;
      RECT  894600.0 738000.0 904800.0 724200.0 ;
      RECT  894600.0 738000.0 904800.0 751800.0 ;
      RECT  894600.0 765600.0 904800.0 751800.0 ;
      RECT  894600.0 765600.0 904800.0 779400.0 ;
      RECT  894600.0 793200.0 904800.0 779400.0 ;
      RECT  894600.0 793200.0 904800.0 807000.0 ;
      RECT  894600.0 820800.0 904800.0 807000.0 ;
      RECT  894600.0 820800.0 904800.0 834600.0 ;
      RECT  894600.0 848400.0 904800.0 834600.0 ;
      RECT  894600.0 848400.0 904800.0 862200.0 ;
      RECT  894600.0 876000.0 904800.0 862200.0 ;
      RECT  894600.0 876000.0 904800.0 889800.0 ;
      RECT  894600.0 903600.0 904800.0 889800.0 ;
      RECT  894600.0 903600.0 904800.0 917400.0 ;
      RECT  894600.0 931200.0 904800.0 917400.0 ;
      RECT  894600.0 931200.0 904800.0 945000.0 ;
      RECT  894600.0 958800.0 904800.0 945000.0 ;
      RECT  894600.0 958800.0 904800.0 972600.0 ;
      RECT  894600.0 986400.0 904800.0 972600.0 ;
      RECT  894600.0 986400.0 904800.0 1000200.0 ;
      RECT  894600.0 1014000.0 904800.0 1000200.0 ;
      RECT  894600.0 1014000.0 904800.0 1027800.0 ;
      RECT  894600.0 1041600.0 904800.0 1027800.0 ;
      RECT  894600.0 1041600.0 904800.0 1055400.0 ;
      RECT  894600.0 1069200.0 904800.0 1055400.0 ;
      RECT  894600.0 1069200.0 904800.0 1083000.0 ;
      RECT  894600.0 1096800.0 904800.0 1083000.0 ;
      RECT  894600.0 1096800.0 904800.0 1110600.0 ;
      RECT  894600.0 1124400.0 904800.0 1110600.0 ;
      RECT  894600.0 1124400.0 904800.0 1138200.0 ;
      RECT  894600.0 1152000.0 904800.0 1138200.0 ;
      RECT  894600.0 1152000.0 904800.0 1165800.0 ;
      RECT  894600.0 1179600.0 904800.0 1165800.0 ;
      RECT  894600.0 1179600.0 904800.0 1193400.0 ;
      RECT  894600.0 1207200.0 904800.0 1193400.0 ;
      RECT  894600.0 1207200.0 904800.0 1221000.0 ;
      RECT  894600.0 1234800.0 904800.0 1221000.0 ;
      RECT  894600.0 1234800.0 904800.0 1248600.0 ;
      RECT  894600.0 1262400.0 904800.0 1248600.0 ;
      RECT  894600.0 1262400.0 904800.0 1276200.0 ;
      RECT  894600.0 1290000.0 904800.0 1276200.0 ;
      RECT  894600.0 1290000.0 904800.0 1303800.0 ;
      RECT  894600.0 1317600.0 904800.0 1303800.0 ;
      RECT  894600.0 1317600.0 904800.0 1331400.0 ;
      RECT  894600.0 1345200.0 904800.0 1331400.0 ;
      RECT  894600.0 1345200.0 904800.0 1359000.0 ;
      RECT  894600.0 1372800.0 904800.0 1359000.0 ;
      RECT  894600.0 1372800.0 904800.0 1386600.0 ;
      RECT  894600.0 1400400.0 904800.0 1386600.0 ;
      RECT  894600.0 1400400.0 904800.0 1414200.0 ;
      RECT  894600.0 1428000.0 904800.0 1414200.0 ;
      RECT  894600.0 1428000.0 904800.0 1441800.0 ;
      RECT  894600.0 1455600.0 904800.0 1441800.0 ;
      RECT  894600.0 1455600.0 904800.0 1469400.0 ;
      RECT  894600.0 1483200.0 904800.0 1469400.0 ;
      RECT  894600.0 1483200.0 904800.0 1497000.0 ;
      RECT  894600.0 1510800.0 904800.0 1497000.0 ;
      RECT  894600.0 1510800.0 904800.0 1524600.0 ;
      RECT  894600.0 1538400.0 904800.0 1524600.0 ;
      RECT  894600.0 1538400.0 904800.0 1552200.0 ;
      RECT  894600.0 1566000.0 904800.0 1552200.0 ;
      RECT  894600.0 1566000.0 904800.0 1579800.0 ;
      RECT  894600.0 1593600.0 904800.0 1579800.0 ;
      RECT  894600.0 1593600.0 904800.0 1607400.0 ;
      RECT  894600.0 1621200.0 904800.0 1607400.0 ;
      RECT  894600.0 1621200.0 904800.0 1635000.0 ;
      RECT  894600.0 1648800.0 904800.0 1635000.0 ;
      RECT  894600.0 1648800.0 904800.0 1662600.0 ;
      RECT  894600.0 1676400.0 904800.0 1662600.0 ;
      RECT  894600.0 1676400.0 904800.0 1690200.0 ;
      RECT  894600.0 1704000.0 904800.0 1690200.0 ;
      RECT  894600.0 1704000.0 904800.0 1717800.0 ;
      RECT  894600.0 1731600.0 904800.0 1717800.0 ;
      RECT  894600.0 1731600.0 904800.0 1745400.0 ;
      RECT  894600.0 1759200.0 904800.0 1745400.0 ;
      RECT  894600.0 1759200.0 904800.0 1773000.0 ;
      RECT  894600.0 1786800.0 904800.0 1773000.0 ;
      RECT  894600.0 1786800.0 904800.0 1800600.0 ;
      RECT  894600.0 1814400.0 904800.0 1800600.0 ;
      RECT  894600.0 1814400.0 904800.0 1828200.0 ;
      RECT  894600.0 1842000.0 904800.0 1828200.0 ;
      RECT  894600.0 1842000.0 904800.0 1855800.0 ;
      RECT  894600.0 1869600.0 904800.0 1855800.0 ;
      RECT  894600.0 1869600.0 904800.0 1883400.0 ;
      RECT  894600.0 1897200.0 904800.0 1883400.0 ;
      RECT  894600.0 1897200.0 904800.0 1911000.0 ;
      RECT  894600.0 1924800.0 904800.0 1911000.0 ;
      RECT  894600.0 1924800.0 904800.0 1938600.0 ;
      RECT  894600.0 1952400.0 904800.0 1938600.0 ;
      RECT  894600.0 1952400.0 904800.0 1966200.0 ;
      RECT  894600.0 1980000.0 904800.0 1966200.0 ;
      RECT  894600.0 1980000.0 904800.0 1993800.0 ;
      RECT  894600.0 2007600.0 904800.0 1993800.0 ;
      RECT  894600.0 2007600.0 904800.0 2021400.0 ;
      RECT  894600.0 2035200.0 904800.0 2021400.0 ;
      RECT  894600.0 2035200.0 904800.0 2049000.0 ;
      RECT  894600.0 2062800.0 904800.0 2049000.0 ;
      RECT  894600.0 2062800.0 904800.0 2076600.0 ;
      RECT  894600.0 2090400.0 904800.0 2076600.0 ;
      RECT  894600.0 2090400.0 904800.0 2104200.0 ;
      RECT  894600.0 2118000.0 904800.0 2104200.0 ;
      RECT  894600.0 2118000.0 904800.0 2131800.0 ;
      RECT  894600.0 2145600.0 904800.0 2131800.0 ;
      RECT  904800.0 379200.0 915000.0 393000.0 ;
      RECT  904800.0 406800.0 915000.0 393000.0 ;
      RECT  904800.0 406800.0 915000.0 420600.0 ;
      RECT  904800.0 434400.0 915000.0 420600.0 ;
      RECT  904800.0 434400.0 915000.0 448200.0 ;
      RECT  904800.0 462000.0 915000.0 448200.0 ;
      RECT  904800.0 462000.0 915000.0 475800.0 ;
      RECT  904800.0 489600.0 915000.0 475800.0 ;
      RECT  904800.0 489600.0 915000.0 503400.0 ;
      RECT  904800.0 517200.0 915000.0 503400.0 ;
      RECT  904800.0 517200.0 915000.0 531000.0 ;
      RECT  904800.0 544800.0 915000.0 531000.0 ;
      RECT  904800.0 544800.0 915000.0 558600.0 ;
      RECT  904800.0 572400.0 915000.0 558600.0 ;
      RECT  904800.0 572400.0 915000.0 586200.0 ;
      RECT  904800.0 600000.0 915000.0 586200.0 ;
      RECT  904800.0 600000.0 915000.0 613800.0 ;
      RECT  904800.0 627600.0 915000.0 613800.0 ;
      RECT  904800.0 627600.0 915000.0 641400.0 ;
      RECT  904800.0 655200.0 915000.0 641400.0 ;
      RECT  904800.0 655200.0 915000.0 669000.0 ;
      RECT  904800.0 682800.0 915000.0 669000.0 ;
      RECT  904800.0 682800.0 915000.0 696600.0 ;
      RECT  904800.0 710400.0 915000.0 696600.0 ;
      RECT  904800.0 710400.0 915000.0 724200.0 ;
      RECT  904800.0 738000.0 915000.0 724200.0 ;
      RECT  904800.0 738000.0 915000.0 751800.0 ;
      RECT  904800.0 765600.0 915000.0 751800.0 ;
      RECT  904800.0 765600.0 915000.0 779400.0 ;
      RECT  904800.0 793200.0 915000.0 779400.0 ;
      RECT  904800.0 793200.0 915000.0 807000.0 ;
      RECT  904800.0 820800.0 915000.0 807000.0 ;
      RECT  904800.0 820800.0 915000.0 834600.0 ;
      RECT  904800.0 848400.0 915000.0 834600.0 ;
      RECT  904800.0 848400.0 915000.0 862200.0 ;
      RECT  904800.0 876000.0 915000.0 862200.0 ;
      RECT  904800.0 876000.0 915000.0 889800.0 ;
      RECT  904800.0 903600.0 915000.0 889800.0 ;
      RECT  904800.0 903600.0 915000.0 917400.0 ;
      RECT  904800.0 931200.0 915000.0 917400.0 ;
      RECT  904800.0 931200.0 915000.0 945000.0 ;
      RECT  904800.0 958800.0 915000.0 945000.0 ;
      RECT  904800.0 958800.0 915000.0 972600.0 ;
      RECT  904800.0 986400.0 915000.0 972600.0 ;
      RECT  904800.0 986400.0 915000.0 1000200.0 ;
      RECT  904800.0 1014000.0 915000.0 1000200.0 ;
      RECT  904800.0 1014000.0 915000.0 1027800.0 ;
      RECT  904800.0 1041600.0 915000.0 1027800.0 ;
      RECT  904800.0 1041600.0 915000.0 1055400.0 ;
      RECT  904800.0 1069200.0 915000.0 1055400.0 ;
      RECT  904800.0 1069200.0 915000.0 1083000.0 ;
      RECT  904800.0 1096800.0 915000.0 1083000.0 ;
      RECT  904800.0 1096800.0 915000.0 1110600.0 ;
      RECT  904800.0 1124400.0 915000.0 1110600.0 ;
      RECT  904800.0 1124400.0 915000.0 1138200.0 ;
      RECT  904800.0 1152000.0 915000.0 1138200.0 ;
      RECT  904800.0 1152000.0 915000.0 1165800.0 ;
      RECT  904800.0 1179600.0 915000.0 1165800.0 ;
      RECT  904800.0 1179600.0 915000.0 1193400.0 ;
      RECT  904800.0 1207200.0 915000.0 1193400.0 ;
      RECT  904800.0 1207200.0 915000.0 1221000.0 ;
      RECT  904800.0 1234800.0 915000.0 1221000.0 ;
      RECT  904800.0 1234800.0 915000.0 1248600.0 ;
      RECT  904800.0 1262400.0 915000.0 1248600.0 ;
      RECT  904800.0 1262400.0 915000.0 1276200.0 ;
      RECT  904800.0 1290000.0 915000.0 1276200.0 ;
      RECT  904800.0 1290000.0 915000.0 1303800.0 ;
      RECT  904800.0 1317600.0 915000.0 1303800.0 ;
      RECT  904800.0 1317600.0 915000.0 1331400.0 ;
      RECT  904800.0 1345200.0 915000.0 1331400.0 ;
      RECT  904800.0 1345200.0 915000.0 1359000.0 ;
      RECT  904800.0 1372800.0 915000.0 1359000.0 ;
      RECT  904800.0 1372800.0 915000.0 1386600.0 ;
      RECT  904800.0 1400400.0 915000.0 1386600.0 ;
      RECT  904800.0 1400400.0 915000.0 1414200.0 ;
      RECT  904800.0 1428000.0 915000.0 1414200.0 ;
      RECT  904800.0 1428000.0 915000.0 1441800.0 ;
      RECT  904800.0 1455600.0 915000.0 1441800.0 ;
      RECT  904800.0 1455600.0 915000.0 1469400.0 ;
      RECT  904800.0 1483200.0 915000.0 1469400.0 ;
      RECT  904800.0 1483200.0 915000.0 1497000.0 ;
      RECT  904800.0 1510800.0 915000.0 1497000.0 ;
      RECT  904800.0 1510800.0 915000.0 1524600.0 ;
      RECT  904800.0 1538400.0 915000.0 1524600.0 ;
      RECT  904800.0 1538400.0 915000.0 1552200.0 ;
      RECT  904800.0 1566000.0 915000.0 1552200.0 ;
      RECT  904800.0 1566000.0 915000.0 1579800.0 ;
      RECT  904800.0 1593600.0 915000.0 1579800.0 ;
      RECT  904800.0 1593600.0 915000.0 1607400.0 ;
      RECT  904800.0 1621200.0 915000.0 1607400.0 ;
      RECT  904800.0 1621200.0 915000.0 1635000.0 ;
      RECT  904800.0 1648800.0 915000.0 1635000.0 ;
      RECT  904800.0 1648800.0 915000.0 1662600.0 ;
      RECT  904800.0 1676400.0 915000.0 1662600.0 ;
      RECT  904800.0 1676400.0 915000.0 1690200.0 ;
      RECT  904800.0 1704000.0 915000.0 1690200.0 ;
      RECT  904800.0 1704000.0 915000.0 1717800.0 ;
      RECT  904800.0 1731600.0 915000.0 1717800.0 ;
      RECT  904800.0 1731600.0 915000.0 1745400.0 ;
      RECT  904800.0 1759200.0 915000.0 1745400.0 ;
      RECT  904800.0 1759200.0 915000.0 1773000.0 ;
      RECT  904800.0 1786800.0 915000.0 1773000.0 ;
      RECT  904800.0 1786800.0 915000.0 1800600.0 ;
      RECT  904800.0 1814400.0 915000.0 1800600.0 ;
      RECT  904800.0 1814400.0 915000.0 1828200.0 ;
      RECT  904800.0 1842000.0 915000.0 1828200.0 ;
      RECT  904800.0 1842000.0 915000.0 1855800.0 ;
      RECT  904800.0 1869600.0 915000.0 1855800.0 ;
      RECT  904800.0 1869600.0 915000.0 1883400.0 ;
      RECT  904800.0 1897200.0 915000.0 1883400.0 ;
      RECT  904800.0 1897200.0 915000.0 1911000.0 ;
      RECT  904800.0 1924800.0 915000.0 1911000.0 ;
      RECT  904800.0 1924800.0 915000.0 1938600.0 ;
      RECT  904800.0 1952400.0 915000.0 1938600.0 ;
      RECT  904800.0 1952400.0 915000.0 1966200.0 ;
      RECT  904800.0 1980000.0 915000.0 1966200.0 ;
      RECT  904800.0 1980000.0 915000.0 1993800.0 ;
      RECT  904800.0 2007600.0 915000.0 1993800.0 ;
      RECT  904800.0 2007600.0 915000.0 2021400.0 ;
      RECT  904800.0 2035200.0 915000.0 2021400.0 ;
      RECT  904800.0 2035200.0 915000.0 2049000.0 ;
      RECT  904800.0 2062800.0 915000.0 2049000.0 ;
      RECT  904800.0 2062800.0 915000.0 2076600.0 ;
      RECT  904800.0 2090400.0 915000.0 2076600.0 ;
      RECT  904800.0 2090400.0 915000.0 2104200.0 ;
      RECT  904800.0 2118000.0 915000.0 2104200.0 ;
      RECT  904800.0 2118000.0 915000.0 2131800.0 ;
      RECT  904800.0 2145600.0 915000.0 2131800.0 ;
      RECT  915000.0 379200.0 925200.0 393000.0 ;
      RECT  915000.0 406800.0 925200.0 393000.0 ;
      RECT  915000.0 406800.0 925200.0 420600.0 ;
      RECT  915000.0 434400.0 925200.0 420600.0 ;
      RECT  915000.0 434400.0 925200.0 448200.0 ;
      RECT  915000.0 462000.0 925200.0 448200.0 ;
      RECT  915000.0 462000.0 925200.0 475800.0 ;
      RECT  915000.0 489600.0 925200.0 475800.0 ;
      RECT  915000.0 489600.0 925200.0 503400.0 ;
      RECT  915000.0 517200.0 925200.0 503400.0 ;
      RECT  915000.0 517200.0 925200.0 531000.0 ;
      RECT  915000.0 544800.0 925200.0 531000.0 ;
      RECT  915000.0 544800.0 925200.0 558600.0 ;
      RECT  915000.0 572400.0 925200.0 558600.0 ;
      RECT  915000.0 572400.0 925200.0 586200.0 ;
      RECT  915000.0 600000.0 925200.0 586200.0 ;
      RECT  915000.0 600000.0 925200.0 613800.0 ;
      RECT  915000.0 627600.0 925200.0 613800.0 ;
      RECT  915000.0 627600.0 925200.0 641400.0 ;
      RECT  915000.0 655200.0 925200.0 641400.0 ;
      RECT  915000.0 655200.0 925200.0 669000.0 ;
      RECT  915000.0 682800.0 925200.0 669000.0 ;
      RECT  915000.0 682800.0 925200.0 696600.0 ;
      RECT  915000.0 710400.0 925200.0 696600.0 ;
      RECT  915000.0 710400.0 925200.0 724200.0 ;
      RECT  915000.0 738000.0 925200.0 724200.0 ;
      RECT  915000.0 738000.0 925200.0 751800.0 ;
      RECT  915000.0 765600.0 925200.0 751800.0 ;
      RECT  915000.0 765600.0 925200.0 779400.0 ;
      RECT  915000.0 793200.0 925200.0 779400.0 ;
      RECT  915000.0 793200.0 925200.0 807000.0 ;
      RECT  915000.0 820800.0 925200.0 807000.0 ;
      RECT  915000.0 820800.0 925200.0 834600.0 ;
      RECT  915000.0 848400.0 925200.0 834600.0 ;
      RECT  915000.0 848400.0 925200.0 862200.0 ;
      RECT  915000.0 876000.0 925200.0 862200.0 ;
      RECT  915000.0 876000.0 925200.0 889800.0 ;
      RECT  915000.0 903600.0 925200.0 889800.0 ;
      RECT  915000.0 903600.0 925200.0 917400.0 ;
      RECT  915000.0 931200.0 925200.0 917400.0 ;
      RECT  915000.0 931200.0 925200.0 945000.0 ;
      RECT  915000.0 958800.0 925200.0 945000.0 ;
      RECT  915000.0 958800.0 925200.0 972600.0 ;
      RECT  915000.0 986400.0 925200.0 972600.0 ;
      RECT  915000.0 986400.0 925200.0 1000200.0 ;
      RECT  915000.0 1014000.0 925200.0 1000200.0 ;
      RECT  915000.0 1014000.0 925200.0 1027800.0 ;
      RECT  915000.0 1041600.0 925200.0 1027800.0 ;
      RECT  915000.0 1041600.0 925200.0 1055400.0 ;
      RECT  915000.0 1069200.0 925200.0 1055400.0 ;
      RECT  915000.0 1069200.0 925200.0 1083000.0 ;
      RECT  915000.0 1096800.0 925200.0 1083000.0 ;
      RECT  915000.0 1096800.0 925200.0 1110600.0 ;
      RECT  915000.0 1124400.0 925200.0 1110600.0 ;
      RECT  915000.0 1124400.0 925200.0 1138200.0 ;
      RECT  915000.0 1152000.0 925200.0 1138200.0 ;
      RECT  915000.0 1152000.0 925200.0 1165800.0 ;
      RECT  915000.0 1179600.0 925200.0 1165800.0 ;
      RECT  915000.0 1179600.0 925200.0 1193400.0 ;
      RECT  915000.0 1207200.0 925200.0 1193400.0 ;
      RECT  915000.0 1207200.0 925200.0 1221000.0 ;
      RECT  915000.0 1234800.0 925200.0 1221000.0 ;
      RECT  915000.0 1234800.0 925200.0 1248600.0 ;
      RECT  915000.0 1262400.0 925200.0 1248600.0 ;
      RECT  915000.0 1262400.0 925200.0 1276200.0 ;
      RECT  915000.0 1290000.0 925200.0 1276200.0 ;
      RECT  915000.0 1290000.0 925200.0 1303800.0 ;
      RECT  915000.0 1317600.0 925200.0 1303800.0 ;
      RECT  915000.0 1317600.0 925200.0 1331400.0 ;
      RECT  915000.0 1345200.0 925200.0 1331400.0 ;
      RECT  915000.0 1345200.0 925200.0 1359000.0 ;
      RECT  915000.0 1372800.0 925200.0 1359000.0 ;
      RECT  915000.0 1372800.0 925200.0 1386600.0 ;
      RECT  915000.0 1400400.0 925200.0 1386600.0 ;
      RECT  915000.0 1400400.0 925200.0 1414200.0 ;
      RECT  915000.0 1428000.0 925200.0 1414200.0 ;
      RECT  915000.0 1428000.0 925200.0 1441800.0 ;
      RECT  915000.0 1455600.0 925200.0 1441800.0 ;
      RECT  915000.0 1455600.0 925200.0 1469400.0 ;
      RECT  915000.0 1483200.0 925200.0 1469400.0 ;
      RECT  915000.0 1483200.0 925200.0 1497000.0 ;
      RECT  915000.0 1510800.0 925200.0 1497000.0 ;
      RECT  915000.0 1510800.0 925200.0 1524600.0 ;
      RECT  915000.0 1538400.0 925200.0 1524600.0 ;
      RECT  915000.0 1538400.0 925200.0 1552200.0 ;
      RECT  915000.0 1566000.0 925200.0 1552200.0 ;
      RECT  915000.0 1566000.0 925200.0 1579800.0 ;
      RECT  915000.0 1593600.0 925200.0 1579800.0 ;
      RECT  915000.0 1593600.0 925200.0 1607400.0 ;
      RECT  915000.0 1621200.0 925200.0 1607400.0 ;
      RECT  915000.0 1621200.0 925200.0 1635000.0 ;
      RECT  915000.0 1648800.0 925200.0 1635000.0 ;
      RECT  915000.0 1648800.0 925200.0 1662600.0 ;
      RECT  915000.0 1676400.0 925200.0 1662600.0 ;
      RECT  915000.0 1676400.0 925200.0 1690200.0 ;
      RECT  915000.0 1704000.0 925200.0 1690200.0 ;
      RECT  915000.0 1704000.0 925200.0 1717800.0 ;
      RECT  915000.0 1731600.0 925200.0 1717800.0 ;
      RECT  915000.0 1731600.0 925200.0 1745400.0 ;
      RECT  915000.0 1759200.0 925200.0 1745400.0 ;
      RECT  915000.0 1759200.0 925200.0 1773000.0 ;
      RECT  915000.0 1786800.0 925200.0 1773000.0 ;
      RECT  915000.0 1786800.0 925200.0 1800600.0 ;
      RECT  915000.0 1814400.0 925200.0 1800600.0 ;
      RECT  915000.0 1814400.0 925200.0 1828200.0 ;
      RECT  915000.0 1842000.0 925200.0 1828200.0 ;
      RECT  915000.0 1842000.0 925200.0 1855800.0 ;
      RECT  915000.0 1869600.0 925200.0 1855800.0 ;
      RECT  915000.0 1869600.0 925200.0 1883400.0 ;
      RECT  915000.0 1897200.0 925200.0 1883400.0 ;
      RECT  915000.0 1897200.0 925200.0 1911000.0 ;
      RECT  915000.0 1924800.0 925200.0 1911000.0 ;
      RECT  915000.0 1924800.0 925200.0 1938600.0 ;
      RECT  915000.0 1952400.0 925200.0 1938600.0 ;
      RECT  915000.0 1952400.0 925200.0 1966200.0 ;
      RECT  915000.0 1980000.0 925200.0 1966200.0 ;
      RECT  915000.0 1980000.0 925200.0 1993800.0 ;
      RECT  915000.0 2007600.0 925200.0 1993800.0 ;
      RECT  915000.0 2007600.0 925200.0 2021400.0 ;
      RECT  915000.0 2035200.0 925200.0 2021400.0 ;
      RECT  915000.0 2035200.0 925200.0 2049000.0 ;
      RECT  915000.0 2062800.0 925200.0 2049000.0 ;
      RECT  915000.0 2062800.0 925200.0 2076600.0 ;
      RECT  915000.0 2090400.0 925200.0 2076600.0 ;
      RECT  915000.0 2090400.0 925200.0 2104200.0 ;
      RECT  915000.0 2118000.0 925200.0 2104200.0 ;
      RECT  915000.0 2118000.0 925200.0 2131800.0 ;
      RECT  915000.0 2145600.0 925200.0 2131800.0 ;
      RECT  925200.0 379200.0 935400.0 393000.0 ;
      RECT  925200.0 406800.0 935400.0 393000.0 ;
      RECT  925200.0 406800.0 935400.0 420600.0 ;
      RECT  925200.0 434400.0 935400.0 420600.0 ;
      RECT  925200.0 434400.0 935400.0 448200.0 ;
      RECT  925200.0 462000.0 935400.0 448200.0 ;
      RECT  925200.0 462000.0 935400.0 475800.0 ;
      RECT  925200.0 489600.0 935400.0 475800.0 ;
      RECT  925200.0 489600.0 935400.0 503400.0 ;
      RECT  925200.0 517200.0 935400.0 503400.0 ;
      RECT  925200.0 517200.0 935400.0 531000.0 ;
      RECT  925200.0 544800.0 935400.0 531000.0 ;
      RECT  925200.0 544800.0 935400.0 558600.0 ;
      RECT  925200.0 572400.0 935400.0 558600.0 ;
      RECT  925200.0 572400.0 935400.0 586200.0 ;
      RECT  925200.0 600000.0 935400.0 586200.0 ;
      RECT  925200.0 600000.0 935400.0 613800.0 ;
      RECT  925200.0 627600.0 935400.0 613800.0 ;
      RECT  925200.0 627600.0 935400.0 641400.0 ;
      RECT  925200.0 655200.0 935400.0 641400.0 ;
      RECT  925200.0 655200.0 935400.0 669000.0 ;
      RECT  925200.0 682800.0 935400.0 669000.0 ;
      RECT  925200.0 682800.0 935400.0 696600.0 ;
      RECT  925200.0 710400.0 935400.0 696600.0 ;
      RECT  925200.0 710400.0 935400.0 724200.0 ;
      RECT  925200.0 738000.0 935400.0 724200.0 ;
      RECT  925200.0 738000.0 935400.0 751800.0 ;
      RECT  925200.0 765600.0 935400.0 751800.0 ;
      RECT  925200.0 765600.0 935400.0 779400.0 ;
      RECT  925200.0 793200.0 935400.0 779400.0 ;
      RECT  925200.0 793200.0 935400.0 807000.0 ;
      RECT  925200.0 820800.0 935400.0 807000.0 ;
      RECT  925200.0 820800.0 935400.0 834600.0 ;
      RECT  925200.0 848400.0 935400.0 834600.0 ;
      RECT  925200.0 848400.0 935400.0 862200.0 ;
      RECT  925200.0 876000.0 935400.0 862200.0 ;
      RECT  925200.0 876000.0 935400.0 889800.0 ;
      RECT  925200.0 903600.0 935400.0 889800.0 ;
      RECT  925200.0 903600.0 935400.0 917400.0 ;
      RECT  925200.0 931200.0 935400.0 917400.0 ;
      RECT  925200.0 931200.0 935400.0 945000.0 ;
      RECT  925200.0 958800.0 935400.0 945000.0 ;
      RECT  925200.0 958800.0 935400.0 972600.0 ;
      RECT  925200.0 986400.0 935400.0 972600.0 ;
      RECT  925200.0 986400.0 935400.0 1000200.0 ;
      RECT  925200.0 1014000.0 935400.0 1000200.0 ;
      RECT  925200.0 1014000.0 935400.0 1027800.0 ;
      RECT  925200.0 1041600.0 935400.0 1027800.0 ;
      RECT  925200.0 1041600.0 935400.0 1055400.0 ;
      RECT  925200.0 1069200.0 935400.0 1055400.0 ;
      RECT  925200.0 1069200.0 935400.0 1083000.0 ;
      RECT  925200.0 1096800.0 935400.0 1083000.0 ;
      RECT  925200.0 1096800.0 935400.0 1110600.0 ;
      RECT  925200.0 1124400.0 935400.0 1110600.0 ;
      RECT  925200.0 1124400.0 935400.0 1138200.0 ;
      RECT  925200.0 1152000.0 935400.0 1138200.0 ;
      RECT  925200.0 1152000.0 935400.0 1165800.0 ;
      RECT  925200.0 1179600.0 935400.0 1165800.0 ;
      RECT  925200.0 1179600.0 935400.0 1193400.0 ;
      RECT  925200.0 1207200.0 935400.0 1193400.0 ;
      RECT  925200.0 1207200.0 935400.0 1221000.0 ;
      RECT  925200.0 1234800.0 935400.0 1221000.0 ;
      RECT  925200.0 1234800.0 935400.0 1248600.0 ;
      RECT  925200.0 1262400.0 935400.0 1248600.0 ;
      RECT  925200.0 1262400.0 935400.0 1276200.0 ;
      RECT  925200.0 1290000.0 935400.0 1276200.0 ;
      RECT  925200.0 1290000.0 935400.0 1303800.0 ;
      RECT  925200.0 1317600.0 935400.0 1303800.0 ;
      RECT  925200.0 1317600.0 935400.0 1331400.0 ;
      RECT  925200.0 1345200.0 935400.0 1331400.0 ;
      RECT  925200.0 1345200.0 935400.0 1359000.0 ;
      RECT  925200.0 1372800.0 935400.0 1359000.0 ;
      RECT  925200.0 1372800.0 935400.0 1386600.0 ;
      RECT  925200.0 1400400.0 935400.0 1386600.0 ;
      RECT  925200.0 1400400.0 935400.0 1414200.0 ;
      RECT  925200.0 1428000.0 935400.0 1414200.0 ;
      RECT  925200.0 1428000.0 935400.0 1441800.0 ;
      RECT  925200.0 1455600.0 935400.0 1441800.0 ;
      RECT  925200.0 1455600.0 935400.0 1469400.0 ;
      RECT  925200.0 1483200.0 935400.0 1469400.0 ;
      RECT  925200.0 1483200.0 935400.0 1497000.0 ;
      RECT  925200.0 1510800.0 935400.0 1497000.0 ;
      RECT  925200.0 1510800.0 935400.0 1524600.0 ;
      RECT  925200.0 1538400.0 935400.0 1524600.0 ;
      RECT  925200.0 1538400.0 935400.0 1552200.0 ;
      RECT  925200.0 1566000.0 935400.0 1552200.0 ;
      RECT  925200.0 1566000.0 935400.0 1579800.0 ;
      RECT  925200.0 1593600.0 935400.0 1579800.0 ;
      RECT  925200.0 1593600.0 935400.0 1607400.0 ;
      RECT  925200.0 1621200.0 935400.0 1607400.0 ;
      RECT  925200.0 1621200.0 935400.0 1635000.0 ;
      RECT  925200.0 1648800.0 935400.0 1635000.0 ;
      RECT  925200.0 1648800.0 935400.0 1662600.0 ;
      RECT  925200.0 1676400.0 935400.0 1662600.0 ;
      RECT  925200.0 1676400.0 935400.0 1690200.0 ;
      RECT  925200.0 1704000.0 935400.0 1690200.0 ;
      RECT  925200.0 1704000.0 935400.0 1717800.0 ;
      RECT  925200.0 1731600.0 935400.0 1717800.0 ;
      RECT  925200.0 1731600.0 935400.0 1745400.0 ;
      RECT  925200.0 1759200.0 935400.0 1745400.0 ;
      RECT  925200.0 1759200.0 935400.0 1773000.0 ;
      RECT  925200.0 1786800.0 935400.0 1773000.0 ;
      RECT  925200.0 1786800.0 935400.0 1800600.0 ;
      RECT  925200.0 1814400.0 935400.0 1800600.0 ;
      RECT  925200.0 1814400.0 935400.0 1828200.0 ;
      RECT  925200.0 1842000.0 935400.0 1828200.0 ;
      RECT  925200.0 1842000.0 935400.0 1855800.0 ;
      RECT  925200.0 1869600.0 935400.0 1855800.0 ;
      RECT  925200.0 1869600.0 935400.0 1883400.0 ;
      RECT  925200.0 1897200.0 935400.0 1883400.0 ;
      RECT  925200.0 1897200.0 935400.0 1911000.0 ;
      RECT  925200.0 1924800.0 935400.0 1911000.0 ;
      RECT  925200.0 1924800.0 935400.0 1938600.0 ;
      RECT  925200.0 1952400.0 935400.0 1938600.0 ;
      RECT  925200.0 1952400.0 935400.0 1966200.0 ;
      RECT  925200.0 1980000.0 935400.0 1966200.0 ;
      RECT  925200.0 1980000.0 935400.0 1993800.0 ;
      RECT  925200.0 2007600.0 935400.0 1993800.0 ;
      RECT  925200.0 2007600.0 935400.0 2021400.0 ;
      RECT  925200.0 2035200.0 935400.0 2021400.0 ;
      RECT  925200.0 2035200.0 935400.0 2049000.0 ;
      RECT  925200.0 2062800.0 935400.0 2049000.0 ;
      RECT  925200.0 2062800.0 935400.0 2076600.0 ;
      RECT  925200.0 2090400.0 935400.0 2076600.0 ;
      RECT  925200.0 2090400.0 935400.0 2104200.0 ;
      RECT  925200.0 2118000.0 935400.0 2104200.0 ;
      RECT  925200.0 2118000.0 935400.0 2131800.0 ;
      RECT  925200.0 2145600.0 935400.0 2131800.0 ;
      RECT  935400.0 379200.0 945600.0 393000.0 ;
      RECT  935400.0 406800.0 945600.0 393000.0 ;
      RECT  935400.0 406800.0 945600.0 420600.0 ;
      RECT  935400.0 434400.0 945600.0 420600.0 ;
      RECT  935400.0 434400.0 945600.0 448200.0 ;
      RECT  935400.0 462000.0 945600.0 448200.0 ;
      RECT  935400.0 462000.0 945600.0 475800.0 ;
      RECT  935400.0 489600.0 945600.0 475800.0 ;
      RECT  935400.0 489600.0 945600.0 503400.0 ;
      RECT  935400.0 517200.0 945600.0 503400.0 ;
      RECT  935400.0 517200.0 945600.0 531000.0 ;
      RECT  935400.0 544800.0 945600.0 531000.0 ;
      RECT  935400.0 544800.0 945600.0 558600.0 ;
      RECT  935400.0 572400.0 945600.0 558600.0 ;
      RECT  935400.0 572400.0 945600.0 586200.0 ;
      RECT  935400.0 600000.0 945600.0 586200.0 ;
      RECT  935400.0 600000.0 945600.0 613800.0 ;
      RECT  935400.0 627600.0 945600.0 613800.0 ;
      RECT  935400.0 627600.0 945600.0 641400.0 ;
      RECT  935400.0 655200.0 945600.0 641400.0 ;
      RECT  935400.0 655200.0 945600.0 669000.0 ;
      RECT  935400.0 682800.0 945600.0 669000.0 ;
      RECT  935400.0 682800.0 945600.0 696600.0 ;
      RECT  935400.0 710400.0 945600.0 696600.0 ;
      RECT  935400.0 710400.0 945600.0 724200.0 ;
      RECT  935400.0 738000.0 945600.0 724200.0 ;
      RECT  935400.0 738000.0 945600.0 751800.0 ;
      RECT  935400.0 765600.0 945600.0 751800.0 ;
      RECT  935400.0 765600.0 945600.0 779400.0 ;
      RECT  935400.0 793200.0 945600.0 779400.0 ;
      RECT  935400.0 793200.0 945600.0 807000.0 ;
      RECT  935400.0 820800.0 945600.0 807000.0 ;
      RECT  935400.0 820800.0 945600.0 834600.0 ;
      RECT  935400.0 848400.0 945600.0 834600.0 ;
      RECT  935400.0 848400.0 945600.0 862200.0 ;
      RECT  935400.0 876000.0 945600.0 862200.0 ;
      RECT  935400.0 876000.0 945600.0 889800.0 ;
      RECT  935400.0 903600.0 945600.0 889800.0 ;
      RECT  935400.0 903600.0 945600.0 917400.0 ;
      RECT  935400.0 931200.0 945600.0 917400.0 ;
      RECT  935400.0 931200.0 945600.0 945000.0 ;
      RECT  935400.0 958800.0 945600.0 945000.0 ;
      RECT  935400.0 958800.0 945600.0 972600.0 ;
      RECT  935400.0 986400.0 945600.0 972600.0 ;
      RECT  935400.0 986400.0 945600.0 1000200.0 ;
      RECT  935400.0 1014000.0 945600.0 1000200.0 ;
      RECT  935400.0 1014000.0 945600.0 1027800.0 ;
      RECT  935400.0 1041600.0 945600.0 1027800.0 ;
      RECT  935400.0 1041600.0 945600.0 1055400.0 ;
      RECT  935400.0 1069200.0 945600.0 1055400.0 ;
      RECT  935400.0 1069200.0 945600.0 1083000.0 ;
      RECT  935400.0 1096800.0 945600.0 1083000.0 ;
      RECT  935400.0 1096800.0 945600.0 1110600.0 ;
      RECT  935400.0 1124400.0 945600.0 1110600.0 ;
      RECT  935400.0 1124400.0 945600.0 1138200.0 ;
      RECT  935400.0 1152000.0 945600.0 1138200.0 ;
      RECT  935400.0 1152000.0 945600.0 1165800.0 ;
      RECT  935400.0 1179600.0 945600.0 1165800.0 ;
      RECT  935400.0 1179600.0 945600.0 1193400.0 ;
      RECT  935400.0 1207200.0 945600.0 1193400.0 ;
      RECT  935400.0 1207200.0 945600.0 1221000.0 ;
      RECT  935400.0 1234800.0 945600.0 1221000.0 ;
      RECT  935400.0 1234800.0 945600.0 1248600.0 ;
      RECT  935400.0 1262400.0 945600.0 1248600.0 ;
      RECT  935400.0 1262400.0 945600.0 1276200.0 ;
      RECT  935400.0 1290000.0 945600.0 1276200.0 ;
      RECT  935400.0 1290000.0 945600.0 1303800.0 ;
      RECT  935400.0 1317600.0 945600.0 1303800.0 ;
      RECT  935400.0 1317600.0 945600.0 1331400.0 ;
      RECT  935400.0 1345200.0 945600.0 1331400.0 ;
      RECT  935400.0 1345200.0 945600.0 1359000.0 ;
      RECT  935400.0 1372800.0 945600.0 1359000.0 ;
      RECT  935400.0 1372800.0 945600.0 1386600.0 ;
      RECT  935400.0 1400400.0 945600.0 1386600.0 ;
      RECT  935400.0 1400400.0 945600.0 1414200.0 ;
      RECT  935400.0 1428000.0 945600.0 1414200.0 ;
      RECT  935400.0 1428000.0 945600.0 1441800.0 ;
      RECT  935400.0 1455600.0 945600.0 1441800.0 ;
      RECT  935400.0 1455600.0 945600.0 1469400.0 ;
      RECT  935400.0 1483200.0 945600.0 1469400.0 ;
      RECT  935400.0 1483200.0 945600.0 1497000.0 ;
      RECT  935400.0 1510800.0 945600.0 1497000.0 ;
      RECT  935400.0 1510800.0 945600.0 1524600.0 ;
      RECT  935400.0 1538400.0 945600.0 1524600.0 ;
      RECT  935400.0 1538400.0 945600.0 1552200.0 ;
      RECT  935400.0 1566000.0 945600.0 1552200.0 ;
      RECT  935400.0 1566000.0 945600.0 1579800.0 ;
      RECT  935400.0 1593600.0 945600.0 1579800.0 ;
      RECT  935400.0 1593600.0 945600.0 1607400.0 ;
      RECT  935400.0 1621200.0 945600.0 1607400.0 ;
      RECT  935400.0 1621200.0 945600.0 1635000.0 ;
      RECT  935400.0 1648800.0 945600.0 1635000.0 ;
      RECT  935400.0 1648800.0 945600.0 1662600.0 ;
      RECT  935400.0 1676400.0 945600.0 1662600.0 ;
      RECT  935400.0 1676400.0 945600.0 1690200.0 ;
      RECT  935400.0 1704000.0 945600.0 1690200.0 ;
      RECT  935400.0 1704000.0 945600.0 1717800.0 ;
      RECT  935400.0 1731600.0 945600.0 1717800.0 ;
      RECT  935400.0 1731600.0 945600.0 1745400.0 ;
      RECT  935400.0 1759200.0 945600.0 1745400.0 ;
      RECT  935400.0 1759200.0 945600.0 1773000.0 ;
      RECT  935400.0 1786800.0 945600.0 1773000.0 ;
      RECT  935400.0 1786800.0 945600.0 1800600.0 ;
      RECT  935400.0 1814400.0 945600.0 1800600.0 ;
      RECT  935400.0 1814400.0 945600.0 1828200.0 ;
      RECT  935400.0 1842000.0 945600.0 1828200.0 ;
      RECT  935400.0 1842000.0 945600.0 1855800.0 ;
      RECT  935400.0 1869600.0 945600.0 1855800.0 ;
      RECT  935400.0 1869600.0 945600.0 1883400.0 ;
      RECT  935400.0 1897200.0 945600.0 1883400.0 ;
      RECT  935400.0 1897200.0 945600.0 1911000.0 ;
      RECT  935400.0 1924800.0 945600.0 1911000.0 ;
      RECT  935400.0 1924800.0 945600.0 1938600.0 ;
      RECT  935400.0 1952400.0 945600.0 1938600.0 ;
      RECT  935400.0 1952400.0 945600.0 1966200.0 ;
      RECT  935400.0 1980000.0 945600.0 1966200.0 ;
      RECT  935400.0 1980000.0 945600.0 1993800.0 ;
      RECT  935400.0 2007600.0 945600.0 1993800.0 ;
      RECT  935400.0 2007600.0 945600.0 2021400.0 ;
      RECT  935400.0 2035200.0 945600.0 2021400.0 ;
      RECT  935400.0 2035200.0 945600.0 2049000.0 ;
      RECT  935400.0 2062800.0 945600.0 2049000.0 ;
      RECT  935400.0 2062800.0 945600.0 2076600.0 ;
      RECT  935400.0 2090400.0 945600.0 2076600.0 ;
      RECT  935400.0 2090400.0 945600.0 2104200.0 ;
      RECT  935400.0 2118000.0 945600.0 2104200.0 ;
      RECT  935400.0 2118000.0 945600.0 2131800.0 ;
      RECT  935400.0 2145600.0 945600.0 2131800.0 ;
      RECT  945600.0 379200.0 955800.0 393000.0 ;
      RECT  945600.0 406800.0 955800.0 393000.0 ;
      RECT  945600.0 406800.0 955800.0 420600.0 ;
      RECT  945600.0 434400.0 955800.0 420600.0 ;
      RECT  945600.0 434400.0 955800.0 448200.0 ;
      RECT  945600.0 462000.0 955800.0 448200.0 ;
      RECT  945600.0 462000.0 955800.0 475800.0 ;
      RECT  945600.0 489600.0 955800.0 475800.0 ;
      RECT  945600.0 489600.0 955800.0 503400.0 ;
      RECT  945600.0 517200.0 955800.0 503400.0 ;
      RECT  945600.0 517200.0 955800.0 531000.0 ;
      RECT  945600.0 544800.0 955800.0 531000.0 ;
      RECT  945600.0 544800.0 955800.0 558600.0 ;
      RECT  945600.0 572400.0 955800.0 558600.0 ;
      RECT  945600.0 572400.0 955800.0 586200.0 ;
      RECT  945600.0 600000.0 955800.0 586200.0 ;
      RECT  945600.0 600000.0 955800.0 613800.0 ;
      RECT  945600.0 627600.0 955800.0 613800.0 ;
      RECT  945600.0 627600.0 955800.0 641400.0 ;
      RECT  945600.0 655200.0 955800.0 641400.0 ;
      RECT  945600.0 655200.0 955800.0 669000.0 ;
      RECT  945600.0 682800.0 955800.0 669000.0 ;
      RECT  945600.0 682800.0 955800.0 696600.0 ;
      RECT  945600.0 710400.0 955800.0 696600.0 ;
      RECT  945600.0 710400.0 955800.0 724200.0 ;
      RECT  945600.0 738000.0 955800.0 724200.0 ;
      RECT  945600.0 738000.0 955800.0 751800.0 ;
      RECT  945600.0 765600.0 955800.0 751800.0 ;
      RECT  945600.0 765600.0 955800.0 779400.0 ;
      RECT  945600.0 793200.0 955800.0 779400.0 ;
      RECT  945600.0 793200.0 955800.0 807000.0 ;
      RECT  945600.0 820800.0 955800.0 807000.0 ;
      RECT  945600.0 820800.0 955800.0 834600.0 ;
      RECT  945600.0 848400.0 955800.0 834600.0 ;
      RECT  945600.0 848400.0 955800.0 862200.0 ;
      RECT  945600.0 876000.0 955800.0 862200.0 ;
      RECT  945600.0 876000.0 955800.0 889800.0 ;
      RECT  945600.0 903600.0 955800.0 889800.0 ;
      RECT  945600.0 903600.0 955800.0 917400.0 ;
      RECT  945600.0 931200.0 955800.0 917400.0 ;
      RECT  945600.0 931200.0 955800.0 945000.0 ;
      RECT  945600.0 958800.0 955800.0 945000.0 ;
      RECT  945600.0 958800.0 955800.0 972600.0 ;
      RECT  945600.0 986400.0 955800.0 972600.0 ;
      RECT  945600.0 986400.0 955800.0 1000200.0 ;
      RECT  945600.0 1014000.0 955800.0 1000200.0 ;
      RECT  945600.0 1014000.0 955800.0 1027800.0 ;
      RECT  945600.0 1041600.0 955800.0 1027800.0 ;
      RECT  945600.0 1041600.0 955800.0 1055400.0 ;
      RECT  945600.0 1069200.0 955800.0 1055400.0 ;
      RECT  945600.0 1069200.0 955800.0 1083000.0 ;
      RECT  945600.0 1096800.0 955800.0 1083000.0 ;
      RECT  945600.0 1096800.0 955800.0 1110600.0 ;
      RECT  945600.0 1124400.0 955800.0 1110600.0 ;
      RECT  945600.0 1124400.0 955800.0 1138200.0 ;
      RECT  945600.0 1152000.0 955800.0 1138200.0 ;
      RECT  945600.0 1152000.0 955800.0 1165800.0 ;
      RECT  945600.0 1179600.0 955800.0 1165800.0 ;
      RECT  945600.0 1179600.0 955800.0 1193400.0 ;
      RECT  945600.0 1207200.0 955800.0 1193400.0 ;
      RECT  945600.0 1207200.0 955800.0 1221000.0 ;
      RECT  945600.0 1234800.0 955800.0 1221000.0 ;
      RECT  945600.0 1234800.0 955800.0 1248600.0 ;
      RECT  945600.0 1262400.0 955800.0 1248600.0 ;
      RECT  945600.0 1262400.0 955800.0 1276200.0 ;
      RECT  945600.0 1290000.0 955800.0 1276200.0 ;
      RECT  945600.0 1290000.0 955800.0 1303800.0 ;
      RECT  945600.0 1317600.0 955800.0 1303800.0 ;
      RECT  945600.0 1317600.0 955800.0 1331400.0 ;
      RECT  945600.0 1345200.0 955800.0 1331400.0 ;
      RECT  945600.0 1345200.0 955800.0 1359000.0 ;
      RECT  945600.0 1372800.0 955800.0 1359000.0 ;
      RECT  945600.0 1372800.0 955800.0 1386600.0 ;
      RECT  945600.0 1400400.0 955800.0 1386600.0 ;
      RECT  945600.0 1400400.0 955800.0 1414200.0 ;
      RECT  945600.0 1428000.0 955800.0 1414200.0 ;
      RECT  945600.0 1428000.0 955800.0 1441800.0 ;
      RECT  945600.0 1455600.0 955800.0 1441800.0 ;
      RECT  945600.0 1455600.0 955800.0 1469400.0 ;
      RECT  945600.0 1483200.0 955800.0 1469400.0 ;
      RECT  945600.0 1483200.0 955800.0 1497000.0 ;
      RECT  945600.0 1510800.0 955800.0 1497000.0 ;
      RECT  945600.0 1510800.0 955800.0 1524600.0 ;
      RECT  945600.0 1538400.0 955800.0 1524600.0 ;
      RECT  945600.0 1538400.0 955800.0 1552200.0 ;
      RECT  945600.0 1566000.0 955800.0 1552200.0 ;
      RECT  945600.0 1566000.0 955800.0 1579800.0 ;
      RECT  945600.0 1593600.0 955800.0 1579800.0 ;
      RECT  945600.0 1593600.0 955800.0 1607400.0 ;
      RECT  945600.0 1621200.0 955800.0 1607400.0 ;
      RECT  945600.0 1621200.0 955800.0 1635000.0 ;
      RECT  945600.0 1648800.0 955800.0 1635000.0 ;
      RECT  945600.0 1648800.0 955800.0 1662600.0 ;
      RECT  945600.0 1676400.0 955800.0 1662600.0 ;
      RECT  945600.0 1676400.0 955800.0 1690200.0 ;
      RECT  945600.0 1704000.0 955800.0 1690200.0 ;
      RECT  945600.0 1704000.0 955800.0 1717800.0 ;
      RECT  945600.0 1731600.0 955800.0 1717800.0 ;
      RECT  945600.0 1731600.0 955800.0 1745400.0 ;
      RECT  945600.0 1759200.0 955800.0 1745400.0 ;
      RECT  945600.0 1759200.0 955800.0 1773000.0 ;
      RECT  945600.0 1786800.0 955800.0 1773000.0 ;
      RECT  945600.0 1786800.0 955800.0 1800600.0 ;
      RECT  945600.0 1814400.0 955800.0 1800600.0 ;
      RECT  945600.0 1814400.0 955800.0 1828200.0 ;
      RECT  945600.0 1842000.0 955800.0 1828200.0 ;
      RECT  945600.0 1842000.0 955800.0 1855800.0 ;
      RECT  945600.0 1869600.0 955800.0 1855800.0 ;
      RECT  945600.0 1869600.0 955800.0 1883400.0 ;
      RECT  945600.0 1897200.0 955800.0 1883400.0 ;
      RECT  945600.0 1897200.0 955800.0 1911000.0 ;
      RECT  945600.0 1924800.0 955800.0 1911000.0 ;
      RECT  945600.0 1924800.0 955800.0 1938600.0 ;
      RECT  945600.0 1952400.0 955800.0 1938600.0 ;
      RECT  945600.0 1952400.0 955800.0 1966200.0 ;
      RECT  945600.0 1980000.0 955800.0 1966200.0 ;
      RECT  945600.0 1980000.0 955800.0 1993800.0 ;
      RECT  945600.0 2007600.0 955800.0 1993800.0 ;
      RECT  945600.0 2007600.0 955800.0 2021400.0 ;
      RECT  945600.0 2035200.0 955800.0 2021400.0 ;
      RECT  945600.0 2035200.0 955800.0 2049000.0 ;
      RECT  945600.0 2062800.0 955800.0 2049000.0 ;
      RECT  945600.0 2062800.0 955800.0 2076600.0 ;
      RECT  945600.0 2090400.0 955800.0 2076600.0 ;
      RECT  945600.0 2090400.0 955800.0 2104200.0 ;
      RECT  945600.0 2118000.0 955800.0 2104200.0 ;
      RECT  945600.0 2118000.0 955800.0 2131800.0 ;
      RECT  945600.0 2145600.0 955800.0 2131800.0 ;
      RECT  955800.0 379200.0 966000.0 393000.0 ;
      RECT  955800.0 406800.0 966000.0 393000.0 ;
      RECT  955800.0 406800.0 966000.0 420600.0 ;
      RECT  955800.0 434400.0 966000.0 420600.0 ;
      RECT  955800.0 434400.0 966000.0 448200.0 ;
      RECT  955800.0 462000.0 966000.0 448200.0 ;
      RECT  955800.0 462000.0 966000.0 475800.0 ;
      RECT  955800.0 489600.0 966000.0 475800.0 ;
      RECT  955800.0 489600.0 966000.0 503400.0 ;
      RECT  955800.0 517200.0 966000.0 503400.0 ;
      RECT  955800.0 517200.0 966000.0 531000.0 ;
      RECT  955800.0 544800.0 966000.0 531000.0 ;
      RECT  955800.0 544800.0 966000.0 558600.0 ;
      RECT  955800.0 572400.0 966000.0 558600.0 ;
      RECT  955800.0 572400.0 966000.0 586200.0 ;
      RECT  955800.0 600000.0 966000.0 586200.0 ;
      RECT  955800.0 600000.0 966000.0 613800.0 ;
      RECT  955800.0 627600.0 966000.0 613800.0 ;
      RECT  955800.0 627600.0 966000.0 641400.0 ;
      RECT  955800.0 655200.0 966000.0 641400.0 ;
      RECT  955800.0 655200.0 966000.0 669000.0 ;
      RECT  955800.0 682800.0 966000.0 669000.0 ;
      RECT  955800.0 682800.0 966000.0 696600.0 ;
      RECT  955800.0 710400.0 966000.0 696600.0 ;
      RECT  955800.0 710400.0 966000.0 724200.0 ;
      RECT  955800.0 738000.0 966000.0 724200.0 ;
      RECT  955800.0 738000.0 966000.0 751800.0 ;
      RECT  955800.0 765600.0 966000.0 751800.0 ;
      RECT  955800.0 765600.0 966000.0 779400.0 ;
      RECT  955800.0 793200.0 966000.0 779400.0 ;
      RECT  955800.0 793200.0 966000.0 807000.0 ;
      RECT  955800.0 820800.0 966000.0 807000.0 ;
      RECT  955800.0 820800.0 966000.0 834600.0 ;
      RECT  955800.0 848400.0 966000.0 834600.0 ;
      RECT  955800.0 848400.0 966000.0 862200.0 ;
      RECT  955800.0 876000.0 966000.0 862200.0 ;
      RECT  955800.0 876000.0 966000.0 889800.0 ;
      RECT  955800.0 903600.0 966000.0 889800.0 ;
      RECT  955800.0 903600.0 966000.0 917400.0 ;
      RECT  955800.0 931200.0 966000.0 917400.0 ;
      RECT  955800.0 931200.0 966000.0 945000.0 ;
      RECT  955800.0 958800.0 966000.0 945000.0 ;
      RECT  955800.0 958800.0 966000.0 972600.0 ;
      RECT  955800.0 986400.0 966000.0 972600.0 ;
      RECT  955800.0 986400.0 966000.0 1000200.0 ;
      RECT  955800.0 1014000.0 966000.0 1000200.0 ;
      RECT  955800.0 1014000.0 966000.0 1027800.0 ;
      RECT  955800.0 1041600.0 966000.0 1027800.0 ;
      RECT  955800.0 1041600.0 966000.0 1055400.0 ;
      RECT  955800.0 1069200.0 966000.0 1055400.0 ;
      RECT  955800.0 1069200.0 966000.0 1083000.0 ;
      RECT  955800.0 1096800.0 966000.0 1083000.0 ;
      RECT  955800.0 1096800.0 966000.0 1110600.0 ;
      RECT  955800.0 1124400.0 966000.0 1110600.0 ;
      RECT  955800.0 1124400.0 966000.0 1138200.0 ;
      RECT  955800.0 1152000.0 966000.0 1138200.0 ;
      RECT  955800.0 1152000.0 966000.0 1165800.0 ;
      RECT  955800.0 1179600.0 966000.0 1165800.0 ;
      RECT  955800.0 1179600.0 966000.0 1193400.0 ;
      RECT  955800.0 1207200.0 966000.0 1193400.0 ;
      RECT  955800.0 1207200.0 966000.0 1221000.0 ;
      RECT  955800.0 1234800.0 966000.0 1221000.0 ;
      RECT  955800.0 1234800.0 966000.0 1248600.0 ;
      RECT  955800.0 1262400.0 966000.0 1248600.0 ;
      RECT  955800.0 1262400.0 966000.0 1276200.0 ;
      RECT  955800.0 1290000.0 966000.0 1276200.0 ;
      RECT  955800.0 1290000.0 966000.0 1303800.0 ;
      RECT  955800.0 1317600.0 966000.0 1303800.0 ;
      RECT  955800.0 1317600.0 966000.0 1331400.0 ;
      RECT  955800.0 1345200.0 966000.0 1331400.0 ;
      RECT  955800.0 1345200.0 966000.0 1359000.0 ;
      RECT  955800.0 1372800.0 966000.0 1359000.0 ;
      RECT  955800.0 1372800.0 966000.0 1386600.0 ;
      RECT  955800.0 1400400.0 966000.0 1386600.0 ;
      RECT  955800.0 1400400.0 966000.0 1414200.0 ;
      RECT  955800.0 1428000.0 966000.0 1414200.0 ;
      RECT  955800.0 1428000.0 966000.0 1441800.0 ;
      RECT  955800.0 1455600.0 966000.0 1441800.0 ;
      RECT  955800.0 1455600.0 966000.0 1469400.0 ;
      RECT  955800.0 1483200.0 966000.0 1469400.0 ;
      RECT  955800.0 1483200.0 966000.0 1497000.0 ;
      RECT  955800.0 1510800.0 966000.0 1497000.0 ;
      RECT  955800.0 1510800.0 966000.0 1524600.0 ;
      RECT  955800.0 1538400.0 966000.0 1524600.0 ;
      RECT  955800.0 1538400.0 966000.0 1552200.0 ;
      RECT  955800.0 1566000.0 966000.0 1552200.0 ;
      RECT  955800.0 1566000.0 966000.0 1579800.0 ;
      RECT  955800.0 1593600.0 966000.0 1579800.0 ;
      RECT  955800.0 1593600.0 966000.0 1607400.0 ;
      RECT  955800.0 1621200.0 966000.0 1607400.0 ;
      RECT  955800.0 1621200.0 966000.0 1635000.0 ;
      RECT  955800.0 1648800.0 966000.0 1635000.0 ;
      RECT  955800.0 1648800.0 966000.0 1662600.0 ;
      RECT  955800.0 1676400.0 966000.0 1662600.0 ;
      RECT  955800.0 1676400.0 966000.0 1690200.0 ;
      RECT  955800.0 1704000.0 966000.0 1690200.0 ;
      RECT  955800.0 1704000.0 966000.0 1717800.0 ;
      RECT  955800.0 1731600.0 966000.0 1717800.0 ;
      RECT  955800.0 1731600.0 966000.0 1745400.0 ;
      RECT  955800.0 1759200.0 966000.0 1745400.0 ;
      RECT  955800.0 1759200.0 966000.0 1773000.0 ;
      RECT  955800.0 1786800.0 966000.0 1773000.0 ;
      RECT  955800.0 1786800.0 966000.0 1800600.0 ;
      RECT  955800.0 1814400.0 966000.0 1800600.0 ;
      RECT  955800.0 1814400.0 966000.0 1828200.0 ;
      RECT  955800.0 1842000.0 966000.0 1828200.0 ;
      RECT  955800.0 1842000.0 966000.0 1855800.0 ;
      RECT  955800.0 1869600.0 966000.0 1855800.0 ;
      RECT  955800.0 1869600.0 966000.0 1883400.0 ;
      RECT  955800.0 1897200.0 966000.0 1883400.0 ;
      RECT  955800.0 1897200.0 966000.0 1911000.0 ;
      RECT  955800.0 1924800.0 966000.0 1911000.0 ;
      RECT  955800.0 1924800.0 966000.0 1938600.0 ;
      RECT  955800.0 1952400.0 966000.0 1938600.0 ;
      RECT  955800.0 1952400.0 966000.0 1966200.0 ;
      RECT  955800.0 1980000.0 966000.0 1966200.0 ;
      RECT  955800.0 1980000.0 966000.0 1993800.0 ;
      RECT  955800.0 2007600.0 966000.0 1993800.0 ;
      RECT  955800.0 2007600.0 966000.0 2021400.0 ;
      RECT  955800.0 2035200.0 966000.0 2021400.0 ;
      RECT  955800.0 2035200.0 966000.0 2049000.0 ;
      RECT  955800.0 2062800.0 966000.0 2049000.0 ;
      RECT  955800.0 2062800.0 966000.0 2076600.0 ;
      RECT  955800.0 2090400.0 966000.0 2076600.0 ;
      RECT  955800.0 2090400.0 966000.0 2104200.0 ;
      RECT  955800.0 2118000.0 966000.0 2104200.0 ;
      RECT  955800.0 2118000.0 966000.0 2131800.0 ;
      RECT  955800.0 2145600.0 966000.0 2131800.0 ;
      RECT  966000.0 379200.0 976200.0 393000.0 ;
      RECT  966000.0 406800.0 976200.0 393000.0 ;
      RECT  966000.0 406800.0 976200.0 420600.0 ;
      RECT  966000.0 434400.0 976200.0 420600.0 ;
      RECT  966000.0 434400.0 976200.0 448200.0 ;
      RECT  966000.0 462000.0 976200.0 448200.0 ;
      RECT  966000.0 462000.0 976200.0 475800.0 ;
      RECT  966000.0 489600.0 976200.0 475800.0 ;
      RECT  966000.0 489600.0 976200.0 503400.0 ;
      RECT  966000.0 517200.0 976200.0 503400.0 ;
      RECT  966000.0 517200.0 976200.0 531000.0 ;
      RECT  966000.0 544800.0 976200.0 531000.0 ;
      RECT  966000.0 544800.0 976200.0 558600.0 ;
      RECT  966000.0 572400.0 976200.0 558600.0 ;
      RECT  966000.0 572400.0 976200.0 586200.0 ;
      RECT  966000.0 600000.0 976200.0 586200.0 ;
      RECT  966000.0 600000.0 976200.0 613800.0 ;
      RECT  966000.0 627600.0 976200.0 613800.0 ;
      RECT  966000.0 627600.0 976200.0 641400.0 ;
      RECT  966000.0 655200.0 976200.0 641400.0 ;
      RECT  966000.0 655200.0 976200.0 669000.0 ;
      RECT  966000.0 682800.0 976200.0 669000.0 ;
      RECT  966000.0 682800.0 976200.0 696600.0 ;
      RECT  966000.0 710400.0 976200.0 696600.0 ;
      RECT  966000.0 710400.0 976200.0 724200.0 ;
      RECT  966000.0 738000.0 976200.0 724200.0 ;
      RECT  966000.0 738000.0 976200.0 751800.0 ;
      RECT  966000.0 765600.0 976200.0 751800.0 ;
      RECT  966000.0 765600.0 976200.0 779400.0 ;
      RECT  966000.0 793200.0 976200.0 779400.0 ;
      RECT  966000.0 793200.0 976200.0 807000.0 ;
      RECT  966000.0 820800.0 976200.0 807000.0 ;
      RECT  966000.0 820800.0 976200.0 834600.0 ;
      RECT  966000.0 848400.0 976200.0 834600.0 ;
      RECT  966000.0 848400.0 976200.0 862200.0 ;
      RECT  966000.0 876000.0 976200.0 862200.0 ;
      RECT  966000.0 876000.0 976200.0 889800.0 ;
      RECT  966000.0 903600.0 976200.0 889800.0 ;
      RECT  966000.0 903600.0 976200.0 917400.0 ;
      RECT  966000.0 931200.0 976200.0 917400.0 ;
      RECT  966000.0 931200.0 976200.0 945000.0 ;
      RECT  966000.0 958800.0 976200.0 945000.0 ;
      RECT  966000.0 958800.0 976200.0 972600.0 ;
      RECT  966000.0 986400.0 976200.0 972600.0 ;
      RECT  966000.0 986400.0 976200.0 1000200.0 ;
      RECT  966000.0 1014000.0 976200.0 1000200.0 ;
      RECT  966000.0 1014000.0 976200.0 1027800.0 ;
      RECT  966000.0 1041600.0 976200.0 1027800.0 ;
      RECT  966000.0 1041600.0 976200.0 1055400.0 ;
      RECT  966000.0 1069200.0 976200.0 1055400.0 ;
      RECT  966000.0 1069200.0 976200.0 1083000.0 ;
      RECT  966000.0 1096800.0 976200.0 1083000.0 ;
      RECT  966000.0 1096800.0 976200.0 1110600.0 ;
      RECT  966000.0 1124400.0 976200.0 1110600.0 ;
      RECT  966000.0 1124400.0 976200.0 1138200.0 ;
      RECT  966000.0 1152000.0 976200.0 1138200.0 ;
      RECT  966000.0 1152000.0 976200.0 1165800.0 ;
      RECT  966000.0 1179600.0 976200.0 1165800.0 ;
      RECT  966000.0 1179600.0 976200.0 1193400.0 ;
      RECT  966000.0 1207200.0 976200.0 1193400.0 ;
      RECT  966000.0 1207200.0 976200.0 1221000.0 ;
      RECT  966000.0 1234800.0 976200.0 1221000.0 ;
      RECT  966000.0 1234800.0 976200.0 1248600.0 ;
      RECT  966000.0 1262400.0 976200.0 1248600.0 ;
      RECT  966000.0 1262400.0 976200.0 1276200.0 ;
      RECT  966000.0 1290000.0 976200.0 1276200.0 ;
      RECT  966000.0 1290000.0 976200.0 1303800.0 ;
      RECT  966000.0 1317600.0 976200.0 1303800.0 ;
      RECT  966000.0 1317600.0 976200.0 1331400.0 ;
      RECT  966000.0 1345200.0 976200.0 1331400.0 ;
      RECT  966000.0 1345200.0 976200.0 1359000.0 ;
      RECT  966000.0 1372800.0 976200.0 1359000.0 ;
      RECT  966000.0 1372800.0 976200.0 1386600.0 ;
      RECT  966000.0 1400400.0 976200.0 1386600.0 ;
      RECT  966000.0 1400400.0 976200.0 1414200.0 ;
      RECT  966000.0 1428000.0 976200.0 1414200.0 ;
      RECT  966000.0 1428000.0 976200.0 1441800.0 ;
      RECT  966000.0 1455600.0 976200.0 1441800.0 ;
      RECT  966000.0 1455600.0 976200.0 1469400.0 ;
      RECT  966000.0 1483200.0 976200.0 1469400.0 ;
      RECT  966000.0 1483200.0 976200.0 1497000.0 ;
      RECT  966000.0 1510800.0 976200.0 1497000.0 ;
      RECT  966000.0 1510800.0 976200.0 1524600.0 ;
      RECT  966000.0 1538400.0 976200.0 1524600.0 ;
      RECT  966000.0 1538400.0 976200.0 1552200.0 ;
      RECT  966000.0 1566000.0 976200.0 1552200.0 ;
      RECT  966000.0 1566000.0 976200.0 1579800.0 ;
      RECT  966000.0 1593600.0 976200.0 1579800.0 ;
      RECT  966000.0 1593600.0 976200.0 1607400.0 ;
      RECT  966000.0 1621200.0 976200.0 1607400.0 ;
      RECT  966000.0 1621200.0 976200.0 1635000.0 ;
      RECT  966000.0 1648800.0 976200.0 1635000.0 ;
      RECT  966000.0 1648800.0 976200.0 1662600.0 ;
      RECT  966000.0 1676400.0 976200.0 1662600.0 ;
      RECT  966000.0 1676400.0 976200.0 1690200.0 ;
      RECT  966000.0 1704000.0 976200.0 1690200.0 ;
      RECT  966000.0 1704000.0 976200.0 1717800.0 ;
      RECT  966000.0 1731600.0 976200.0 1717800.0 ;
      RECT  966000.0 1731600.0 976200.0 1745400.0 ;
      RECT  966000.0 1759200.0 976200.0 1745400.0 ;
      RECT  966000.0 1759200.0 976200.0 1773000.0 ;
      RECT  966000.0 1786800.0 976200.0 1773000.0 ;
      RECT  966000.0 1786800.0 976200.0 1800600.0 ;
      RECT  966000.0 1814400.0 976200.0 1800600.0 ;
      RECT  966000.0 1814400.0 976200.0 1828200.0 ;
      RECT  966000.0 1842000.0 976200.0 1828200.0 ;
      RECT  966000.0 1842000.0 976200.0 1855800.0 ;
      RECT  966000.0 1869600.0 976200.0 1855800.0 ;
      RECT  966000.0 1869600.0 976200.0 1883400.0 ;
      RECT  966000.0 1897200.0 976200.0 1883400.0 ;
      RECT  966000.0 1897200.0 976200.0 1911000.0 ;
      RECT  966000.0 1924800.0 976200.0 1911000.0 ;
      RECT  966000.0 1924800.0 976200.0 1938600.0 ;
      RECT  966000.0 1952400.0 976200.0 1938600.0 ;
      RECT  966000.0 1952400.0 976200.0 1966200.0 ;
      RECT  966000.0 1980000.0 976200.0 1966200.0 ;
      RECT  966000.0 1980000.0 976200.0 1993800.0 ;
      RECT  966000.0 2007600.0 976200.0 1993800.0 ;
      RECT  966000.0 2007600.0 976200.0 2021400.0 ;
      RECT  966000.0 2035200.0 976200.0 2021400.0 ;
      RECT  966000.0 2035200.0 976200.0 2049000.0 ;
      RECT  966000.0 2062800.0 976200.0 2049000.0 ;
      RECT  966000.0 2062800.0 976200.0 2076600.0 ;
      RECT  966000.0 2090400.0 976200.0 2076600.0 ;
      RECT  966000.0 2090400.0 976200.0 2104200.0 ;
      RECT  966000.0 2118000.0 976200.0 2104200.0 ;
      RECT  966000.0 2118000.0 976200.0 2131800.0 ;
      RECT  966000.0 2145600.0 976200.0 2131800.0 ;
      RECT  976200.0 379200.0 986400.0 393000.0 ;
      RECT  976200.0 406800.0 986400.0 393000.0 ;
      RECT  976200.0 406800.0 986400.0 420600.0 ;
      RECT  976200.0 434400.0 986400.0 420600.0 ;
      RECT  976200.0 434400.0 986400.0 448200.0 ;
      RECT  976200.0 462000.0 986400.0 448200.0 ;
      RECT  976200.0 462000.0 986400.0 475800.0 ;
      RECT  976200.0 489600.0 986400.0 475800.0 ;
      RECT  976200.0 489600.0 986400.0 503400.0 ;
      RECT  976200.0 517200.0 986400.0 503400.0 ;
      RECT  976200.0 517200.0 986400.0 531000.0 ;
      RECT  976200.0 544800.0 986400.0 531000.0 ;
      RECT  976200.0 544800.0 986400.0 558600.0 ;
      RECT  976200.0 572400.0 986400.0 558600.0 ;
      RECT  976200.0 572400.0 986400.0 586200.0 ;
      RECT  976200.0 600000.0 986400.0 586200.0 ;
      RECT  976200.0 600000.0 986400.0 613800.0 ;
      RECT  976200.0 627600.0 986400.0 613800.0 ;
      RECT  976200.0 627600.0 986400.0 641400.0 ;
      RECT  976200.0 655200.0 986400.0 641400.0 ;
      RECT  976200.0 655200.0 986400.0 669000.0 ;
      RECT  976200.0 682800.0 986400.0 669000.0 ;
      RECT  976200.0 682800.0 986400.0 696600.0 ;
      RECT  976200.0 710400.0 986400.0 696600.0 ;
      RECT  976200.0 710400.0 986400.0 724200.0 ;
      RECT  976200.0 738000.0 986400.0 724200.0 ;
      RECT  976200.0 738000.0 986400.0 751800.0 ;
      RECT  976200.0 765600.0 986400.0 751800.0 ;
      RECT  976200.0 765600.0 986400.0 779400.0 ;
      RECT  976200.0 793200.0 986400.0 779400.0 ;
      RECT  976200.0 793200.0 986400.0 807000.0 ;
      RECT  976200.0 820800.0 986400.0 807000.0 ;
      RECT  976200.0 820800.0 986400.0 834600.0 ;
      RECT  976200.0 848400.0 986400.0 834600.0 ;
      RECT  976200.0 848400.0 986400.0 862200.0 ;
      RECT  976200.0 876000.0 986400.0 862200.0 ;
      RECT  976200.0 876000.0 986400.0 889800.0 ;
      RECT  976200.0 903600.0 986400.0 889800.0 ;
      RECT  976200.0 903600.0 986400.0 917400.0 ;
      RECT  976200.0 931200.0 986400.0 917400.0 ;
      RECT  976200.0 931200.0 986400.0 945000.0 ;
      RECT  976200.0 958800.0 986400.0 945000.0 ;
      RECT  976200.0 958800.0 986400.0 972600.0 ;
      RECT  976200.0 986400.0 986400.0 972600.0 ;
      RECT  976200.0 986400.0 986400.0 1000200.0 ;
      RECT  976200.0 1014000.0 986400.0 1000200.0 ;
      RECT  976200.0 1014000.0 986400.0 1027800.0 ;
      RECT  976200.0 1041600.0 986400.0 1027800.0 ;
      RECT  976200.0 1041600.0 986400.0 1055400.0 ;
      RECT  976200.0 1069200.0 986400.0 1055400.0 ;
      RECT  976200.0 1069200.0 986400.0 1083000.0 ;
      RECT  976200.0 1096800.0 986400.0 1083000.0 ;
      RECT  976200.0 1096800.0 986400.0 1110600.0 ;
      RECT  976200.0 1124400.0 986400.0 1110600.0 ;
      RECT  976200.0 1124400.0 986400.0 1138200.0 ;
      RECT  976200.0 1152000.0 986400.0 1138200.0 ;
      RECT  976200.0 1152000.0 986400.0 1165800.0 ;
      RECT  976200.0 1179600.0 986400.0 1165800.0 ;
      RECT  976200.0 1179600.0 986400.0 1193400.0 ;
      RECT  976200.0 1207200.0 986400.0 1193400.0 ;
      RECT  976200.0 1207200.0 986400.0 1221000.0 ;
      RECT  976200.0 1234800.0 986400.0 1221000.0 ;
      RECT  976200.0 1234800.0 986400.0 1248600.0 ;
      RECT  976200.0 1262400.0 986400.0 1248600.0 ;
      RECT  976200.0 1262400.0 986400.0 1276200.0 ;
      RECT  976200.0 1290000.0 986400.0 1276200.0 ;
      RECT  976200.0 1290000.0 986400.0 1303800.0 ;
      RECT  976200.0 1317600.0 986400.0 1303800.0 ;
      RECT  976200.0 1317600.0 986400.0 1331400.0 ;
      RECT  976200.0 1345200.0 986400.0 1331400.0 ;
      RECT  976200.0 1345200.0 986400.0 1359000.0 ;
      RECT  976200.0 1372800.0 986400.0 1359000.0 ;
      RECT  976200.0 1372800.0 986400.0 1386600.0 ;
      RECT  976200.0 1400400.0 986400.0 1386600.0 ;
      RECT  976200.0 1400400.0 986400.0 1414200.0 ;
      RECT  976200.0 1428000.0 986400.0 1414200.0 ;
      RECT  976200.0 1428000.0 986400.0 1441800.0 ;
      RECT  976200.0 1455600.0 986400.0 1441800.0 ;
      RECT  976200.0 1455600.0 986400.0 1469400.0 ;
      RECT  976200.0 1483200.0 986400.0 1469400.0 ;
      RECT  976200.0 1483200.0 986400.0 1497000.0 ;
      RECT  976200.0 1510800.0 986400.0 1497000.0 ;
      RECT  976200.0 1510800.0 986400.0 1524600.0 ;
      RECT  976200.0 1538400.0 986400.0 1524600.0 ;
      RECT  976200.0 1538400.0 986400.0 1552200.0 ;
      RECT  976200.0 1566000.0 986400.0 1552200.0 ;
      RECT  976200.0 1566000.0 986400.0 1579800.0 ;
      RECT  976200.0 1593600.0 986400.0 1579800.0 ;
      RECT  976200.0 1593600.0 986400.0 1607400.0 ;
      RECT  976200.0 1621200.0 986400.0 1607400.0 ;
      RECT  976200.0 1621200.0 986400.0 1635000.0 ;
      RECT  976200.0 1648800.0 986400.0 1635000.0 ;
      RECT  976200.0 1648800.0 986400.0 1662600.0 ;
      RECT  976200.0 1676400.0 986400.0 1662600.0 ;
      RECT  976200.0 1676400.0 986400.0 1690200.0 ;
      RECT  976200.0 1704000.0 986400.0 1690200.0 ;
      RECT  976200.0 1704000.0 986400.0 1717800.0 ;
      RECT  976200.0 1731600.0 986400.0 1717800.0 ;
      RECT  976200.0 1731600.0 986400.0 1745400.0 ;
      RECT  976200.0 1759200.0 986400.0 1745400.0 ;
      RECT  976200.0 1759200.0 986400.0 1773000.0 ;
      RECT  976200.0 1786800.0 986400.0 1773000.0 ;
      RECT  976200.0 1786800.0 986400.0 1800600.0 ;
      RECT  976200.0 1814400.0 986400.0 1800600.0 ;
      RECT  976200.0 1814400.0 986400.0 1828200.0 ;
      RECT  976200.0 1842000.0 986400.0 1828200.0 ;
      RECT  976200.0 1842000.0 986400.0 1855800.0 ;
      RECT  976200.0 1869600.0 986400.0 1855800.0 ;
      RECT  976200.0 1869600.0 986400.0 1883400.0 ;
      RECT  976200.0 1897200.0 986400.0 1883400.0 ;
      RECT  976200.0 1897200.0 986400.0 1911000.0 ;
      RECT  976200.0 1924800.0 986400.0 1911000.0 ;
      RECT  976200.0 1924800.0 986400.0 1938600.0 ;
      RECT  976200.0 1952400.0 986400.0 1938600.0 ;
      RECT  976200.0 1952400.0 986400.0 1966200.0 ;
      RECT  976200.0 1980000.0 986400.0 1966200.0 ;
      RECT  976200.0 1980000.0 986400.0 1993800.0 ;
      RECT  976200.0 2007600.0 986400.0 1993800.0 ;
      RECT  976200.0 2007600.0 986400.0 2021400.0 ;
      RECT  976200.0 2035200.0 986400.0 2021400.0 ;
      RECT  976200.0 2035200.0 986400.0 2049000.0 ;
      RECT  976200.0 2062800.0 986400.0 2049000.0 ;
      RECT  976200.0 2062800.0 986400.0 2076600.0 ;
      RECT  976200.0 2090400.0 986400.0 2076600.0 ;
      RECT  976200.0 2090400.0 986400.0 2104200.0 ;
      RECT  976200.0 2118000.0 986400.0 2104200.0 ;
      RECT  976200.0 2118000.0 986400.0 2131800.0 ;
      RECT  976200.0 2145600.0 986400.0 2131800.0 ;
      RECT  986400.0 379200.0 996600.0 393000.0 ;
      RECT  986400.0 406800.0 996600.0 393000.0 ;
      RECT  986400.0 406800.0 996600.0 420600.0 ;
      RECT  986400.0 434400.0 996600.0 420600.0 ;
      RECT  986400.0 434400.0 996600.0 448200.0 ;
      RECT  986400.0 462000.0 996600.0 448200.0 ;
      RECT  986400.0 462000.0 996600.0 475800.0 ;
      RECT  986400.0 489600.0 996600.0 475800.0 ;
      RECT  986400.0 489600.0 996600.0 503400.0 ;
      RECT  986400.0 517200.0 996600.0 503400.0 ;
      RECT  986400.0 517200.0 996600.0 531000.0 ;
      RECT  986400.0 544800.0 996600.0 531000.0 ;
      RECT  986400.0 544800.0 996600.0 558600.0 ;
      RECT  986400.0 572400.0 996600.0 558600.0 ;
      RECT  986400.0 572400.0 996600.0 586200.0 ;
      RECT  986400.0 600000.0 996600.0 586200.0 ;
      RECT  986400.0 600000.0 996600.0 613800.0 ;
      RECT  986400.0 627600.0 996600.0 613800.0 ;
      RECT  986400.0 627600.0 996600.0 641400.0 ;
      RECT  986400.0 655200.0 996600.0 641400.0 ;
      RECT  986400.0 655200.0 996600.0 669000.0 ;
      RECT  986400.0 682800.0 996600.0 669000.0 ;
      RECT  986400.0 682800.0 996600.0 696600.0 ;
      RECT  986400.0 710400.0 996600.0 696600.0 ;
      RECT  986400.0 710400.0 996600.0 724200.0 ;
      RECT  986400.0 738000.0 996600.0 724200.0 ;
      RECT  986400.0 738000.0 996600.0 751800.0 ;
      RECT  986400.0 765600.0 996600.0 751800.0 ;
      RECT  986400.0 765600.0 996600.0 779400.0 ;
      RECT  986400.0 793200.0 996600.0 779400.0 ;
      RECT  986400.0 793200.0 996600.0 807000.0 ;
      RECT  986400.0 820800.0 996600.0 807000.0 ;
      RECT  986400.0 820800.0 996600.0 834600.0 ;
      RECT  986400.0 848400.0 996600.0 834600.0 ;
      RECT  986400.0 848400.0 996600.0 862200.0 ;
      RECT  986400.0 876000.0 996600.0 862200.0 ;
      RECT  986400.0 876000.0 996600.0 889800.0 ;
      RECT  986400.0 903600.0 996600.0 889800.0 ;
      RECT  986400.0 903600.0 996600.0 917400.0 ;
      RECT  986400.0 931200.0 996600.0 917400.0 ;
      RECT  986400.0 931200.0 996600.0 945000.0 ;
      RECT  986400.0 958800.0 996600.0 945000.0 ;
      RECT  986400.0 958800.0 996600.0 972600.0 ;
      RECT  986400.0 986400.0 996600.0 972600.0 ;
      RECT  986400.0 986400.0 996600.0 1000200.0 ;
      RECT  986400.0 1014000.0 996600.0 1000200.0 ;
      RECT  986400.0 1014000.0 996600.0 1027800.0 ;
      RECT  986400.0 1041600.0 996600.0 1027800.0 ;
      RECT  986400.0 1041600.0 996600.0 1055400.0 ;
      RECT  986400.0 1069200.0 996600.0 1055400.0 ;
      RECT  986400.0 1069200.0 996600.0 1083000.0 ;
      RECT  986400.0 1096800.0 996600.0 1083000.0 ;
      RECT  986400.0 1096800.0 996600.0 1110600.0 ;
      RECT  986400.0 1124400.0 996600.0 1110600.0 ;
      RECT  986400.0 1124400.0 996600.0 1138200.0 ;
      RECT  986400.0 1152000.0 996600.0 1138200.0 ;
      RECT  986400.0 1152000.0 996600.0 1165800.0 ;
      RECT  986400.0 1179600.0 996600.0 1165800.0 ;
      RECT  986400.0 1179600.0 996600.0 1193400.0 ;
      RECT  986400.0 1207200.0 996600.0 1193400.0 ;
      RECT  986400.0 1207200.0 996600.0 1221000.0 ;
      RECT  986400.0 1234800.0 996600.0 1221000.0 ;
      RECT  986400.0 1234800.0 996600.0 1248600.0 ;
      RECT  986400.0 1262400.0 996600.0 1248600.0 ;
      RECT  986400.0 1262400.0 996600.0 1276200.0 ;
      RECT  986400.0 1290000.0 996600.0 1276200.0 ;
      RECT  986400.0 1290000.0 996600.0 1303800.0 ;
      RECT  986400.0 1317600.0 996600.0 1303800.0 ;
      RECT  986400.0 1317600.0 996600.0 1331400.0 ;
      RECT  986400.0 1345200.0 996600.0 1331400.0 ;
      RECT  986400.0 1345200.0 996600.0 1359000.0 ;
      RECT  986400.0 1372800.0 996600.0 1359000.0 ;
      RECT  986400.0 1372800.0 996600.0 1386600.0 ;
      RECT  986400.0 1400400.0 996600.0 1386600.0 ;
      RECT  986400.0 1400400.0 996600.0 1414200.0 ;
      RECT  986400.0 1428000.0 996600.0 1414200.0 ;
      RECT  986400.0 1428000.0 996600.0 1441800.0 ;
      RECT  986400.0 1455600.0 996600.0 1441800.0 ;
      RECT  986400.0 1455600.0 996600.0 1469400.0 ;
      RECT  986400.0 1483200.0 996600.0 1469400.0 ;
      RECT  986400.0 1483200.0 996600.0 1497000.0 ;
      RECT  986400.0 1510800.0 996600.0 1497000.0 ;
      RECT  986400.0 1510800.0 996600.0 1524600.0 ;
      RECT  986400.0 1538400.0 996600.0 1524600.0 ;
      RECT  986400.0 1538400.0 996600.0 1552200.0 ;
      RECT  986400.0 1566000.0 996600.0 1552200.0 ;
      RECT  986400.0 1566000.0 996600.0 1579800.0 ;
      RECT  986400.0 1593600.0 996600.0 1579800.0 ;
      RECT  986400.0 1593600.0 996600.0 1607400.0 ;
      RECT  986400.0 1621200.0 996600.0 1607400.0 ;
      RECT  986400.0 1621200.0 996600.0 1635000.0 ;
      RECT  986400.0 1648800.0 996600.0 1635000.0 ;
      RECT  986400.0 1648800.0 996600.0 1662600.0 ;
      RECT  986400.0 1676400.0 996600.0 1662600.0 ;
      RECT  986400.0 1676400.0 996600.0 1690200.0 ;
      RECT  986400.0 1704000.0 996600.0 1690200.0 ;
      RECT  986400.0 1704000.0 996600.0 1717800.0 ;
      RECT  986400.0 1731600.0 996600.0 1717800.0 ;
      RECT  986400.0 1731600.0 996600.0 1745400.0 ;
      RECT  986400.0 1759200.0 996600.0 1745400.0 ;
      RECT  986400.0 1759200.0 996600.0 1773000.0 ;
      RECT  986400.0 1786800.0 996600.0 1773000.0 ;
      RECT  986400.0 1786800.0 996600.0 1800600.0 ;
      RECT  986400.0 1814400.0 996600.0 1800600.0 ;
      RECT  986400.0 1814400.0 996600.0 1828200.0 ;
      RECT  986400.0 1842000.0 996600.0 1828200.0 ;
      RECT  986400.0 1842000.0 996600.0 1855800.0 ;
      RECT  986400.0 1869600.0 996600.0 1855800.0 ;
      RECT  986400.0 1869600.0 996600.0 1883400.0 ;
      RECT  986400.0 1897200.0 996600.0 1883400.0 ;
      RECT  986400.0 1897200.0 996600.0 1911000.0 ;
      RECT  986400.0 1924800.0 996600.0 1911000.0 ;
      RECT  986400.0 1924800.0 996600.0 1938600.0 ;
      RECT  986400.0 1952400.0 996600.0 1938600.0 ;
      RECT  986400.0 1952400.0 996600.0 1966200.0 ;
      RECT  986400.0 1980000.0 996600.0 1966200.0 ;
      RECT  986400.0 1980000.0 996600.0 1993800.0 ;
      RECT  986400.0 2007600.0 996600.0 1993800.0 ;
      RECT  986400.0 2007600.0 996600.0 2021400.0 ;
      RECT  986400.0 2035200.0 996600.0 2021400.0 ;
      RECT  986400.0 2035200.0 996600.0 2049000.0 ;
      RECT  986400.0 2062800.0 996600.0 2049000.0 ;
      RECT  986400.0 2062800.0 996600.0 2076600.0 ;
      RECT  986400.0 2090400.0 996600.0 2076600.0 ;
      RECT  986400.0 2090400.0 996600.0 2104200.0 ;
      RECT  986400.0 2118000.0 996600.0 2104200.0 ;
      RECT  986400.0 2118000.0 996600.0 2131800.0 ;
      RECT  986400.0 2145600.0 996600.0 2131800.0 ;
      RECT  996600.0 379200.0 1006800.0 393000.0 ;
      RECT  996600.0 406800.0 1006800.0 393000.0 ;
      RECT  996600.0 406800.0 1006800.0 420600.0 ;
      RECT  996600.0 434400.0 1006800.0 420600.0 ;
      RECT  996600.0 434400.0 1006800.0 448200.0 ;
      RECT  996600.0 462000.0 1006800.0 448200.0 ;
      RECT  996600.0 462000.0 1006800.0 475800.0 ;
      RECT  996600.0 489600.0 1006800.0 475800.0 ;
      RECT  996600.0 489600.0 1006800.0 503400.0 ;
      RECT  996600.0 517200.0 1006800.0 503400.0 ;
      RECT  996600.0 517200.0 1006800.0 531000.0 ;
      RECT  996600.0 544800.0 1006800.0 531000.0 ;
      RECT  996600.0 544800.0 1006800.0 558600.0 ;
      RECT  996600.0 572400.0 1006800.0 558600.0 ;
      RECT  996600.0 572400.0 1006800.0 586200.0 ;
      RECT  996600.0 600000.0 1006800.0 586200.0 ;
      RECT  996600.0 600000.0 1006800.0 613800.0 ;
      RECT  996600.0 627600.0 1006800.0 613800.0 ;
      RECT  996600.0 627600.0 1006800.0 641400.0 ;
      RECT  996600.0 655200.0 1006800.0 641400.0 ;
      RECT  996600.0 655200.0 1006800.0 669000.0 ;
      RECT  996600.0 682800.0 1006800.0 669000.0 ;
      RECT  996600.0 682800.0 1006800.0 696600.0 ;
      RECT  996600.0 710400.0 1006800.0 696600.0 ;
      RECT  996600.0 710400.0 1006800.0 724200.0 ;
      RECT  996600.0 738000.0 1006800.0 724200.0 ;
      RECT  996600.0 738000.0 1006800.0 751800.0 ;
      RECT  996600.0 765600.0 1006800.0 751800.0 ;
      RECT  996600.0 765600.0 1006800.0 779400.0 ;
      RECT  996600.0 793200.0 1006800.0 779400.0 ;
      RECT  996600.0 793200.0 1006800.0 807000.0 ;
      RECT  996600.0 820800.0 1006800.0 807000.0 ;
      RECT  996600.0 820800.0 1006800.0 834600.0 ;
      RECT  996600.0 848400.0 1006800.0 834600.0 ;
      RECT  996600.0 848400.0 1006800.0 862200.0 ;
      RECT  996600.0 876000.0 1006800.0 862200.0 ;
      RECT  996600.0 876000.0 1006800.0 889800.0 ;
      RECT  996600.0 903600.0 1006800.0 889800.0 ;
      RECT  996600.0 903600.0 1006800.0 917400.0 ;
      RECT  996600.0 931200.0 1006800.0 917400.0 ;
      RECT  996600.0 931200.0 1006800.0 945000.0 ;
      RECT  996600.0 958800.0 1006800.0 945000.0 ;
      RECT  996600.0 958800.0 1006800.0 972600.0 ;
      RECT  996600.0 986400.0 1006800.0 972600.0 ;
      RECT  996600.0 986400.0 1006800.0 1000200.0 ;
      RECT  996600.0 1014000.0 1006800.0 1000200.0 ;
      RECT  996600.0 1014000.0 1006800.0 1027800.0 ;
      RECT  996600.0 1041600.0 1006800.0 1027800.0 ;
      RECT  996600.0 1041600.0 1006800.0 1055400.0 ;
      RECT  996600.0 1069200.0 1006800.0 1055400.0 ;
      RECT  996600.0 1069200.0 1006800.0 1083000.0 ;
      RECT  996600.0 1096800.0 1006800.0 1083000.0 ;
      RECT  996600.0 1096800.0 1006800.0 1110600.0 ;
      RECT  996600.0 1124400.0 1006800.0 1110600.0 ;
      RECT  996600.0 1124400.0 1006800.0 1138200.0 ;
      RECT  996600.0 1152000.0 1006800.0 1138200.0 ;
      RECT  996600.0 1152000.0 1006800.0 1165800.0 ;
      RECT  996600.0 1179600.0 1006800.0 1165800.0 ;
      RECT  996600.0 1179600.0 1006800.0 1193400.0 ;
      RECT  996600.0 1207200.0 1006800.0 1193400.0 ;
      RECT  996600.0 1207200.0 1006800.0 1221000.0 ;
      RECT  996600.0 1234800.0 1006800.0 1221000.0 ;
      RECT  996600.0 1234800.0 1006800.0 1248600.0 ;
      RECT  996600.0 1262400.0 1006800.0 1248600.0 ;
      RECT  996600.0 1262400.0 1006800.0 1276200.0 ;
      RECT  996600.0 1290000.0 1006800.0 1276200.0 ;
      RECT  996600.0 1290000.0 1006800.0 1303800.0 ;
      RECT  996600.0 1317600.0 1006800.0 1303800.0 ;
      RECT  996600.0 1317600.0 1006800.0 1331400.0 ;
      RECT  996600.0 1345200.0 1006800.0 1331400.0 ;
      RECT  996600.0 1345200.0 1006800.0 1359000.0 ;
      RECT  996600.0 1372800.0 1006800.0 1359000.0 ;
      RECT  996600.0 1372800.0 1006800.0 1386600.0 ;
      RECT  996600.0 1400400.0 1006800.0 1386600.0 ;
      RECT  996600.0 1400400.0 1006800.0 1414200.0 ;
      RECT  996600.0 1428000.0 1006800.0 1414200.0 ;
      RECT  996600.0 1428000.0 1006800.0 1441800.0 ;
      RECT  996600.0 1455600.0 1006800.0 1441800.0 ;
      RECT  996600.0 1455600.0 1006800.0 1469400.0 ;
      RECT  996600.0 1483200.0 1006800.0 1469400.0 ;
      RECT  996600.0 1483200.0 1006800.0 1497000.0 ;
      RECT  996600.0 1510800.0 1006800.0 1497000.0 ;
      RECT  996600.0 1510800.0 1006800.0 1524600.0 ;
      RECT  996600.0 1538400.0 1006800.0 1524600.0 ;
      RECT  996600.0 1538400.0 1006800.0 1552200.0 ;
      RECT  996600.0 1566000.0 1006800.0 1552200.0 ;
      RECT  996600.0 1566000.0 1006800.0 1579800.0 ;
      RECT  996600.0 1593600.0 1006800.0 1579800.0 ;
      RECT  996600.0 1593600.0 1006800.0 1607400.0 ;
      RECT  996600.0 1621200.0 1006800.0 1607400.0 ;
      RECT  996600.0 1621200.0 1006800.0 1635000.0 ;
      RECT  996600.0 1648800.0 1006800.0 1635000.0 ;
      RECT  996600.0 1648800.0 1006800.0 1662600.0 ;
      RECT  996600.0 1676400.0 1006800.0 1662600.0 ;
      RECT  996600.0 1676400.0 1006800.0 1690200.0 ;
      RECT  996600.0 1704000.0 1006800.0 1690200.0 ;
      RECT  996600.0 1704000.0 1006800.0 1717800.0 ;
      RECT  996600.0 1731600.0 1006800.0 1717800.0 ;
      RECT  996600.0 1731600.0 1006800.0 1745400.0 ;
      RECT  996600.0 1759200.0 1006800.0 1745400.0 ;
      RECT  996600.0 1759200.0 1006800.0 1773000.0 ;
      RECT  996600.0 1786800.0 1006800.0 1773000.0 ;
      RECT  996600.0 1786800.0 1006800.0 1800600.0 ;
      RECT  996600.0 1814400.0 1006800.0 1800600.0 ;
      RECT  996600.0 1814400.0 1006800.0 1828200.0 ;
      RECT  996600.0 1842000.0 1006800.0 1828200.0 ;
      RECT  996600.0 1842000.0 1006800.0 1855800.0 ;
      RECT  996600.0 1869600.0 1006800.0 1855800.0 ;
      RECT  996600.0 1869600.0 1006800.0 1883400.0 ;
      RECT  996600.0 1897200.0 1006800.0 1883400.0 ;
      RECT  996600.0 1897200.0 1006800.0 1911000.0 ;
      RECT  996600.0 1924800.0 1006800.0 1911000.0 ;
      RECT  996600.0 1924800.0 1006800.0 1938600.0 ;
      RECT  996600.0 1952400.0 1006800.0 1938600.0 ;
      RECT  996600.0 1952400.0 1006800.0 1966200.0 ;
      RECT  996600.0 1980000.0 1006800.0 1966200.0 ;
      RECT  996600.0 1980000.0 1006800.0 1993800.0 ;
      RECT  996600.0 2007600.0 1006800.0 1993800.0 ;
      RECT  996600.0 2007600.0 1006800.0 2021400.0 ;
      RECT  996600.0 2035200.0 1006800.0 2021400.0 ;
      RECT  996600.0 2035200.0 1006800.0 2049000.0 ;
      RECT  996600.0 2062800.0 1006800.0 2049000.0 ;
      RECT  996600.0 2062800.0 1006800.0 2076600.0 ;
      RECT  996600.0 2090400.0 1006800.0 2076600.0 ;
      RECT  996600.0 2090400.0 1006800.0 2104200.0 ;
      RECT  996600.0 2118000.0 1006800.0 2104200.0 ;
      RECT  996600.0 2118000.0 1006800.0 2131800.0 ;
      RECT  996600.0 2145600.0 1006800.0 2131800.0 ;
      RECT  1006800.0 379200.0 1017000.0 393000.0 ;
      RECT  1006800.0 406800.0 1017000.0 393000.0 ;
      RECT  1006800.0 406800.0 1017000.0 420600.0 ;
      RECT  1006800.0 434400.0 1017000.0 420600.0 ;
      RECT  1006800.0 434400.0 1017000.0 448200.0 ;
      RECT  1006800.0 462000.0 1017000.0 448200.0 ;
      RECT  1006800.0 462000.0 1017000.0 475800.0 ;
      RECT  1006800.0 489600.0 1017000.0 475800.0 ;
      RECT  1006800.0 489600.0 1017000.0 503400.0 ;
      RECT  1006800.0 517200.0 1017000.0 503400.0 ;
      RECT  1006800.0 517200.0 1017000.0 531000.0 ;
      RECT  1006800.0 544800.0 1017000.0 531000.0 ;
      RECT  1006800.0 544800.0 1017000.0 558600.0 ;
      RECT  1006800.0 572400.0 1017000.0 558600.0 ;
      RECT  1006800.0 572400.0 1017000.0 586200.0 ;
      RECT  1006800.0 600000.0 1017000.0 586200.0 ;
      RECT  1006800.0 600000.0 1017000.0 613800.0 ;
      RECT  1006800.0 627600.0 1017000.0 613800.0 ;
      RECT  1006800.0 627600.0 1017000.0 641400.0 ;
      RECT  1006800.0 655200.0 1017000.0 641400.0 ;
      RECT  1006800.0 655200.0 1017000.0 669000.0 ;
      RECT  1006800.0 682800.0 1017000.0 669000.0 ;
      RECT  1006800.0 682800.0 1017000.0 696600.0 ;
      RECT  1006800.0 710400.0 1017000.0 696600.0 ;
      RECT  1006800.0 710400.0 1017000.0 724200.0 ;
      RECT  1006800.0 738000.0 1017000.0 724200.0 ;
      RECT  1006800.0 738000.0 1017000.0 751800.0 ;
      RECT  1006800.0 765600.0 1017000.0 751800.0 ;
      RECT  1006800.0 765600.0 1017000.0 779400.0 ;
      RECT  1006800.0 793200.0 1017000.0 779400.0 ;
      RECT  1006800.0 793200.0 1017000.0 807000.0 ;
      RECT  1006800.0 820800.0 1017000.0 807000.0 ;
      RECT  1006800.0 820800.0 1017000.0 834600.0 ;
      RECT  1006800.0 848400.0 1017000.0 834600.0 ;
      RECT  1006800.0 848400.0 1017000.0 862200.0 ;
      RECT  1006800.0 876000.0 1017000.0 862200.0 ;
      RECT  1006800.0 876000.0 1017000.0 889800.0 ;
      RECT  1006800.0 903600.0 1017000.0 889800.0 ;
      RECT  1006800.0 903600.0 1017000.0 917400.0 ;
      RECT  1006800.0 931200.0 1017000.0 917400.0 ;
      RECT  1006800.0 931200.0 1017000.0 945000.0 ;
      RECT  1006800.0 958800.0 1017000.0 945000.0 ;
      RECT  1006800.0 958800.0 1017000.0 972600.0 ;
      RECT  1006800.0 986400.0 1017000.0 972600.0 ;
      RECT  1006800.0 986400.0 1017000.0 1000200.0 ;
      RECT  1006800.0 1014000.0 1017000.0 1000200.0 ;
      RECT  1006800.0 1014000.0 1017000.0 1027800.0 ;
      RECT  1006800.0 1041600.0 1017000.0 1027800.0 ;
      RECT  1006800.0 1041600.0 1017000.0 1055400.0 ;
      RECT  1006800.0 1069200.0 1017000.0 1055400.0 ;
      RECT  1006800.0 1069200.0 1017000.0 1083000.0 ;
      RECT  1006800.0 1096800.0 1017000.0 1083000.0 ;
      RECT  1006800.0 1096800.0 1017000.0 1110600.0 ;
      RECT  1006800.0 1124400.0 1017000.0 1110600.0 ;
      RECT  1006800.0 1124400.0 1017000.0 1138200.0 ;
      RECT  1006800.0 1152000.0 1017000.0 1138200.0 ;
      RECT  1006800.0 1152000.0 1017000.0 1165800.0 ;
      RECT  1006800.0 1179600.0 1017000.0 1165800.0 ;
      RECT  1006800.0 1179600.0 1017000.0 1193400.0 ;
      RECT  1006800.0 1207200.0 1017000.0 1193400.0 ;
      RECT  1006800.0 1207200.0 1017000.0 1221000.0 ;
      RECT  1006800.0 1234800.0 1017000.0 1221000.0 ;
      RECT  1006800.0 1234800.0 1017000.0 1248600.0 ;
      RECT  1006800.0 1262400.0 1017000.0 1248600.0 ;
      RECT  1006800.0 1262400.0 1017000.0 1276200.0 ;
      RECT  1006800.0 1290000.0 1017000.0 1276200.0 ;
      RECT  1006800.0 1290000.0 1017000.0 1303800.0 ;
      RECT  1006800.0 1317600.0 1017000.0 1303800.0 ;
      RECT  1006800.0 1317600.0 1017000.0 1331400.0 ;
      RECT  1006800.0 1345200.0 1017000.0 1331400.0 ;
      RECT  1006800.0 1345200.0 1017000.0 1359000.0 ;
      RECT  1006800.0 1372800.0 1017000.0 1359000.0 ;
      RECT  1006800.0 1372800.0 1017000.0 1386600.0 ;
      RECT  1006800.0 1400400.0 1017000.0 1386600.0 ;
      RECT  1006800.0 1400400.0 1017000.0 1414200.0 ;
      RECT  1006800.0 1428000.0 1017000.0 1414200.0 ;
      RECT  1006800.0 1428000.0 1017000.0 1441800.0 ;
      RECT  1006800.0 1455600.0 1017000.0 1441800.0 ;
      RECT  1006800.0 1455600.0 1017000.0 1469400.0 ;
      RECT  1006800.0 1483200.0 1017000.0 1469400.0 ;
      RECT  1006800.0 1483200.0 1017000.0 1497000.0 ;
      RECT  1006800.0 1510800.0 1017000.0 1497000.0 ;
      RECT  1006800.0 1510800.0 1017000.0 1524600.0 ;
      RECT  1006800.0 1538400.0 1017000.0 1524600.0 ;
      RECT  1006800.0 1538400.0 1017000.0 1552200.0 ;
      RECT  1006800.0 1566000.0 1017000.0 1552200.0 ;
      RECT  1006800.0 1566000.0 1017000.0 1579800.0 ;
      RECT  1006800.0 1593600.0 1017000.0 1579800.0 ;
      RECT  1006800.0 1593600.0 1017000.0 1607400.0 ;
      RECT  1006800.0 1621200.0 1017000.0 1607400.0 ;
      RECT  1006800.0 1621200.0 1017000.0 1635000.0 ;
      RECT  1006800.0 1648800.0 1017000.0 1635000.0 ;
      RECT  1006800.0 1648800.0 1017000.0 1662600.0 ;
      RECT  1006800.0 1676400.0 1017000.0 1662600.0 ;
      RECT  1006800.0 1676400.0 1017000.0 1690200.0 ;
      RECT  1006800.0 1704000.0 1017000.0 1690200.0 ;
      RECT  1006800.0 1704000.0 1017000.0 1717800.0 ;
      RECT  1006800.0 1731600.0 1017000.0 1717800.0 ;
      RECT  1006800.0 1731600.0 1017000.0 1745400.0 ;
      RECT  1006800.0 1759200.0 1017000.0 1745400.0 ;
      RECT  1006800.0 1759200.0 1017000.0 1773000.0 ;
      RECT  1006800.0 1786800.0 1017000.0 1773000.0 ;
      RECT  1006800.0 1786800.0 1017000.0 1800600.0 ;
      RECT  1006800.0 1814400.0 1017000.0 1800600.0 ;
      RECT  1006800.0 1814400.0 1017000.0 1828200.0 ;
      RECT  1006800.0 1842000.0 1017000.0 1828200.0 ;
      RECT  1006800.0 1842000.0 1017000.0 1855800.0 ;
      RECT  1006800.0 1869600.0 1017000.0 1855800.0 ;
      RECT  1006800.0 1869600.0 1017000.0 1883400.0 ;
      RECT  1006800.0 1897200.0 1017000.0 1883400.0 ;
      RECT  1006800.0 1897200.0 1017000.0 1911000.0 ;
      RECT  1006800.0 1924800.0 1017000.0 1911000.0 ;
      RECT  1006800.0 1924800.0 1017000.0 1938600.0 ;
      RECT  1006800.0 1952400.0 1017000.0 1938600.0 ;
      RECT  1006800.0 1952400.0 1017000.0 1966200.0 ;
      RECT  1006800.0 1980000.0 1017000.0 1966200.0 ;
      RECT  1006800.0 1980000.0 1017000.0 1993800.0 ;
      RECT  1006800.0 2007600.0 1017000.0 1993800.0 ;
      RECT  1006800.0 2007600.0 1017000.0 2021400.0 ;
      RECT  1006800.0 2035200.0 1017000.0 2021400.0 ;
      RECT  1006800.0 2035200.0 1017000.0 2049000.0 ;
      RECT  1006800.0 2062800.0 1017000.0 2049000.0 ;
      RECT  1006800.0 2062800.0 1017000.0 2076600.0 ;
      RECT  1006800.0 2090400.0 1017000.0 2076600.0 ;
      RECT  1006800.0 2090400.0 1017000.0 2104200.0 ;
      RECT  1006800.0 2118000.0 1017000.0 2104200.0 ;
      RECT  1006800.0 2118000.0 1017000.0 2131800.0 ;
      RECT  1006800.0 2145600.0 1017000.0 2131800.0 ;
      RECT  1017000.0 379200.0 1027200.0 393000.0 ;
      RECT  1017000.0 406800.0 1027200.0 393000.0 ;
      RECT  1017000.0 406800.0 1027200.0 420600.0 ;
      RECT  1017000.0 434400.0 1027200.0 420600.0 ;
      RECT  1017000.0 434400.0 1027200.0 448200.0 ;
      RECT  1017000.0 462000.0 1027200.0 448200.0 ;
      RECT  1017000.0 462000.0 1027200.0 475800.0 ;
      RECT  1017000.0 489600.0 1027200.0 475800.0 ;
      RECT  1017000.0 489600.0 1027200.0 503400.0 ;
      RECT  1017000.0 517200.0 1027200.0 503400.0 ;
      RECT  1017000.0 517200.0 1027200.0 531000.0 ;
      RECT  1017000.0 544800.0 1027200.0 531000.0 ;
      RECT  1017000.0 544800.0 1027200.0 558600.0 ;
      RECT  1017000.0 572400.0 1027200.0 558600.0 ;
      RECT  1017000.0 572400.0 1027200.0 586200.0 ;
      RECT  1017000.0 600000.0 1027200.0 586200.0 ;
      RECT  1017000.0 600000.0 1027200.0 613800.0 ;
      RECT  1017000.0 627600.0 1027200.0 613800.0 ;
      RECT  1017000.0 627600.0 1027200.0 641400.0 ;
      RECT  1017000.0 655200.0 1027200.0 641400.0 ;
      RECT  1017000.0 655200.0 1027200.0 669000.0 ;
      RECT  1017000.0 682800.0 1027200.0 669000.0 ;
      RECT  1017000.0 682800.0 1027200.0 696600.0 ;
      RECT  1017000.0 710400.0 1027200.0 696600.0 ;
      RECT  1017000.0 710400.0 1027200.0 724200.0 ;
      RECT  1017000.0 738000.0 1027200.0 724200.0 ;
      RECT  1017000.0 738000.0 1027200.0 751800.0 ;
      RECT  1017000.0 765600.0 1027200.0 751800.0 ;
      RECT  1017000.0 765600.0 1027200.0 779400.0 ;
      RECT  1017000.0 793200.0 1027200.0 779400.0 ;
      RECT  1017000.0 793200.0 1027200.0 807000.0 ;
      RECT  1017000.0 820800.0 1027200.0 807000.0 ;
      RECT  1017000.0 820800.0 1027200.0 834600.0 ;
      RECT  1017000.0 848400.0 1027200.0 834600.0 ;
      RECT  1017000.0 848400.0 1027200.0 862200.0 ;
      RECT  1017000.0 876000.0 1027200.0 862200.0 ;
      RECT  1017000.0 876000.0 1027200.0 889800.0 ;
      RECT  1017000.0 903600.0 1027200.0 889800.0 ;
      RECT  1017000.0 903600.0 1027200.0 917400.0 ;
      RECT  1017000.0 931200.0 1027200.0 917400.0 ;
      RECT  1017000.0 931200.0 1027200.0 945000.0 ;
      RECT  1017000.0 958800.0 1027200.0 945000.0 ;
      RECT  1017000.0 958800.0 1027200.0 972600.0 ;
      RECT  1017000.0 986400.0 1027200.0 972600.0 ;
      RECT  1017000.0 986400.0 1027200.0 1000200.0 ;
      RECT  1017000.0 1014000.0 1027200.0 1000200.0 ;
      RECT  1017000.0 1014000.0 1027200.0 1027800.0 ;
      RECT  1017000.0 1041600.0 1027200.0 1027800.0 ;
      RECT  1017000.0 1041600.0 1027200.0 1055400.0 ;
      RECT  1017000.0 1069200.0 1027200.0 1055400.0 ;
      RECT  1017000.0 1069200.0 1027200.0 1083000.0 ;
      RECT  1017000.0 1096800.0 1027200.0 1083000.0 ;
      RECT  1017000.0 1096800.0 1027200.0 1110600.0 ;
      RECT  1017000.0 1124400.0 1027200.0 1110600.0 ;
      RECT  1017000.0 1124400.0 1027200.0 1138200.0 ;
      RECT  1017000.0 1152000.0 1027200.0 1138200.0 ;
      RECT  1017000.0 1152000.0 1027200.0 1165800.0 ;
      RECT  1017000.0 1179600.0 1027200.0 1165800.0 ;
      RECT  1017000.0 1179600.0 1027200.0 1193400.0 ;
      RECT  1017000.0 1207200.0 1027200.0 1193400.0 ;
      RECT  1017000.0 1207200.0 1027200.0 1221000.0 ;
      RECT  1017000.0 1234800.0 1027200.0 1221000.0 ;
      RECT  1017000.0 1234800.0 1027200.0 1248600.0 ;
      RECT  1017000.0 1262400.0 1027200.0 1248600.0 ;
      RECT  1017000.0 1262400.0 1027200.0 1276200.0 ;
      RECT  1017000.0 1290000.0 1027200.0 1276200.0 ;
      RECT  1017000.0 1290000.0 1027200.0 1303800.0 ;
      RECT  1017000.0 1317600.0 1027200.0 1303800.0 ;
      RECT  1017000.0 1317600.0 1027200.0 1331400.0 ;
      RECT  1017000.0 1345200.0 1027200.0 1331400.0 ;
      RECT  1017000.0 1345200.0 1027200.0 1359000.0 ;
      RECT  1017000.0 1372800.0 1027200.0 1359000.0 ;
      RECT  1017000.0 1372800.0 1027200.0 1386600.0 ;
      RECT  1017000.0 1400400.0 1027200.0 1386600.0 ;
      RECT  1017000.0 1400400.0 1027200.0 1414200.0 ;
      RECT  1017000.0 1428000.0 1027200.0 1414200.0 ;
      RECT  1017000.0 1428000.0 1027200.0 1441800.0 ;
      RECT  1017000.0 1455600.0 1027200.0 1441800.0 ;
      RECT  1017000.0 1455600.0 1027200.0 1469400.0 ;
      RECT  1017000.0 1483200.0 1027200.0 1469400.0 ;
      RECT  1017000.0 1483200.0 1027200.0 1497000.0 ;
      RECT  1017000.0 1510800.0 1027200.0 1497000.0 ;
      RECT  1017000.0 1510800.0 1027200.0 1524600.0 ;
      RECT  1017000.0 1538400.0 1027200.0 1524600.0 ;
      RECT  1017000.0 1538400.0 1027200.0 1552200.0 ;
      RECT  1017000.0 1566000.0 1027200.0 1552200.0 ;
      RECT  1017000.0 1566000.0 1027200.0 1579800.0 ;
      RECT  1017000.0 1593600.0 1027200.0 1579800.0 ;
      RECT  1017000.0 1593600.0 1027200.0 1607400.0 ;
      RECT  1017000.0 1621200.0 1027200.0 1607400.0 ;
      RECT  1017000.0 1621200.0 1027200.0 1635000.0 ;
      RECT  1017000.0 1648800.0 1027200.0 1635000.0 ;
      RECT  1017000.0 1648800.0 1027200.0 1662600.0 ;
      RECT  1017000.0 1676400.0 1027200.0 1662600.0 ;
      RECT  1017000.0 1676400.0 1027200.0 1690200.0 ;
      RECT  1017000.0 1704000.0 1027200.0 1690200.0 ;
      RECT  1017000.0 1704000.0 1027200.0 1717800.0 ;
      RECT  1017000.0 1731600.0 1027200.0 1717800.0 ;
      RECT  1017000.0 1731600.0 1027200.0 1745400.0 ;
      RECT  1017000.0 1759200.0 1027200.0 1745400.0 ;
      RECT  1017000.0 1759200.0 1027200.0 1773000.0 ;
      RECT  1017000.0 1786800.0 1027200.0 1773000.0 ;
      RECT  1017000.0 1786800.0 1027200.0 1800600.0 ;
      RECT  1017000.0 1814400.0 1027200.0 1800600.0 ;
      RECT  1017000.0 1814400.0 1027200.0 1828200.0 ;
      RECT  1017000.0 1842000.0 1027200.0 1828200.0 ;
      RECT  1017000.0 1842000.0 1027200.0 1855800.0 ;
      RECT  1017000.0 1869600.0 1027200.0 1855800.0 ;
      RECT  1017000.0 1869600.0 1027200.0 1883400.0 ;
      RECT  1017000.0 1897200.0 1027200.0 1883400.0 ;
      RECT  1017000.0 1897200.0 1027200.0 1911000.0 ;
      RECT  1017000.0 1924800.0 1027200.0 1911000.0 ;
      RECT  1017000.0 1924800.0 1027200.0 1938600.0 ;
      RECT  1017000.0 1952400.0 1027200.0 1938600.0 ;
      RECT  1017000.0 1952400.0 1027200.0 1966200.0 ;
      RECT  1017000.0 1980000.0 1027200.0 1966200.0 ;
      RECT  1017000.0 1980000.0 1027200.0 1993800.0 ;
      RECT  1017000.0 2007600.0 1027200.0 1993800.0 ;
      RECT  1017000.0 2007600.0 1027200.0 2021400.0 ;
      RECT  1017000.0 2035200.0 1027200.0 2021400.0 ;
      RECT  1017000.0 2035200.0 1027200.0 2049000.0 ;
      RECT  1017000.0 2062800.0 1027200.0 2049000.0 ;
      RECT  1017000.0 2062800.0 1027200.0 2076600.0 ;
      RECT  1017000.0 2090400.0 1027200.0 2076600.0 ;
      RECT  1017000.0 2090400.0 1027200.0 2104200.0 ;
      RECT  1017000.0 2118000.0 1027200.0 2104200.0 ;
      RECT  1017000.0 2118000.0 1027200.0 2131800.0 ;
      RECT  1017000.0 2145600.0 1027200.0 2131800.0 ;
      RECT  1027200.0 379200.0 1037400.0 393000.0 ;
      RECT  1027200.0 406800.0 1037400.0 393000.0 ;
      RECT  1027200.0 406800.0 1037400.0 420600.0 ;
      RECT  1027200.0 434400.0 1037400.0 420600.0 ;
      RECT  1027200.0 434400.0 1037400.0 448200.0 ;
      RECT  1027200.0 462000.0 1037400.0 448200.0 ;
      RECT  1027200.0 462000.0 1037400.0 475800.0 ;
      RECT  1027200.0 489600.0 1037400.0 475800.0 ;
      RECT  1027200.0 489600.0 1037400.0 503400.0 ;
      RECT  1027200.0 517200.0 1037400.0 503400.0 ;
      RECT  1027200.0 517200.0 1037400.0 531000.0 ;
      RECT  1027200.0 544800.0 1037400.0 531000.0 ;
      RECT  1027200.0 544800.0 1037400.0 558600.0 ;
      RECT  1027200.0 572400.0 1037400.0 558600.0 ;
      RECT  1027200.0 572400.0 1037400.0 586200.0 ;
      RECT  1027200.0 600000.0 1037400.0 586200.0 ;
      RECT  1027200.0 600000.0 1037400.0 613800.0 ;
      RECT  1027200.0 627600.0 1037400.0 613800.0 ;
      RECT  1027200.0 627600.0 1037400.0 641400.0 ;
      RECT  1027200.0 655200.0 1037400.0 641400.0 ;
      RECT  1027200.0 655200.0 1037400.0 669000.0 ;
      RECT  1027200.0 682800.0 1037400.0 669000.0 ;
      RECT  1027200.0 682800.0 1037400.0 696600.0 ;
      RECT  1027200.0 710400.0 1037400.0 696600.0 ;
      RECT  1027200.0 710400.0 1037400.0 724200.0 ;
      RECT  1027200.0 738000.0 1037400.0 724200.0 ;
      RECT  1027200.0 738000.0 1037400.0 751800.0 ;
      RECT  1027200.0 765600.0 1037400.0 751800.0 ;
      RECT  1027200.0 765600.0 1037400.0 779400.0 ;
      RECT  1027200.0 793200.0 1037400.0 779400.0 ;
      RECT  1027200.0 793200.0 1037400.0 807000.0 ;
      RECT  1027200.0 820800.0 1037400.0 807000.0 ;
      RECT  1027200.0 820800.0 1037400.0 834600.0 ;
      RECT  1027200.0 848400.0 1037400.0 834600.0 ;
      RECT  1027200.0 848400.0 1037400.0 862200.0 ;
      RECT  1027200.0 876000.0 1037400.0 862200.0 ;
      RECT  1027200.0 876000.0 1037400.0 889800.0 ;
      RECT  1027200.0 903600.0 1037400.0 889800.0 ;
      RECT  1027200.0 903600.0 1037400.0 917400.0 ;
      RECT  1027200.0 931200.0 1037400.0 917400.0 ;
      RECT  1027200.0 931200.0 1037400.0 945000.0 ;
      RECT  1027200.0 958800.0 1037400.0 945000.0 ;
      RECT  1027200.0 958800.0 1037400.0 972600.0 ;
      RECT  1027200.0 986400.0 1037400.0 972600.0 ;
      RECT  1027200.0 986400.0 1037400.0 1000200.0 ;
      RECT  1027200.0 1014000.0 1037400.0 1000200.0 ;
      RECT  1027200.0 1014000.0 1037400.0 1027800.0 ;
      RECT  1027200.0 1041600.0 1037400.0 1027800.0 ;
      RECT  1027200.0 1041600.0 1037400.0 1055400.0 ;
      RECT  1027200.0 1069200.0 1037400.0 1055400.0 ;
      RECT  1027200.0 1069200.0 1037400.0 1083000.0 ;
      RECT  1027200.0 1096800.0 1037400.0 1083000.0 ;
      RECT  1027200.0 1096800.0 1037400.0 1110600.0 ;
      RECT  1027200.0 1124400.0 1037400.0 1110600.0 ;
      RECT  1027200.0 1124400.0 1037400.0 1138200.0 ;
      RECT  1027200.0 1152000.0 1037400.0 1138200.0 ;
      RECT  1027200.0 1152000.0 1037400.0 1165800.0 ;
      RECT  1027200.0 1179600.0 1037400.0 1165800.0 ;
      RECT  1027200.0 1179600.0 1037400.0 1193400.0 ;
      RECT  1027200.0 1207200.0 1037400.0 1193400.0 ;
      RECT  1027200.0 1207200.0 1037400.0 1221000.0 ;
      RECT  1027200.0 1234800.0 1037400.0 1221000.0 ;
      RECT  1027200.0 1234800.0 1037400.0 1248600.0 ;
      RECT  1027200.0 1262400.0 1037400.0 1248600.0 ;
      RECT  1027200.0 1262400.0 1037400.0 1276200.0 ;
      RECT  1027200.0 1290000.0 1037400.0 1276200.0 ;
      RECT  1027200.0 1290000.0 1037400.0 1303800.0 ;
      RECT  1027200.0 1317600.0 1037400.0 1303800.0 ;
      RECT  1027200.0 1317600.0 1037400.0 1331400.0 ;
      RECT  1027200.0 1345200.0 1037400.0 1331400.0 ;
      RECT  1027200.0 1345200.0 1037400.0 1359000.0 ;
      RECT  1027200.0 1372800.0 1037400.0 1359000.0 ;
      RECT  1027200.0 1372800.0 1037400.0 1386600.0 ;
      RECT  1027200.0 1400400.0 1037400.0 1386600.0 ;
      RECT  1027200.0 1400400.0 1037400.0 1414200.0 ;
      RECT  1027200.0 1428000.0 1037400.0 1414200.0 ;
      RECT  1027200.0 1428000.0 1037400.0 1441800.0 ;
      RECT  1027200.0 1455600.0 1037400.0 1441800.0 ;
      RECT  1027200.0 1455600.0 1037400.0 1469400.0 ;
      RECT  1027200.0 1483200.0 1037400.0 1469400.0 ;
      RECT  1027200.0 1483200.0 1037400.0 1497000.0 ;
      RECT  1027200.0 1510800.0 1037400.0 1497000.0 ;
      RECT  1027200.0 1510800.0 1037400.0 1524600.0 ;
      RECT  1027200.0 1538400.0 1037400.0 1524600.0 ;
      RECT  1027200.0 1538400.0 1037400.0 1552200.0 ;
      RECT  1027200.0 1566000.0 1037400.0 1552200.0 ;
      RECT  1027200.0 1566000.0 1037400.0 1579800.0 ;
      RECT  1027200.0 1593600.0 1037400.0 1579800.0 ;
      RECT  1027200.0 1593600.0 1037400.0 1607400.0 ;
      RECT  1027200.0 1621200.0 1037400.0 1607400.0 ;
      RECT  1027200.0 1621200.0 1037400.0 1635000.0 ;
      RECT  1027200.0 1648800.0 1037400.0 1635000.0 ;
      RECT  1027200.0 1648800.0 1037400.0 1662600.0 ;
      RECT  1027200.0 1676400.0 1037400.0 1662600.0 ;
      RECT  1027200.0 1676400.0 1037400.0 1690200.0 ;
      RECT  1027200.0 1704000.0 1037400.0 1690200.0 ;
      RECT  1027200.0 1704000.0 1037400.0 1717800.0 ;
      RECT  1027200.0 1731600.0 1037400.0 1717800.0 ;
      RECT  1027200.0 1731600.0 1037400.0 1745400.0 ;
      RECT  1027200.0 1759200.0 1037400.0 1745400.0 ;
      RECT  1027200.0 1759200.0 1037400.0 1773000.0 ;
      RECT  1027200.0 1786800.0 1037400.0 1773000.0 ;
      RECT  1027200.0 1786800.0 1037400.0 1800600.0 ;
      RECT  1027200.0 1814400.0 1037400.0 1800600.0 ;
      RECT  1027200.0 1814400.0 1037400.0 1828200.0 ;
      RECT  1027200.0 1842000.0 1037400.0 1828200.0 ;
      RECT  1027200.0 1842000.0 1037400.0 1855800.0 ;
      RECT  1027200.0 1869600.0 1037400.0 1855800.0 ;
      RECT  1027200.0 1869600.0 1037400.0 1883400.0 ;
      RECT  1027200.0 1897200.0 1037400.0 1883400.0 ;
      RECT  1027200.0 1897200.0 1037400.0 1911000.0 ;
      RECT  1027200.0 1924800.0 1037400.0 1911000.0 ;
      RECT  1027200.0 1924800.0 1037400.0 1938600.0 ;
      RECT  1027200.0 1952400.0 1037400.0 1938600.0 ;
      RECT  1027200.0 1952400.0 1037400.0 1966200.0 ;
      RECT  1027200.0 1980000.0 1037400.0 1966200.0 ;
      RECT  1027200.0 1980000.0 1037400.0 1993800.0 ;
      RECT  1027200.0 2007600.0 1037400.0 1993800.0 ;
      RECT  1027200.0 2007600.0 1037400.0 2021400.0 ;
      RECT  1027200.0 2035200.0 1037400.0 2021400.0 ;
      RECT  1027200.0 2035200.0 1037400.0 2049000.0 ;
      RECT  1027200.0 2062800.0 1037400.0 2049000.0 ;
      RECT  1027200.0 2062800.0 1037400.0 2076600.0 ;
      RECT  1027200.0 2090400.0 1037400.0 2076600.0 ;
      RECT  1027200.0 2090400.0 1037400.0 2104200.0 ;
      RECT  1027200.0 2118000.0 1037400.0 2104200.0 ;
      RECT  1027200.0 2118000.0 1037400.0 2131800.0 ;
      RECT  1027200.0 2145600.0 1037400.0 2131800.0 ;
      RECT  1037400.0 379200.0 1047600.0 393000.0 ;
      RECT  1037400.0 406800.0 1047600.0 393000.0 ;
      RECT  1037400.0 406800.0 1047600.0 420600.0 ;
      RECT  1037400.0 434400.0 1047600.0 420600.0 ;
      RECT  1037400.0 434400.0 1047600.0 448200.0 ;
      RECT  1037400.0 462000.0 1047600.0 448200.0 ;
      RECT  1037400.0 462000.0 1047600.0 475800.0 ;
      RECT  1037400.0 489600.0 1047600.0 475800.0 ;
      RECT  1037400.0 489600.0 1047600.0 503400.0 ;
      RECT  1037400.0 517200.0 1047600.0 503400.0 ;
      RECT  1037400.0 517200.0 1047600.0 531000.0 ;
      RECT  1037400.0 544800.0 1047600.0 531000.0 ;
      RECT  1037400.0 544800.0 1047600.0 558600.0 ;
      RECT  1037400.0 572400.0 1047600.0 558600.0 ;
      RECT  1037400.0 572400.0 1047600.0 586200.0 ;
      RECT  1037400.0 600000.0 1047600.0 586200.0 ;
      RECT  1037400.0 600000.0 1047600.0 613800.0 ;
      RECT  1037400.0 627600.0 1047600.0 613800.0 ;
      RECT  1037400.0 627600.0 1047600.0 641400.0 ;
      RECT  1037400.0 655200.0 1047600.0 641400.0 ;
      RECT  1037400.0 655200.0 1047600.0 669000.0 ;
      RECT  1037400.0 682800.0 1047600.0 669000.0 ;
      RECT  1037400.0 682800.0 1047600.0 696600.0 ;
      RECT  1037400.0 710400.0 1047600.0 696600.0 ;
      RECT  1037400.0 710400.0 1047600.0 724200.0 ;
      RECT  1037400.0 738000.0 1047600.0 724200.0 ;
      RECT  1037400.0 738000.0 1047600.0 751800.0 ;
      RECT  1037400.0 765600.0 1047600.0 751800.0 ;
      RECT  1037400.0 765600.0 1047600.0 779400.0 ;
      RECT  1037400.0 793200.0 1047600.0 779400.0 ;
      RECT  1037400.0 793200.0 1047600.0 807000.0 ;
      RECT  1037400.0 820800.0 1047600.0 807000.0 ;
      RECT  1037400.0 820800.0 1047600.0 834600.0 ;
      RECT  1037400.0 848400.0 1047600.0 834600.0 ;
      RECT  1037400.0 848400.0 1047600.0 862200.0 ;
      RECT  1037400.0 876000.0 1047600.0 862200.0 ;
      RECT  1037400.0 876000.0 1047600.0 889800.0 ;
      RECT  1037400.0 903600.0 1047600.0 889800.0 ;
      RECT  1037400.0 903600.0 1047600.0 917400.0 ;
      RECT  1037400.0 931200.0 1047600.0 917400.0 ;
      RECT  1037400.0 931200.0 1047600.0 945000.0 ;
      RECT  1037400.0 958800.0 1047600.0 945000.0 ;
      RECT  1037400.0 958800.0 1047600.0 972600.0 ;
      RECT  1037400.0 986400.0 1047600.0 972600.0 ;
      RECT  1037400.0 986400.0 1047600.0 1000200.0 ;
      RECT  1037400.0 1014000.0 1047600.0 1000200.0 ;
      RECT  1037400.0 1014000.0 1047600.0 1027800.0 ;
      RECT  1037400.0 1041600.0 1047600.0 1027800.0 ;
      RECT  1037400.0 1041600.0 1047600.0 1055400.0 ;
      RECT  1037400.0 1069200.0 1047600.0 1055400.0 ;
      RECT  1037400.0 1069200.0 1047600.0 1083000.0 ;
      RECT  1037400.0 1096800.0 1047600.0 1083000.0 ;
      RECT  1037400.0 1096800.0 1047600.0 1110600.0 ;
      RECT  1037400.0 1124400.0 1047600.0 1110600.0 ;
      RECT  1037400.0 1124400.0 1047600.0 1138200.0 ;
      RECT  1037400.0 1152000.0 1047600.0 1138200.0 ;
      RECT  1037400.0 1152000.0 1047600.0 1165800.0 ;
      RECT  1037400.0 1179600.0 1047600.0 1165800.0 ;
      RECT  1037400.0 1179600.0 1047600.0 1193400.0 ;
      RECT  1037400.0 1207200.0 1047600.0 1193400.0 ;
      RECT  1037400.0 1207200.0 1047600.0 1221000.0 ;
      RECT  1037400.0 1234800.0 1047600.0 1221000.0 ;
      RECT  1037400.0 1234800.0 1047600.0 1248600.0 ;
      RECT  1037400.0 1262400.0 1047600.0 1248600.0 ;
      RECT  1037400.0 1262400.0 1047600.0 1276200.0 ;
      RECT  1037400.0 1290000.0 1047600.0 1276200.0 ;
      RECT  1037400.0 1290000.0 1047600.0 1303800.0 ;
      RECT  1037400.0 1317600.0 1047600.0 1303800.0 ;
      RECT  1037400.0 1317600.0 1047600.0 1331400.0 ;
      RECT  1037400.0 1345200.0 1047600.0 1331400.0 ;
      RECT  1037400.0 1345200.0 1047600.0 1359000.0 ;
      RECT  1037400.0 1372800.0 1047600.0 1359000.0 ;
      RECT  1037400.0 1372800.0 1047600.0 1386600.0 ;
      RECT  1037400.0 1400400.0 1047600.0 1386600.0 ;
      RECT  1037400.0 1400400.0 1047600.0 1414200.0 ;
      RECT  1037400.0 1428000.0 1047600.0 1414200.0 ;
      RECT  1037400.0 1428000.0 1047600.0 1441800.0 ;
      RECT  1037400.0 1455600.0 1047600.0 1441800.0 ;
      RECT  1037400.0 1455600.0 1047600.0 1469400.0 ;
      RECT  1037400.0 1483200.0 1047600.0 1469400.0 ;
      RECT  1037400.0 1483200.0 1047600.0 1497000.0 ;
      RECT  1037400.0 1510800.0 1047600.0 1497000.0 ;
      RECT  1037400.0 1510800.0 1047600.0 1524600.0 ;
      RECT  1037400.0 1538400.0 1047600.0 1524600.0 ;
      RECT  1037400.0 1538400.0 1047600.0 1552200.0 ;
      RECT  1037400.0 1566000.0 1047600.0 1552200.0 ;
      RECT  1037400.0 1566000.0 1047600.0 1579800.0 ;
      RECT  1037400.0 1593600.0 1047600.0 1579800.0 ;
      RECT  1037400.0 1593600.0 1047600.0 1607400.0 ;
      RECT  1037400.0 1621200.0 1047600.0 1607400.0 ;
      RECT  1037400.0 1621200.0 1047600.0 1635000.0 ;
      RECT  1037400.0 1648800.0 1047600.0 1635000.0 ;
      RECT  1037400.0 1648800.0 1047600.0 1662600.0 ;
      RECT  1037400.0 1676400.0 1047600.0 1662600.0 ;
      RECT  1037400.0 1676400.0 1047600.0 1690200.0 ;
      RECT  1037400.0 1704000.0 1047600.0 1690200.0 ;
      RECT  1037400.0 1704000.0 1047600.0 1717800.0 ;
      RECT  1037400.0 1731600.0 1047600.0 1717800.0 ;
      RECT  1037400.0 1731600.0 1047600.0 1745400.0 ;
      RECT  1037400.0 1759200.0 1047600.0 1745400.0 ;
      RECT  1037400.0 1759200.0 1047600.0 1773000.0 ;
      RECT  1037400.0 1786800.0 1047600.0 1773000.0 ;
      RECT  1037400.0 1786800.0 1047600.0 1800600.0 ;
      RECT  1037400.0 1814400.0 1047600.0 1800600.0 ;
      RECT  1037400.0 1814400.0 1047600.0 1828200.0 ;
      RECT  1037400.0 1842000.0 1047600.0 1828200.0 ;
      RECT  1037400.0 1842000.0 1047600.0 1855800.0 ;
      RECT  1037400.0 1869600.0 1047600.0 1855800.0 ;
      RECT  1037400.0 1869600.0 1047600.0 1883400.0 ;
      RECT  1037400.0 1897200.0 1047600.0 1883400.0 ;
      RECT  1037400.0 1897200.0 1047600.0 1911000.0 ;
      RECT  1037400.0 1924800.0 1047600.0 1911000.0 ;
      RECT  1037400.0 1924800.0 1047600.0 1938600.0 ;
      RECT  1037400.0 1952400.0 1047600.0 1938600.0 ;
      RECT  1037400.0 1952400.0 1047600.0 1966200.0 ;
      RECT  1037400.0 1980000.0 1047600.0 1966200.0 ;
      RECT  1037400.0 1980000.0 1047600.0 1993800.0 ;
      RECT  1037400.0 2007600.0 1047600.0 1993800.0 ;
      RECT  1037400.0 2007600.0 1047600.0 2021400.0 ;
      RECT  1037400.0 2035200.0 1047600.0 2021400.0 ;
      RECT  1037400.0 2035200.0 1047600.0 2049000.0 ;
      RECT  1037400.0 2062800.0 1047600.0 2049000.0 ;
      RECT  1037400.0 2062800.0 1047600.0 2076600.0 ;
      RECT  1037400.0 2090400.0 1047600.0 2076600.0 ;
      RECT  1037400.0 2090400.0 1047600.0 2104200.0 ;
      RECT  1037400.0 2118000.0 1047600.0 2104200.0 ;
      RECT  1037400.0 2118000.0 1047600.0 2131800.0 ;
      RECT  1037400.0 2145600.0 1047600.0 2131800.0 ;
      RECT  1047600.0 379200.0 1057800.0 393000.0 ;
      RECT  1047600.0 406800.0 1057800.0 393000.0 ;
      RECT  1047600.0 406800.0 1057800.0 420600.0 ;
      RECT  1047600.0 434400.0 1057800.0 420600.0 ;
      RECT  1047600.0 434400.0 1057800.0 448200.0 ;
      RECT  1047600.0 462000.0 1057800.0 448200.0 ;
      RECT  1047600.0 462000.0 1057800.0 475800.0 ;
      RECT  1047600.0 489600.0 1057800.0 475800.0 ;
      RECT  1047600.0 489600.0 1057800.0 503400.0 ;
      RECT  1047600.0 517200.0 1057800.0 503400.0 ;
      RECT  1047600.0 517200.0 1057800.0 531000.0 ;
      RECT  1047600.0 544800.0 1057800.0 531000.0 ;
      RECT  1047600.0 544800.0 1057800.0 558600.0 ;
      RECT  1047600.0 572400.0 1057800.0 558600.0 ;
      RECT  1047600.0 572400.0 1057800.0 586200.0 ;
      RECT  1047600.0 600000.0 1057800.0 586200.0 ;
      RECT  1047600.0 600000.0 1057800.0 613800.0 ;
      RECT  1047600.0 627600.0 1057800.0 613800.0 ;
      RECT  1047600.0 627600.0 1057800.0 641400.0 ;
      RECT  1047600.0 655200.0 1057800.0 641400.0 ;
      RECT  1047600.0 655200.0 1057800.0 669000.0 ;
      RECT  1047600.0 682800.0 1057800.0 669000.0 ;
      RECT  1047600.0 682800.0 1057800.0 696600.0 ;
      RECT  1047600.0 710400.0 1057800.0 696600.0 ;
      RECT  1047600.0 710400.0 1057800.0 724200.0 ;
      RECT  1047600.0 738000.0 1057800.0 724200.0 ;
      RECT  1047600.0 738000.0 1057800.0 751800.0 ;
      RECT  1047600.0 765600.0 1057800.0 751800.0 ;
      RECT  1047600.0 765600.0 1057800.0 779400.0 ;
      RECT  1047600.0 793200.0 1057800.0 779400.0 ;
      RECT  1047600.0 793200.0 1057800.0 807000.0 ;
      RECT  1047600.0 820800.0 1057800.0 807000.0 ;
      RECT  1047600.0 820800.0 1057800.0 834600.0 ;
      RECT  1047600.0 848400.0 1057800.0 834600.0 ;
      RECT  1047600.0 848400.0 1057800.0 862200.0 ;
      RECT  1047600.0 876000.0 1057800.0 862200.0 ;
      RECT  1047600.0 876000.0 1057800.0 889800.0 ;
      RECT  1047600.0 903600.0 1057800.0 889800.0 ;
      RECT  1047600.0 903600.0 1057800.0 917400.0 ;
      RECT  1047600.0 931200.0 1057800.0 917400.0 ;
      RECT  1047600.0 931200.0 1057800.0 945000.0 ;
      RECT  1047600.0 958800.0 1057800.0 945000.0 ;
      RECT  1047600.0 958800.0 1057800.0 972600.0 ;
      RECT  1047600.0 986400.0 1057800.0 972600.0 ;
      RECT  1047600.0 986400.0 1057800.0 1000200.0 ;
      RECT  1047600.0 1014000.0 1057800.0 1000200.0 ;
      RECT  1047600.0 1014000.0 1057800.0 1027800.0 ;
      RECT  1047600.0 1041600.0 1057800.0 1027800.0 ;
      RECT  1047600.0 1041600.0 1057800.0 1055400.0 ;
      RECT  1047600.0 1069200.0 1057800.0 1055400.0 ;
      RECT  1047600.0 1069200.0 1057800.0 1083000.0 ;
      RECT  1047600.0 1096800.0 1057800.0 1083000.0 ;
      RECT  1047600.0 1096800.0 1057800.0 1110600.0 ;
      RECT  1047600.0 1124400.0 1057800.0 1110600.0 ;
      RECT  1047600.0 1124400.0 1057800.0 1138200.0 ;
      RECT  1047600.0 1152000.0 1057800.0 1138200.0 ;
      RECT  1047600.0 1152000.0 1057800.0 1165800.0 ;
      RECT  1047600.0 1179600.0 1057800.0 1165800.0 ;
      RECT  1047600.0 1179600.0 1057800.0 1193400.0 ;
      RECT  1047600.0 1207200.0 1057800.0 1193400.0 ;
      RECT  1047600.0 1207200.0 1057800.0 1221000.0 ;
      RECT  1047600.0 1234800.0 1057800.0 1221000.0 ;
      RECT  1047600.0 1234800.0 1057800.0 1248600.0 ;
      RECT  1047600.0 1262400.0 1057800.0 1248600.0 ;
      RECT  1047600.0 1262400.0 1057800.0 1276200.0 ;
      RECT  1047600.0 1290000.0 1057800.0 1276200.0 ;
      RECT  1047600.0 1290000.0 1057800.0 1303800.0 ;
      RECT  1047600.0 1317600.0 1057800.0 1303800.0 ;
      RECT  1047600.0 1317600.0 1057800.0 1331400.0 ;
      RECT  1047600.0 1345200.0 1057800.0 1331400.0 ;
      RECT  1047600.0 1345200.0 1057800.0 1359000.0 ;
      RECT  1047600.0 1372800.0 1057800.0 1359000.0 ;
      RECT  1047600.0 1372800.0 1057800.0 1386600.0 ;
      RECT  1047600.0 1400400.0 1057800.0 1386600.0 ;
      RECT  1047600.0 1400400.0 1057800.0 1414200.0 ;
      RECT  1047600.0 1428000.0 1057800.0 1414200.0 ;
      RECT  1047600.0 1428000.0 1057800.0 1441800.0 ;
      RECT  1047600.0 1455600.0 1057800.0 1441800.0 ;
      RECT  1047600.0 1455600.0 1057800.0 1469400.0 ;
      RECT  1047600.0 1483200.0 1057800.0 1469400.0 ;
      RECT  1047600.0 1483200.0 1057800.0 1497000.0 ;
      RECT  1047600.0 1510800.0 1057800.0 1497000.0 ;
      RECT  1047600.0 1510800.0 1057800.0 1524600.0 ;
      RECT  1047600.0 1538400.0 1057800.0 1524600.0 ;
      RECT  1047600.0 1538400.0 1057800.0 1552200.0 ;
      RECT  1047600.0 1566000.0 1057800.0 1552200.0 ;
      RECT  1047600.0 1566000.0 1057800.0 1579800.0 ;
      RECT  1047600.0 1593600.0 1057800.0 1579800.0 ;
      RECT  1047600.0 1593600.0 1057800.0 1607400.0 ;
      RECT  1047600.0 1621200.0 1057800.0 1607400.0 ;
      RECT  1047600.0 1621200.0 1057800.0 1635000.0 ;
      RECT  1047600.0 1648800.0 1057800.0 1635000.0 ;
      RECT  1047600.0 1648800.0 1057800.0 1662600.0 ;
      RECT  1047600.0 1676400.0 1057800.0 1662600.0 ;
      RECT  1047600.0 1676400.0 1057800.0 1690200.0 ;
      RECT  1047600.0 1704000.0 1057800.0 1690200.0 ;
      RECT  1047600.0 1704000.0 1057800.0 1717800.0 ;
      RECT  1047600.0 1731600.0 1057800.0 1717800.0 ;
      RECT  1047600.0 1731600.0 1057800.0 1745400.0 ;
      RECT  1047600.0 1759200.0 1057800.0 1745400.0 ;
      RECT  1047600.0 1759200.0 1057800.0 1773000.0 ;
      RECT  1047600.0 1786800.0 1057800.0 1773000.0 ;
      RECT  1047600.0 1786800.0 1057800.0 1800600.0 ;
      RECT  1047600.0 1814400.0 1057800.0 1800600.0 ;
      RECT  1047600.0 1814400.0 1057800.0 1828200.0 ;
      RECT  1047600.0 1842000.0 1057800.0 1828200.0 ;
      RECT  1047600.0 1842000.0 1057800.0 1855800.0 ;
      RECT  1047600.0 1869600.0 1057800.0 1855800.0 ;
      RECT  1047600.0 1869600.0 1057800.0 1883400.0 ;
      RECT  1047600.0 1897200.0 1057800.0 1883400.0 ;
      RECT  1047600.0 1897200.0 1057800.0 1911000.0 ;
      RECT  1047600.0 1924800.0 1057800.0 1911000.0 ;
      RECT  1047600.0 1924800.0 1057800.0 1938600.0 ;
      RECT  1047600.0 1952400.0 1057800.0 1938600.0 ;
      RECT  1047600.0 1952400.0 1057800.0 1966200.0 ;
      RECT  1047600.0 1980000.0 1057800.0 1966200.0 ;
      RECT  1047600.0 1980000.0 1057800.0 1993800.0 ;
      RECT  1047600.0 2007600.0 1057800.0 1993800.0 ;
      RECT  1047600.0 2007600.0 1057800.0 2021400.0 ;
      RECT  1047600.0 2035200.0 1057800.0 2021400.0 ;
      RECT  1047600.0 2035200.0 1057800.0 2049000.0 ;
      RECT  1047600.0 2062800.0 1057800.0 2049000.0 ;
      RECT  1047600.0 2062800.0 1057800.0 2076600.0 ;
      RECT  1047600.0 2090400.0 1057800.0 2076600.0 ;
      RECT  1047600.0 2090400.0 1057800.0 2104200.0 ;
      RECT  1047600.0 2118000.0 1057800.0 2104200.0 ;
      RECT  1047600.0 2118000.0 1057800.0 2131800.0 ;
      RECT  1047600.0 2145600.0 1057800.0 2131800.0 ;
      RECT  1057800.0 379200.0 1068000.0 393000.0 ;
      RECT  1057800.0 406800.0 1068000.0 393000.0 ;
      RECT  1057800.0 406800.0 1068000.0 420600.0 ;
      RECT  1057800.0 434400.0 1068000.0 420600.0 ;
      RECT  1057800.0 434400.0 1068000.0 448200.0 ;
      RECT  1057800.0 462000.0 1068000.0 448200.0 ;
      RECT  1057800.0 462000.0 1068000.0 475800.0 ;
      RECT  1057800.0 489600.0 1068000.0 475800.0 ;
      RECT  1057800.0 489600.0 1068000.0 503400.0 ;
      RECT  1057800.0 517200.0 1068000.0 503400.0 ;
      RECT  1057800.0 517200.0 1068000.0 531000.0 ;
      RECT  1057800.0 544800.0 1068000.0 531000.0 ;
      RECT  1057800.0 544800.0 1068000.0 558600.0 ;
      RECT  1057800.0 572400.0 1068000.0 558600.0 ;
      RECT  1057800.0 572400.0 1068000.0 586200.0 ;
      RECT  1057800.0 600000.0 1068000.0 586200.0 ;
      RECT  1057800.0 600000.0 1068000.0 613800.0 ;
      RECT  1057800.0 627600.0 1068000.0 613800.0 ;
      RECT  1057800.0 627600.0 1068000.0 641400.0 ;
      RECT  1057800.0 655200.0 1068000.0 641400.0 ;
      RECT  1057800.0 655200.0 1068000.0 669000.0 ;
      RECT  1057800.0 682800.0 1068000.0 669000.0 ;
      RECT  1057800.0 682800.0 1068000.0 696600.0 ;
      RECT  1057800.0 710400.0 1068000.0 696600.0 ;
      RECT  1057800.0 710400.0 1068000.0 724200.0 ;
      RECT  1057800.0 738000.0 1068000.0 724200.0 ;
      RECT  1057800.0 738000.0 1068000.0 751800.0 ;
      RECT  1057800.0 765600.0 1068000.0 751800.0 ;
      RECT  1057800.0 765600.0 1068000.0 779400.0 ;
      RECT  1057800.0 793200.0 1068000.0 779400.0 ;
      RECT  1057800.0 793200.0 1068000.0 807000.0 ;
      RECT  1057800.0 820800.0 1068000.0 807000.0 ;
      RECT  1057800.0 820800.0 1068000.0 834600.0 ;
      RECT  1057800.0 848400.0 1068000.0 834600.0 ;
      RECT  1057800.0 848400.0 1068000.0 862200.0 ;
      RECT  1057800.0 876000.0 1068000.0 862200.0 ;
      RECT  1057800.0 876000.0 1068000.0 889800.0 ;
      RECT  1057800.0 903600.0 1068000.0 889800.0 ;
      RECT  1057800.0 903600.0 1068000.0 917400.0 ;
      RECT  1057800.0 931200.0 1068000.0 917400.0 ;
      RECT  1057800.0 931200.0 1068000.0 945000.0 ;
      RECT  1057800.0 958800.0 1068000.0 945000.0 ;
      RECT  1057800.0 958800.0 1068000.0 972600.0 ;
      RECT  1057800.0 986400.0 1068000.0 972600.0 ;
      RECT  1057800.0 986400.0 1068000.0 1000200.0 ;
      RECT  1057800.0 1014000.0 1068000.0 1000200.0 ;
      RECT  1057800.0 1014000.0 1068000.0 1027800.0 ;
      RECT  1057800.0 1041600.0 1068000.0 1027800.0 ;
      RECT  1057800.0 1041600.0 1068000.0 1055400.0 ;
      RECT  1057800.0 1069200.0 1068000.0 1055400.0 ;
      RECT  1057800.0 1069200.0 1068000.0 1083000.0 ;
      RECT  1057800.0 1096800.0 1068000.0 1083000.0 ;
      RECT  1057800.0 1096800.0 1068000.0 1110600.0 ;
      RECT  1057800.0 1124400.0 1068000.0 1110600.0 ;
      RECT  1057800.0 1124400.0 1068000.0 1138200.0 ;
      RECT  1057800.0 1152000.0 1068000.0 1138200.0 ;
      RECT  1057800.0 1152000.0 1068000.0 1165800.0 ;
      RECT  1057800.0 1179600.0 1068000.0 1165800.0 ;
      RECT  1057800.0 1179600.0 1068000.0 1193400.0 ;
      RECT  1057800.0 1207200.0 1068000.0 1193400.0 ;
      RECT  1057800.0 1207200.0 1068000.0 1221000.0 ;
      RECT  1057800.0 1234800.0 1068000.0 1221000.0 ;
      RECT  1057800.0 1234800.0 1068000.0 1248600.0 ;
      RECT  1057800.0 1262400.0 1068000.0 1248600.0 ;
      RECT  1057800.0 1262400.0 1068000.0 1276200.0 ;
      RECT  1057800.0 1290000.0 1068000.0 1276200.0 ;
      RECT  1057800.0 1290000.0 1068000.0 1303800.0 ;
      RECT  1057800.0 1317600.0 1068000.0 1303800.0 ;
      RECT  1057800.0 1317600.0 1068000.0 1331400.0 ;
      RECT  1057800.0 1345200.0 1068000.0 1331400.0 ;
      RECT  1057800.0 1345200.0 1068000.0 1359000.0 ;
      RECT  1057800.0 1372800.0 1068000.0 1359000.0 ;
      RECT  1057800.0 1372800.0 1068000.0 1386600.0 ;
      RECT  1057800.0 1400400.0 1068000.0 1386600.0 ;
      RECT  1057800.0 1400400.0 1068000.0 1414200.0 ;
      RECT  1057800.0 1428000.0 1068000.0 1414200.0 ;
      RECT  1057800.0 1428000.0 1068000.0 1441800.0 ;
      RECT  1057800.0 1455600.0 1068000.0 1441800.0 ;
      RECT  1057800.0 1455600.0 1068000.0 1469400.0 ;
      RECT  1057800.0 1483200.0 1068000.0 1469400.0 ;
      RECT  1057800.0 1483200.0 1068000.0 1497000.0 ;
      RECT  1057800.0 1510800.0 1068000.0 1497000.0 ;
      RECT  1057800.0 1510800.0 1068000.0 1524600.0 ;
      RECT  1057800.0 1538400.0 1068000.0 1524600.0 ;
      RECT  1057800.0 1538400.0 1068000.0 1552200.0 ;
      RECT  1057800.0 1566000.0 1068000.0 1552200.0 ;
      RECT  1057800.0 1566000.0 1068000.0 1579800.0 ;
      RECT  1057800.0 1593600.0 1068000.0 1579800.0 ;
      RECT  1057800.0 1593600.0 1068000.0 1607400.0 ;
      RECT  1057800.0 1621200.0 1068000.0 1607400.0 ;
      RECT  1057800.0 1621200.0 1068000.0 1635000.0 ;
      RECT  1057800.0 1648800.0 1068000.0 1635000.0 ;
      RECT  1057800.0 1648800.0 1068000.0 1662600.0 ;
      RECT  1057800.0 1676400.0 1068000.0 1662600.0 ;
      RECT  1057800.0 1676400.0 1068000.0 1690200.0 ;
      RECT  1057800.0 1704000.0 1068000.0 1690200.0 ;
      RECT  1057800.0 1704000.0 1068000.0 1717800.0 ;
      RECT  1057800.0 1731600.0 1068000.0 1717800.0 ;
      RECT  1057800.0 1731600.0 1068000.0 1745400.0 ;
      RECT  1057800.0 1759200.0 1068000.0 1745400.0 ;
      RECT  1057800.0 1759200.0 1068000.0 1773000.0 ;
      RECT  1057800.0 1786800.0 1068000.0 1773000.0 ;
      RECT  1057800.0 1786800.0 1068000.0 1800600.0 ;
      RECT  1057800.0 1814400.0 1068000.0 1800600.0 ;
      RECT  1057800.0 1814400.0 1068000.0 1828200.0 ;
      RECT  1057800.0 1842000.0 1068000.0 1828200.0 ;
      RECT  1057800.0 1842000.0 1068000.0 1855800.0 ;
      RECT  1057800.0 1869600.0 1068000.0 1855800.0 ;
      RECT  1057800.0 1869600.0 1068000.0 1883400.0 ;
      RECT  1057800.0 1897200.0 1068000.0 1883400.0 ;
      RECT  1057800.0 1897200.0 1068000.0 1911000.0 ;
      RECT  1057800.0 1924800.0 1068000.0 1911000.0 ;
      RECT  1057800.0 1924800.0 1068000.0 1938600.0 ;
      RECT  1057800.0 1952400.0 1068000.0 1938600.0 ;
      RECT  1057800.0 1952400.0 1068000.0 1966200.0 ;
      RECT  1057800.0 1980000.0 1068000.0 1966200.0 ;
      RECT  1057800.0 1980000.0 1068000.0 1993800.0 ;
      RECT  1057800.0 2007600.0 1068000.0 1993800.0 ;
      RECT  1057800.0 2007600.0 1068000.0 2021400.0 ;
      RECT  1057800.0 2035200.0 1068000.0 2021400.0 ;
      RECT  1057800.0 2035200.0 1068000.0 2049000.0 ;
      RECT  1057800.0 2062800.0 1068000.0 2049000.0 ;
      RECT  1057800.0 2062800.0 1068000.0 2076600.0 ;
      RECT  1057800.0 2090400.0 1068000.0 2076600.0 ;
      RECT  1057800.0 2090400.0 1068000.0 2104200.0 ;
      RECT  1057800.0 2118000.0 1068000.0 2104200.0 ;
      RECT  1057800.0 2118000.0 1068000.0 2131800.0 ;
      RECT  1057800.0 2145600.0 1068000.0 2131800.0 ;
      RECT  1068000.0 379200.0 1078200.0 393000.0 ;
      RECT  1068000.0 406800.0 1078200.0 393000.0 ;
      RECT  1068000.0 406800.0 1078200.0 420600.0 ;
      RECT  1068000.0 434400.0 1078200.0 420600.0 ;
      RECT  1068000.0 434400.0 1078200.0 448200.0 ;
      RECT  1068000.0 462000.0 1078200.0 448200.0 ;
      RECT  1068000.0 462000.0 1078200.0 475800.0 ;
      RECT  1068000.0 489600.0 1078200.0 475800.0 ;
      RECT  1068000.0 489600.0 1078200.0 503400.0 ;
      RECT  1068000.0 517200.0 1078200.0 503400.0 ;
      RECT  1068000.0 517200.0 1078200.0 531000.0 ;
      RECT  1068000.0 544800.0 1078200.0 531000.0 ;
      RECT  1068000.0 544800.0 1078200.0 558600.0 ;
      RECT  1068000.0 572400.0 1078200.0 558600.0 ;
      RECT  1068000.0 572400.0 1078200.0 586200.0 ;
      RECT  1068000.0 600000.0 1078200.0 586200.0 ;
      RECT  1068000.0 600000.0 1078200.0 613800.0 ;
      RECT  1068000.0 627600.0 1078200.0 613800.0 ;
      RECT  1068000.0 627600.0 1078200.0 641400.0 ;
      RECT  1068000.0 655200.0 1078200.0 641400.0 ;
      RECT  1068000.0 655200.0 1078200.0 669000.0 ;
      RECT  1068000.0 682800.0 1078200.0 669000.0 ;
      RECT  1068000.0 682800.0 1078200.0 696600.0 ;
      RECT  1068000.0 710400.0 1078200.0 696600.0 ;
      RECT  1068000.0 710400.0 1078200.0 724200.0 ;
      RECT  1068000.0 738000.0 1078200.0 724200.0 ;
      RECT  1068000.0 738000.0 1078200.0 751800.0 ;
      RECT  1068000.0 765600.0 1078200.0 751800.0 ;
      RECT  1068000.0 765600.0 1078200.0 779400.0 ;
      RECT  1068000.0 793200.0 1078200.0 779400.0 ;
      RECT  1068000.0 793200.0 1078200.0 807000.0 ;
      RECT  1068000.0 820800.0 1078200.0 807000.0 ;
      RECT  1068000.0 820800.0 1078200.0 834600.0 ;
      RECT  1068000.0 848400.0 1078200.0 834600.0 ;
      RECT  1068000.0 848400.0 1078200.0 862200.0 ;
      RECT  1068000.0 876000.0 1078200.0 862200.0 ;
      RECT  1068000.0 876000.0 1078200.0 889800.0 ;
      RECT  1068000.0 903600.0 1078200.0 889800.0 ;
      RECT  1068000.0 903600.0 1078200.0 917400.0 ;
      RECT  1068000.0 931200.0 1078200.0 917400.0 ;
      RECT  1068000.0 931200.0 1078200.0 945000.0 ;
      RECT  1068000.0 958800.0 1078200.0 945000.0 ;
      RECT  1068000.0 958800.0 1078200.0 972600.0 ;
      RECT  1068000.0 986400.0 1078200.0 972600.0 ;
      RECT  1068000.0 986400.0 1078200.0 1000200.0 ;
      RECT  1068000.0 1014000.0 1078200.0 1000200.0 ;
      RECT  1068000.0 1014000.0 1078200.0 1027800.0 ;
      RECT  1068000.0 1041600.0 1078200.0 1027800.0 ;
      RECT  1068000.0 1041600.0 1078200.0 1055400.0 ;
      RECT  1068000.0 1069200.0 1078200.0 1055400.0 ;
      RECT  1068000.0 1069200.0 1078200.0 1083000.0 ;
      RECT  1068000.0 1096800.0 1078200.0 1083000.0 ;
      RECT  1068000.0 1096800.0 1078200.0 1110600.0 ;
      RECT  1068000.0 1124400.0 1078200.0 1110600.0 ;
      RECT  1068000.0 1124400.0 1078200.0 1138200.0 ;
      RECT  1068000.0 1152000.0 1078200.0 1138200.0 ;
      RECT  1068000.0 1152000.0 1078200.0 1165800.0 ;
      RECT  1068000.0 1179600.0 1078200.0 1165800.0 ;
      RECT  1068000.0 1179600.0 1078200.0 1193400.0 ;
      RECT  1068000.0 1207200.0 1078200.0 1193400.0 ;
      RECT  1068000.0 1207200.0 1078200.0 1221000.0 ;
      RECT  1068000.0 1234800.0 1078200.0 1221000.0 ;
      RECT  1068000.0 1234800.0 1078200.0 1248600.0 ;
      RECT  1068000.0 1262400.0 1078200.0 1248600.0 ;
      RECT  1068000.0 1262400.0 1078200.0 1276200.0 ;
      RECT  1068000.0 1290000.0 1078200.0 1276200.0 ;
      RECT  1068000.0 1290000.0 1078200.0 1303800.0 ;
      RECT  1068000.0 1317600.0 1078200.0 1303800.0 ;
      RECT  1068000.0 1317600.0 1078200.0 1331400.0 ;
      RECT  1068000.0 1345200.0 1078200.0 1331400.0 ;
      RECT  1068000.0 1345200.0 1078200.0 1359000.0 ;
      RECT  1068000.0 1372800.0 1078200.0 1359000.0 ;
      RECT  1068000.0 1372800.0 1078200.0 1386600.0 ;
      RECT  1068000.0 1400400.0 1078200.0 1386600.0 ;
      RECT  1068000.0 1400400.0 1078200.0 1414200.0 ;
      RECT  1068000.0 1428000.0 1078200.0 1414200.0 ;
      RECT  1068000.0 1428000.0 1078200.0 1441800.0 ;
      RECT  1068000.0 1455600.0 1078200.0 1441800.0 ;
      RECT  1068000.0 1455600.0 1078200.0 1469400.0 ;
      RECT  1068000.0 1483200.0 1078200.0 1469400.0 ;
      RECT  1068000.0 1483200.0 1078200.0 1497000.0 ;
      RECT  1068000.0 1510800.0 1078200.0 1497000.0 ;
      RECT  1068000.0 1510800.0 1078200.0 1524600.0 ;
      RECT  1068000.0 1538400.0 1078200.0 1524600.0 ;
      RECT  1068000.0 1538400.0 1078200.0 1552200.0 ;
      RECT  1068000.0 1566000.0 1078200.0 1552200.0 ;
      RECT  1068000.0 1566000.0 1078200.0 1579800.0 ;
      RECT  1068000.0 1593600.0 1078200.0 1579800.0 ;
      RECT  1068000.0 1593600.0 1078200.0 1607400.0 ;
      RECT  1068000.0 1621200.0 1078200.0 1607400.0 ;
      RECT  1068000.0 1621200.0 1078200.0 1635000.0 ;
      RECT  1068000.0 1648800.0 1078200.0 1635000.0 ;
      RECT  1068000.0 1648800.0 1078200.0 1662600.0 ;
      RECT  1068000.0 1676400.0 1078200.0 1662600.0 ;
      RECT  1068000.0 1676400.0 1078200.0 1690200.0 ;
      RECT  1068000.0 1704000.0 1078200.0 1690200.0 ;
      RECT  1068000.0 1704000.0 1078200.0 1717800.0 ;
      RECT  1068000.0 1731600.0 1078200.0 1717800.0 ;
      RECT  1068000.0 1731600.0 1078200.0 1745400.0 ;
      RECT  1068000.0 1759200.0 1078200.0 1745400.0 ;
      RECT  1068000.0 1759200.0 1078200.0 1773000.0 ;
      RECT  1068000.0 1786800.0 1078200.0 1773000.0 ;
      RECT  1068000.0 1786800.0 1078200.0 1800600.0 ;
      RECT  1068000.0 1814400.0 1078200.0 1800600.0 ;
      RECT  1068000.0 1814400.0 1078200.0 1828200.0 ;
      RECT  1068000.0 1842000.0 1078200.0 1828200.0 ;
      RECT  1068000.0 1842000.0 1078200.0 1855800.0 ;
      RECT  1068000.0 1869600.0 1078200.0 1855800.0 ;
      RECT  1068000.0 1869600.0 1078200.0 1883400.0 ;
      RECT  1068000.0 1897200.0 1078200.0 1883400.0 ;
      RECT  1068000.0 1897200.0 1078200.0 1911000.0 ;
      RECT  1068000.0 1924800.0 1078200.0 1911000.0 ;
      RECT  1068000.0 1924800.0 1078200.0 1938600.0 ;
      RECT  1068000.0 1952400.0 1078200.0 1938600.0 ;
      RECT  1068000.0 1952400.0 1078200.0 1966200.0 ;
      RECT  1068000.0 1980000.0 1078200.0 1966200.0 ;
      RECT  1068000.0 1980000.0 1078200.0 1993800.0 ;
      RECT  1068000.0 2007600.0 1078200.0 1993800.0 ;
      RECT  1068000.0 2007600.0 1078200.0 2021400.0 ;
      RECT  1068000.0 2035200.0 1078200.0 2021400.0 ;
      RECT  1068000.0 2035200.0 1078200.0 2049000.0 ;
      RECT  1068000.0 2062800.0 1078200.0 2049000.0 ;
      RECT  1068000.0 2062800.0 1078200.0 2076600.0 ;
      RECT  1068000.0 2090400.0 1078200.0 2076600.0 ;
      RECT  1068000.0 2090400.0 1078200.0 2104200.0 ;
      RECT  1068000.0 2118000.0 1078200.0 2104200.0 ;
      RECT  1068000.0 2118000.0 1078200.0 2131800.0 ;
      RECT  1068000.0 2145600.0 1078200.0 2131800.0 ;
      RECT  1078200.0 379200.0 1088400.0 393000.0 ;
      RECT  1078200.0 406800.0 1088400.0 393000.0 ;
      RECT  1078200.0 406800.0 1088400.0 420600.0 ;
      RECT  1078200.0 434400.0 1088400.0 420600.0 ;
      RECT  1078200.0 434400.0 1088400.0 448200.0 ;
      RECT  1078200.0 462000.0 1088400.0 448200.0 ;
      RECT  1078200.0 462000.0 1088400.0 475800.0 ;
      RECT  1078200.0 489600.0 1088400.0 475800.0 ;
      RECT  1078200.0 489600.0 1088400.0 503400.0 ;
      RECT  1078200.0 517200.0 1088400.0 503400.0 ;
      RECT  1078200.0 517200.0 1088400.0 531000.0 ;
      RECT  1078200.0 544800.0 1088400.0 531000.0 ;
      RECT  1078200.0 544800.0 1088400.0 558600.0 ;
      RECT  1078200.0 572400.0 1088400.0 558600.0 ;
      RECT  1078200.0 572400.0 1088400.0 586200.0 ;
      RECT  1078200.0 600000.0 1088400.0 586200.0 ;
      RECT  1078200.0 600000.0 1088400.0 613800.0 ;
      RECT  1078200.0 627600.0 1088400.0 613800.0 ;
      RECT  1078200.0 627600.0 1088400.0 641400.0 ;
      RECT  1078200.0 655200.0 1088400.0 641400.0 ;
      RECT  1078200.0 655200.0 1088400.0 669000.0 ;
      RECT  1078200.0 682800.0 1088400.0 669000.0 ;
      RECT  1078200.0 682800.0 1088400.0 696600.0 ;
      RECT  1078200.0 710400.0 1088400.0 696600.0 ;
      RECT  1078200.0 710400.0 1088400.0 724200.0 ;
      RECT  1078200.0 738000.0 1088400.0 724200.0 ;
      RECT  1078200.0 738000.0 1088400.0 751800.0 ;
      RECT  1078200.0 765600.0 1088400.0 751800.0 ;
      RECT  1078200.0 765600.0 1088400.0 779400.0 ;
      RECT  1078200.0 793200.0 1088400.0 779400.0 ;
      RECT  1078200.0 793200.0 1088400.0 807000.0 ;
      RECT  1078200.0 820800.0 1088400.0 807000.0 ;
      RECT  1078200.0 820800.0 1088400.0 834600.0 ;
      RECT  1078200.0 848400.0 1088400.0 834600.0 ;
      RECT  1078200.0 848400.0 1088400.0 862200.0 ;
      RECT  1078200.0 876000.0 1088400.0 862200.0 ;
      RECT  1078200.0 876000.0 1088400.0 889800.0 ;
      RECT  1078200.0 903600.0 1088400.0 889800.0 ;
      RECT  1078200.0 903600.0 1088400.0 917400.0 ;
      RECT  1078200.0 931200.0 1088400.0 917400.0 ;
      RECT  1078200.0 931200.0 1088400.0 945000.0 ;
      RECT  1078200.0 958800.0 1088400.0 945000.0 ;
      RECT  1078200.0 958800.0 1088400.0 972600.0 ;
      RECT  1078200.0 986400.0 1088400.0 972600.0 ;
      RECT  1078200.0 986400.0 1088400.0 1000200.0 ;
      RECT  1078200.0 1014000.0 1088400.0 1000200.0 ;
      RECT  1078200.0 1014000.0 1088400.0 1027800.0 ;
      RECT  1078200.0 1041600.0 1088400.0 1027800.0 ;
      RECT  1078200.0 1041600.0 1088400.0 1055400.0 ;
      RECT  1078200.0 1069200.0 1088400.0 1055400.0 ;
      RECT  1078200.0 1069200.0 1088400.0 1083000.0 ;
      RECT  1078200.0 1096800.0 1088400.0 1083000.0 ;
      RECT  1078200.0 1096800.0 1088400.0 1110600.0 ;
      RECT  1078200.0 1124400.0 1088400.0 1110600.0 ;
      RECT  1078200.0 1124400.0 1088400.0 1138200.0 ;
      RECT  1078200.0 1152000.0 1088400.0 1138200.0 ;
      RECT  1078200.0 1152000.0 1088400.0 1165800.0 ;
      RECT  1078200.0 1179600.0 1088400.0 1165800.0 ;
      RECT  1078200.0 1179600.0 1088400.0 1193400.0 ;
      RECT  1078200.0 1207200.0 1088400.0 1193400.0 ;
      RECT  1078200.0 1207200.0 1088400.0 1221000.0 ;
      RECT  1078200.0 1234800.0 1088400.0 1221000.0 ;
      RECT  1078200.0 1234800.0 1088400.0 1248600.0 ;
      RECT  1078200.0 1262400.0 1088400.0 1248600.0 ;
      RECT  1078200.0 1262400.0 1088400.0 1276200.0 ;
      RECT  1078200.0 1290000.0 1088400.0 1276200.0 ;
      RECT  1078200.0 1290000.0 1088400.0 1303800.0 ;
      RECT  1078200.0 1317600.0 1088400.0 1303800.0 ;
      RECT  1078200.0 1317600.0 1088400.0 1331400.0 ;
      RECT  1078200.0 1345200.0 1088400.0 1331400.0 ;
      RECT  1078200.0 1345200.0 1088400.0 1359000.0 ;
      RECT  1078200.0 1372800.0 1088400.0 1359000.0 ;
      RECT  1078200.0 1372800.0 1088400.0 1386600.0 ;
      RECT  1078200.0 1400400.0 1088400.0 1386600.0 ;
      RECT  1078200.0 1400400.0 1088400.0 1414200.0 ;
      RECT  1078200.0 1428000.0 1088400.0 1414200.0 ;
      RECT  1078200.0 1428000.0 1088400.0 1441800.0 ;
      RECT  1078200.0 1455600.0 1088400.0 1441800.0 ;
      RECT  1078200.0 1455600.0 1088400.0 1469400.0 ;
      RECT  1078200.0 1483200.0 1088400.0 1469400.0 ;
      RECT  1078200.0 1483200.0 1088400.0 1497000.0 ;
      RECT  1078200.0 1510800.0 1088400.0 1497000.0 ;
      RECT  1078200.0 1510800.0 1088400.0 1524600.0 ;
      RECT  1078200.0 1538400.0 1088400.0 1524600.0 ;
      RECT  1078200.0 1538400.0 1088400.0 1552200.0 ;
      RECT  1078200.0 1566000.0 1088400.0 1552200.0 ;
      RECT  1078200.0 1566000.0 1088400.0 1579800.0 ;
      RECT  1078200.0 1593600.0 1088400.0 1579800.0 ;
      RECT  1078200.0 1593600.0 1088400.0 1607400.0 ;
      RECT  1078200.0 1621200.0 1088400.0 1607400.0 ;
      RECT  1078200.0 1621200.0 1088400.0 1635000.0 ;
      RECT  1078200.0 1648800.0 1088400.0 1635000.0 ;
      RECT  1078200.0 1648800.0 1088400.0 1662600.0 ;
      RECT  1078200.0 1676400.0 1088400.0 1662600.0 ;
      RECT  1078200.0 1676400.0 1088400.0 1690200.0 ;
      RECT  1078200.0 1704000.0 1088400.0 1690200.0 ;
      RECT  1078200.0 1704000.0 1088400.0 1717800.0 ;
      RECT  1078200.0 1731600.0 1088400.0 1717800.0 ;
      RECT  1078200.0 1731600.0 1088400.0 1745400.0 ;
      RECT  1078200.0 1759200.0 1088400.0 1745400.0 ;
      RECT  1078200.0 1759200.0 1088400.0 1773000.0 ;
      RECT  1078200.0 1786800.0 1088400.0 1773000.0 ;
      RECT  1078200.0 1786800.0 1088400.0 1800600.0 ;
      RECT  1078200.0 1814400.0 1088400.0 1800600.0 ;
      RECT  1078200.0 1814400.0 1088400.0 1828200.0 ;
      RECT  1078200.0 1842000.0 1088400.0 1828200.0 ;
      RECT  1078200.0 1842000.0 1088400.0 1855800.0 ;
      RECT  1078200.0 1869600.0 1088400.0 1855800.0 ;
      RECT  1078200.0 1869600.0 1088400.0 1883400.0 ;
      RECT  1078200.0 1897200.0 1088400.0 1883400.0 ;
      RECT  1078200.0 1897200.0 1088400.0 1911000.0 ;
      RECT  1078200.0 1924800.0 1088400.0 1911000.0 ;
      RECT  1078200.0 1924800.0 1088400.0 1938600.0 ;
      RECT  1078200.0 1952400.0 1088400.0 1938600.0 ;
      RECT  1078200.0 1952400.0 1088400.0 1966200.0 ;
      RECT  1078200.0 1980000.0 1088400.0 1966200.0 ;
      RECT  1078200.0 1980000.0 1088400.0 1993800.0 ;
      RECT  1078200.0 2007600.0 1088400.0 1993800.0 ;
      RECT  1078200.0 2007600.0 1088400.0 2021400.0 ;
      RECT  1078200.0 2035200.0 1088400.0 2021400.0 ;
      RECT  1078200.0 2035200.0 1088400.0 2049000.0 ;
      RECT  1078200.0 2062800.0 1088400.0 2049000.0 ;
      RECT  1078200.0 2062800.0 1088400.0 2076600.0 ;
      RECT  1078200.0 2090400.0 1088400.0 2076600.0 ;
      RECT  1078200.0 2090400.0 1088400.0 2104200.0 ;
      RECT  1078200.0 2118000.0 1088400.0 2104200.0 ;
      RECT  1078200.0 2118000.0 1088400.0 2131800.0 ;
      RECT  1078200.0 2145600.0 1088400.0 2131800.0 ;
      RECT  1088400.0 379200.0 1098600.0 393000.0 ;
      RECT  1088400.0 406800.0 1098600.0 393000.0 ;
      RECT  1088400.0 406800.0 1098600.0 420600.0 ;
      RECT  1088400.0 434400.0 1098600.0 420600.0 ;
      RECT  1088400.0 434400.0 1098600.0 448200.0 ;
      RECT  1088400.0 462000.0 1098600.0 448200.0 ;
      RECT  1088400.0 462000.0 1098600.0 475800.0 ;
      RECT  1088400.0 489600.0 1098600.0 475800.0 ;
      RECT  1088400.0 489600.0 1098600.0 503400.0 ;
      RECT  1088400.0 517200.0 1098600.0 503400.0 ;
      RECT  1088400.0 517200.0 1098600.0 531000.0 ;
      RECT  1088400.0 544800.0 1098600.0 531000.0 ;
      RECT  1088400.0 544800.0 1098600.0 558600.0 ;
      RECT  1088400.0 572400.0 1098600.0 558600.0 ;
      RECT  1088400.0 572400.0 1098600.0 586200.0 ;
      RECT  1088400.0 600000.0 1098600.0 586200.0 ;
      RECT  1088400.0 600000.0 1098600.0 613800.0 ;
      RECT  1088400.0 627600.0 1098600.0 613800.0 ;
      RECT  1088400.0 627600.0 1098600.0 641400.0 ;
      RECT  1088400.0 655200.0 1098600.0 641400.0 ;
      RECT  1088400.0 655200.0 1098600.0 669000.0 ;
      RECT  1088400.0 682800.0 1098600.0 669000.0 ;
      RECT  1088400.0 682800.0 1098600.0 696600.0 ;
      RECT  1088400.0 710400.0 1098600.0 696600.0 ;
      RECT  1088400.0 710400.0 1098600.0 724200.0 ;
      RECT  1088400.0 738000.0 1098600.0 724200.0 ;
      RECT  1088400.0 738000.0 1098600.0 751800.0 ;
      RECT  1088400.0 765600.0 1098600.0 751800.0 ;
      RECT  1088400.0 765600.0 1098600.0 779400.0 ;
      RECT  1088400.0 793200.0 1098600.0 779400.0 ;
      RECT  1088400.0 793200.0 1098600.0 807000.0 ;
      RECT  1088400.0 820800.0 1098600.0 807000.0 ;
      RECT  1088400.0 820800.0 1098600.0 834600.0 ;
      RECT  1088400.0 848400.0 1098600.0 834600.0 ;
      RECT  1088400.0 848400.0 1098600.0 862200.0 ;
      RECT  1088400.0 876000.0 1098600.0 862200.0 ;
      RECT  1088400.0 876000.0 1098600.0 889800.0 ;
      RECT  1088400.0 903600.0 1098600.0 889800.0 ;
      RECT  1088400.0 903600.0 1098600.0 917400.0 ;
      RECT  1088400.0 931200.0 1098600.0 917400.0 ;
      RECT  1088400.0 931200.0 1098600.0 945000.0 ;
      RECT  1088400.0 958800.0 1098600.0 945000.0 ;
      RECT  1088400.0 958800.0 1098600.0 972600.0 ;
      RECT  1088400.0 986400.0 1098600.0 972600.0 ;
      RECT  1088400.0 986400.0 1098600.0 1000200.0 ;
      RECT  1088400.0 1014000.0 1098600.0 1000200.0 ;
      RECT  1088400.0 1014000.0 1098600.0 1027800.0 ;
      RECT  1088400.0 1041600.0 1098600.0 1027800.0 ;
      RECT  1088400.0 1041600.0 1098600.0 1055400.0 ;
      RECT  1088400.0 1069200.0 1098600.0 1055400.0 ;
      RECT  1088400.0 1069200.0 1098600.0 1083000.0 ;
      RECT  1088400.0 1096800.0 1098600.0 1083000.0 ;
      RECT  1088400.0 1096800.0 1098600.0 1110600.0 ;
      RECT  1088400.0 1124400.0 1098600.0 1110600.0 ;
      RECT  1088400.0 1124400.0 1098600.0 1138200.0 ;
      RECT  1088400.0 1152000.0 1098600.0 1138200.0 ;
      RECT  1088400.0 1152000.0 1098600.0 1165800.0 ;
      RECT  1088400.0 1179600.0 1098600.0 1165800.0 ;
      RECT  1088400.0 1179600.0 1098600.0 1193400.0 ;
      RECT  1088400.0 1207200.0 1098600.0 1193400.0 ;
      RECT  1088400.0 1207200.0 1098600.0 1221000.0 ;
      RECT  1088400.0 1234800.0 1098600.0 1221000.0 ;
      RECT  1088400.0 1234800.0 1098600.0 1248600.0 ;
      RECT  1088400.0 1262400.0 1098600.0 1248600.0 ;
      RECT  1088400.0 1262400.0 1098600.0 1276200.0 ;
      RECT  1088400.0 1290000.0 1098600.0 1276200.0 ;
      RECT  1088400.0 1290000.0 1098600.0 1303800.0 ;
      RECT  1088400.0 1317600.0 1098600.0 1303800.0 ;
      RECT  1088400.0 1317600.0 1098600.0 1331400.0 ;
      RECT  1088400.0 1345200.0 1098600.0 1331400.0 ;
      RECT  1088400.0 1345200.0 1098600.0 1359000.0 ;
      RECT  1088400.0 1372800.0 1098600.0 1359000.0 ;
      RECT  1088400.0 1372800.0 1098600.0 1386600.0 ;
      RECT  1088400.0 1400400.0 1098600.0 1386600.0 ;
      RECT  1088400.0 1400400.0 1098600.0 1414200.0 ;
      RECT  1088400.0 1428000.0 1098600.0 1414200.0 ;
      RECT  1088400.0 1428000.0 1098600.0 1441800.0 ;
      RECT  1088400.0 1455600.0 1098600.0 1441800.0 ;
      RECT  1088400.0 1455600.0 1098600.0 1469400.0 ;
      RECT  1088400.0 1483200.0 1098600.0 1469400.0 ;
      RECT  1088400.0 1483200.0 1098600.0 1497000.0 ;
      RECT  1088400.0 1510800.0 1098600.0 1497000.0 ;
      RECT  1088400.0 1510800.0 1098600.0 1524600.0 ;
      RECT  1088400.0 1538400.0 1098600.0 1524600.0 ;
      RECT  1088400.0 1538400.0 1098600.0 1552200.0 ;
      RECT  1088400.0 1566000.0 1098600.0 1552200.0 ;
      RECT  1088400.0 1566000.0 1098600.0 1579800.0 ;
      RECT  1088400.0 1593600.0 1098600.0 1579800.0 ;
      RECT  1088400.0 1593600.0 1098600.0 1607400.0 ;
      RECT  1088400.0 1621200.0 1098600.0 1607400.0 ;
      RECT  1088400.0 1621200.0 1098600.0 1635000.0 ;
      RECT  1088400.0 1648800.0 1098600.0 1635000.0 ;
      RECT  1088400.0 1648800.0 1098600.0 1662600.0 ;
      RECT  1088400.0 1676400.0 1098600.0 1662600.0 ;
      RECT  1088400.0 1676400.0 1098600.0 1690200.0 ;
      RECT  1088400.0 1704000.0 1098600.0 1690200.0 ;
      RECT  1088400.0 1704000.0 1098600.0 1717800.0 ;
      RECT  1088400.0 1731600.0 1098600.0 1717800.0 ;
      RECT  1088400.0 1731600.0 1098600.0 1745400.0 ;
      RECT  1088400.0 1759200.0 1098600.0 1745400.0 ;
      RECT  1088400.0 1759200.0 1098600.0 1773000.0 ;
      RECT  1088400.0 1786800.0 1098600.0 1773000.0 ;
      RECT  1088400.0 1786800.0 1098600.0 1800600.0 ;
      RECT  1088400.0 1814400.0 1098600.0 1800600.0 ;
      RECT  1088400.0 1814400.0 1098600.0 1828200.0 ;
      RECT  1088400.0 1842000.0 1098600.0 1828200.0 ;
      RECT  1088400.0 1842000.0 1098600.0 1855800.0 ;
      RECT  1088400.0 1869600.0 1098600.0 1855800.0 ;
      RECT  1088400.0 1869600.0 1098600.0 1883400.0 ;
      RECT  1088400.0 1897200.0 1098600.0 1883400.0 ;
      RECT  1088400.0 1897200.0 1098600.0 1911000.0 ;
      RECT  1088400.0 1924800.0 1098600.0 1911000.0 ;
      RECT  1088400.0 1924800.0 1098600.0 1938600.0 ;
      RECT  1088400.0 1952400.0 1098600.0 1938600.0 ;
      RECT  1088400.0 1952400.0 1098600.0 1966200.0 ;
      RECT  1088400.0 1980000.0 1098600.0 1966200.0 ;
      RECT  1088400.0 1980000.0 1098600.0 1993800.0 ;
      RECT  1088400.0 2007600.0 1098600.0 1993800.0 ;
      RECT  1088400.0 2007600.0 1098600.0 2021400.0 ;
      RECT  1088400.0 2035200.0 1098600.0 2021400.0 ;
      RECT  1088400.0 2035200.0 1098600.0 2049000.0 ;
      RECT  1088400.0 2062800.0 1098600.0 2049000.0 ;
      RECT  1088400.0 2062800.0 1098600.0 2076600.0 ;
      RECT  1088400.0 2090400.0 1098600.0 2076600.0 ;
      RECT  1088400.0 2090400.0 1098600.0 2104200.0 ;
      RECT  1088400.0 2118000.0 1098600.0 2104200.0 ;
      RECT  1088400.0 2118000.0 1098600.0 2131800.0 ;
      RECT  1088400.0 2145600.0 1098600.0 2131800.0 ;
      RECT  1098600.0 379200.0 1108800.0 393000.0 ;
      RECT  1098600.0 406800.0 1108800.0 393000.0 ;
      RECT  1098600.0 406800.0 1108800.0 420600.0 ;
      RECT  1098600.0 434400.0 1108800.0 420600.0 ;
      RECT  1098600.0 434400.0 1108800.0 448200.0 ;
      RECT  1098600.0 462000.0 1108800.0 448200.0 ;
      RECT  1098600.0 462000.0 1108800.0 475800.0 ;
      RECT  1098600.0 489600.0 1108800.0 475800.0 ;
      RECT  1098600.0 489600.0 1108800.0 503400.0 ;
      RECT  1098600.0 517200.0 1108800.0 503400.0 ;
      RECT  1098600.0 517200.0 1108800.0 531000.0 ;
      RECT  1098600.0 544800.0 1108800.0 531000.0 ;
      RECT  1098600.0 544800.0 1108800.0 558600.0 ;
      RECT  1098600.0 572400.0 1108800.0 558600.0 ;
      RECT  1098600.0 572400.0 1108800.0 586200.0 ;
      RECT  1098600.0 600000.0 1108800.0 586200.0 ;
      RECT  1098600.0 600000.0 1108800.0 613800.0 ;
      RECT  1098600.0 627600.0 1108800.0 613800.0 ;
      RECT  1098600.0 627600.0 1108800.0 641400.0 ;
      RECT  1098600.0 655200.0 1108800.0 641400.0 ;
      RECT  1098600.0 655200.0 1108800.0 669000.0 ;
      RECT  1098600.0 682800.0 1108800.0 669000.0 ;
      RECT  1098600.0 682800.0 1108800.0 696600.0 ;
      RECT  1098600.0 710400.0 1108800.0 696600.0 ;
      RECT  1098600.0 710400.0 1108800.0 724200.0 ;
      RECT  1098600.0 738000.0 1108800.0 724200.0 ;
      RECT  1098600.0 738000.0 1108800.0 751800.0 ;
      RECT  1098600.0 765600.0 1108800.0 751800.0 ;
      RECT  1098600.0 765600.0 1108800.0 779400.0 ;
      RECT  1098600.0 793200.0 1108800.0 779400.0 ;
      RECT  1098600.0 793200.0 1108800.0 807000.0 ;
      RECT  1098600.0 820800.0 1108800.0 807000.0 ;
      RECT  1098600.0 820800.0 1108800.0 834600.0 ;
      RECT  1098600.0 848400.0 1108800.0 834600.0 ;
      RECT  1098600.0 848400.0 1108800.0 862200.0 ;
      RECT  1098600.0 876000.0 1108800.0 862200.0 ;
      RECT  1098600.0 876000.0 1108800.0 889800.0 ;
      RECT  1098600.0 903600.0 1108800.0 889800.0 ;
      RECT  1098600.0 903600.0 1108800.0 917400.0 ;
      RECT  1098600.0 931200.0 1108800.0 917400.0 ;
      RECT  1098600.0 931200.0 1108800.0 945000.0 ;
      RECT  1098600.0 958800.0 1108800.0 945000.0 ;
      RECT  1098600.0 958800.0 1108800.0 972600.0 ;
      RECT  1098600.0 986400.0 1108800.0 972600.0 ;
      RECT  1098600.0 986400.0 1108800.0 1000200.0 ;
      RECT  1098600.0 1014000.0 1108800.0 1000200.0 ;
      RECT  1098600.0 1014000.0 1108800.0 1027800.0 ;
      RECT  1098600.0 1041600.0 1108800.0 1027800.0 ;
      RECT  1098600.0 1041600.0 1108800.0 1055400.0 ;
      RECT  1098600.0 1069200.0 1108800.0 1055400.0 ;
      RECT  1098600.0 1069200.0 1108800.0 1083000.0 ;
      RECT  1098600.0 1096800.0 1108800.0 1083000.0 ;
      RECT  1098600.0 1096800.0 1108800.0 1110600.0 ;
      RECT  1098600.0 1124400.0 1108800.0 1110600.0 ;
      RECT  1098600.0 1124400.0 1108800.0 1138200.0 ;
      RECT  1098600.0 1152000.0 1108800.0 1138200.0 ;
      RECT  1098600.0 1152000.0 1108800.0 1165800.0 ;
      RECT  1098600.0 1179600.0 1108800.0 1165800.0 ;
      RECT  1098600.0 1179600.0 1108800.0 1193400.0 ;
      RECT  1098600.0 1207200.0 1108800.0 1193400.0 ;
      RECT  1098600.0 1207200.0 1108800.0 1221000.0 ;
      RECT  1098600.0 1234800.0 1108800.0 1221000.0 ;
      RECT  1098600.0 1234800.0 1108800.0 1248600.0 ;
      RECT  1098600.0 1262400.0 1108800.0 1248600.0 ;
      RECT  1098600.0 1262400.0 1108800.0 1276200.0 ;
      RECT  1098600.0 1290000.0 1108800.0 1276200.0 ;
      RECT  1098600.0 1290000.0 1108800.0 1303800.0 ;
      RECT  1098600.0 1317600.0 1108800.0 1303800.0 ;
      RECT  1098600.0 1317600.0 1108800.0 1331400.0 ;
      RECT  1098600.0 1345200.0 1108800.0 1331400.0 ;
      RECT  1098600.0 1345200.0 1108800.0 1359000.0 ;
      RECT  1098600.0 1372800.0 1108800.0 1359000.0 ;
      RECT  1098600.0 1372800.0 1108800.0 1386600.0 ;
      RECT  1098600.0 1400400.0 1108800.0 1386600.0 ;
      RECT  1098600.0 1400400.0 1108800.0 1414200.0 ;
      RECT  1098600.0 1428000.0 1108800.0 1414200.0 ;
      RECT  1098600.0 1428000.0 1108800.0 1441800.0 ;
      RECT  1098600.0 1455600.0 1108800.0 1441800.0 ;
      RECT  1098600.0 1455600.0 1108800.0 1469400.0 ;
      RECT  1098600.0 1483200.0 1108800.0 1469400.0 ;
      RECT  1098600.0 1483200.0 1108800.0 1497000.0 ;
      RECT  1098600.0 1510800.0 1108800.0 1497000.0 ;
      RECT  1098600.0 1510800.0 1108800.0 1524600.0 ;
      RECT  1098600.0 1538400.0 1108800.0 1524600.0 ;
      RECT  1098600.0 1538400.0 1108800.0 1552200.0 ;
      RECT  1098600.0 1566000.0 1108800.0 1552200.0 ;
      RECT  1098600.0 1566000.0 1108800.0 1579800.0 ;
      RECT  1098600.0 1593600.0 1108800.0 1579800.0 ;
      RECT  1098600.0 1593600.0 1108800.0 1607400.0 ;
      RECT  1098600.0 1621200.0 1108800.0 1607400.0 ;
      RECT  1098600.0 1621200.0 1108800.0 1635000.0 ;
      RECT  1098600.0 1648800.0 1108800.0 1635000.0 ;
      RECT  1098600.0 1648800.0 1108800.0 1662600.0 ;
      RECT  1098600.0 1676400.0 1108800.0 1662600.0 ;
      RECT  1098600.0 1676400.0 1108800.0 1690200.0 ;
      RECT  1098600.0 1704000.0 1108800.0 1690200.0 ;
      RECT  1098600.0 1704000.0 1108800.0 1717800.0 ;
      RECT  1098600.0 1731600.0 1108800.0 1717800.0 ;
      RECT  1098600.0 1731600.0 1108800.0 1745400.0 ;
      RECT  1098600.0 1759200.0 1108800.0 1745400.0 ;
      RECT  1098600.0 1759200.0 1108800.0 1773000.0 ;
      RECT  1098600.0 1786800.0 1108800.0 1773000.0 ;
      RECT  1098600.0 1786800.0 1108800.0 1800600.0 ;
      RECT  1098600.0 1814400.0 1108800.0 1800600.0 ;
      RECT  1098600.0 1814400.0 1108800.0 1828200.0 ;
      RECT  1098600.0 1842000.0 1108800.0 1828200.0 ;
      RECT  1098600.0 1842000.0 1108800.0 1855800.0 ;
      RECT  1098600.0 1869600.0 1108800.0 1855800.0 ;
      RECT  1098600.0 1869600.0 1108800.0 1883400.0 ;
      RECT  1098600.0 1897200.0 1108800.0 1883400.0 ;
      RECT  1098600.0 1897200.0 1108800.0 1911000.0 ;
      RECT  1098600.0 1924800.0 1108800.0 1911000.0 ;
      RECT  1098600.0 1924800.0 1108800.0 1938600.0 ;
      RECT  1098600.0 1952400.0 1108800.0 1938600.0 ;
      RECT  1098600.0 1952400.0 1108800.0 1966200.0 ;
      RECT  1098600.0 1980000.0 1108800.0 1966200.0 ;
      RECT  1098600.0 1980000.0 1108800.0 1993800.0 ;
      RECT  1098600.0 2007600.0 1108800.0 1993800.0 ;
      RECT  1098600.0 2007600.0 1108800.0 2021400.0 ;
      RECT  1098600.0 2035200.0 1108800.0 2021400.0 ;
      RECT  1098600.0 2035200.0 1108800.0 2049000.0 ;
      RECT  1098600.0 2062800.0 1108800.0 2049000.0 ;
      RECT  1098600.0 2062800.0 1108800.0 2076600.0 ;
      RECT  1098600.0 2090400.0 1108800.0 2076600.0 ;
      RECT  1098600.0 2090400.0 1108800.0 2104200.0 ;
      RECT  1098600.0 2118000.0 1108800.0 2104200.0 ;
      RECT  1098600.0 2118000.0 1108800.0 2131800.0 ;
      RECT  1098600.0 2145600.0 1108800.0 2131800.0 ;
      RECT  1108800.0 379200.0 1119000.0 393000.0 ;
      RECT  1108800.0 406800.0 1119000.0 393000.0 ;
      RECT  1108800.0 406800.0 1119000.0 420600.0 ;
      RECT  1108800.0 434400.0 1119000.0 420600.0 ;
      RECT  1108800.0 434400.0 1119000.0 448200.0 ;
      RECT  1108800.0 462000.0 1119000.0 448200.0 ;
      RECT  1108800.0 462000.0 1119000.0 475800.0 ;
      RECT  1108800.0 489600.0 1119000.0 475800.0 ;
      RECT  1108800.0 489600.0 1119000.0 503400.0 ;
      RECT  1108800.0 517200.0 1119000.0 503400.0 ;
      RECT  1108800.0 517200.0 1119000.0 531000.0 ;
      RECT  1108800.0 544800.0 1119000.0 531000.0 ;
      RECT  1108800.0 544800.0 1119000.0 558600.0 ;
      RECT  1108800.0 572400.0 1119000.0 558600.0 ;
      RECT  1108800.0 572400.0 1119000.0 586200.0 ;
      RECT  1108800.0 600000.0 1119000.0 586200.0 ;
      RECT  1108800.0 600000.0 1119000.0 613800.0 ;
      RECT  1108800.0 627600.0 1119000.0 613800.0 ;
      RECT  1108800.0 627600.0 1119000.0 641400.0 ;
      RECT  1108800.0 655200.0 1119000.0 641400.0 ;
      RECT  1108800.0 655200.0 1119000.0 669000.0 ;
      RECT  1108800.0 682800.0 1119000.0 669000.0 ;
      RECT  1108800.0 682800.0 1119000.0 696600.0 ;
      RECT  1108800.0 710400.0 1119000.0 696600.0 ;
      RECT  1108800.0 710400.0 1119000.0 724200.0 ;
      RECT  1108800.0 738000.0 1119000.0 724200.0 ;
      RECT  1108800.0 738000.0 1119000.0 751800.0 ;
      RECT  1108800.0 765600.0 1119000.0 751800.0 ;
      RECT  1108800.0 765600.0 1119000.0 779400.0 ;
      RECT  1108800.0 793200.0 1119000.0 779400.0 ;
      RECT  1108800.0 793200.0 1119000.0 807000.0 ;
      RECT  1108800.0 820800.0 1119000.0 807000.0 ;
      RECT  1108800.0 820800.0 1119000.0 834600.0 ;
      RECT  1108800.0 848400.0 1119000.0 834600.0 ;
      RECT  1108800.0 848400.0 1119000.0 862200.0 ;
      RECT  1108800.0 876000.0 1119000.0 862200.0 ;
      RECT  1108800.0 876000.0 1119000.0 889800.0 ;
      RECT  1108800.0 903600.0 1119000.0 889800.0 ;
      RECT  1108800.0 903600.0 1119000.0 917400.0 ;
      RECT  1108800.0 931200.0 1119000.0 917400.0 ;
      RECT  1108800.0 931200.0 1119000.0 945000.0 ;
      RECT  1108800.0 958800.0 1119000.0 945000.0 ;
      RECT  1108800.0 958800.0 1119000.0 972600.0 ;
      RECT  1108800.0 986400.0 1119000.0 972600.0 ;
      RECT  1108800.0 986400.0 1119000.0 1000200.0 ;
      RECT  1108800.0 1014000.0 1119000.0 1000200.0 ;
      RECT  1108800.0 1014000.0 1119000.0 1027800.0 ;
      RECT  1108800.0 1041600.0 1119000.0 1027800.0 ;
      RECT  1108800.0 1041600.0 1119000.0 1055400.0 ;
      RECT  1108800.0 1069200.0 1119000.0 1055400.0 ;
      RECT  1108800.0 1069200.0 1119000.0 1083000.0 ;
      RECT  1108800.0 1096800.0 1119000.0 1083000.0 ;
      RECT  1108800.0 1096800.0 1119000.0 1110600.0 ;
      RECT  1108800.0 1124400.0 1119000.0 1110600.0 ;
      RECT  1108800.0 1124400.0 1119000.0 1138200.0 ;
      RECT  1108800.0 1152000.0 1119000.0 1138200.0 ;
      RECT  1108800.0 1152000.0 1119000.0 1165800.0 ;
      RECT  1108800.0 1179600.0 1119000.0 1165800.0 ;
      RECT  1108800.0 1179600.0 1119000.0 1193400.0 ;
      RECT  1108800.0 1207200.0 1119000.0 1193400.0 ;
      RECT  1108800.0 1207200.0 1119000.0 1221000.0 ;
      RECT  1108800.0 1234800.0 1119000.0 1221000.0 ;
      RECT  1108800.0 1234800.0 1119000.0 1248600.0 ;
      RECT  1108800.0 1262400.0 1119000.0 1248600.0 ;
      RECT  1108800.0 1262400.0 1119000.0 1276200.0 ;
      RECT  1108800.0 1290000.0 1119000.0 1276200.0 ;
      RECT  1108800.0 1290000.0 1119000.0 1303800.0 ;
      RECT  1108800.0 1317600.0 1119000.0 1303800.0 ;
      RECT  1108800.0 1317600.0 1119000.0 1331400.0 ;
      RECT  1108800.0 1345200.0 1119000.0 1331400.0 ;
      RECT  1108800.0 1345200.0 1119000.0 1359000.0 ;
      RECT  1108800.0 1372800.0 1119000.0 1359000.0 ;
      RECT  1108800.0 1372800.0 1119000.0 1386600.0 ;
      RECT  1108800.0 1400400.0 1119000.0 1386600.0 ;
      RECT  1108800.0 1400400.0 1119000.0 1414200.0 ;
      RECT  1108800.0 1428000.0 1119000.0 1414200.0 ;
      RECT  1108800.0 1428000.0 1119000.0 1441800.0 ;
      RECT  1108800.0 1455600.0 1119000.0 1441800.0 ;
      RECT  1108800.0 1455600.0 1119000.0 1469400.0 ;
      RECT  1108800.0 1483200.0 1119000.0 1469400.0 ;
      RECT  1108800.0 1483200.0 1119000.0 1497000.0 ;
      RECT  1108800.0 1510800.0 1119000.0 1497000.0 ;
      RECT  1108800.0 1510800.0 1119000.0 1524600.0 ;
      RECT  1108800.0 1538400.0 1119000.0 1524600.0 ;
      RECT  1108800.0 1538400.0 1119000.0 1552200.0 ;
      RECT  1108800.0 1566000.0 1119000.0 1552200.0 ;
      RECT  1108800.0 1566000.0 1119000.0 1579800.0 ;
      RECT  1108800.0 1593600.0 1119000.0 1579800.0 ;
      RECT  1108800.0 1593600.0 1119000.0 1607400.0 ;
      RECT  1108800.0 1621200.0 1119000.0 1607400.0 ;
      RECT  1108800.0 1621200.0 1119000.0 1635000.0 ;
      RECT  1108800.0 1648800.0 1119000.0 1635000.0 ;
      RECT  1108800.0 1648800.0 1119000.0 1662600.0 ;
      RECT  1108800.0 1676400.0 1119000.0 1662600.0 ;
      RECT  1108800.0 1676400.0 1119000.0 1690200.0 ;
      RECT  1108800.0 1704000.0 1119000.0 1690200.0 ;
      RECT  1108800.0 1704000.0 1119000.0 1717800.0 ;
      RECT  1108800.0 1731600.0 1119000.0 1717800.0 ;
      RECT  1108800.0 1731600.0 1119000.0 1745400.0 ;
      RECT  1108800.0 1759200.0 1119000.0 1745400.0 ;
      RECT  1108800.0 1759200.0 1119000.0 1773000.0 ;
      RECT  1108800.0 1786800.0 1119000.0 1773000.0 ;
      RECT  1108800.0 1786800.0 1119000.0 1800600.0 ;
      RECT  1108800.0 1814400.0 1119000.0 1800600.0 ;
      RECT  1108800.0 1814400.0 1119000.0 1828200.0 ;
      RECT  1108800.0 1842000.0 1119000.0 1828200.0 ;
      RECT  1108800.0 1842000.0 1119000.0 1855800.0 ;
      RECT  1108800.0 1869600.0 1119000.0 1855800.0 ;
      RECT  1108800.0 1869600.0 1119000.0 1883400.0 ;
      RECT  1108800.0 1897200.0 1119000.0 1883400.0 ;
      RECT  1108800.0 1897200.0 1119000.0 1911000.0 ;
      RECT  1108800.0 1924800.0 1119000.0 1911000.0 ;
      RECT  1108800.0 1924800.0 1119000.0 1938600.0 ;
      RECT  1108800.0 1952400.0 1119000.0 1938600.0 ;
      RECT  1108800.0 1952400.0 1119000.0 1966200.0 ;
      RECT  1108800.0 1980000.0 1119000.0 1966200.0 ;
      RECT  1108800.0 1980000.0 1119000.0 1993800.0 ;
      RECT  1108800.0 2007600.0 1119000.0 1993800.0 ;
      RECT  1108800.0 2007600.0 1119000.0 2021400.0 ;
      RECT  1108800.0 2035200.0 1119000.0 2021400.0 ;
      RECT  1108800.0 2035200.0 1119000.0 2049000.0 ;
      RECT  1108800.0 2062800.0 1119000.0 2049000.0 ;
      RECT  1108800.0 2062800.0 1119000.0 2076600.0 ;
      RECT  1108800.0 2090400.0 1119000.0 2076600.0 ;
      RECT  1108800.0 2090400.0 1119000.0 2104200.0 ;
      RECT  1108800.0 2118000.0 1119000.0 2104200.0 ;
      RECT  1108800.0 2118000.0 1119000.0 2131800.0 ;
      RECT  1108800.0 2145600.0 1119000.0 2131800.0 ;
      RECT  1119000.0 379200.0 1129200.0 393000.0 ;
      RECT  1119000.0 406800.0 1129200.0 393000.0 ;
      RECT  1119000.0 406800.0 1129200.0 420600.0 ;
      RECT  1119000.0 434400.0 1129200.0 420600.0 ;
      RECT  1119000.0 434400.0 1129200.0 448200.0 ;
      RECT  1119000.0 462000.0 1129200.0 448200.0 ;
      RECT  1119000.0 462000.0 1129200.0 475800.0 ;
      RECT  1119000.0 489600.0 1129200.0 475800.0 ;
      RECT  1119000.0 489600.0 1129200.0 503400.0 ;
      RECT  1119000.0 517200.0 1129200.0 503400.0 ;
      RECT  1119000.0 517200.0 1129200.0 531000.0 ;
      RECT  1119000.0 544800.0 1129200.0 531000.0 ;
      RECT  1119000.0 544800.0 1129200.0 558600.0 ;
      RECT  1119000.0 572400.0 1129200.0 558600.0 ;
      RECT  1119000.0 572400.0 1129200.0 586200.0 ;
      RECT  1119000.0 600000.0 1129200.0 586200.0 ;
      RECT  1119000.0 600000.0 1129200.0 613800.0 ;
      RECT  1119000.0 627600.0 1129200.0 613800.0 ;
      RECT  1119000.0 627600.0 1129200.0 641400.0 ;
      RECT  1119000.0 655200.0 1129200.0 641400.0 ;
      RECT  1119000.0 655200.0 1129200.0 669000.0 ;
      RECT  1119000.0 682800.0 1129200.0 669000.0 ;
      RECT  1119000.0 682800.0 1129200.0 696600.0 ;
      RECT  1119000.0 710400.0 1129200.0 696600.0 ;
      RECT  1119000.0 710400.0 1129200.0 724200.0 ;
      RECT  1119000.0 738000.0 1129200.0 724200.0 ;
      RECT  1119000.0 738000.0 1129200.0 751800.0 ;
      RECT  1119000.0 765600.0 1129200.0 751800.0 ;
      RECT  1119000.0 765600.0 1129200.0 779400.0 ;
      RECT  1119000.0 793200.0 1129200.0 779400.0 ;
      RECT  1119000.0 793200.0 1129200.0 807000.0 ;
      RECT  1119000.0 820800.0 1129200.0 807000.0 ;
      RECT  1119000.0 820800.0 1129200.0 834600.0 ;
      RECT  1119000.0 848400.0 1129200.0 834600.0 ;
      RECT  1119000.0 848400.0 1129200.0 862200.0 ;
      RECT  1119000.0 876000.0 1129200.0 862200.0 ;
      RECT  1119000.0 876000.0 1129200.0 889800.0 ;
      RECT  1119000.0 903600.0 1129200.0 889800.0 ;
      RECT  1119000.0 903600.0 1129200.0 917400.0 ;
      RECT  1119000.0 931200.0 1129200.0 917400.0 ;
      RECT  1119000.0 931200.0 1129200.0 945000.0 ;
      RECT  1119000.0 958800.0 1129200.0 945000.0 ;
      RECT  1119000.0 958800.0 1129200.0 972600.0 ;
      RECT  1119000.0 986400.0 1129200.0 972600.0 ;
      RECT  1119000.0 986400.0 1129200.0 1000200.0 ;
      RECT  1119000.0 1014000.0 1129200.0 1000200.0 ;
      RECT  1119000.0 1014000.0 1129200.0 1027800.0 ;
      RECT  1119000.0 1041600.0 1129200.0 1027800.0 ;
      RECT  1119000.0 1041600.0 1129200.0 1055400.0 ;
      RECT  1119000.0 1069200.0 1129200.0 1055400.0 ;
      RECT  1119000.0 1069200.0 1129200.0 1083000.0 ;
      RECT  1119000.0 1096800.0 1129200.0 1083000.0 ;
      RECT  1119000.0 1096800.0 1129200.0 1110600.0 ;
      RECT  1119000.0 1124400.0 1129200.0 1110600.0 ;
      RECT  1119000.0 1124400.0 1129200.0 1138200.0 ;
      RECT  1119000.0 1152000.0 1129200.0 1138200.0 ;
      RECT  1119000.0 1152000.0 1129200.0 1165800.0 ;
      RECT  1119000.0 1179600.0 1129200.0 1165800.0 ;
      RECT  1119000.0 1179600.0 1129200.0 1193400.0 ;
      RECT  1119000.0 1207200.0 1129200.0 1193400.0 ;
      RECT  1119000.0 1207200.0 1129200.0 1221000.0 ;
      RECT  1119000.0 1234800.0 1129200.0 1221000.0 ;
      RECT  1119000.0 1234800.0 1129200.0 1248600.0 ;
      RECT  1119000.0 1262400.0 1129200.0 1248600.0 ;
      RECT  1119000.0 1262400.0 1129200.0 1276200.0 ;
      RECT  1119000.0 1290000.0 1129200.0 1276200.0 ;
      RECT  1119000.0 1290000.0 1129200.0 1303800.0 ;
      RECT  1119000.0 1317600.0 1129200.0 1303800.0 ;
      RECT  1119000.0 1317600.0 1129200.0 1331400.0 ;
      RECT  1119000.0 1345200.0 1129200.0 1331400.0 ;
      RECT  1119000.0 1345200.0 1129200.0 1359000.0 ;
      RECT  1119000.0 1372800.0 1129200.0 1359000.0 ;
      RECT  1119000.0 1372800.0 1129200.0 1386600.0 ;
      RECT  1119000.0 1400400.0 1129200.0 1386600.0 ;
      RECT  1119000.0 1400400.0 1129200.0 1414200.0 ;
      RECT  1119000.0 1428000.0 1129200.0 1414200.0 ;
      RECT  1119000.0 1428000.0 1129200.0 1441800.0 ;
      RECT  1119000.0 1455600.0 1129200.0 1441800.0 ;
      RECT  1119000.0 1455600.0 1129200.0 1469400.0 ;
      RECT  1119000.0 1483200.0 1129200.0 1469400.0 ;
      RECT  1119000.0 1483200.0 1129200.0 1497000.0 ;
      RECT  1119000.0 1510800.0 1129200.0 1497000.0 ;
      RECT  1119000.0 1510800.0 1129200.0 1524600.0 ;
      RECT  1119000.0 1538400.0 1129200.0 1524600.0 ;
      RECT  1119000.0 1538400.0 1129200.0 1552200.0 ;
      RECT  1119000.0 1566000.0 1129200.0 1552200.0 ;
      RECT  1119000.0 1566000.0 1129200.0 1579800.0 ;
      RECT  1119000.0 1593600.0 1129200.0 1579800.0 ;
      RECT  1119000.0 1593600.0 1129200.0 1607400.0 ;
      RECT  1119000.0 1621200.0 1129200.0 1607400.0 ;
      RECT  1119000.0 1621200.0 1129200.0 1635000.0 ;
      RECT  1119000.0 1648800.0 1129200.0 1635000.0 ;
      RECT  1119000.0 1648800.0 1129200.0 1662600.0 ;
      RECT  1119000.0 1676400.0 1129200.0 1662600.0 ;
      RECT  1119000.0 1676400.0 1129200.0 1690200.0 ;
      RECT  1119000.0 1704000.0 1129200.0 1690200.0 ;
      RECT  1119000.0 1704000.0 1129200.0 1717800.0 ;
      RECT  1119000.0 1731600.0 1129200.0 1717800.0 ;
      RECT  1119000.0 1731600.0 1129200.0 1745400.0 ;
      RECT  1119000.0 1759200.0 1129200.0 1745400.0 ;
      RECT  1119000.0 1759200.0 1129200.0 1773000.0 ;
      RECT  1119000.0 1786800.0 1129200.0 1773000.0 ;
      RECT  1119000.0 1786800.0 1129200.0 1800600.0 ;
      RECT  1119000.0 1814400.0 1129200.0 1800600.0 ;
      RECT  1119000.0 1814400.0 1129200.0 1828200.0 ;
      RECT  1119000.0 1842000.0 1129200.0 1828200.0 ;
      RECT  1119000.0 1842000.0 1129200.0 1855800.0 ;
      RECT  1119000.0 1869600.0 1129200.0 1855800.0 ;
      RECT  1119000.0 1869600.0 1129200.0 1883400.0 ;
      RECT  1119000.0 1897200.0 1129200.0 1883400.0 ;
      RECT  1119000.0 1897200.0 1129200.0 1911000.0 ;
      RECT  1119000.0 1924800.0 1129200.0 1911000.0 ;
      RECT  1119000.0 1924800.0 1129200.0 1938600.0 ;
      RECT  1119000.0 1952400.0 1129200.0 1938600.0 ;
      RECT  1119000.0 1952400.0 1129200.0 1966200.0 ;
      RECT  1119000.0 1980000.0 1129200.0 1966200.0 ;
      RECT  1119000.0 1980000.0 1129200.0 1993800.0 ;
      RECT  1119000.0 2007600.0 1129200.0 1993800.0 ;
      RECT  1119000.0 2007600.0 1129200.0 2021400.0 ;
      RECT  1119000.0 2035200.0 1129200.0 2021400.0 ;
      RECT  1119000.0 2035200.0 1129200.0 2049000.0 ;
      RECT  1119000.0 2062800.0 1129200.0 2049000.0 ;
      RECT  1119000.0 2062800.0 1129200.0 2076600.0 ;
      RECT  1119000.0 2090400.0 1129200.0 2076600.0 ;
      RECT  1119000.0 2090400.0 1129200.0 2104200.0 ;
      RECT  1119000.0 2118000.0 1129200.0 2104200.0 ;
      RECT  1119000.0 2118000.0 1129200.0 2131800.0 ;
      RECT  1119000.0 2145600.0 1129200.0 2131800.0 ;
      RECT  1129200.0 379200.0 1139400.0 393000.0 ;
      RECT  1129200.0 406800.0 1139400.0 393000.0 ;
      RECT  1129200.0 406800.0 1139400.0 420600.0 ;
      RECT  1129200.0 434400.0 1139400.0 420600.0 ;
      RECT  1129200.0 434400.0 1139400.0 448200.0 ;
      RECT  1129200.0 462000.0 1139400.0 448200.0 ;
      RECT  1129200.0 462000.0 1139400.0 475800.0 ;
      RECT  1129200.0 489600.0 1139400.0 475800.0 ;
      RECT  1129200.0 489600.0 1139400.0 503400.0 ;
      RECT  1129200.0 517200.0 1139400.0 503400.0 ;
      RECT  1129200.0 517200.0 1139400.0 531000.0 ;
      RECT  1129200.0 544800.0 1139400.0 531000.0 ;
      RECT  1129200.0 544800.0 1139400.0 558600.0 ;
      RECT  1129200.0 572400.0 1139400.0 558600.0 ;
      RECT  1129200.0 572400.0 1139400.0 586200.0 ;
      RECT  1129200.0 600000.0 1139400.0 586200.0 ;
      RECT  1129200.0 600000.0 1139400.0 613800.0 ;
      RECT  1129200.0 627600.0 1139400.0 613800.0 ;
      RECT  1129200.0 627600.0 1139400.0 641400.0 ;
      RECT  1129200.0 655200.0 1139400.0 641400.0 ;
      RECT  1129200.0 655200.0 1139400.0 669000.0 ;
      RECT  1129200.0 682800.0 1139400.0 669000.0 ;
      RECT  1129200.0 682800.0 1139400.0 696600.0 ;
      RECT  1129200.0 710400.0 1139400.0 696600.0 ;
      RECT  1129200.0 710400.0 1139400.0 724200.0 ;
      RECT  1129200.0 738000.0 1139400.0 724200.0 ;
      RECT  1129200.0 738000.0 1139400.0 751800.0 ;
      RECT  1129200.0 765600.0 1139400.0 751800.0 ;
      RECT  1129200.0 765600.0 1139400.0 779400.0 ;
      RECT  1129200.0 793200.0 1139400.0 779400.0 ;
      RECT  1129200.0 793200.0 1139400.0 807000.0 ;
      RECT  1129200.0 820800.0 1139400.0 807000.0 ;
      RECT  1129200.0 820800.0 1139400.0 834600.0 ;
      RECT  1129200.0 848400.0 1139400.0 834600.0 ;
      RECT  1129200.0 848400.0 1139400.0 862200.0 ;
      RECT  1129200.0 876000.0 1139400.0 862200.0 ;
      RECT  1129200.0 876000.0 1139400.0 889800.0 ;
      RECT  1129200.0 903600.0 1139400.0 889800.0 ;
      RECT  1129200.0 903600.0 1139400.0 917400.0 ;
      RECT  1129200.0 931200.0 1139400.0 917400.0 ;
      RECT  1129200.0 931200.0 1139400.0 945000.0 ;
      RECT  1129200.0 958800.0 1139400.0 945000.0 ;
      RECT  1129200.0 958800.0 1139400.0 972600.0 ;
      RECT  1129200.0 986400.0 1139400.0 972600.0 ;
      RECT  1129200.0 986400.0 1139400.0 1000200.0 ;
      RECT  1129200.0 1014000.0 1139400.0 1000200.0 ;
      RECT  1129200.0 1014000.0 1139400.0 1027800.0 ;
      RECT  1129200.0 1041600.0 1139400.0 1027800.0 ;
      RECT  1129200.0 1041600.0 1139400.0 1055400.0 ;
      RECT  1129200.0 1069200.0 1139400.0 1055400.0 ;
      RECT  1129200.0 1069200.0 1139400.0 1083000.0 ;
      RECT  1129200.0 1096800.0 1139400.0 1083000.0 ;
      RECT  1129200.0 1096800.0 1139400.0 1110600.0 ;
      RECT  1129200.0 1124400.0 1139400.0 1110600.0 ;
      RECT  1129200.0 1124400.0 1139400.0 1138200.0 ;
      RECT  1129200.0 1152000.0 1139400.0 1138200.0 ;
      RECT  1129200.0 1152000.0 1139400.0 1165800.0 ;
      RECT  1129200.0 1179600.0 1139400.0 1165800.0 ;
      RECT  1129200.0 1179600.0 1139400.0 1193400.0 ;
      RECT  1129200.0 1207200.0 1139400.0 1193400.0 ;
      RECT  1129200.0 1207200.0 1139400.0 1221000.0 ;
      RECT  1129200.0 1234800.0 1139400.0 1221000.0 ;
      RECT  1129200.0 1234800.0 1139400.0 1248600.0 ;
      RECT  1129200.0 1262400.0 1139400.0 1248600.0 ;
      RECT  1129200.0 1262400.0 1139400.0 1276200.0 ;
      RECT  1129200.0 1290000.0 1139400.0 1276200.0 ;
      RECT  1129200.0 1290000.0 1139400.0 1303800.0 ;
      RECT  1129200.0 1317600.0 1139400.0 1303800.0 ;
      RECT  1129200.0 1317600.0 1139400.0 1331400.0 ;
      RECT  1129200.0 1345200.0 1139400.0 1331400.0 ;
      RECT  1129200.0 1345200.0 1139400.0 1359000.0 ;
      RECT  1129200.0 1372800.0 1139400.0 1359000.0 ;
      RECT  1129200.0 1372800.0 1139400.0 1386600.0 ;
      RECT  1129200.0 1400400.0 1139400.0 1386600.0 ;
      RECT  1129200.0 1400400.0 1139400.0 1414200.0 ;
      RECT  1129200.0 1428000.0 1139400.0 1414200.0 ;
      RECT  1129200.0 1428000.0 1139400.0 1441800.0 ;
      RECT  1129200.0 1455600.0 1139400.0 1441800.0 ;
      RECT  1129200.0 1455600.0 1139400.0 1469400.0 ;
      RECT  1129200.0 1483200.0 1139400.0 1469400.0 ;
      RECT  1129200.0 1483200.0 1139400.0 1497000.0 ;
      RECT  1129200.0 1510800.0 1139400.0 1497000.0 ;
      RECT  1129200.0 1510800.0 1139400.0 1524600.0 ;
      RECT  1129200.0 1538400.0 1139400.0 1524600.0 ;
      RECT  1129200.0 1538400.0 1139400.0 1552200.0 ;
      RECT  1129200.0 1566000.0 1139400.0 1552200.0 ;
      RECT  1129200.0 1566000.0 1139400.0 1579800.0 ;
      RECT  1129200.0 1593600.0 1139400.0 1579800.0 ;
      RECT  1129200.0 1593600.0 1139400.0 1607400.0 ;
      RECT  1129200.0 1621200.0 1139400.0 1607400.0 ;
      RECT  1129200.0 1621200.0 1139400.0 1635000.0 ;
      RECT  1129200.0 1648800.0 1139400.0 1635000.0 ;
      RECT  1129200.0 1648800.0 1139400.0 1662600.0 ;
      RECT  1129200.0 1676400.0 1139400.0 1662600.0 ;
      RECT  1129200.0 1676400.0 1139400.0 1690200.0 ;
      RECT  1129200.0 1704000.0 1139400.0 1690200.0 ;
      RECT  1129200.0 1704000.0 1139400.0 1717800.0 ;
      RECT  1129200.0 1731600.0 1139400.0 1717800.0 ;
      RECT  1129200.0 1731600.0 1139400.0 1745400.0 ;
      RECT  1129200.0 1759200.0 1139400.0 1745400.0 ;
      RECT  1129200.0 1759200.0 1139400.0 1773000.0 ;
      RECT  1129200.0 1786800.0 1139400.0 1773000.0 ;
      RECT  1129200.0 1786800.0 1139400.0 1800600.0 ;
      RECT  1129200.0 1814400.0 1139400.0 1800600.0 ;
      RECT  1129200.0 1814400.0 1139400.0 1828200.0 ;
      RECT  1129200.0 1842000.0 1139400.0 1828200.0 ;
      RECT  1129200.0 1842000.0 1139400.0 1855800.0 ;
      RECT  1129200.0 1869600.0 1139400.0 1855800.0 ;
      RECT  1129200.0 1869600.0 1139400.0 1883400.0 ;
      RECT  1129200.0 1897200.0 1139400.0 1883400.0 ;
      RECT  1129200.0 1897200.0 1139400.0 1911000.0 ;
      RECT  1129200.0 1924800.0 1139400.0 1911000.0 ;
      RECT  1129200.0 1924800.0 1139400.0 1938600.0 ;
      RECT  1129200.0 1952400.0 1139400.0 1938600.0 ;
      RECT  1129200.0 1952400.0 1139400.0 1966200.0 ;
      RECT  1129200.0 1980000.0 1139400.0 1966200.0 ;
      RECT  1129200.0 1980000.0 1139400.0 1993800.0 ;
      RECT  1129200.0 2007600.0 1139400.0 1993800.0 ;
      RECT  1129200.0 2007600.0 1139400.0 2021400.0 ;
      RECT  1129200.0 2035200.0 1139400.0 2021400.0 ;
      RECT  1129200.0 2035200.0 1139400.0 2049000.0 ;
      RECT  1129200.0 2062800.0 1139400.0 2049000.0 ;
      RECT  1129200.0 2062800.0 1139400.0 2076600.0 ;
      RECT  1129200.0 2090400.0 1139400.0 2076600.0 ;
      RECT  1129200.0 2090400.0 1139400.0 2104200.0 ;
      RECT  1129200.0 2118000.0 1139400.0 2104200.0 ;
      RECT  1129200.0 2118000.0 1139400.0 2131800.0 ;
      RECT  1129200.0 2145600.0 1139400.0 2131800.0 ;
      RECT  1139400.0 379200.0 1149600.0 393000.0 ;
      RECT  1139400.0 406800.0 1149600.0 393000.0 ;
      RECT  1139400.0 406800.0 1149600.0 420600.0 ;
      RECT  1139400.0 434400.0 1149600.0 420600.0 ;
      RECT  1139400.0 434400.0 1149600.0 448200.0 ;
      RECT  1139400.0 462000.0 1149600.0 448200.0 ;
      RECT  1139400.0 462000.0 1149600.0 475800.0 ;
      RECT  1139400.0 489600.0 1149600.0 475800.0 ;
      RECT  1139400.0 489600.0 1149600.0 503400.0 ;
      RECT  1139400.0 517200.0 1149600.0 503400.0 ;
      RECT  1139400.0 517200.0 1149600.0 531000.0 ;
      RECT  1139400.0 544800.0 1149600.0 531000.0 ;
      RECT  1139400.0 544800.0 1149600.0 558600.0 ;
      RECT  1139400.0 572400.0 1149600.0 558600.0 ;
      RECT  1139400.0 572400.0 1149600.0 586200.0 ;
      RECT  1139400.0 600000.0 1149600.0 586200.0 ;
      RECT  1139400.0 600000.0 1149600.0 613800.0 ;
      RECT  1139400.0 627600.0 1149600.0 613800.0 ;
      RECT  1139400.0 627600.0 1149600.0 641400.0 ;
      RECT  1139400.0 655200.0 1149600.0 641400.0 ;
      RECT  1139400.0 655200.0 1149600.0 669000.0 ;
      RECT  1139400.0 682800.0 1149600.0 669000.0 ;
      RECT  1139400.0 682800.0 1149600.0 696600.0 ;
      RECT  1139400.0 710400.0 1149600.0 696600.0 ;
      RECT  1139400.0 710400.0 1149600.0 724200.0 ;
      RECT  1139400.0 738000.0 1149600.0 724200.0 ;
      RECT  1139400.0 738000.0 1149600.0 751800.0 ;
      RECT  1139400.0 765600.0 1149600.0 751800.0 ;
      RECT  1139400.0 765600.0 1149600.0 779400.0 ;
      RECT  1139400.0 793200.0 1149600.0 779400.0 ;
      RECT  1139400.0 793200.0 1149600.0 807000.0 ;
      RECT  1139400.0 820800.0 1149600.0 807000.0 ;
      RECT  1139400.0 820800.0 1149600.0 834600.0 ;
      RECT  1139400.0 848400.0 1149600.0 834600.0 ;
      RECT  1139400.0 848400.0 1149600.0 862200.0 ;
      RECT  1139400.0 876000.0 1149600.0 862200.0 ;
      RECT  1139400.0 876000.0 1149600.0 889800.0 ;
      RECT  1139400.0 903600.0 1149600.0 889800.0 ;
      RECT  1139400.0 903600.0 1149600.0 917400.0 ;
      RECT  1139400.0 931200.0 1149600.0 917400.0 ;
      RECT  1139400.0 931200.0 1149600.0 945000.0 ;
      RECT  1139400.0 958800.0 1149600.0 945000.0 ;
      RECT  1139400.0 958800.0 1149600.0 972600.0 ;
      RECT  1139400.0 986400.0 1149600.0 972600.0 ;
      RECT  1139400.0 986400.0 1149600.0 1000200.0 ;
      RECT  1139400.0 1014000.0 1149600.0 1000200.0 ;
      RECT  1139400.0 1014000.0 1149600.0 1027800.0 ;
      RECT  1139400.0 1041600.0 1149600.0 1027800.0 ;
      RECT  1139400.0 1041600.0 1149600.0 1055400.0 ;
      RECT  1139400.0 1069200.0 1149600.0 1055400.0 ;
      RECT  1139400.0 1069200.0 1149600.0 1083000.0 ;
      RECT  1139400.0 1096800.0 1149600.0 1083000.0 ;
      RECT  1139400.0 1096800.0 1149600.0 1110600.0 ;
      RECT  1139400.0 1124400.0 1149600.0 1110600.0 ;
      RECT  1139400.0 1124400.0 1149600.0 1138200.0 ;
      RECT  1139400.0 1152000.0 1149600.0 1138200.0 ;
      RECT  1139400.0 1152000.0 1149600.0 1165800.0 ;
      RECT  1139400.0 1179600.0 1149600.0 1165800.0 ;
      RECT  1139400.0 1179600.0 1149600.0 1193400.0 ;
      RECT  1139400.0 1207200.0 1149600.0 1193400.0 ;
      RECT  1139400.0 1207200.0 1149600.0 1221000.0 ;
      RECT  1139400.0 1234800.0 1149600.0 1221000.0 ;
      RECT  1139400.0 1234800.0 1149600.0 1248600.0 ;
      RECT  1139400.0 1262400.0 1149600.0 1248600.0 ;
      RECT  1139400.0 1262400.0 1149600.0 1276200.0 ;
      RECT  1139400.0 1290000.0 1149600.0 1276200.0 ;
      RECT  1139400.0 1290000.0 1149600.0 1303800.0 ;
      RECT  1139400.0 1317600.0 1149600.0 1303800.0 ;
      RECT  1139400.0 1317600.0 1149600.0 1331400.0 ;
      RECT  1139400.0 1345200.0 1149600.0 1331400.0 ;
      RECT  1139400.0 1345200.0 1149600.0 1359000.0 ;
      RECT  1139400.0 1372800.0 1149600.0 1359000.0 ;
      RECT  1139400.0 1372800.0 1149600.0 1386600.0 ;
      RECT  1139400.0 1400400.0 1149600.0 1386600.0 ;
      RECT  1139400.0 1400400.0 1149600.0 1414200.0 ;
      RECT  1139400.0 1428000.0 1149600.0 1414200.0 ;
      RECT  1139400.0 1428000.0 1149600.0 1441800.0 ;
      RECT  1139400.0 1455600.0 1149600.0 1441800.0 ;
      RECT  1139400.0 1455600.0 1149600.0 1469400.0 ;
      RECT  1139400.0 1483200.0 1149600.0 1469400.0 ;
      RECT  1139400.0 1483200.0 1149600.0 1497000.0 ;
      RECT  1139400.0 1510800.0 1149600.0 1497000.0 ;
      RECT  1139400.0 1510800.0 1149600.0 1524600.0 ;
      RECT  1139400.0 1538400.0 1149600.0 1524600.0 ;
      RECT  1139400.0 1538400.0 1149600.0 1552200.0 ;
      RECT  1139400.0 1566000.0 1149600.0 1552200.0 ;
      RECT  1139400.0 1566000.0 1149600.0 1579800.0 ;
      RECT  1139400.0 1593600.0 1149600.0 1579800.0 ;
      RECT  1139400.0 1593600.0 1149600.0 1607400.0 ;
      RECT  1139400.0 1621200.0 1149600.0 1607400.0 ;
      RECT  1139400.0 1621200.0 1149600.0 1635000.0 ;
      RECT  1139400.0 1648800.0 1149600.0 1635000.0 ;
      RECT  1139400.0 1648800.0 1149600.0 1662600.0 ;
      RECT  1139400.0 1676400.0 1149600.0 1662600.0 ;
      RECT  1139400.0 1676400.0 1149600.0 1690200.0 ;
      RECT  1139400.0 1704000.0 1149600.0 1690200.0 ;
      RECT  1139400.0 1704000.0 1149600.0 1717800.0 ;
      RECT  1139400.0 1731600.0 1149600.0 1717800.0 ;
      RECT  1139400.0 1731600.0 1149600.0 1745400.0 ;
      RECT  1139400.0 1759200.0 1149600.0 1745400.0 ;
      RECT  1139400.0 1759200.0 1149600.0 1773000.0 ;
      RECT  1139400.0 1786800.0 1149600.0 1773000.0 ;
      RECT  1139400.0 1786800.0 1149600.0 1800600.0 ;
      RECT  1139400.0 1814400.0 1149600.0 1800600.0 ;
      RECT  1139400.0 1814400.0 1149600.0 1828200.0 ;
      RECT  1139400.0 1842000.0 1149600.0 1828200.0 ;
      RECT  1139400.0 1842000.0 1149600.0 1855800.0 ;
      RECT  1139400.0 1869600.0 1149600.0 1855800.0 ;
      RECT  1139400.0 1869600.0 1149600.0 1883400.0 ;
      RECT  1139400.0 1897200.0 1149600.0 1883400.0 ;
      RECT  1139400.0 1897200.0 1149600.0 1911000.0 ;
      RECT  1139400.0 1924800.0 1149600.0 1911000.0 ;
      RECT  1139400.0 1924800.0 1149600.0 1938600.0 ;
      RECT  1139400.0 1952400.0 1149600.0 1938600.0 ;
      RECT  1139400.0 1952400.0 1149600.0 1966200.0 ;
      RECT  1139400.0 1980000.0 1149600.0 1966200.0 ;
      RECT  1139400.0 1980000.0 1149600.0 1993800.0 ;
      RECT  1139400.0 2007600.0 1149600.0 1993800.0 ;
      RECT  1139400.0 2007600.0 1149600.0 2021400.0 ;
      RECT  1139400.0 2035200.0 1149600.0 2021400.0 ;
      RECT  1139400.0 2035200.0 1149600.0 2049000.0 ;
      RECT  1139400.0 2062800.0 1149600.0 2049000.0 ;
      RECT  1139400.0 2062800.0 1149600.0 2076600.0 ;
      RECT  1139400.0 2090400.0 1149600.0 2076600.0 ;
      RECT  1139400.0 2090400.0 1149600.0 2104200.0 ;
      RECT  1139400.0 2118000.0 1149600.0 2104200.0 ;
      RECT  1139400.0 2118000.0 1149600.0 2131800.0 ;
      RECT  1139400.0 2145600.0 1149600.0 2131800.0 ;
      RECT  1149600.0 379200.0 1159800.0 393000.0 ;
      RECT  1149600.0 406800.0 1159800.0 393000.0 ;
      RECT  1149600.0 406800.0 1159800.0 420600.0 ;
      RECT  1149600.0 434400.0 1159800.0 420600.0 ;
      RECT  1149600.0 434400.0 1159800.0 448200.0 ;
      RECT  1149600.0 462000.0 1159800.0 448200.0 ;
      RECT  1149600.0 462000.0 1159800.0 475800.0 ;
      RECT  1149600.0 489600.0 1159800.0 475800.0 ;
      RECT  1149600.0 489600.0 1159800.0 503400.0 ;
      RECT  1149600.0 517200.0 1159800.0 503400.0 ;
      RECT  1149600.0 517200.0 1159800.0 531000.0 ;
      RECT  1149600.0 544800.0 1159800.0 531000.0 ;
      RECT  1149600.0 544800.0 1159800.0 558600.0 ;
      RECT  1149600.0 572400.0 1159800.0 558600.0 ;
      RECT  1149600.0 572400.0 1159800.0 586200.0 ;
      RECT  1149600.0 600000.0 1159800.0 586200.0 ;
      RECT  1149600.0 600000.0 1159800.0 613800.0 ;
      RECT  1149600.0 627600.0 1159800.0 613800.0 ;
      RECT  1149600.0 627600.0 1159800.0 641400.0 ;
      RECT  1149600.0 655200.0 1159800.0 641400.0 ;
      RECT  1149600.0 655200.0 1159800.0 669000.0 ;
      RECT  1149600.0 682800.0 1159800.0 669000.0 ;
      RECT  1149600.0 682800.0 1159800.0 696600.0 ;
      RECT  1149600.0 710400.0 1159800.0 696600.0 ;
      RECT  1149600.0 710400.0 1159800.0 724200.0 ;
      RECT  1149600.0 738000.0 1159800.0 724200.0 ;
      RECT  1149600.0 738000.0 1159800.0 751800.0 ;
      RECT  1149600.0 765600.0 1159800.0 751800.0 ;
      RECT  1149600.0 765600.0 1159800.0 779400.0 ;
      RECT  1149600.0 793200.0 1159800.0 779400.0 ;
      RECT  1149600.0 793200.0 1159800.0 807000.0 ;
      RECT  1149600.0 820800.0 1159800.0 807000.0 ;
      RECT  1149600.0 820800.0 1159800.0 834600.0 ;
      RECT  1149600.0 848400.0 1159800.0 834600.0 ;
      RECT  1149600.0 848400.0 1159800.0 862200.0 ;
      RECT  1149600.0 876000.0 1159800.0 862200.0 ;
      RECT  1149600.0 876000.0 1159800.0 889800.0 ;
      RECT  1149600.0 903600.0 1159800.0 889800.0 ;
      RECT  1149600.0 903600.0 1159800.0 917400.0 ;
      RECT  1149600.0 931200.0 1159800.0 917400.0 ;
      RECT  1149600.0 931200.0 1159800.0 945000.0 ;
      RECT  1149600.0 958800.0 1159800.0 945000.0 ;
      RECT  1149600.0 958800.0 1159800.0 972600.0 ;
      RECT  1149600.0 986400.0 1159800.0 972600.0 ;
      RECT  1149600.0 986400.0 1159800.0 1000200.0 ;
      RECT  1149600.0 1014000.0 1159800.0 1000200.0 ;
      RECT  1149600.0 1014000.0 1159800.0 1027800.0 ;
      RECT  1149600.0 1041600.0 1159800.0 1027800.0 ;
      RECT  1149600.0 1041600.0 1159800.0 1055400.0 ;
      RECT  1149600.0 1069200.0 1159800.0 1055400.0 ;
      RECT  1149600.0 1069200.0 1159800.0 1083000.0 ;
      RECT  1149600.0 1096800.0 1159800.0 1083000.0 ;
      RECT  1149600.0 1096800.0 1159800.0 1110600.0 ;
      RECT  1149600.0 1124400.0 1159800.0 1110600.0 ;
      RECT  1149600.0 1124400.0 1159800.0 1138200.0 ;
      RECT  1149600.0 1152000.0 1159800.0 1138200.0 ;
      RECT  1149600.0 1152000.0 1159800.0 1165800.0 ;
      RECT  1149600.0 1179600.0 1159800.0 1165800.0 ;
      RECT  1149600.0 1179600.0 1159800.0 1193400.0 ;
      RECT  1149600.0 1207200.0 1159800.0 1193400.0 ;
      RECT  1149600.0 1207200.0 1159800.0 1221000.0 ;
      RECT  1149600.0 1234800.0 1159800.0 1221000.0 ;
      RECT  1149600.0 1234800.0 1159800.0 1248600.0 ;
      RECT  1149600.0 1262400.0 1159800.0 1248600.0 ;
      RECT  1149600.0 1262400.0 1159800.0 1276200.0 ;
      RECT  1149600.0 1290000.0 1159800.0 1276200.0 ;
      RECT  1149600.0 1290000.0 1159800.0 1303800.0 ;
      RECT  1149600.0 1317600.0 1159800.0 1303800.0 ;
      RECT  1149600.0 1317600.0 1159800.0 1331400.0 ;
      RECT  1149600.0 1345200.0 1159800.0 1331400.0 ;
      RECT  1149600.0 1345200.0 1159800.0 1359000.0 ;
      RECT  1149600.0 1372800.0 1159800.0 1359000.0 ;
      RECT  1149600.0 1372800.0 1159800.0 1386600.0 ;
      RECT  1149600.0 1400400.0 1159800.0 1386600.0 ;
      RECT  1149600.0 1400400.0 1159800.0 1414200.0 ;
      RECT  1149600.0 1428000.0 1159800.0 1414200.0 ;
      RECT  1149600.0 1428000.0 1159800.0 1441800.0 ;
      RECT  1149600.0 1455600.0 1159800.0 1441800.0 ;
      RECT  1149600.0 1455600.0 1159800.0 1469400.0 ;
      RECT  1149600.0 1483200.0 1159800.0 1469400.0 ;
      RECT  1149600.0 1483200.0 1159800.0 1497000.0 ;
      RECT  1149600.0 1510800.0 1159800.0 1497000.0 ;
      RECT  1149600.0 1510800.0 1159800.0 1524600.0 ;
      RECT  1149600.0 1538400.0 1159800.0 1524600.0 ;
      RECT  1149600.0 1538400.0 1159800.0 1552200.0 ;
      RECT  1149600.0 1566000.0 1159800.0 1552200.0 ;
      RECT  1149600.0 1566000.0 1159800.0 1579800.0 ;
      RECT  1149600.0 1593600.0 1159800.0 1579800.0 ;
      RECT  1149600.0 1593600.0 1159800.0 1607400.0 ;
      RECT  1149600.0 1621200.0 1159800.0 1607400.0 ;
      RECT  1149600.0 1621200.0 1159800.0 1635000.0 ;
      RECT  1149600.0 1648800.0 1159800.0 1635000.0 ;
      RECT  1149600.0 1648800.0 1159800.0 1662600.0 ;
      RECT  1149600.0 1676400.0 1159800.0 1662600.0 ;
      RECT  1149600.0 1676400.0 1159800.0 1690200.0 ;
      RECT  1149600.0 1704000.0 1159800.0 1690200.0 ;
      RECT  1149600.0 1704000.0 1159800.0 1717800.0 ;
      RECT  1149600.0 1731600.0 1159800.0 1717800.0 ;
      RECT  1149600.0 1731600.0 1159800.0 1745400.0 ;
      RECT  1149600.0 1759200.0 1159800.0 1745400.0 ;
      RECT  1149600.0 1759200.0 1159800.0 1773000.0 ;
      RECT  1149600.0 1786800.0 1159800.0 1773000.0 ;
      RECT  1149600.0 1786800.0 1159800.0 1800600.0 ;
      RECT  1149600.0 1814400.0 1159800.0 1800600.0 ;
      RECT  1149600.0 1814400.0 1159800.0 1828200.0 ;
      RECT  1149600.0 1842000.0 1159800.0 1828200.0 ;
      RECT  1149600.0 1842000.0 1159800.0 1855800.0 ;
      RECT  1149600.0 1869600.0 1159800.0 1855800.0 ;
      RECT  1149600.0 1869600.0 1159800.0 1883400.0 ;
      RECT  1149600.0 1897200.0 1159800.0 1883400.0 ;
      RECT  1149600.0 1897200.0 1159800.0 1911000.0 ;
      RECT  1149600.0 1924800.0 1159800.0 1911000.0 ;
      RECT  1149600.0 1924800.0 1159800.0 1938600.0 ;
      RECT  1149600.0 1952400.0 1159800.0 1938600.0 ;
      RECT  1149600.0 1952400.0 1159800.0 1966200.0 ;
      RECT  1149600.0 1980000.0 1159800.0 1966200.0 ;
      RECT  1149600.0 1980000.0 1159800.0 1993800.0 ;
      RECT  1149600.0 2007600.0 1159800.0 1993800.0 ;
      RECT  1149600.0 2007600.0 1159800.0 2021400.0 ;
      RECT  1149600.0 2035200.0 1159800.0 2021400.0 ;
      RECT  1149600.0 2035200.0 1159800.0 2049000.0 ;
      RECT  1149600.0 2062800.0 1159800.0 2049000.0 ;
      RECT  1149600.0 2062800.0 1159800.0 2076600.0 ;
      RECT  1149600.0 2090400.0 1159800.0 2076600.0 ;
      RECT  1149600.0 2090400.0 1159800.0 2104200.0 ;
      RECT  1149600.0 2118000.0 1159800.0 2104200.0 ;
      RECT  1149600.0 2118000.0 1159800.0 2131800.0 ;
      RECT  1149600.0 2145600.0 1159800.0 2131800.0 ;
      RECT  1159800.0 379200.0 1170000.0 393000.0 ;
      RECT  1159800.0 406800.0 1170000.0 393000.0 ;
      RECT  1159800.0 406800.0 1170000.0 420600.0 ;
      RECT  1159800.0 434400.0 1170000.0 420600.0 ;
      RECT  1159800.0 434400.0 1170000.0 448200.0 ;
      RECT  1159800.0 462000.0 1170000.0 448200.0 ;
      RECT  1159800.0 462000.0 1170000.0 475800.0 ;
      RECT  1159800.0 489600.0 1170000.0 475800.0 ;
      RECT  1159800.0 489600.0 1170000.0 503400.0 ;
      RECT  1159800.0 517200.0 1170000.0 503400.0 ;
      RECT  1159800.0 517200.0 1170000.0 531000.0 ;
      RECT  1159800.0 544800.0 1170000.0 531000.0 ;
      RECT  1159800.0 544800.0 1170000.0 558600.0 ;
      RECT  1159800.0 572400.0 1170000.0 558600.0 ;
      RECT  1159800.0 572400.0 1170000.0 586200.0 ;
      RECT  1159800.0 600000.0 1170000.0 586200.0 ;
      RECT  1159800.0 600000.0 1170000.0 613800.0 ;
      RECT  1159800.0 627600.0 1170000.0 613800.0 ;
      RECT  1159800.0 627600.0 1170000.0 641400.0 ;
      RECT  1159800.0 655200.0 1170000.0 641400.0 ;
      RECT  1159800.0 655200.0 1170000.0 669000.0 ;
      RECT  1159800.0 682800.0 1170000.0 669000.0 ;
      RECT  1159800.0 682800.0 1170000.0 696600.0 ;
      RECT  1159800.0 710400.0 1170000.0 696600.0 ;
      RECT  1159800.0 710400.0 1170000.0 724200.0 ;
      RECT  1159800.0 738000.0 1170000.0 724200.0 ;
      RECT  1159800.0 738000.0 1170000.0 751800.0 ;
      RECT  1159800.0 765600.0 1170000.0 751800.0 ;
      RECT  1159800.0 765600.0 1170000.0 779400.0 ;
      RECT  1159800.0 793200.0 1170000.0 779400.0 ;
      RECT  1159800.0 793200.0 1170000.0 807000.0 ;
      RECT  1159800.0 820800.0 1170000.0 807000.0 ;
      RECT  1159800.0 820800.0 1170000.0 834600.0 ;
      RECT  1159800.0 848400.0 1170000.0 834600.0 ;
      RECT  1159800.0 848400.0 1170000.0 862200.0 ;
      RECT  1159800.0 876000.0 1170000.0 862200.0 ;
      RECT  1159800.0 876000.0 1170000.0 889800.0 ;
      RECT  1159800.0 903600.0 1170000.0 889800.0 ;
      RECT  1159800.0 903600.0 1170000.0 917400.0 ;
      RECT  1159800.0 931200.0 1170000.0 917400.0 ;
      RECT  1159800.0 931200.0 1170000.0 945000.0 ;
      RECT  1159800.0 958800.0 1170000.0 945000.0 ;
      RECT  1159800.0 958800.0 1170000.0 972600.0 ;
      RECT  1159800.0 986400.0 1170000.0 972600.0 ;
      RECT  1159800.0 986400.0 1170000.0 1000200.0 ;
      RECT  1159800.0 1014000.0 1170000.0 1000200.0 ;
      RECT  1159800.0 1014000.0 1170000.0 1027800.0 ;
      RECT  1159800.0 1041600.0 1170000.0 1027800.0 ;
      RECT  1159800.0 1041600.0 1170000.0 1055400.0 ;
      RECT  1159800.0 1069200.0 1170000.0 1055400.0 ;
      RECT  1159800.0 1069200.0 1170000.0 1083000.0 ;
      RECT  1159800.0 1096800.0 1170000.0 1083000.0 ;
      RECT  1159800.0 1096800.0 1170000.0 1110600.0 ;
      RECT  1159800.0 1124400.0 1170000.0 1110600.0 ;
      RECT  1159800.0 1124400.0 1170000.0 1138200.0 ;
      RECT  1159800.0 1152000.0 1170000.0 1138200.0 ;
      RECT  1159800.0 1152000.0 1170000.0 1165800.0 ;
      RECT  1159800.0 1179600.0 1170000.0 1165800.0 ;
      RECT  1159800.0 1179600.0 1170000.0 1193400.0 ;
      RECT  1159800.0 1207200.0 1170000.0 1193400.0 ;
      RECT  1159800.0 1207200.0 1170000.0 1221000.0 ;
      RECT  1159800.0 1234800.0 1170000.0 1221000.0 ;
      RECT  1159800.0 1234800.0 1170000.0 1248600.0 ;
      RECT  1159800.0 1262400.0 1170000.0 1248600.0 ;
      RECT  1159800.0 1262400.0 1170000.0 1276200.0 ;
      RECT  1159800.0 1290000.0 1170000.0 1276200.0 ;
      RECT  1159800.0 1290000.0 1170000.0 1303800.0 ;
      RECT  1159800.0 1317600.0 1170000.0 1303800.0 ;
      RECT  1159800.0 1317600.0 1170000.0 1331400.0 ;
      RECT  1159800.0 1345200.0 1170000.0 1331400.0 ;
      RECT  1159800.0 1345200.0 1170000.0 1359000.0 ;
      RECT  1159800.0 1372800.0 1170000.0 1359000.0 ;
      RECT  1159800.0 1372800.0 1170000.0 1386600.0 ;
      RECT  1159800.0 1400400.0 1170000.0 1386600.0 ;
      RECT  1159800.0 1400400.0 1170000.0 1414200.0 ;
      RECT  1159800.0 1428000.0 1170000.0 1414200.0 ;
      RECT  1159800.0 1428000.0 1170000.0 1441800.0 ;
      RECT  1159800.0 1455600.0 1170000.0 1441800.0 ;
      RECT  1159800.0 1455600.0 1170000.0 1469400.0 ;
      RECT  1159800.0 1483200.0 1170000.0 1469400.0 ;
      RECT  1159800.0 1483200.0 1170000.0 1497000.0 ;
      RECT  1159800.0 1510800.0 1170000.0 1497000.0 ;
      RECT  1159800.0 1510800.0 1170000.0 1524600.0 ;
      RECT  1159800.0 1538400.0 1170000.0 1524600.0 ;
      RECT  1159800.0 1538400.0 1170000.0 1552200.0 ;
      RECT  1159800.0 1566000.0 1170000.0 1552200.0 ;
      RECT  1159800.0 1566000.0 1170000.0 1579800.0 ;
      RECT  1159800.0 1593600.0 1170000.0 1579800.0 ;
      RECT  1159800.0 1593600.0 1170000.0 1607400.0 ;
      RECT  1159800.0 1621200.0 1170000.0 1607400.0 ;
      RECT  1159800.0 1621200.0 1170000.0 1635000.0 ;
      RECT  1159800.0 1648800.0 1170000.0 1635000.0 ;
      RECT  1159800.0 1648800.0 1170000.0 1662600.0 ;
      RECT  1159800.0 1676400.0 1170000.0 1662600.0 ;
      RECT  1159800.0 1676400.0 1170000.0 1690200.0 ;
      RECT  1159800.0 1704000.0 1170000.0 1690200.0 ;
      RECT  1159800.0 1704000.0 1170000.0 1717800.0 ;
      RECT  1159800.0 1731600.0 1170000.0 1717800.0 ;
      RECT  1159800.0 1731600.0 1170000.0 1745400.0 ;
      RECT  1159800.0 1759200.0 1170000.0 1745400.0 ;
      RECT  1159800.0 1759200.0 1170000.0 1773000.0 ;
      RECT  1159800.0 1786800.0 1170000.0 1773000.0 ;
      RECT  1159800.0 1786800.0 1170000.0 1800600.0 ;
      RECT  1159800.0 1814400.0 1170000.0 1800600.0 ;
      RECT  1159800.0 1814400.0 1170000.0 1828200.0 ;
      RECT  1159800.0 1842000.0 1170000.0 1828200.0 ;
      RECT  1159800.0 1842000.0 1170000.0 1855800.0 ;
      RECT  1159800.0 1869600.0 1170000.0 1855800.0 ;
      RECT  1159800.0 1869600.0 1170000.0 1883400.0 ;
      RECT  1159800.0 1897200.0 1170000.0 1883400.0 ;
      RECT  1159800.0 1897200.0 1170000.0 1911000.0 ;
      RECT  1159800.0 1924800.0 1170000.0 1911000.0 ;
      RECT  1159800.0 1924800.0 1170000.0 1938600.0 ;
      RECT  1159800.0 1952400.0 1170000.0 1938600.0 ;
      RECT  1159800.0 1952400.0 1170000.0 1966200.0 ;
      RECT  1159800.0 1980000.0 1170000.0 1966200.0 ;
      RECT  1159800.0 1980000.0 1170000.0 1993800.0 ;
      RECT  1159800.0 2007600.0 1170000.0 1993800.0 ;
      RECT  1159800.0 2007600.0 1170000.0 2021400.0 ;
      RECT  1159800.0 2035200.0 1170000.0 2021400.0 ;
      RECT  1159800.0 2035200.0 1170000.0 2049000.0 ;
      RECT  1159800.0 2062800.0 1170000.0 2049000.0 ;
      RECT  1159800.0 2062800.0 1170000.0 2076600.0 ;
      RECT  1159800.0 2090400.0 1170000.0 2076600.0 ;
      RECT  1159800.0 2090400.0 1170000.0 2104200.0 ;
      RECT  1159800.0 2118000.0 1170000.0 2104200.0 ;
      RECT  1159800.0 2118000.0 1170000.0 2131800.0 ;
      RECT  1159800.0 2145600.0 1170000.0 2131800.0 ;
      RECT  1170000.0 379200.0 1180200.0 393000.0 ;
      RECT  1170000.0 406800.0 1180200.0 393000.0 ;
      RECT  1170000.0 406800.0 1180200.0 420600.0 ;
      RECT  1170000.0 434400.0 1180200.0 420600.0 ;
      RECT  1170000.0 434400.0 1180200.0 448200.0 ;
      RECT  1170000.0 462000.0 1180200.0 448200.0 ;
      RECT  1170000.0 462000.0 1180200.0 475800.0 ;
      RECT  1170000.0 489600.0 1180200.0 475800.0 ;
      RECT  1170000.0 489600.0 1180200.0 503400.0 ;
      RECT  1170000.0 517200.0 1180200.0 503400.0 ;
      RECT  1170000.0 517200.0 1180200.0 531000.0 ;
      RECT  1170000.0 544800.0 1180200.0 531000.0 ;
      RECT  1170000.0 544800.0 1180200.0 558600.0 ;
      RECT  1170000.0 572400.0 1180200.0 558600.0 ;
      RECT  1170000.0 572400.0 1180200.0 586200.0 ;
      RECT  1170000.0 600000.0 1180200.0 586200.0 ;
      RECT  1170000.0 600000.0 1180200.0 613800.0 ;
      RECT  1170000.0 627600.0 1180200.0 613800.0 ;
      RECT  1170000.0 627600.0 1180200.0 641400.0 ;
      RECT  1170000.0 655200.0 1180200.0 641400.0 ;
      RECT  1170000.0 655200.0 1180200.0 669000.0 ;
      RECT  1170000.0 682800.0 1180200.0 669000.0 ;
      RECT  1170000.0 682800.0 1180200.0 696600.0 ;
      RECT  1170000.0 710400.0 1180200.0 696600.0 ;
      RECT  1170000.0 710400.0 1180200.0 724200.0 ;
      RECT  1170000.0 738000.0 1180200.0 724200.0 ;
      RECT  1170000.0 738000.0 1180200.0 751800.0 ;
      RECT  1170000.0 765600.0 1180200.0 751800.0 ;
      RECT  1170000.0 765600.0 1180200.0 779400.0 ;
      RECT  1170000.0 793200.0 1180200.0 779400.0 ;
      RECT  1170000.0 793200.0 1180200.0 807000.0 ;
      RECT  1170000.0 820800.0 1180200.0 807000.0 ;
      RECT  1170000.0 820800.0 1180200.0 834600.0 ;
      RECT  1170000.0 848400.0 1180200.0 834600.0 ;
      RECT  1170000.0 848400.0 1180200.0 862200.0 ;
      RECT  1170000.0 876000.0 1180200.0 862200.0 ;
      RECT  1170000.0 876000.0 1180200.0 889800.0 ;
      RECT  1170000.0 903600.0 1180200.0 889800.0 ;
      RECT  1170000.0 903600.0 1180200.0 917400.0 ;
      RECT  1170000.0 931200.0 1180200.0 917400.0 ;
      RECT  1170000.0 931200.0 1180200.0 945000.0 ;
      RECT  1170000.0 958800.0 1180200.0 945000.0 ;
      RECT  1170000.0 958800.0 1180200.0 972600.0 ;
      RECT  1170000.0 986400.0 1180200.0 972600.0 ;
      RECT  1170000.0 986400.0 1180200.0 1000200.0 ;
      RECT  1170000.0 1014000.0 1180200.0 1000200.0 ;
      RECT  1170000.0 1014000.0 1180200.0 1027800.0 ;
      RECT  1170000.0 1041600.0 1180200.0 1027800.0 ;
      RECT  1170000.0 1041600.0 1180200.0 1055400.0 ;
      RECT  1170000.0 1069200.0 1180200.0 1055400.0 ;
      RECT  1170000.0 1069200.0 1180200.0 1083000.0 ;
      RECT  1170000.0 1096800.0 1180200.0 1083000.0 ;
      RECT  1170000.0 1096800.0 1180200.0 1110600.0 ;
      RECT  1170000.0 1124400.0 1180200.0 1110600.0 ;
      RECT  1170000.0 1124400.0 1180200.0 1138200.0 ;
      RECT  1170000.0 1152000.0 1180200.0 1138200.0 ;
      RECT  1170000.0 1152000.0 1180200.0 1165800.0 ;
      RECT  1170000.0 1179600.0 1180200.0 1165800.0 ;
      RECT  1170000.0 1179600.0 1180200.0 1193400.0 ;
      RECT  1170000.0 1207200.0 1180200.0 1193400.0 ;
      RECT  1170000.0 1207200.0 1180200.0 1221000.0 ;
      RECT  1170000.0 1234800.0 1180200.0 1221000.0 ;
      RECT  1170000.0 1234800.0 1180200.0 1248600.0 ;
      RECT  1170000.0 1262400.0 1180200.0 1248600.0 ;
      RECT  1170000.0 1262400.0 1180200.0 1276200.0 ;
      RECT  1170000.0 1290000.0 1180200.0 1276200.0 ;
      RECT  1170000.0 1290000.0 1180200.0 1303800.0 ;
      RECT  1170000.0 1317600.0 1180200.0 1303800.0 ;
      RECT  1170000.0 1317600.0 1180200.0 1331400.0 ;
      RECT  1170000.0 1345200.0 1180200.0 1331400.0 ;
      RECT  1170000.0 1345200.0 1180200.0 1359000.0 ;
      RECT  1170000.0 1372800.0 1180200.0 1359000.0 ;
      RECT  1170000.0 1372800.0 1180200.0 1386600.0 ;
      RECT  1170000.0 1400400.0 1180200.0 1386600.0 ;
      RECT  1170000.0 1400400.0 1180200.0 1414200.0 ;
      RECT  1170000.0 1428000.0 1180200.0 1414200.0 ;
      RECT  1170000.0 1428000.0 1180200.0 1441800.0 ;
      RECT  1170000.0 1455600.0 1180200.0 1441800.0 ;
      RECT  1170000.0 1455600.0 1180200.0 1469400.0 ;
      RECT  1170000.0 1483200.0 1180200.0 1469400.0 ;
      RECT  1170000.0 1483200.0 1180200.0 1497000.0 ;
      RECT  1170000.0 1510800.0 1180200.0 1497000.0 ;
      RECT  1170000.0 1510800.0 1180200.0 1524600.0 ;
      RECT  1170000.0 1538400.0 1180200.0 1524600.0 ;
      RECT  1170000.0 1538400.0 1180200.0 1552200.0 ;
      RECT  1170000.0 1566000.0 1180200.0 1552200.0 ;
      RECT  1170000.0 1566000.0 1180200.0 1579800.0 ;
      RECT  1170000.0 1593600.0 1180200.0 1579800.0 ;
      RECT  1170000.0 1593600.0 1180200.0 1607400.0 ;
      RECT  1170000.0 1621200.0 1180200.0 1607400.0 ;
      RECT  1170000.0 1621200.0 1180200.0 1635000.0 ;
      RECT  1170000.0 1648800.0 1180200.0 1635000.0 ;
      RECT  1170000.0 1648800.0 1180200.0 1662600.0 ;
      RECT  1170000.0 1676400.0 1180200.0 1662600.0 ;
      RECT  1170000.0 1676400.0 1180200.0 1690200.0 ;
      RECT  1170000.0 1704000.0 1180200.0 1690200.0 ;
      RECT  1170000.0 1704000.0 1180200.0 1717800.0 ;
      RECT  1170000.0 1731600.0 1180200.0 1717800.0 ;
      RECT  1170000.0 1731600.0 1180200.0 1745400.0 ;
      RECT  1170000.0 1759200.0 1180200.0 1745400.0 ;
      RECT  1170000.0 1759200.0 1180200.0 1773000.0 ;
      RECT  1170000.0 1786800.0 1180200.0 1773000.0 ;
      RECT  1170000.0 1786800.0 1180200.0 1800600.0 ;
      RECT  1170000.0 1814400.0 1180200.0 1800600.0 ;
      RECT  1170000.0 1814400.0 1180200.0 1828200.0 ;
      RECT  1170000.0 1842000.0 1180200.0 1828200.0 ;
      RECT  1170000.0 1842000.0 1180200.0 1855800.0 ;
      RECT  1170000.0 1869600.0 1180200.0 1855800.0 ;
      RECT  1170000.0 1869600.0 1180200.0 1883400.0 ;
      RECT  1170000.0 1897200.0 1180200.0 1883400.0 ;
      RECT  1170000.0 1897200.0 1180200.0 1911000.0 ;
      RECT  1170000.0 1924800.0 1180200.0 1911000.0 ;
      RECT  1170000.0 1924800.0 1180200.0 1938600.0 ;
      RECT  1170000.0 1952400.0 1180200.0 1938600.0 ;
      RECT  1170000.0 1952400.0 1180200.0 1966200.0 ;
      RECT  1170000.0 1980000.0 1180200.0 1966200.0 ;
      RECT  1170000.0 1980000.0 1180200.0 1993800.0 ;
      RECT  1170000.0 2007600.0 1180200.0 1993800.0 ;
      RECT  1170000.0 2007600.0 1180200.0 2021400.0 ;
      RECT  1170000.0 2035200.0 1180200.0 2021400.0 ;
      RECT  1170000.0 2035200.0 1180200.0 2049000.0 ;
      RECT  1170000.0 2062800.0 1180200.0 2049000.0 ;
      RECT  1170000.0 2062800.0 1180200.0 2076600.0 ;
      RECT  1170000.0 2090400.0 1180200.0 2076600.0 ;
      RECT  1170000.0 2090400.0 1180200.0 2104200.0 ;
      RECT  1170000.0 2118000.0 1180200.0 2104200.0 ;
      RECT  1170000.0 2118000.0 1180200.0 2131800.0 ;
      RECT  1170000.0 2145600.0 1180200.0 2131800.0 ;
      RECT  1180200.0 379200.0 1190400.0 393000.0 ;
      RECT  1180200.0 406800.0 1190400.0 393000.0 ;
      RECT  1180200.0 406800.0 1190400.0 420600.0 ;
      RECT  1180200.0 434400.0 1190400.0 420600.0 ;
      RECT  1180200.0 434400.0 1190400.0 448200.0 ;
      RECT  1180200.0 462000.0 1190400.0 448200.0 ;
      RECT  1180200.0 462000.0 1190400.0 475800.0 ;
      RECT  1180200.0 489600.0 1190400.0 475800.0 ;
      RECT  1180200.0 489600.0 1190400.0 503400.0 ;
      RECT  1180200.0 517200.0 1190400.0 503400.0 ;
      RECT  1180200.0 517200.0 1190400.0 531000.0 ;
      RECT  1180200.0 544800.0 1190400.0 531000.0 ;
      RECT  1180200.0 544800.0 1190400.0 558600.0 ;
      RECT  1180200.0 572400.0 1190400.0 558600.0 ;
      RECT  1180200.0 572400.0 1190400.0 586200.0 ;
      RECT  1180200.0 600000.0 1190400.0 586200.0 ;
      RECT  1180200.0 600000.0 1190400.0 613800.0 ;
      RECT  1180200.0 627600.0 1190400.0 613800.0 ;
      RECT  1180200.0 627600.0 1190400.0 641400.0 ;
      RECT  1180200.0 655200.0 1190400.0 641400.0 ;
      RECT  1180200.0 655200.0 1190400.0 669000.0 ;
      RECT  1180200.0 682800.0 1190400.0 669000.0 ;
      RECT  1180200.0 682800.0 1190400.0 696600.0 ;
      RECT  1180200.0 710400.0 1190400.0 696600.0 ;
      RECT  1180200.0 710400.0 1190400.0 724200.0 ;
      RECT  1180200.0 738000.0 1190400.0 724200.0 ;
      RECT  1180200.0 738000.0 1190400.0 751800.0 ;
      RECT  1180200.0 765600.0 1190400.0 751800.0 ;
      RECT  1180200.0 765600.0 1190400.0 779400.0 ;
      RECT  1180200.0 793200.0 1190400.0 779400.0 ;
      RECT  1180200.0 793200.0 1190400.0 807000.0 ;
      RECT  1180200.0 820800.0 1190400.0 807000.0 ;
      RECT  1180200.0 820800.0 1190400.0 834600.0 ;
      RECT  1180200.0 848400.0 1190400.0 834600.0 ;
      RECT  1180200.0 848400.0 1190400.0 862200.0 ;
      RECT  1180200.0 876000.0 1190400.0 862200.0 ;
      RECT  1180200.0 876000.0 1190400.0 889800.0 ;
      RECT  1180200.0 903600.0 1190400.0 889800.0 ;
      RECT  1180200.0 903600.0 1190400.0 917400.0 ;
      RECT  1180200.0 931200.0 1190400.0 917400.0 ;
      RECT  1180200.0 931200.0 1190400.0 945000.0 ;
      RECT  1180200.0 958800.0 1190400.0 945000.0 ;
      RECT  1180200.0 958800.0 1190400.0 972600.0 ;
      RECT  1180200.0 986400.0 1190400.0 972600.0 ;
      RECT  1180200.0 986400.0 1190400.0 1000200.0 ;
      RECT  1180200.0 1014000.0 1190400.0 1000200.0 ;
      RECT  1180200.0 1014000.0 1190400.0 1027800.0 ;
      RECT  1180200.0 1041600.0 1190400.0 1027800.0 ;
      RECT  1180200.0 1041600.0 1190400.0 1055400.0 ;
      RECT  1180200.0 1069200.0 1190400.0 1055400.0 ;
      RECT  1180200.0 1069200.0 1190400.0 1083000.0 ;
      RECT  1180200.0 1096800.0 1190400.0 1083000.0 ;
      RECT  1180200.0 1096800.0 1190400.0 1110600.0 ;
      RECT  1180200.0 1124400.0 1190400.0 1110600.0 ;
      RECT  1180200.0 1124400.0 1190400.0 1138200.0 ;
      RECT  1180200.0 1152000.0 1190400.0 1138200.0 ;
      RECT  1180200.0 1152000.0 1190400.0 1165800.0 ;
      RECT  1180200.0 1179600.0 1190400.0 1165800.0 ;
      RECT  1180200.0 1179600.0 1190400.0 1193400.0 ;
      RECT  1180200.0 1207200.0 1190400.0 1193400.0 ;
      RECT  1180200.0 1207200.0 1190400.0 1221000.0 ;
      RECT  1180200.0 1234800.0 1190400.0 1221000.0 ;
      RECT  1180200.0 1234800.0 1190400.0 1248600.0 ;
      RECT  1180200.0 1262400.0 1190400.0 1248600.0 ;
      RECT  1180200.0 1262400.0 1190400.0 1276200.0 ;
      RECT  1180200.0 1290000.0 1190400.0 1276200.0 ;
      RECT  1180200.0 1290000.0 1190400.0 1303800.0 ;
      RECT  1180200.0 1317600.0 1190400.0 1303800.0 ;
      RECT  1180200.0 1317600.0 1190400.0 1331400.0 ;
      RECT  1180200.0 1345200.0 1190400.0 1331400.0 ;
      RECT  1180200.0 1345200.0 1190400.0 1359000.0 ;
      RECT  1180200.0 1372800.0 1190400.0 1359000.0 ;
      RECT  1180200.0 1372800.0 1190400.0 1386600.0 ;
      RECT  1180200.0 1400400.0 1190400.0 1386600.0 ;
      RECT  1180200.0 1400400.0 1190400.0 1414200.0 ;
      RECT  1180200.0 1428000.0 1190400.0 1414200.0 ;
      RECT  1180200.0 1428000.0 1190400.0 1441800.0 ;
      RECT  1180200.0 1455600.0 1190400.0 1441800.0 ;
      RECT  1180200.0 1455600.0 1190400.0 1469400.0 ;
      RECT  1180200.0 1483200.0 1190400.0 1469400.0 ;
      RECT  1180200.0 1483200.0 1190400.0 1497000.0 ;
      RECT  1180200.0 1510800.0 1190400.0 1497000.0 ;
      RECT  1180200.0 1510800.0 1190400.0 1524600.0 ;
      RECT  1180200.0 1538400.0 1190400.0 1524600.0 ;
      RECT  1180200.0 1538400.0 1190400.0 1552200.0 ;
      RECT  1180200.0 1566000.0 1190400.0 1552200.0 ;
      RECT  1180200.0 1566000.0 1190400.0 1579800.0 ;
      RECT  1180200.0 1593600.0 1190400.0 1579800.0 ;
      RECT  1180200.0 1593600.0 1190400.0 1607400.0 ;
      RECT  1180200.0 1621200.0 1190400.0 1607400.0 ;
      RECT  1180200.0 1621200.0 1190400.0 1635000.0 ;
      RECT  1180200.0 1648800.0 1190400.0 1635000.0 ;
      RECT  1180200.0 1648800.0 1190400.0 1662600.0 ;
      RECT  1180200.0 1676400.0 1190400.0 1662600.0 ;
      RECT  1180200.0 1676400.0 1190400.0 1690200.0 ;
      RECT  1180200.0 1704000.0 1190400.0 1690200.0 ;
      RECT  1180200.0 1704000.0 1190400.0 1717800.0 ;
      RECT  1180200.0 1731600.0 1190400.0 1717800.0 ;
      RECT  1180200.0 1731600.0 1190400.0 1745400.0 ;
      RECT  1180200.0 1759200.0 1190400.0 1745400.0 ;
      RECT  1180200.0 1759200.0 1190400.0 1773000.0 ;
      RECT  1180200.0 1786800.0 1190400.0 1773000.0 ;
      RECT  1180200.0 1786800.0 1190400.0 1800600.0 ;
      RECT  1180200.0 1814400.0 1190400.0 1800600.0 ;
      RECT  1180200.0 1814400.0 1190400.0 1828200.0 ;
      RECT  1180200.0 1842000.0 1190400.0 1828200.0 ;
      RECT  1180200.0 1842000.0 1190400.0 1855800.0 ;
      RECT  1180200.0 1869600.0 1190400.0 1855800.0 ;
      RECT  1180200.0 1869600.0 1190400.0 1883400.0 ;
      RECT  1180200.0 1897200.0 1190400.0 1883400.0 ;
      RECT  1180200.0 1897200.0 1190400.0 1911000.0 ;
      RECT  1180200.0 1924800.0 1190400.0 1911000.0 ;
      RECT  1180200.0 1924800.0 1190400.0 1938600.0 ;
      RECT  1180200.0 1952400.0 1190400.0 1938600.0 ;
      RECT  1180200.0 1952400.0 1190400.0 1966200.0 ;
      RECT  1180200.0 1980000.0 1190400.0 1966200.0 ;
      RECT  1180200.0 1980000.0 1190400.0 1993800.0 ;
      RECT  1180200.0 2007600.0 1190400.0 1993800.0 ;
      RECT  1180200.0 2007600.0 1190400.0 2021400.0 ;
      RECT  1180200.0 2035200.0 1190400.0 2021400.0 ;
      RECT  1180200.0 2035200.0 1190400.0 2049000.0 ;
      RECT  1180200.0 2062800.0 1190400.0 2049000.0 ;
      RECT  1180200.0 2062800.0 1190400.0 2076600.0 ;
      RECT  1180200.0 2090400.0 1190400.0 2076600.0 ;
      RECT  1180200.0 2090400.0 1190400.0 2104200.0 ;
      RECT  1180200.0 2118000.0 1190400.0 2104200.0 ;
      RECT  1180200.0 2118000.0 1190400.0 2131800.0 ;
      RECT  1180200.0 2145600.0 1190400.0 2131800.0 ;
      RECT  1190400.0 379200.0 1200600.0 393000.0 ;
      RECT  1190400.0 406800.0 1200600.0 393000.0 ;
      RECT  1190400.0 406800.0 1200600.0 420600.0 ;
      RECT  1190400.0 434400.0 1200600.0 420600.0 ;
      RECT  1190400.0 434400.0 1200600.0 448200.0 ;
      RECT  1190400.0 462000.0 1200600.0 448200.0 ;
      RECT  1190400.0 462000.0 1200600.0 475800.0 ;
      RECT  1190400.0 489600.0 1200600.0 475800.0 ;
      RECT  1190400.0 489600.0 1200600.0 503400.0 ;
      RECT  1190400.0 517200.0 1200600.0 503400.0 ;
      RECT  1190400.0 517200.0 1200600.0 531000.0 ;
      RECT  1190400.0 544800.0 1200600.0 531000.0 ;
      RECT  1190400.0 544800.0 1200600.0 558600.0 ;
      RECT  1190400.0 572400.0 1200600.0 558600.0 ;
      RECT  1190400.0 572400.0 1200600.0 586200.0 ;
      RECT  1190400.0 600000.0 1200600.0 586200.0 ;
      RECT  1190400.0 600000.0 1200600.0 613800.0 ;
      RECT  1190400.0 627600.0 1200600.0 613800.0 ;
      RECT  1190400.0 627600.0 1200600.0 641400.0 ;
      RECT  1190400.0 655200.0 1200600.0 641400.0 ;
      RECT  1190400.0 655200.0 1200600.0 669000.0 ;
      RECT  1190400.0 682800.0 1200600.0 669000.0 ;
      RECT  1190400.0 682800.0 1200600.0 696600.0 ;
      RECT  1190400.0 710400.0 1200600.0 696600.0 ;
      RECT  1190400.0 710400.0 1200600.0 724200.0 ;
      RECT  1190400.0 738000.0 1200600.0 724200.0 ;
      RECT  1190400.0 738000.0 1200600.0 751800.0 ;
      RECT  1190400.0 765600.0 1200600.0 751800.0 ;
      RECT  1190400.0 765600.0 1200600.0 779400.0 ;
      RECT  1190400.0 793200.0 1200600.0 779400.0 ;
      RECT  1190400.0 793200.0 1200600.0 807000.0 ;
      RECT  1190400.0 820800.0 1200600.0 807000.0 ;
      RECT  1190400.0 820800.0 1200600.0 834600.0 ;
      RECT  1190400.0 848400.0 1200600.0 834600.0 ;
      RECT  1190400.0 848400.0 1200600.0 862200.0 ;
      RECT  1190400.0 876000.0 1200600.0 862200.0 ;
      RECT  1190400.0 876000.0 1200600.0 889800.0 ;
      RECT  1190400.0 903600.0 1200600.0 889800.0 ;
      RECT  1190400.0 903600.0 1200600.0 917400.0 ;
      RECT  1190400.0 931200.0 1200600.0 917400.0 ;
      RECT  1190400.0 931200.0 1200600.0 945000.0 ;
      RECT  1190400.0 958800.0 1200600.0 945000.0 ;
      RECT  1190400.0 958800.0 1200600.0 972600.0 ;
      RECT  1190400.0 986400.0 1200600.0 972600.0 ;
      RECT  1190400.0 986400.0 1200600.0 1000200.0 ;
      RECT  1190400.0 1014000.0 1200600.0 1000200.0 ;
      RECT  1190400.0 1014000.0 1200600.0 1027800.0 ;
      RECT  1190400.0 1041600.0 1200600.0 1027800.0 ;
      RECT  1190400.0 1041600.0 1200600.0 1055400.0 ;
      RECT  1190400.0 1069200.0 1200600.0 1055400.0 ;
      RECT  1190400.0 1069200.0 1200600.0 1083000.0 ;
      RECT  1190400.0 1096800.0 1200600.0 1083000.0 ;
      RECT  1190400.0 1096800.0 1200600.0 1110600.0 ;
      RECT  1190400.0 1124400.0 1200600.0 1110600.0 ;
      RECT  1190400.0 1124400.0 1200600.0 1138200.0 ;
      RECT  1190400.0 1152000.0 1200600.0 1138200.0 ;
      RECT  1190400.0 1152000.0 1200600.0 1165800.0 ;
      RECT  1190400.0 1179600.0 1200600.0 1165800.0 ;
      RECT  1190400.0 1179600.0 1200600.0 1193400.0 ;
      RECT  1190400.0 1207200.0 1200600.0 1193400.0 ;
      RECT  1190400.0 1207200.0 1200600.0 1221000.0 ;
      RECT  1190400.0 1234800.0 1200600.0 1221000.0 ;
      RECT  1190400.0 1234800.0 1200600.0 1248600.0 ;
      RECT  1190400.0 1262400.0 1200600.0 1248600.0 ;
      RECT  1190400.0 1262400.0 1200600.0 1276200.0 ;
      RECT  1190400.0 1290000.0 1200600.0 1276200.0 ;
      RECT  1190400.0 1290000.0 1200600.0 1303800.0 ;
      RECT  1190400.0 1317600.0 1200600.0 1303800.0 ;
      RECT  1190400.0 1317600.0 1200600.0 1331400.0 ;
      RECT  1190400.0 1345200.0 1200600.0 1331400.0 ;
      RECT  1190400.0 1345200.0 1200600.0 1359000.0 ;
      RECT  1190400.0 1372800.0 1200600.0 1359000.0 ;
      RECT  1190400.0 1372800.0 1200600.0 1386600.0 ;
      RECT  1190400.0 1400400.0 1200600.0 1386600.0 ;
      RECT  1190400.0 1400400.0 1200600.0 1414200.0 ;
      RECT  1190400.0 1428000.0 1200600.0 1414200.0 ;
      RECT  1190400.0 1428000.0 1200600.0 1441800.0 ;
      RECT  1190400.0 1455600.0 1200600.0 1441800.0 ;
      RECT  1190400.0 1455600.0 1200600.0 1469400.0 ;
      RECT  1190400.0 1483200.0 1200600.0 1469400.0 ;
      RECT  1190400.0 1483200.0 1200600.0 1497000.0 ;
      RECT  1190400.0 1510800.0 1200600.0 1497000.0 ;
      RECT  1190400.0 1510800.0 1200600.0 1524600.0 ;
      RECT  1190400.0 1538400.0 1200600.0 1524600.0 ;
      RECT  1190400.0 1538400.0 1200600.0 1552200.0 ;
      RECT  1190400.0 1566000.0 1200600.0 1552200.0 ;
      RECT  1190400.0 1566000.0 1200600.0 1579800.0 ;
      RECT  1190400.0 1593600.0 1200600.0 1579800.0 ;
      RECT  1190400.0 1593600.0 1200600.0 1607400.0 ;
      RECT  1190400.0 1621200.0 1200600.0 1607400.0 ;
      RECT  1190400.0 1621200.0 1200600.0 1635000.0 ;
      RECT  1190400.0 1648800.0 1200600.0 1635000.0 ;
      RECT  1190400.0 1648800.0 1200600.0 1662600.0 ;
      RECT  1190400.0 1676400.0 1200600.0 1662600.0 ;
      RECT  1190400.0 1676400.0 1200600.0 1690200.0 ;
      RECT  1190400.0 1704000.0 1200600.0 1690200.0 ;
      RECT  1190400.0 1704000.0 1200600.0 1717800.0 ;
      RECT  1190400.0 1731600.0 1200600.0 1717800.0 ;
      RECT  1190400.0 1731600.0 1200600.0 1745400.0 ;
      RECT  1190400.0 1759200.0 1200600.0 1745400.0 ;
      RECT  1190400.0 1759200.0 1200600.0 1773000.0 ;
      RECT  1190400.0 1786800.0 1200600.0 1773000.0 ;
      RECT  1190400.0 1786800.0 1200600.0 1800600.0 ;
      RECT  1190400.0 1814400.0 1200600.0 1800600.0 ;
      RECT  1190400.0 1814400.0 1200600.0 1828200.0 ;
      RECT  1190400.0 1842000.0 1200600.0 1828200.0 ;
      RECT  1190400.0 1842000.0 1200600.0 1855800.0 ;
      RECT  1190400.0 1869600.0 1200600.0 1855800.0 ;
      RECT  1190400.0 1869600.0 1200600.0 1883400.0 ;
      RECT  1190400.0 1897200.0 1200600.0 1883400.0 ;
      RECT  1190400.0 1897200.0 1200600.0 1911000.0 ;
      RECT  1190400.0 1924800.0 1200600.0 1911000.0 ;
      RECT  1190400.0 1924800.0 1200600.0 1938600.0 ;
      RECT  1190400.0 1952400.0 1200600.0 1938600.0 ;
      RECT  1190400.0 1952400.0 1200600.0 1966200.0 ;
      RECT  1190400.0 1980000.0 1200600.0 1966200.0 ;
      RECT  1190400.0 1980000.0 1200600.0 1993800.0 ;
      RECT  1190400.0 2007600.0 1200600.0 1993800.0 ;
      RECT  1190400.0 2007600.0 1200600.0 2021400.0 ;
      RECT  1190400.0 2035200.0 1200600.0 2021400.0 ;
      RECT  1190400.0 2035200.0 1200600.0 2049000.0 ;
      RECT  1190400.0 2062800.0 1200600.0 2049000.0 ;
      RECT  1190400.0 2062800.0 1200600.0 2076600.0 ;
      RECT  1190400.0 2090400.0 1200600.0 2076600.0 ;
      RECT  1190400.0 2090400.0 1200600.0 2104200.0 ;
      RECT  1190400.0 2118000.0 1200600.0 2104200.0 ;
      RECT  1190400.0 2118000.0 1200600.0 2131800.0 ;
      RECT  1190400.0 2145600.0 1200600.0 2131800.0 ;
      RECT  1200600.0 379200.0 1210800.0 393000.0 ;
      RECT  1200600.0 406800.0 1210800.0 393000.0 ;
      RECT  1200600.0 406800.0 1210800.0 420600.0 ;
      RECT  1200600.0 434400.0 1210800.0 420600.0 ;
      RECT  1200600.0 434400.0 1210800.0 448200.0 ;
      RECT  1200600.0 462000.0 1210800.0 448200.0 ;
      RECT  1200600.0 462000.0 1210800.0 475800.0 ;
      RECT  1200600.0 489600.0 1210800.0 475800.0 ;
      RECT  1200600.0 489600.0 1210800.0 503400.0 ;
      RECT  1200600.0 517200.0 1210800.0 503400.0 ;
      RECT  1200600.0 517200.0 1210800.0 531000.0 ;
      RECT  1200600.0 544800.0 1210800.0 531000.0 ;
      RECT  1200600.0 544800.0 1210800.0 558600.0 ;
      RECT  1200600.0 572400.0 1210800.0 558600.0 ;
      RECT  1200600.0 572400.0 1210800.0 586200.0 ;
      RECT  1200600.0 600000.0 1210800.0 586200.0 ;
      RECT  1200600.0 600000.0 1210800.0 613800.0 ;
      RECT  1200600.0 627600.0 1210800.0 613800.0 ;
      RECT  1200600.0 627600.0 1210800.0 641400.0 ;
      RECT  1200600.0 655200.0 1210800.0 641400.0 ;
      RECT  1200600.0 655200.0 1210800.0 669000.0 ;
      RECT  1200600.0 682800.0 1210800.0 669000.0 ;
      RECT  1200600.0 682800.0 1210800.0 696600.0 ;
      RECT  1200600.0 710400.0 1210800.0 696600.0 ;
      RECT  1200600.0 710400.0 1210800.0 724200.0 ;
      RECT  1200600.0 738000.0 1210800.0 724200.0 ;
      RECT  1200600.0 738000.0 1210800.0 751800.0 ;
      RECT  1200600.0 765600.0 1210800.0 751800.0 ;
      RECT  1200600.0 765600.0 1210800.0 779400.0 ;
      RECT  1200600.0 793200.0 1210800.0 779400.0 ;
      RECT  1200600.0 793200.0 1210800.0 807000.0 ;
      RECT  1200600.0 820800.0 1210800.0 807000.0 ;
      RECT  1200600.0 820800.0 1210800.0 834600.0 ;
      RECT  1200600.0 848400.0 1210800.0 834600.0 ;
      RECT  1200600.0 848400.0 1210800.0 862200.0 ;
      RECT  1200600.0 876000.0 1210800.0 862200.0 ;
      RECT  1200600.0 876000.0 1210800.0 889800.0 ;
      RECT  1200600.0 903600.0 1210800.0 889800.0 ;
      RECT  1200600.0 903600.0 1210800.0 917400.0 ;
      RECT  1200600.0 931200.0 1210800.0 917400.0 ;
      RECT  1200600.0 931200.0 1210800.0 945000.0 ;
      RECT  1200600.0 958800.0 1210800.0 945000.0 ;
      RECT  1200600.0 958800.0 1210800.0 972600.0 ;
      RECT  1200600.0 986400.0 1210800.0 972600.0 ;
      RECT  1200600.0 986400.0 1210800.0 1000200.0 ;
      RECT  1200600.0 1014000.0 1210800.0 1000200.0 ;
      RECT  1200600.0 1014000.0 1210800.0 1027800.0 ;
      RECT  1200600.0 1041600.0 1210800.0 1027800.0 ;
      RECT  1200600.0 1041600.0 1210800.0 1055400.0 ;
      RECT  1200600.0 1069200.0 1210800.0 1055400.0 ;
      RECT  1200600.0 1069200.0 1210800.0 1083000.0 ;
      RECT  1200600.0 1096800.0 1210800.0 1083000.0 ;
      RECT  1200600.0 1096800.0 1210800.0 1110600.0 ;
      RECT  1200600.0 1124400.0 1210800.0 1110600.0 ;
      RECT  1200600.0 1124400.0 1210800.0 1138200.0 ;
      RECT  1200600.0 1152000.0 1210800.0 1138200.0 ;
      RECT  1200600.0 1152000.0 1210800.0 1165800.0 ;
      RECT  1200600.0 1179600.0 1210800.0 1165800.0 ;
      RECT  1200600.0 1179600.0 1210800.0 1193400.0 ;
      RECT  1200600.0 1207200.0 1210800.0 1193400.0 ;
      RECT  1200600.0 1207200.0 1210800.0 1221000.0 ;
      RECT  1200600.0 1234800.0 1210800.0 1221000.0 ;
      RECT  1200600.0 1234800.0 1210800.0 1248600.0 ;
      RECT  1200600.0 1262400.0 1210800.0 1248600.0 ;
      RECT  1200600.0 1262400.0 1210800.0 1276200.0 ;
      RECT  1200600.0 1290000.0 1210800.0 1276200.0 ;
      RECT  1200600.0 1290000.0 1210800.0 1303800.0 ;
      RECT  1200600.0 1317600.0 1210800.0 1303800.0 ;
      RECT  1200600.0 1317600.0 1210800.0 1331400.0 ;
      RECT  1200600.0 1345200.0 1210800.0 1331400.0 ;
      RECT  1200600.0 1345200.0 1210800.0 1359000.0 ;
      RECT  1200600.0 1372800.0 1210800.0 1359000.0 ;
      RECT  1200600.0 1372800.0 1210800.0 1386600.0 ;
      RECT  1200600.0 1400400.0 1210800.0 1386600.0 ;
      RECT  1200600.0 1400400.0 1210800.0 1414200.0 ;
      RECT  1200600.0 1428000.0 1210800.0 1414200.0 ;
      RECT  1200600.0 1428000.0 1210800.0 1441800.0 ;
      RECT  1200600.0 1455600.0 1210800.0 1441800.0 ;
      RECT  1200600.0 1455600.0 1210800.0 1469400.0 ;
      RECT  1200600.0 1483200.0 1210800.0 1469400.0 ;
      RECT  1200600.0 1483200.0 1210800.0 1497000.0 ;
      RECT  1200600.0 1510800.0 1210800.0 1497000.0 ;
      RECT  1200600.0 1510800.0 1210800.0 1524600.0 ;
      RECT  1200600.0 1538400.0 1210800.0 1524600.0 ;
      RECT  1200600.0 1538400.0 1210800.0 1552200.0 ;
      RECT  1200600.0 1566000.0 1210800.0 1552200.0 ;
      RECT  1200600.0 1566000.0 1210800.0 1579800.0 ;
      RECT  1200600.0 1593600.0 1210800.0 1579800.0 ;
      RECT  1200600.0 1593600.0 1210800.0 1607400.0 ;
      RECT  1200600.0 1621200.0 1210800.0 1607400.0 ;
      RECT  1200600.0 1621200.0 1210800.0 1635000.0 ;
      RECT  1200600.0 1648800.0 1210800.0 1635000.0 ;
      RECT  1200600.0 1648800.0 1210800.0 1662600.0 ;
      RECT  1200600.0 1676400.0 1210800.0 1662600.0 ;
      RECT  1200600.0 1676400.0 1210800.0 1690200.0 ;
      RECT  1200600.0 1704000.0 1210800.0 1690200.0 ;
      RECT  1200600.0 1704000.0 1210800.0 1717800.0 ;
      RECT  1200600.0 1731600.0 1210800.0 1717800.0 ;
      RECT  1200600.0 1731600.0 1210800.0 1745400.0 ;
      RECT  1200600.0 1759200.0 1210800.0 1745400.0 ;
      RECT  1200600.0 1759200.0 1210800.0 1773000.0 ;
      RECT  1200600.0 1786800.0 1210800.0 1773000.0 ;
      RECT  1200600.0 1786800.0 1210800.0 1800600.0 ;
      RECT  1200600.0 1814400.0 1210800.0 1800600.0 ;
      RECT  1200600.0 1814400.0 1210800.0 1828200.0 ;
      RECT  1200600.0 1842000.0 1210800.0 1828200.0 ;
      RECT  1200600.0 1842000.0 1210800.0 1855800.0 ;
      RECT  1200600.0 1869600.0 1210800.0 1855800.0 ;
      RECT  1200600.0 1869600.0 1210800.0 1883400.0 ;
      RECT  1200600.0 1897200.0 1210800.0 1883400.0 ;
      RECT  1200600.0 1897200.0 1210800.0 1911000.0 ;
      RECT  1200600.0 1924800.0 1210800.0 1911000.0 ;
      RECT  1200600.0 1924800.0 1210800.0 1938600.0 ;
      RECT  1200600.0 1952400.0 1210800.0 1938600.0 ;
      RECT  1200600.0 1952400.0 1210800.0 1966200.0 ;
      RECT  1200600.0 1980000.0 1210800.0 1966200.0 ;
      RECT  1200600.0 1980000.0 1210800.0 1993800.0 ;
      RECT  1200600.0 2007600.0 1210800.0 1993800.0 ;
      RECT  1200600.0 2007600.0 1210800.0 2021400.0 ;
      RECT  1200600.0 2035200.0 1210800.0 2021400.0 ;
      RECT  1200600.0 2035200.0 1210800.0 2049000.0 ;
      RECT  1200600.0 2062800.0 1210800.0 2049000.0 ;
      RECT  1200600.0 2062800.0 1210800.0 2076600.0 ;
      RECT  1200600.0 2090400.0 1210800.0 2076600.0 ;
      RECT  1200600.0 2090400.0 1210800.0 2104200.0 ;
      RECT  1200600.0 2118000.0 1210800.0 2104200.0 ;
      RECT  1200600.0 2118000.0 1210800.0 2131800.0 ;
      RECT  1200600.0 2145600.0 1210800.0 2131800.0 ;
      RECT  1210800.0 379200.0 1221000.0 393000.0 ;
      RECT  1210800.0 406800.0 1221000.0 393000.0 ;
      RECT  1210800.0 406800.0 1221000.0 420600.0 ;
      RECT  1210800.0 434400.0 1221000.0 420600.0 ;
      RECT  1210800.0 434400.0 1221000.0 448200.0 ;
      RECT  1210800.0 462000.0 1221000.0 448200.0 ;
      RECT  1210800.0 462000.0 1221000.0 475800.0 ;
      RECT  1210800.0 489600.0 1221000.0 475800.0 ;
      RECT  1210800.0 489600.0 1221000.0 503400.0 ;
      RECT  1210800.0 517200.0 1221000.0 503400.0 ;
      RECT  1210800.0 517200.0 1221000.0 531000.0 ;
      RECT  1210800.0 544800.0 1221000.0 531000.0 ;
      RECT  1210800.0 544800.0 1221000.0 558600.0 ;
      RECT  1210800.0 572400.0 1221000.0 558600.0 ;
      RECT  1210800.0 572400.0 1221000.0 586200.0 ;
      RECT  1210800.0 600000.0 1221000.0 586200.0 ;
      RECT  1210800.0 600000.0 1221000.0 613800.0 ;
      RECT  1210800.0 627600.0 1221000.0 613800.0 ;
      RECT  1210800.0 627600.0 1221000.0 641400.0 ;
      RECT  1210800.0 655200.0 1221000.0 641400.0 ;
      RECT  1210800.0 655200.0 1221000.0 669000.0 ;
      RECT  1210800.0 682800.0 1221000.0 669000.0 ;
      RECT  1210800.0 682800.0 1221000.0 696600.0 ;
      RECT  1210800.0 710400.0 1221000.0 696600.0 ;
      RECT  1210800.0 710400.0 1221000.0 724200.0 ;
      RECT  1210800.0 738000.0 1221000.0 724200.0 ;
      RECT  1210800.0 738000.0 1221000.0 751800.0 ;
      RECT  1210800.0 765600.0 1221000.0 751800.0 ;
      RECT  1210800.0 765600.0 1221000.0 779400.0 ;
      RECT  1210800.0 793200.0 1221000.0 779400.0 ;
      RECT  1210800.0 793200.0 1221000.0 807000.0 ;
      RECT  1210800.0 820800.0 1221000.0 807000.0 ;
      RECT  1210800.0 820800.0 1221000.0 834600.0 ;
      RECT  1210800.0 848400.0 1221000.0 834600.0 ;
      RECT  1210800.0 848400.0 1221000.0 862200.0 ;
      RECT  1210800.0 876000.0 1221000.0 862200.0 ;
      RECT  1210800.0 876000.0 1221000.0 889800.0 ;
      RECT  1210800.0 903600.0 1221000.0 889800.0 ;
      RECT  1210800.0 903600.0 1221000.0 917400.0 ;
      RECT  1210800.0 931200.0 1221000.0 917400.0 ;
      RECT  1210800.0 931200.0 1221000.0 945000.0 ;
      RECT  1210800.0 958800.0 1221000.0 945000.0 ;
      RECT  1210800.0 958800.0 1221000.0 972600.0 ;
      RECT  1210800.0 986400.0 1221000.0 972600.0 ;
      RECT  1210800.0 986400.0 1221000.0 1000200.0 ;
      RECT  1210800.0 1014000.0 1221000.0 1000200.0 ;
      RECT  1210800.0 1014000.0 1221000.0 1027800.0 ;
      RECT  1210800.0 1041600.0 1221000.0 1027800.0 ;
      RECT  1210800.0 1041600.0 1221000.0 1055400.0 ;
      RECT  1210800.0 1069200.0 1221000.0 1055400.0 ;
      RECT  1210800.0 1069200.0 1221000.0 1083000.0 ;
      RECT  1210800.0 1096800.0 1221000.0 1083000.0 ;
      RECT  1210800.0 1096800.0 1221000.0 1110600.0 ;
      RECT  1210800.0 1124400.0 1221000.0 1110600.0 ;
      RECT  1210800.0 1124400.0 1221000.0 1138200.0 ;
      RECT  1210800.0 1152000.0 1221000.0 1138200.0 ;
      RECT  1210800.0 1152000.0 1221000.0 1165800.0 ;
      RECT  1210800.0 1179600.0 1221000.0 1165800.0 ;
      RECT  1210800.0 1179600.0 1221000.0 1193400.0 ;
      RECT  1210800.0 1207200.0 1221000.0 1193400.0 ;
      RECT  1210800.0 1207200.0 1221000.0 1221000.0 ;
      RECT  1210800.0 1234800.0 1221000.0 1221000.0 ;
      RECT  1210800.0 1234800.0 1221000.0 1248600.0 ;
      RECT  1210800.0 1262400.0 1221000.0 1248600.0 ;
      RECT  1210800.0 1262400.0 1221000.0 1276200.0 ;
      RECT  1210800.0 1290000.0 1221000.0 1276200.0 ;
      RECT  1210800.0 1290000.0 1221000.0 1303800.0 ;
      RECT  1210800.0 1317600.0 1221000.0 1303800.0 ;
      RECT  1210800.0 1317600.0 1221000.0 1331400.0 ;
      RECT  1210800.0 1345200.0 1221000.0 1331400.0 ;
      RECT  1210800.0 1345200.0 1221000.0 1359000.0 ;
      RECT  1210800.0 1372800.0 1221000.0 1359000.0 ;
      RECT  1210800.0 1372800.0 1221000.0 1386600.0 ;
      RECT  1210800.0 1400400.0 1221000.0 1386600.0 ;
      RECT  1210800.0 1400400.0 1221000.0 1414200.0 ;
      RECT  1210800.0 1428000.0 1221000.0 1414200.0 ;
      RECT  1210800.0 1428000.0 1221000.0 1441800.0 ;
      RECT  1210800.0 1455600.0 1221000.0 1441800.0 ;
      RECT  1210800.0 1455600.0 1221000.0 1469400.0 ;
      RECT  1210800.0 1483200.0 1221000.0 1469400.0 ;
      RECT  1210800.0 1483200.0 1221000.0 1497000.0 ;
      RECT  1210800.0 1510800.0 1221000.0 1497000.0 ;
      RECT  1210800.0 1510800.0 1221000.0 1524600.0 ;
      RECT  1210800.0 1538400.0 1221000.0 1524600.0 ;
      RECT  1210800.0 1538400.0 1221000.0 1552200.0 ;
      RECT  1210800.0 1566000.0 1221000.0 1552200.0 ;
      RECT  1210800.0 1566000.0 1221000.0 1579800.0 ;
      RECT  1210800.0 1593600.0 1221000.0 1579800.0 ;
      RECT  1210800.0 1593600.0 1221000.0 1607400.0 ;
      RECT  1210800.0 1621200.0 1221000.0 1607400.0 ;
      RECT  1210800.0 1621200.0 1221000.0 1635000.0 ;
      RECT  1210800.0 1648800.0 1221000.0 1635000.0 ;
      RECT  1210800.0 1648800.0 1221000.0 1662600.0 ;
      RECT  1210800.0 1676400.0 1221000.0 1662600.0 ;
      RECT  1210800.0 1676400.0 1221000.0 1690200.0 ;
      RECT  1210800.0 1704000.0 1221000.0 1690200.0 ;
      RECT  1210800.0 1704000.0 1221000.0 1717800.0 ;
      RECT  1210800.0 1731600.0 1221000.0 1717800.0 ;
      RECT  1210800.0 1731600.0 1221000.0 1745400.0 ;
      RECT  1210800.0 1759200.0 1221000.0 1745400.0 ;
      RECT  1210800.0 1759200.0 1221000.0 1773000.0 ;
      RECT  1210800.0 1786800.0 1221000.0 1773000.0 ;
      RECT  1210800.0 1786800.0 1221000.0 1800600.0 ;
      RECT  1210800.0 1814400.0 1221000.0 1800600.0 ;
      RECT  1210800.0 1814400.0 1221000.0 1828200.0 ;
      RECT  1210800.0 1842000.0 1221000.0 1828200.0 ;
      RECT  1210800.0 1842000.0 1221000.0 1855800.0 ;
      RECT  1210800.0 1869600.0 1221000.0 1855800.0 ;
      RECT  1210800.0 1869600.0 1221000.0 1883400.0 ;
      RECT  1210800.0 1897200.0 1221000.0 1883400.0 ;
      RECT  1210800.0 1897200.0 1221000.0 1911000.0 ;
      RECT  1210800.0 1924800.0 1221000.0 1911000.0 ;
      RECT  1210800.0 1924800.0 1221000.0 1938600.0 ;
      RECT  1210800.0 1952400.0 1221000.0 1938600.0 ;
      RECT  1210800.0 1952400.0 1221000.0 1966200.0 ;
      RECT  1210800.0 1980000.0 1221000.0 1966200.0 ;
      RECT  1210800.0 1980000.0 1221000.0 1993800.0 ;
      RECT  1210800.0 2007600.0 1221000.0 1993800.0 ;
      RECT  1210800.0 2007600.0 1221000.0 2021400.0 ;
      RECT  1210800.0 2035200.0 1221000.0 2021400.0 ;
      RECT  1210800.0 2035200.0 1221000.0 2049000.0 ;
      RECT  1210800.0 2062800.0 1221000.0 2049000.0 ;
      RECT  1210800.0 2062800.0 1221000.0 2076600.0 ;
      RECT  1210800.0 2090400.0 1221000.0 2076600.0 ;
      RECT  1210800.0 2090400.0 1221000.0 2104200.0 ;
      RECT  1210800.0 2118000.0 1221000.0 2104200.0 ;
      RECT  1210800.0 2118000.0 1221000.0 2131800.0 ;
      RECT  1210800.0 2145600.0 1221000.0 2131800.0 ;
      RECT  1221000.0 379200.0 1231200.0 393000.0 ;
      RECT  1221000.0 406800.0 1231200.0 393000.0 ;
      RECT  1221000.0 406800.0 1231200.0 420600.0 ;
      RECT  1221000.0 434400.0 1231200.0 420600.0 ;
      RECT  1221000.0 434400.0 1231200.0 448200.0 ;
      RECT  1221000.0 462000.0 1231200.0 448200.0 ;
      RECT  1221000.0 462000.0 1231200.0 475800.0 ;
      RECT  1221000.0 489600.0 1231200.0 475800.0 ;
      RECT  1221000.0 489600.0 1231200.0 503400.0 ;
      RECT  1221000.0 517200.0 1231200.0 503400.0 ;
      RECT  1221000.0 517200.0 1231200.0 531000.0 ;
      RECT  1221000.0 544800.0 1231200.0 531000.0 ;
      RECT  1221000.0 544800.0 1231200.0 558600.0 ;
      RECT  1221000.0 572400.0 1231200.0 558600.0 ;
      RECT  1221000.0 572400.0 1231200.0 586200.0 ;
      RECT  1221000.0 600000.0 1231200.0 586200.0 ;
      RECT  1221000.0 600000.0 1231200.0 613800.0 ;
      RECT  1221000.0 627600.0 1231200.0 613800.0 ;
      RECT  1221000.0 627600.0 1231200.0 641400.0 ;
      RECT  1221000.0 655200.0 1231200.0 641400.0 ;
      RECT  1221000.0 655200.0 1231200.0 669000.0 ;
      RECT  1221000.0 682800.0 1231200.0 669000.0 ;
      RECT  1221000.0 682800.0 1231200.0 696600.0 ;
      RECT  1221000.0 710400.0 1231200.0 696600.0 ;
      RECT  1221000.0 710400.0 1231200.0 724200.0 ;
      RECT  1221000.0 738000.0 1231200.0 724200.0 ;
      RECT  1221000.0 738000.0 1231200.0 751800.0 ;
      RECT  1221000.0 765600.0 1231200.0 751800.0 ;
      RECT  1221000.0 765600.0 1231200.0 779400.0 ;
      RECT  1221000.0 793200.0 1231200.0 779400.0 ;
      RECT  1221000.0 793200.0 1231200.0 807000.0 ;
      RECT  1221000.0 820800.0 1231200.0 807000.0 ;
      RECT  1221000.0 820800.0 1231200.0 834600.0 ;
      RECT  1221000.0 848400.0 1231200.0 834600.0 ;
      RECT  1221000.0 848400.0 1231200.0 862200.0 ;
      RECT  1221000.0 876000.0 1231200.0 862200.0 ;
      RECT  1221000.0 876000.0 1231200.0 889800.0 ;
      RECT  1221000.0 903600.0 1231200.0 889800.0 ;
      RECT  1221000.0 903600.0 1231200.0 917400.0 ;
      RECT  1221000.0 931200.0 1231200.0 917400.0 ;
      RECT  1221000.0 931200.0 1231200.0 945000.0 ;
      RECT  1221000.0 958800.0 1231200.0 945000.0 ;
      RECT  1221000.0 958800.0 1231200.0 972600.0 ;
      RECT  1221000.0 986400.0 1231200.0 972600.0 ;
      RECT  1221000.0 986400.0 1231200.0 1000200.0 ;
      RECT  1221000.0 1014000.0 1231200.0 1000200.0 ;
      RECT  1221000.0 1014000.0 1231200.0 1027800.0 ;
      RECT  1221000.0 1041600.0 1231200.0 1027800.0 ;
      RECT  1221000.0 1041600.0 1231200.0 1055400.0 ;
      RECT  1221000.0 1069200.0 1231200.0 1055400.0 ;
      RECT  1221000.0 1069200.0 1231200.0 1083000.0 ;
      RECT  1221000.0 1096800.0 1231200.0 1083000.0 ;
      RECT  1221000.0 1096800.0 1231200.0 1110600.0 ;
      RECT  1221000.0 1124400.0 1231200.0 1110600.0 ;
      RECT  1221000.0 1124400.0 1231200.0 1138200.0 ;
      RECT  1221000.0 1152000.0 1231200.0 1138200.0 ;
      RECT  1221000.0 1152000.0 1231200.0 1165800.0 ;
      RECT  1221000.0 1179600.0 1231200.0 1165800.0 ;
      RECT  1221000.0 1179600.0 1231200.0 1193400.0 ;
      RECT  1221000.0 1207200.0 1231200.0 1193400.0 ;
      RECT  1221000.0 1207200.0 1231200.0 1221000.0 ;
      RECT  1221000.0 1234800.0 1231200.0 1221000.0 ;
      RECT  1221000.0 1234800.0 1231200.0 1248600.0 ;
      RECT  1221000.0 1262400.0 1231200.0 1248600.0 ;
      RECT  1221000.0 1262400.0 1231200.0 1276200.0 ;
      RECT  1221000.0 1290000.0 1231200.0 1276200.0 ;
      RECT  1221000.0 1290000.0 1231200.0 1303800.0 ;
      RECT  1221000.0 1317600.0 1231200.0 1303800.0 ;
      RECT  1221000.0 1317600.0 1231200.0 1331400.0 ;
      RECT  1221000.0 1345200.0 1231200.0 1331400.0 ;
      RECT  1221000.0 1345200.0 1231200.0 1359000.0 ;
      RECT  1221000.0 1372800.0 1231200.0 1359000.0 ;
      RECT  1221000.0 1372800.0 1231200.0 1386600.0 ;
      RECT  1221000.0 1400400.0 1231200.0 1386600.0 ;
      RECT  1221000.0 1400400.0 1231200.0 1414200.0 ;
      RECT  1221000.0 1428000.0 1231200.0 1414200.0 ;
      RECT  1221000.0 1428000.0 1231200.0 1441800.0 ;
      RECT  1221000.0 1455600.0 1231200.0 1441800.0 ;
      RECT  1221000.0 1455600.0 1231200.0 1469400.0 ;
      RECT  1221000.0 1483200.0 1231200.0 1469400.0 ;
      RECT  1221000.0 1483200.0 1231200.0 1497000.0 ;
      RECT  1221000.0 1510800.0 1231200.0 1497000.0 ;
      RECT  1221000.0 1510800.0 1231200.0 1524600.0 ;
      RECT  1221000.0 1538400.0 1231200.0 1524600.0 ;
      RECT  1221000.0 1538400.0 1231200.0 1552200.0 ;
      RECT  1221000.0 1566000.0 1231200.0 1552200.0 ;
      RECT  1221000.0 1566000.0 1231200.0 1579800.0 ;
      RECT  1221000.0 1593600.0 1231200.0 1579800.0 ;
      RECT  1221000.0 1593600.0 1231200.0 1607400.0 ;
      RECT  1221000.0 1621200.0 1231200.0 1607400.0 ;
      RECT  1221000.0 1621200.0 1231200.0 1635000.0 ;
      RECT  1221000.0 1648800.0 1231200.0 1635000.0 ;
      RECT  1221000.0 1648800.0 1231200.0 1662600.0 ;
      RECT  1221000.0 1676400.0 1231200.0 1662600.0 ;
      RECT  1221000.0 1676400.0 1231200.0 1690200.0 ;
      RECT  1221000.0 1704000.0 1231200.0 1690200.0 ;
      RECT  1221000.0 1704000.0 1231200.0 1717800.0 ;
      RECT  1221000.0 1731600.0 1231200.0 1717800.0 ;
      RECT  1221000.0 1731600.0 1231200.0 1745400.0 ;
      RECT  1221000.0 1759200.0 1231200.0 1745400.0 ;
      RECT  1221000.0 1759200.0 1231200.0 1773000.0 ;
      RECT  1221000.0 1786800.0 1231200.0 1773000.0 ;
      RECT  1221000.0 1786800.0 1231200.0 1800600.0 ;
      RECT  1221000.0 1814400.0 1231200.0 1800600.0 ;
      RECT  1221000.0 1814400.0 1231200.0 1828200.0 ;
      RECT  1221000.0 1842000.0 1231200.0 1828200.0 ;
      RECT  1221000.0 1842000.0 1231200.0 1855800.0 ;
      RECT  1221000.0 1869600.0 1231200.0 1855800.0 ;
      RECT  1221000.0 1869600.0 1231200.0 1883400.0 ;
      RECT  1221000.0 1897200.0 1231200.0 1883400.0 ;
      RECT  1221000.0 1897200.0 1231200.0 1911000.0 ;
      RECT  1221000.0 1924800.0 1231200.0 1911000.0 ;
      RECT  1221000.0 1924800.0 1231200.0 1938600.0 ;
      RECT  1221000.0 1952400.0 1231200.0 1938600.0 ;
      RECT  1221000.0 1952400.0 1231200.0 1966200.0 ;
      RECT  1221000.0 1980000.0 1231200.0 1966200.0 ;
      RECT  1221000.0 1980000.0 1231200.0 1993800.0 ;
      RECT  1221000.0 2007600.0 1231200.0 1993800.0 ;
      RECT  1221000.0 2007600.0 1231200.0 2021400.0 ;
      RECT  1221000.0 2035200.0 1231200.0 2021400.0 ;
      RECT  1221000.0 2035200.0 1231200.0 2049000.0 ;
      RECT  1221000.0 2062800.0 1231200.0 2049000.0 ;
      RECT  1221000.0 2062800.0 1231200.0 2076600.0 ;
      RECT  1221000.0 2090400.0 1231200.0 2076600.0 ;
      RECT  1221000.0 2090400.0 1231200.0 2104200.0 ;
      RECT  1221000.0 2118000.0 1231200.0 2104200.0 ;
      RECT  1221000.0 2118000.0 1231200.0 2131800.0 ;
      RECT  1221000.0 2145600.0 1231200.0 2131800.0 ;
      RECT  1231200.0 379200.0 1241400.0 393000.0 ;
      RECT  1231200.0 406800.0 1241400.0 393000.0 ;
      RECT  1231200.0 406800.0 1241400.0 420600.0 ;
      RECT  1231200.0 434400.0 1241400.0 420600.0 ;
      RECT  1231200.0 434400.0 1241400.0 448200.0 ;
      RECT  1231200.0 462000.0 1241400.0 448200.0 ;
      RECT  1231200.0 462000.0 1241400.0 475800.0 ;
      RECT  1231200.0 489600.0 1241400.0 475800.0 ;
      RECT  1231200.0 489600.0 1241400.0 503400.0 ;
      RECT  1231200.0 517200.0 1241400.0 503400.0 ;
      RECT  1231200.0 517200.0 1241400.0 531000.0 ;
      RECT  1231200.0 544800.0 1241400.0 531000.0 ;
      RECT  1231200.0 544800.0 1241400.0 558600.0 ;
      RECT  1231200.0 572400.0 1241400.0 558600.0 ;
      RECT  1231200.0 572400.0 1241400.0 586200.0 ;
      RECT  1231200.0 600000.0 1241400.0 586200.0 ;
      RECT  1231200.0 600000.0 1241400.0 613800.0 ;
      RECT  1231200.0 627600.0 1241400.0 613800.0 ;
      RECT  1231200.0 627600.0 1241400.0 641400.0 ;
      RECT  1231200.0 655200.0 1241400.0 641400.0 ;
      RECT  1231200.0 655200.0 1241400.0 669000.0 ;
      RECT  1231200.0 682800.0 1241400.0 669000.0 ;
      RECT  1231200.0 682800.0 1241400.0 696600.0 ;
      RECT  1231200.0 710400.0 1241400.0 696600.0 ;
      RECT  1231200.0 710400.0 1241400.0 724200.0 ;
      RECT  1231200.0 738000.0 1241400.0 724200.0 ;
      RECT  1231200.0 738000.0 1241400.0 751800.0 ;
      RECT  1231200.0 765600.0 1241400.0 751800.0 ;
      RECT  1231200.0 765600.0 1241400.0 779400.0 ;
      RECT  1231200.0 793200.0 1241400.0 779400.0 ;
      RECT  1231200.0 793200.0 1241400.0 807000.0 ;
      RECT  1231200.0 820800.0 1241400.0 807000.0 ;
      RECT  1231200.0 820800.0 1241400.0 834600.0 ;
      RECT  1231200.0 848400.0 1241400.0 834600.0 ;
      RECT  1231200.0 848400.0 1241400.0 862200.0 ;
      RECT  1231200.0 876000.0 1241400.0 862200.0 ;
      RECT  1231200.0 876000.0 1241400.0 889800.0 ;
      RECT  1231200.0 903600.0 1241400.0 889800.0 ;
      RECT  1231200.0 903600.0 1241400.0 917400.0 ;
      RECT  1231200.0 931200.0 1241400.0 917400.0 ;
      RECT  1231200.0 931200.0 1241400.0 945000.0 ;
      RECT  1231200.0 958800.0 1241400.0 945000.0 ;
      RECT  1231200.0 958800.0 1241400.0 972600.0 ;
      RECT  1231200.0 986400.0 1241400.0 972600.0 ;
      RECT  1231200.0 986400.0 1241400.0 1000200.0 ;
      RECT  1231200.0 1014000.0 1241400.0 1000200.0 ;
      RECT  1231200.0 1014000.0 1241400.0 1027800.0 ;
      RECT  1231200.0 1041600.0 1241400.0 1027800.0 ;
      RECT  1231200.0 1041600.0 1241400.0 1055400.0 ;
      RECT  1231200.0 1069200.0 1241400.0 1055400.0 ;
      RECT  1231200.0 1069200.0 1241400.0 1083000.0 ;
      RECT  1231200.0 1096800.0 1241400.0 1083000.0 ;
      RECT  1231200.0 1096800.0 1241400.0 1110600.0 ;
      RECT  1231200.0 1124400.0 1241400.0 1110600.0 ;
      RECT  1231200.0 1124400.0 1241400.0 1138200.0 ;
      RECT  1231200.0 1152000.0 1241400.0 1138200.0 ;
      RECT  1231200.0 1152000.0 1241400.0 1165800.0 ;
      RECT  1231200.0 1179600.0 1241400.0 1165800.0 ;
      RECT  1231200.0 1179600.0 1241400.0 1193400.0 ;
      RECT  1231200.0 1207200.0 1241400.0 1193400.0 ;
      RECT  1231200.0 1207200.0 1241400.0 1221000.0 ;
      RECT  1231200.0 1234800.0 1241400.0 1221000.0 ;
      RECT  1231200.0 1234800.0 1241400.0 1248600.0 ;
      RECT  1231200.0 1262400.0 1241400.0 1248600.0 ;
      RECT  1231200.0 1262400.0 1241400.0 1276200.0 ;
      RECT  1231200.0 1290000.0 1241400.0 1276200.0 ;
      RECT  1231200.0 1290000.0 1241400.0 1303800.0 ;
      RECT  1231200.0 1317600.0 1241400.0 1303800.0 ;
      RECT  1231200.0 1317600.0 1241400.0 1331400.0 ;
      RECT  1231200.0 1345200.0 1241400.0 1331400.0 ;
      RECT  1231200.0 1345200.0 1241400.0 1359000.0 ;
      RECT  1231200.0 1372800.0 1241400.0 1359000.0 ;
      RECT  1231200.0 1372800.0 1241400.0 1386600.0 ;
      RECT  1231200.0 1400400.0 1241400.0 1386600.0 ;
      RECT  1231200.0 1400400.0 1241400.0 1414200.0 ;
      RECT  1231200.0 1428000.0 1241400.0 1414200.0 ;
      RECT  1231200.0 1428000.0 1241400.0 1441800.0 ;
      RECT  1231200.0 1455600.0 1241400.0 1441800.0 ;
      RECT  1231200.0 1455600.0 1241400.0 1469400.0 ;
      RECT  1231200.0 1483200.0 1241400.0 1469400.0 ;
      RECT  1231200.0 1483200.0 1241400.0 1497000.0 ;
      RECT  1231200.0 1510800.0 1241400.0 1497000.0 ;
      RECT  1231200.0 1510800.0 1241400.0 1524600.0 ;
      RECT  1231200.0 1538400.0 1241400.0 1524600.0 ;
      RECT  1231200.0 1538400.0 1241400.0 1552200.0 ;
      RECT  1231200.0 1566000.0 1241400.0 1552200.0 ;
      RECT  1231200.0 1566000.0 1241400.0 1579800.0 ;
      RECT  1231200.0 1593600.0 1241400.0 1579800.0 ;
      RECT  1231200.0 1593600.0 1241400.0 1607400.0 ;
      RECT  1231200.0 1621200.0 1241400.0 1607400.0 ;
      RECT  1231200.0 1621200.0 1241400.0 1635000.0 ;
      RECT  1231200.0 1648800.0 1241400.0 1635000.0 ;
      RECT  1231200.0 1648800.0 1241400.0 1662600.0 ;
      RECT  1231200.0 1676400.0 1241400.0 1662600.0 ;
      RECT  1231200.0 1676400.0 1241400.0 1690200.0 ;
      RECT  1231200.0 1704000.0 1241400.0 1690200.0 ;
      RECT  1231200.0 1704000.0 1241400.0 1717800.0 ;
      RECT  1231200.0 1731600.0 1241400.0 1717800.0 ;
      RECT  1231200.0 1731600.0 1241400.0 1745400.0 ;
      RECT  1231200.0 1759200.0 1241400.0 1745400.0 ;
      RECT  1231200.0 1759200.0 1241400.0 1773000.0 ;
      RECT  1231200.0 1786800.0 1241400.0 1773000.0 ;
      RECT  1231200.0 1786800.0 1241400.0 1800600.0 ;
      RECT  1231200.0 1814400.0 1241400.0 1800600.0 ;
      RECT  1231200.0 1814400.0 1241400.0 1828200.0 ;
      RECT  1231200.0 1842000.0 1241400.0 1828200.0 ;
      RECT  1231200.0 1842000.0 1241400.0 1855800.0 ;
      RECT  1231200.0 1869600.0 1241400.0 1855800.0 ;
      RECT  1231200.0 1869600.0 1241400.0 1883400.0 ;
      RECT  1231200.0 1897200.0 1241400.0 1883400.0 ;
      RECT  1231200.0 1897200.0 1241400.0 1911000.0 ;
      RECT  1231200.0 1924800.0 1241400.0 1911000.0 ;
      RECT  1231200.0 1924800.0 1241400.0 1938600.0 ;
      RECT  1231200.0 1952400.0 1241400.0 1938600.0 ;
      RECT  1231200.0 1952400.0 1241400.0 1966200.0 ;
      RECT  1231200.0 1980000.0 1241400.0 1966200.0 ;
      RECT  1231200.0 1980000.0 1241400.0 1993800.0 ;
      RECT  1231200.0 2007600.0 1241400.0 1993800.0 ;
      RECT  1231200.0 2007600.0 1241400.0 2021400.0 ;
      RECT  1231200.0 2035200.0 1241400.0 2021400.0 ;
      RECT  1231200.0 2035200.0 1241400.0 2049000.0 ;
      RECT  1231200.0 2062800.0 1241400.0 2049000.0 ;
      RECT  1231200.0 2062800.0 1241400.0 2076600.0 ;
      RECT  1231200.0 2090400.0 1241400.0 2076600.0 ;
      RECT  1231200.0 2090400.0 1241400.0 2104200.0 ;
      RECT  1231200.0 2118000.0 1241400.0 2104200.0 ;
      RECT  1231200.0 2118000.0 1241400.0 2131800.0 ;
      RECT  1231200.0 2145600.0 1241400.0 2131800.0 ;
      RECT  1241400.0 379200.0 1251600.0 393000.0 ;
      RECT  1241400.0 406800.0 1251600.0 393000.0 ;
      RECT  1241400.0 406800.0 1251600.0 420600.0 ;
      RECT  1241400.0 434400.0 1251600.0 420600.0 ;
      RECT  1241400.0 434400.0 1251600.0 448200.0 ;
      RECT  1241400.0 462000.0 1251600.0 448200.0 ;
      RECT  1241400.0 462000.0 1251600.0 475800.0 ;
      RECT  1241400.0 489600.0 1251600.0 475800.0 ;
      RECT  1241400.0 489600.0 1251600.0 503400.0 ;
      RECT  1241400.0 517200.0 1251600.0 503400.0 ;
      RECT  1241400.0 517200.0 1251600.0 531000.0 ;
      RECT  1241400.0 544800.0 1251600.0 531000.0 ;
      RECT  1241400.0 544800.0 1251600.0 558600.0 ;
      RECT  1241400.0 572400.0 1251600.0 558600.0 ;
      RECT  1241400.0 572400.0 1251600.0 586200.0 ;
      RECT  1241400.0 600000.0 1251600.0 586200.0 ;
      RECT  1241400.0 600000.0 1251600.0 613800.0 ;
      RECT  1241400.0 627600.0 1251600.0 613800.0 ;
      RECT  1241400.0 627600.0 1251600.0 641400.0 ;
      RECT  1241400.0 655200.0 1251600.0 641400.0 ;
      RECT  1241400.0 655200.0 1251600.0 669000.0 ;
      RECT  1241400.0 682800.0 1251600.0 669000.0 ;
      RECT  1241400.0 682800.0 1251600.0 696600.0 ;
      RECT  1241400.0 710400.0 1251600.0 696600.0 ;
      RECT  1241400.0 710400.0 1251600.0 724200.0 ;
      RECT  1241400.0 738000.0 1251600.0 724200.0 ;
      RECT  1241400.0 738000.0 1251600.0 751800.0 ;
      RECT  1241400.0 765600.0 1251600.0 751800.0 ;
      RECT  1241400.0 765600.0 1251600.0 779400.0 ;
      RECT  1241400.0 793200.0 1251600.0 779400.0 ;
      RECT  1241400.0 793200.0 1251600.0 807000.0 ;
      RECT  1241400.0 820800.0 1251600.0 807000.0 ;
      RECT  1241400.0 820800.0 1251600.0 834600.0 ;
      RECT  1241400.0 848400.0 1251600.0 834600.0 ;
      RECT  1241400.0 848400.0 1251600.0 862200.0 ;
      RECT  1241400.0 876000.0 1251600.0 862200.0 ;
      RECT  1241400.0 876000.0 1251600.0 889800.0 ;
      RECT  1241400.0 903600.0 1251600.0 889800.0 ;
      RECT  1241400.0 903600.0 1251600.0 917400.0 ;
      RECT  1241400.0 931200.0 1251600.0 917400.0 ;
      RECT  1241400.0 931200.0 1251600.0 945000.0 ;
      RECT  1241400.0 958800.0 1251600.0 945000.0 ;
      RECT  1241400.0 958800.0 1251600.0 972600.0 ;
      RECT  1241400.0 986400.0 1251600.0 972600.0 ;
      RECT  1241400.0 986400.0 1251600.0 1000200.0 ;
      RECT  1241400.0 1014000.0 1251600.0 1000200.0 ;
      RECT  1241400.0 1014000.0 1251600.0 1027800.0 ;
      RECT  1241400.0 1041600.0 1251600.0 1027800.0 ;
      RECT  1241400.0 1041600.0 1251600.0 1055400.0 ;
      RECT  1241400.0 1069200.0 1251600.0 1055400.0 ;
      RECT  1241400.0 1069200.0 1251600.0 1083000.0 ;
      RECT  1241400.0 1096800.0 1251600.0 1083000.0 ;
      RECT  1241400.0 1096800.0 1251600.0 1110600.0 ;
      RECT  1241400.0 1124400.0 1251600.0 1110600.0 ;
      RECT  1241400.0 1124400.0 1251600.0 1138200.0 ;
      RECT  1241400.0 1152000.0 1251600.0 1138200.0 ;
      RECT  1241400.0 1152000.0 1251600.0 1165800.0 ;
      RECT  1241400.0 1179600.0 1251600.0 1165800.0 ;
      RECT  1241400.0 1179600.0 1251600.0 1193400.0 ;
      RECT  1241400.0 1207200.0 1251600.0 1193400.0 ;
      RECT  1241400.0 1207200.0 1251600.0 1221000.0 ;
      RECT  1241400.0 1234800.0 1251600.0 1221000.0 ;
      RECT  1241400.0 1234800.0 1251600.0 1248600.0 ;
      RECT  1241400.0 1262400.0 1251600.0 1248600.0 ;
      RECT  1241400.0 1262400.0 1251600.0 1276200.0 ;
      RECT  1241400.0 1290000.0 1251600.0 1276200.0 ;
      RECT  1241400.0 1290000.0 1251600.0 1303800.0 ;
      RECT  1241400.0 1317600.0 1251600.0 1303800.0 ;
      RECT  1241400.0 1317600.0 1251600.0 1331400.0 ;
      RECT  1241400.0 1345200.0 1251600.0 1331400.0 ;
      RECT  1241400.0 1345200.0 1251600.0 1359000.0 ;
      RECT  1241400.0 1372800.0 1251600.0 1359000.0 ;
      RECT  1241400.0 1372800.0 1251600.0 1386600.0 ;
      RECT  1241400.0 1400400.0 1251600.0 1386600.0 ;
      RECT  1241400.0 1400400.0 1251600.0 1414200.0 ;
      RECT  1241400.0 1428000.0 1251600.0 1414200.0 ;
      RECT  1241400.0 1428000.0 1251600.0 1441800.0 ;
      RECT  1241400.0 1455600.0 1251600.0 1441800.0 ;
      RECT  1241400.0 1455600.0 1251600.0 1469400.0 ;
      RECT  1241400.0 1483200.0 1251600.0 1469400.0 ;
      RECT  1241400.0 1483200.0 1251600.0 1497000.0 ;
      RECT  1241400.0 1510800.0 1251600.0 1497000.0 ;
      RECT  1241400.0 1510800.0 1251600.0 1524600.0 ;
      RECT  1241400.0 1538400.0 1251600.0 1524600.0 ;
      RECT  1241400.0 1538400.0 1251600.0 1552200.0 ;
      RECT  1241400.0 1566000.0 1251600.0 1552200.0 ;
      RECT  1241400.0 1566000.0 1251600.0 1579800.0 ;
      RECT  1241400.0 1593600.0 1251600.0 1579800.0 ;
      RECT  1241400.0 1593600.0 1251600.0 1607400.0 ;
      RECT  1241400.0 1621200.0 1251600.0 1607400.0 ;
      RECT  1241400.0 1621200.0 1251600.0 1635000.0 ;
      RECT  1241400.0 1648800.0 1251600.0 1635000.0 ;
      RECT  1241400.0 1648800.0 1251600.0 1662600.0 ;
      RECT  1241400.0 1676400.0 1251600.0 1662600.0 ;
      RECT  1241400.0 1676400.0 1251600.0 1690200.0 ;
      RECT  1241400.0 1704000.0 1251600.0 1690200.0 ;
      RECT  1241400.0 1704000.0 1251600.0 1717800.0 ;
      RECT  1241400.0 1731600.0 1251600.0 1717800.0 ;
      RECT  1241400.0 1731600.0 1251600.0 1745400.0 ;
      RECT  1241400.0 1759200.0 1251600.0 1745400.0 ;
      RECT  1241400.0 1759200.0 1251600.0 1773000.0 ;
      RECT  1241400.0 1786800.0 1251600.0 1773000.0 ;
      RECT  1241400.0 1786800.0 1251600.0 1800600.0 ;
      RECT  1241400.0 1814400.0 1251600.0 1800600.0 ;
      RECT  1241400.0 1814400.0 1251600.0 1828200.0 ;
      RECT  1241400.0 1842000.0 1251600.0 1828200.0 ;
      RECT  1241400.0 1842000.0 1251600.0 1855800.0 ;
      RECT  1241400.0 1869600.0 1251600.0 1855800.0 ;
      RECT  1241400.0 1869600.0 1251600.0 1883400.0 ;
      RECT  1241400.0 1897200.0 1251600.0 1883400.0 ;
      RECT  1241400.0 1897200.0 1251600.0 1911000.0 ;
      RECT  1241400.0 1924800.0 1251600.0 1911000.0 ;
      RECT  1241400.0 1924800.0 1251600.0 1938600.0 ;
      RECT  1241400.0 1952400.0 1251600.0 1938600.0 ;
      RECT  1241400.0 1952400.0 1251600.0 1966200.0 ;
      RECT  1241400.0 1980000.0 1251600.0 1966200.0 ;
      RECT  1241400.0 1980000.0 1251600.0 1993800.0 ;
      RECT  1241400.0 2007600.0 1251600.0 1993800.0 ;
      RECT  1241400.0 2007600.0 1251600.0 2021400.0 ;
      RECT  1241400.0 2035200.0 1251600.0 2021400.0 ;
      RECT  1241400.0 2035200.0 1251600.0 2049000.0 ;
      RECT  1241400.0 2062800.0 1251600.0 2049000.0 ;
      RECT  1241400.0 2062800.0 1251600.0 2076600.0 ;
      RECT  1241400.0 2090400.0 1251600.0 2076600.0 ;
      RECT  1241400.0 2090400.0 1251600.0 2104200.0 ;
      RECT  1241400.0 2118000.0 1251600.0 2104200.0 ;
      RECT  1241400.0 2118000.0 1251600.0 2131800.0 ;
      RECT  1241400.0 2145600.0 1251600.0 2131800.0 ;
      RECT  1251600.0 379200.0 1261800.0 393000.0 ;
      RECT  1251600.0 406800.0 1261800.0 393000.0 ;
      RECT  1251600.0 406800.0 1261800.0 420600.0 ;
      RECT  1251600.0 434400.0 1261800.0 420600.0 ;
      RECT  1251600.0 434400.0 1261800.0 448200.0 ;
      RECT  1251600.0 462000.0 1261800.0 448200.0 ;
      RECT  1251600.0 462000.0 1261800.0 475800.0 ;
      RECT  1251600.0 489600.0 1261800.0 475800.0 ;
      RECT  1251600.0 489600.0 1261800.0 503400.0 ;
      RECT  1251600.0 517200.0 1261800.0 503400.0 ;
      RECT  1251600.0 517200.0 1261800.0 531000.0 ;
      RECT  1251600.0 544800.0 1261800.0 531000.0 ;
      RECT  1251600.0 544800.0 1261800.0 558600.0 ;
      RECT  1251600.0 572400.0 1261800.0 558600.0 ;
      RECT  1251600.0 572400.0 1261800.0 586200.0 ;
      RECT  1251600.0 600000.0 1261800.0 586200.0 ;
      RECT  1251600.0 600000.0 1261800.0 613800.0 ;
      RECT  1251600.0 627600.0 1261800.0 613800.0 ;
      RECT  1251600.0 627600.0 1261800.0 641400.0 ;
      RECT  1251600.0 655200.0 1261800.0 641400.0 ;
      RECT  1251600.0 655200.0 1261800.0 669000.0 ;
      RECT  1251600.0 682800.0 1261800.0 669000.0 ;
      RECT  1251600.0 682800.0 1261800.0 696600.0 ;
      RECT  1251600.0 710400.0 1261800.0 696600.0 ;
      RECT  1251600.0 710400.0 1261800.0 724200.0 ;
      RECT  1251600.0 738000.0 1261800.0 724200.0 ;
      RECT  1251600.0 738000.0 1261800.0 751800.0 ;
      RECT  1251600.0 765600.0 1261800.0 751800.0 ;
      RECT  1251600.0 765600.0 1261800.0 779400.0 ;
      RECT  1251600.0 793200.0 1261800.0 779400.0 ;
      RECT  1251600.0 793200.0 1261800.0 807000.0 ;
      RECT  1251600.0 820800.0 1261800.0 807000.0 ;
      RECT  1251600.0 820800.0 1261800.0 834600.0 ;
      RECT  1251600.0 848400.0 1261800.0 834600.0 ;
      RECT  1251600.0 848400.0 1261800.0 862200.0 ;
      RECT  1251600.0 876000.0 1261800.0 862200.0 ;
      RECT  1251600.0 876000.0 1261800.0 889800.0 ;
      RECT  1251600.0 903600.0 1261800.0 889800.0 ;
      RECT  1251600.0 903600.0 1261800.0 917400.0 ;
      RECT  1251600.0 931200.0 1261800.0 917400.0 ;
      RECT  1251600.0 931200.0 1261800.0 945000.0 ;
      RECT  1251600.0 958800.0 1261800.0 945000.0 ;
      RECT  1251600.0 958800.0 1261800.0 972600.0 ;
      RECT  1251600.0 986400.0 1261800.0 972600.0 ;
      RECT  1251600.0 986400.0 1261800.0 1000200.0 ;
      RECT  1251600.0 1014000.0 1261800.0 1000200.0 ;
      RECT  1251600.0 1014000.0 1261800.0 1027800.0 ;
      RECT  1251600.0 1041600.0 1261800.0 1027800.0 ;
      RECT  1251600.0 1041600.0 1261800.0 1055400.0 ;
      RECT  1251600.0 1069200.0 1261800.0 1055400.0 ;
      RECT  1251600.0 1069200.0 1261800.0 1083000.0 ;
      RECT  1251600.0 1096800.0 1261800.0 1083000.0 ;
      RECT  1251600.0 1096800.0 1261800.0 1110600.0 ;
      RECT  1251600.0 1124400.0 1261800.0 1110600.0 ;
      RECT  1251600.0 1124400.0 1261800.0 1138200.0 ;
      RECT  1251600.0 1152000.0 1261800.0 1138200.0 ;
      RECT  1251600.0 1152000.0 1261800.0 1165800.0 ;
      RECT  1251600.0 1179600.0 1261800.0 1165800.0 ;
      RECT  1251600.0 1179600.0 1261800.0 1193400.0 ;
      RECT  1251600.0 1207200.0 1261800.0 1193400.0 ;
      RECT  1251600.0 1207200.0 1261800.0 1221000.0 ;
      RECT  1251600.0 1234800.0 1261800.0 1221000.0 ;
      RECT  1251600.0 1234800.0 1261800.0 1248600.0 ;
      RECT  1251600.0 1262400.0 1261800.0 1248600.0 ;
      RECT  1251600.0 1262400.0 1261800.0 1276200.0 ;
      RECT  1251600.0 1290000.0 1261800.0 1276200.0 ;
      RECT  1251600.0 1290000.0 1261800.0 1303800.0 ;
      RECT  1251600.0 1317600.0 1261800.0 1303800.0 ;
      RECT  1251600.0 1317600.0 1261800.0 1331400.0 ;
      RECT  1251600.0 1345200.0 1261800.0 1331400.0 ;
      RECT  1251600.0 1345200.0 1261800.0 1359000.0 ;
      RECT  1251600.0 1372800.0 1261800.0 1359000.0 ;
      RECT  1251600.0 1372800.0 1261800.0 1386600.0 ;
      RECT  1251600.0 1400400.0 1261800.0 1386600.0 ;
      RECT  1251600.0 1400400.0 1261800.0 1414200.0 ;
      RECT  1251600.0 1428000.0 1261800.0 1414200.0 ;
      RECT  1251600.0 1428000.0 1261800.0 1441800.0 ;
      RECT  1251600.0 1455600.0 1261800.0 1441800.0 ;
      RECT  1251600.0 1455600.0 1261800.0 1469400.0 ;
      RECT  1251600.0 1483200.0 1261800.0 1469400.0 ;
      RECT  1251600.0 1483200.0 1261800.0 1497000.0 ;
      RECT  1251600.0 1510800.0 1261800.0 1497000.0 ;
      RECT  1251600.0 1510800.0 1261800.0 1524600.0 ;
      RECT  1251600.0 1538400.0 1261800.0 1524600.0 ;
      RECT  1251600.0 1538400.0 1261800.0 1552200.0 ;
      RECT  1251600.0 1566000.0 1261800.0 1552200.0 ;
      RECT  1251600.0 1566000.0 1261800.0 1579800.0 ;
      RECT  1251600.0 1593600.0 1261800.0 1579800.0 ;
      RECT  1251600.0 1593600.0 1261800.0 1607400.0 ;
      RECT  1251600.0 1621200.0 1261800.0 1607400.0 ;
      RECT  1251600.0 1621200.0 1261800.0 1635000.0 ;
      RECT  1251600.0 1648800.0 1261800.0 1635000.0 ;
      RECT  1251600.0 1648800.0 1261800.0 1662600.0 ;
      RECT  1251600.0 1676400.0 1261800.0 1662600.0 ;
      RECT  1251600.0 1676400.0 1261800.0 1690200.0 ;
      RECT  1251600.0 1704000.0 1261800.0 1690200.0 ;
      RECT  1251600.0 1704000.0 1261800.0 1717800.0 ;
      RECT  1251600.0 1731600.0 1261800.0 1717800.0 ;
      RECT  1251600.0 1731600.0 1261800.0 1745400.0 ;
      RECT  1251600.0 1759200.0 1261800.0 1745400.0 ;
      RECT  1251600.0 1759200.0 1261800.0 1773000.0 ;
      RECT  1251600.0 1786800.0 1261800.0 1773000.0 ;
      RECT  1251600.0 1786800.0 1261800.0 1800600.0 ;
      RECT  1251600.0 1814400.0 1261800.0 1800600.0 ;
      RECT  1251600.0 1814400.0 1261800.0 1828200.0 ;
      RECT  1251600.0 1842000.0 1261800.0 1828200.0 ;
      RECT  1251600.0 1842000.0 1261800.0 1855800.0 ;
      RECT  1251600.0 1869600.0 1261800.0 1855800.0 ;
      RECT  1251600.0 1869600.0 1261800.0 1883400.0 ;
      RECT  1251600.0 1897200.0 1261800.0 1883400.0 ;
      RECT  1251600.0 1897200.0 1261800.0 1911000.0 ;
      RECT  1251600.0 1924800.0 1261800.0 1911000.0 ;
      RECT  1251600.0 1924800.0 1261800.0 1938600.0 ;
      RECT  1251600.0 1952400.0 1261800.0 1938600.0 ;
      RECT  1251600.0 1952400.0 1261800.0 1966200.0 ;
      RECT  1251600.0 1980000.0 1261800.0 1966200.0 ;
      RECT  1251600.0 1980000.0 1261800.0 1993800.0 ;
      RECT  1251600.0 2007600.0 1261800.0 1993800.0 ;
      RECT  1251600.0 2007600.0 1261800.0 2021400.0 ;
      RECT  1251600.0 2035200.0 1261800.0 2021400.0 ;
      RECT  1251600.0 2035200.0 1261800.0 2049000.0 ;
      RECT  1251600.0 2062800.0 1261800.0 2049000.0 ;
      RECT  1251600.0 2062800.0 1261800.0 2076600.0 ;
      RECT  1251600.0 2090400.0 1261800.0 2076600.0 ;
      RECT  1251600.0 2090400.0 1261800.0 2104200.0 ;
      RECT  1251600.0 2118000.0 1261800.0 2104200.0 ;
      RECT  1251600.0 2118000.0 1261800.0 2131800.0 ;
      RECT  1251600.0 2145600.0 1261800.0 2131800.0 ;
      RECT  1261800.0 379200.0 1272000.0 393000.0 ;
      RECT  1261800.0 406800.0 1272000.0 393000.0 ;
      RECT  1261800.0 406800.0 1272000.0 420600.0 ;
      RECT  1261800.0 434400.0 1272000.0 420600.0 ;
      RECT  1261800.0 434400.0 1272000.0 448200.0 ;
      RECT  1261800.0 462000.0 1272000.0 448200.0 ;
      RECT  1261800.0 462000.0 1272000.0 475800.0 ;
      RECT  1261800.0 489600.0 1272000.0 475800.0 ;
      RECT  1261800.0 489600.0 1272000.0 503400.0 ;
      RECT  1261800.0 517200.0 1272000.0 503400.0 ;
      RECT  1261800.0 517200.0 1272000.0 531000.0 ;
      RECT  1261800.0 544800.0 1272000.0 531000.0 ;
      RECT  1261800.0 544800.0 1272000.0 558600.0 ;
      RECT  1261800.0 572400.0 1272000.0 558600.0 ;
      RECT  1261800.0 572400.0 1272000.0 586200.0 ;
      RECT  1261800.0 600000.0 1272000.0 586200.0 ;
      RECT  1261800.0 600000.0 1272000.0 613800.0 ;
      RECT  1261800.0 627600.0 1272000.0 613800.0 ;
      RECT  1261800.0 627600.0 1272000.0 641400.0 ;
      RECT  1261800.0 655200.0 1272000.0 641400.0 ;
      RECT  1261800.0 655200.0 1272000.0 669000.0 ;
      RECT  1261800.0 682800.0 1272000.0 669000.0 ;
      RECT  1261800.0 682800.0 1272000.0 696600.0 ;
      RECT  1261800.0 710400.0 1272000.0 696600.0 ;
      RECT  1261800.0 710400.0 1272000.0 724200.0 ;
      RECT  1261800.0 738000.0 1272000.0 724200.0 ;
      RECT  1261800.0 738000.0 1272000.0 751800.0 ;
      RECT  1261800.0 765600.0 1272000.0 751800.0 ;
      RECT  1261800.0 765600.0 1272000.0 779400.0 ;
      RECT  1261800.0 793200.0 1272000.0 779400.0 ;
      RECT  1261800.0 793200.0 1272000.0 807000.0 ;
      RECT  1261800.0 820800.0 1272000.0 807000.0 ;
      RECT  1261800.0 820800.0 1272000.0 834600.0 ;
      RECT  1261800.0 848400.0 1272000.0 834600.0 ;
      RECT  1261800.0 848400.0 1272000.0 862200.0 ;
      RECT  1261800.0 876000.0 1272000.0 862200.0 ;
      RECT  1261800.0 876000.0 1272000.0 889800.0 ;
      RECT  1261800.0 903600.0 1272000.0 889800.0 ;
      RECT  1261800.0 903600.0 1272000.0 917400.0 ;
      RECT  1261800.0 931200.0 1272000.0 917400.0 ;
      RECT  1261800.0 931200.0 1272000.0 945000.0 ;
      RECT  1261800.0 958800.0 1272000.0 945000.0 ;
      RECT  1261800.0 958800.0 1272000.0 972600.0 ;
      RECT  1261800.0 986400.0 1272000.0 972600.0 ;
      RECT  1261800.0 986400.0 1272000.0 1000200.0 ;
      RECT  1261800.0 1014000.0 1272000.0 1000200.0 ;
      RECT  1261800.0 1014000.0 1272000.0 1027800.0 ;
      RECT  1261800.0 1041600.0 1272000.0 1027800.0 ;
      RECT  1261800.0 1041600.0 1272000.0 1055400.0 ;
      RECT  1261800.0 1069200.0 1272000.0 1055400.0 ;
      RECT  1261800.0 1069200.0 1272000.0 1083000.0 ;
      RECT  1261800.0 1096800.0 1272000.0 1083000.0 ;
      RECT  1261800.0 1096800.0 1272000.0 1110600.0 ;
      RECT  1261800.0 1124400.0 1272000.0 1110600.0 ;
      RECT  1261800.0 1124400.0 1272000.0 1138200.0 ;
      RECT  1261800.0 1152000.0 1272000.0 1138200.0 ;
      RECT  1261800.0 1152000.0 1272000.0 1165800.0 ;
      RECT  1261800.0 1179600.0 1272000.0 1165800.0 ;
      RECT  1261800.0 1179600.0 1272000.0 1193400.0 ;
      RECT  1261800.0 1207200.0 1272000.0 1193400.0 ;
      RECT  1261800.0 1207200.0 1272000.0 1221000.0 ;
      RECT  1261800.0 1234800.0 1272000.0 1221000.0 ;
      RECT  1261800.0 1234800.0 1272000.0 1248600.0 ;
      RECT  1261800.0 1262400.0 1272000.0 1248600.0 ;
      RECT  1261800.0 1262400.0 1272000.0 1276200.0 ;
      RECT  1261800.0 1290000.0 1272000.0 1276200.0 ;
      RECT  1261800.0 1290000.0 1272000.0 1303800.0 ;
      RECT  1261800.0 1317600.0 1272000.0 1303800.0 ;
      RECT  1261800.0 1317600.0 1272000.0 1331400.0 ;
      RECT  1261800.0 1345200.0 1272000.0 1331400.0 ;
      RECT  1261800.0 1345200.0 1272000.0 1359000.0 ;
      RECT  1261800.0 1372800.0 1272000.0 1359000.0 ;
      RECT  1261800.0 1372800.0 1272000.0 1386600.0 ;
      RECT  1261800.0 1400400.0 1272000.0 1386600.0 ;
      RECT  1261800.0 1400400.0 1272000.0 1414200.0 ;
      RECT  1261800.0 1428000.0 1272000.0 1414200.0 ;
      RECT  1261800.0 1428000.0 1272000.0 1441800.0 ;
      RECT  1261800.0 1455600.0 1272000.0 1441800.0 ;
      RECT  1261800.0 1455600.0 1272000.0 1469400.0 ;
      RECT  1261800.0 1483200.0 1272000.0 1469400.0 ;
      RECT  1261800.0 1483200.0 1272000.0 1497000.0 ;
      RECT  1261800.0 1510800.0 1272000.0 1497000.0 ;
      RECT  1261800.0 1510800.0 1272000.0 1524600.0 ;
      RECT  1261800.0 1538400.0 1272000.0 1524600.0 ;
      RECT  1261800.0 1538400.0 1272000.0 1552200.0 ;
      RECT  1261800.0 1566000.0 1272000.0 1552200.0 ;
      RECT  1261800.0 1566000.0 1272000.0 1579800.0 ;
      RECT  1261800.0 1593600.0 1272000.0 1579800.0 ;
      RECT  1261800.0 1593600.0 1272000.0 1607400.0 ;
      RECT  1261800.0 1621200.0 1272000.0 1607400.0 ;
      RECT  1261800.0 1621200.0 1272000.0 1635000.0 ;
      RECT  1261800.0 1648800.0 1272000.0 1635000.0 ;
      RECT  1261800.0 1648800.0 1272000.0 1662600.0 ;
      RECT  1261800.0 1676400.0 1272000.0 1662600.0 ;
      RECT  1261800.0 1676400.0 1272000.0 1690200.0 ;
      RECT  1261800.0 1704000.0 1272000.0 1690200.0 ;
      RECT  1261800.0 1704000.0 1272000.0 1717800.0 ;
      RECT  1261800.0 1731600.0 1272000.0 1717800.0 ;
      RECT  1261800.0 1731600.0 1272000.0 1745400.0 ;
      RECT  1261800.0 1759200.0 1272000.0 1745400.0 ;
      RECT  1261800.0 1759200.0 1272000.0 1773000.0 ;
      RECT  1261800.0 1786800.0 1272000.0 1773000.0 ;
      RECT  1261800.0 1786800.0 1272000.0 1800600.0 ;
      RECT  1261800.0 1814400.0 1272000.0 1800600.0 ;
      RECT  1261800.0 1814400.0 1272000.0 1828200.0 ;
      RECT  1261800.0 1842000.0 1272000.0 1828200.0 ;
      RECT  1261800.0 1842000.0 1272000.0 1855800.0 ;
      RECT  1261800.0 1869600.0 1272000.0 1855800.0 ;
      RECT  1261800.0 1869600.0 1272000.0 1883400.0 ;
      RECT  1261800.0 1897200.0 1272000.0 1883400.0 ;
      RECT  1261800.0 1897200.0 1272000.0 1911000.0 ;
      RECT  1261800.0 1924800.0 1272000.0 1911000.0 ;
      RECT  1261800.0 1924800.0 1272000.0 1938600.0 ;
      RECT  1261800.0 1952400.0 1272000.0 1938600.0 ;
      RECT  1261800.0 1952400.0 1272000.0 1966200.0 ;
      RECT  1261800.0 1980000.0 1272000.0 1966200.0 ;
      RECT  1261800.0 1980000.0 1272000.0 1993800.0 ;
      RECT  1261800.0 2007600.0 1272000.0 1993800.0 ;
      RECT  1261800.0 2007600.0 1272000.0 2021400.0 ;
      RECT  1261800.0 2035200.0 1272000.0 2021400.0 ;
      RECT  1261800.0 2035200.0 1272000.0 2049000.0 ;
      RECT  1261800.0 2062800.0 1272000.0 2049000.0 ;
      RECT  1261800.0 2062800.0 1272000.0 2076600.0 ;
      RECT  1261800.0 2090400.0 1272000.0 2076600.0 ;
      RECT  1261800.0 2090400.0 1272000.0 2104200.0 ;
      RECT  1261800.0 2118000.0 1272000.0 2104200.0 ;
      RECT  1261800.0 2118000.0 1272000.0 2131800.0 ;
      RECT  1261800.0 2145600.0 1272000.0 2131800.0 ;
      RECT  1272000.0 379200.0 1282200.0 393000.0 ;
      RECT  1272000.0 406800.0 1282200.0 393000.0 ;
      RECT  1272000.0 406800.0 1282200.0 420600.0 ;
      RECT  1272000.0 434400.0 1282200.0 420600.0 ;
      RECT  1272000.0 434400.0 1282200.0 448200.0 ;
      RECT  1272000.0 462000.0 1282200.0 448200.0 ;
      RECT  1272000.0 462000.0 1282200.0 475800.0 ;
      RECT  1272000.0 489600.0 1282200.0 475800.0 ;
      RECT  1272000.0 489600.0 1282200.0 503400.0 ;
      RECT  1272000.0 517200.0 1282200.0 503400.0 ;
      RECT  1272000.0 517200.0 1282200.0 531000.0 ;
      RECT  1272000.0 544800.0 1282200.0 531000.0 ;
      RECT  1272000.0 544800.0 1282200.0 558600.0 ;
      RECT  1272000.0 572400.0 1282200.0 558600.0 ;
      RECT  1272000.0 572400.0 1282200.0 586200.0 ;
      RECT  1272000.0 600000.0 1282200.0 586200.0 ;
      RECT  1272000.0 600000.0 1282200.0 613800.0 ;
      RECT  1272000.0 627600.0 1282200.0 613800.0 ;
      RECT  1272000.0 627600.0 1282200.0 641400.0 ;
      RECT  1272000.0 655200.0 1282200.0 641400.0 ;
      RECT  1272000.0 655200.0 1282200.0 669000.0 ;
      RECT  1272000.0 682800.0 1282200.0 669000.0 ;
      RECT  1272000.0 682800.0 1282200.0 696600.0 ;
      RECT  1272000.0 710400.0 1282200.0 696600.0 ;
      RECT  1272000.0 710400.0 1282200.0 724200.0 ;
      RECT  1272000.0 738000.0 1282200.0 724200.0 ;
      RECT  1272000.0 738000.0 1282200.0 751800.0 ;
      RECT  1272000.0 765600.0 1282200.0 751800.0 ;
      RECT  1272000.0 765600.0 1282200.0 779400.0 ;
      RECT  1272000.0 793200.0 1282200.0 779400.0 ;
      RECT  1272000.0 793200.0 1282200.0 807000.0 ;
      RECT  1272000.0 820800.0 1282200.0 807000.0 ;
      RECT  1272000.0 820800.0 1282200.0 834600.0 ;
      RECT  1272000.0 848400.0 1282200.0 834600.0 ;
      RECT  1272000.0 848400.0 1282200.0 862200.0 ;
      RECT  1272000.0 876000.0 1282200.0 862200.0 ;
      RECT  1272000.0 876000.0 1282200.0 889800.0 ;
      RECT  1272000.0 903600.0 1282200.0 889800.0 ;
      RECT  1272000.0 903600.0 1282200.0 917400.0 ;
      RECT  1272000.0 931200.0 1282200.0 917400.0 ;
      RECT  1272000.0 931200.0 1282200.0 945000.0 ;
      RECT  1272000.0 958800.0 1282200.0 945000.0 ;
      RECT  1272000.0 958800.0 1282200.0 972600.0 ;
      RECT  1272000.0 986400.0 1282200.0 972600.0 ;
      RECT  1272000.0 986400.0 1282200.0 1000200.0 ;
      RECT  1272000.0 1014000.0 1282200.0 1000200.0 ;
      RECT  1272000.0 1014000.0 1282200.0 1027800.0 ;
      RECT  1272000.0 1041600.0 1282200.0 1027800.0 ;
      RECT  1272000.0 1041600.0 1282200.0 1055400.0 ;
      RECT  1272000.0 1069200.0 1282200.0 1055400.0 ;
      RECT  1272000.0 1069200.0 1282200.0 1083000.0 ;
      RECT  1272000.0 1096800.0 1282200.0 1083000.0 ;
      RECT  1272000.0 1096800.0 1282200.0 1110600.0 ;
      RECT  1272000.0 1124400.0 1282200.0 1110600.0 ;
      RECT  1272000.0 1124400.0 1282200.0 1138200.0 ;
      RECT  1272000.0 1152000.0 1282200.0 1138200.0 ;
      RECT  1272000.0 1152000.0 1282200.0 1165800.0 ;
      RECT  1272000.0 1179600.0 1282200.0 1165800.0 ;
      RECT  1272000.0 1179600.0 1282200.0 1193400.0 ;
      RECT  1272000.0 1207200.0 1282200.0 1193400.0 ;
      RECT  1272000.0 1207200.0 1282200.0 1221000.0 ;
      RECT  1272000.0 1234800.0 1282200.0 1221000.0 ;
      RECT  1272000.0 1234800.0 1282200.0 1248600.0 ;
      RECT  1272000.0 1262400.0 1282200.0 1248600.0 ;
      RECT  1272000.0 1262400.0 1282200.0 1276200.0 ;
      RECT  1272000.0 1290000.0 1282200.0 1276200.0 ;
      RECT  1272000.0 1290000.0 1282200.0 1303800.0 ;
      RECT  1272000.0 1317600.0 1282200.0 1303800.0 ;
      RECT  1272000.0 1317600.0 1282200.0 1331400.0 ;
      RECT  1272000.0 1345200.0 1282200.0 1331400.0 ;
      RECT  1272000.0 1345200.0 1282200.0 1359000.0 ;
      RECT  1272000.0 1372800.0 1282200.0 1359000.0 ;
      RECT  1272000.0 1372800.0 1282200.0 1386600.0 ;
      RECT  1272000.0 1400400.0 1282200.0 1386600.0 ;
      RECT  1272000.0 1400400.0 1282200.0 1414200.0 ;
      RECT  1272000.0 1428000.0 1282200.0 1414200.0 ;
      RECT  1272000.0 1428000.0 1282200.0 1441800.0 ;
      RECT  1272000.0 1455600.0 1282200.0 1441800.0 ;
      RECT  1272000.0 1455600.0 1282200.0 1469400.0 ;
      RECT  1272000.0 1483200.0 1282200.0 1469400.0 ;
      RECT  1272000.0 1483200.0 1282200.0 1497000.0 ;
      RECT  1272000.0 1510800.0 1282200.0 1497000.0 ;
      RECT  1272000.0 1510800.0 1282200.0 1524600.0 ;
      RECT  1272000.0 1538400.0 1282200.0 1524600.0 ;
      RECT  1272000.0 1538400.0 1282200.0 1552200.0 ;
      RECT  1272000.0 1566000.0 1282200.0 1552200.0 ;
      RECT  1272000.0 1566000.0 1282200.0 1579800.0 ;
      RECT  1272000.0 1593600.0 1282200.0 1579800.0 ;
      RECT  1272000.0 1593600.0 1282200.0 1607400.0 ;
      RECT  1272000.0 1621200.0 1282200.0 1607400.0 ;
      RECT  1272000.0 1621200.0 1282200.0 1635000.0 ;
      RECT  1272000.0 1648800.0 1282200.0 1635000.0 ;
      RECT  1272000.0 1648800.0 1282200.0 1662600.0 ;
      RECT  1272000.0 1676400.0 1282200.0 1662600.0 ;
      RECT  1272000.0 1676400.0 1282200.0 1690200.0 ;
      RECT  1272000.0 1704000.0 1282200.0 1690200.0 ;
      RECT  1272000.0 1704000.0 1282200.0 1717800.0 ;
      RECT  1272000.0 1731600.0 1282200.0 1717800.0 ;
      RECT  1272000.0 1731600.0 1282200.0 1745400.0 ;
      RECT  1272000.0 1759200.0 1282200.0 1745400.0 ;
      RECT  1272000.0 1759200.0 1282200.0 1773000.0 ;
      RECT  1272000.0 1786800.0 1282200.0 1773000.0 ;
      RECT  1272000.0 1786800.0 1282200.0 1800600.0 ;
      RECT  1272000.0 1814400.0 1282200.0 1800600.0 ;
      RECT  1272000.0 1814400.0 1282200.0 1828200.0 ;
      RECT  1272000.0 1842000.0 1282200.0 1828200.0 ;
      RECT  1272000.0 1842000.0 1282200.0 1855800.0 ;
      RECT  1272000.0 1869600.0 1282200.0 1855800.0 ;
      RECT  1272000.0 1869600.0 1282200.0 1883400.0 ;
      RECT  1272000.0 1897200.0 1282200.0 1883400.0 ;
      RECT  1272000.0 1897200.0 1282200.0 1911000.0 ;
      RECT  1272000.0 1924800.0 1282200.0 1911000.0 ;
      RECT  1272000.0 1924800.0 1282200.0 1938600.0 ;
      RECT  1272000.0 1952400.0 1282200.0 1938600.0 ;
      RECT  1272000.0 1952400.0 1282200.0 1966200.0 ;
      RECT  1272000.0 1980000.0 1282200.0 1966200.0 ;
      RECT  1272000.0 1980000.0 1282200.0 1993800.0 ;
      RECT  1272000.0 2007600.0 1282200.0 1993800.0 ;
      RECT  1272000.0 2007600.0 1282200.0 2021400.0 ;
      RECT  1272000.0 2035200.0 1282200.0 2021400.0 ;
      RECT  1272000.0 2035200.0 1282200.0 2049000.0 ;
      RECT  1272000.0 2062800.0 1282200.0 2049000.0 ;
      RECT  1272000.0 2062800.0 1282200.0 2076600.0 ;
      RECT  1272000.0 2090400.0 1282200.0 2076600.0 ;
      RECT  1272000.0 2090400.0 1282200.0 2104200.0 ;
      RECT  1272000.0 2118000.0 1282200.0 2104200.0 ;
      RECT  1272000.0 2118000.0 1282200.0 2131800.0 ;
      RECT  1272000.0 2145600.0 1282200.0 2131800.0 ;
      RECT  1282200.0 379200.0 1292400.0 393000.0 ;
      RECT  1282200.0 406800.0 1292400.0 393000.0 ;
      RECT  1282200.0 406800.0 1292400.0 420600.0 ;
      RECT  1282200.0 434400.0 1292400.0 420600.0 ;
      RECT  1282200.0 434400.0 1292400.0 448200.0 ;
      RECT  1282200.0 462000.0 1292400.0 448200.0 ;
      RECT  1282200.0 462000.0 1292400.0 475800.0 ;
      RECT  1282200.0 489600.0 1292400.0 475800.0 ;
      RECT  1282200.0 489600.0 1292400.0 503400.0 ;
      RECT  1282200.0 517200.0 1292400.0 503400.0 ;
      RECT  1282200.0 517200.0 1292400.0 531000.0 ;
      RECT  1282200.0 544800.0 1292400.0 531000.0 ;
      RECT  1282200.0 544800.0 1292400.0 558600.0 ;
      RECT  1282200.0 572400.0 1292400.0 558600.0 ;
      RECT  1282200.0 572400.0 1292400.0 586200.0 ;
      RECT  1282200.0 600000.0 1292400.0 586200.0 ;
      RECT  1282200.0 600000.0 1292400.0 613800.0 ;
      RECT  1282200.0 627600.0 1292400.0 613800.0 ;
      RECT  1282200.0 627600.0 1292400.0 641400.0 ;
      RECT  1282200.0 655200.0 1292400.0 641400.0 ;
      RECT  1282200.0 655200.0 1292400.0 669000.0 ;
      RECT  1282200.0 682800.0 1292400.0 669000.0 ;
      RECT  1282200.0 682800.0 1292400.0 696600.0 ;
      RECT  1282200.0 710400.0 1292400.0 696600.0 ;
      RECT  1282200.0 710400.0 1292400.0 724200.0 ;
      RECT  1282200.0 738000.0 1292400.0 724200.0 ;
      RECT  1282200.0 738000.0 1292400.0 751800.0 ;
      RECT  1282200.0 765600.0 1292400.0 751800.0 ;
      RECT  1282200.0 765600.0 1292400.0 779400.0 ;
      RECT  1282200.0 793200.0 1292400.0 779400.0 ;
      RECT  1282200.0 793200.0 1292400.0 807000.0 ;
      RECT  1282200.0 820800.0 1292400.0 807000.0 ;
      RECT  1282200.0 820800.0 1292400.0 834600.0 ;
      RECT  1282200.0 848400.0 1292400.0 834600.0 ;
      RECT  1282200.0 848400.0 1292400.0 862200.0 ;
      RECT  1282200.0 876000.0 1292400.0 862200.0 ;
      RECT  1282200.0 876000.0 1292400.0 889800.0 ;
      RECT  1282200.0 903600.0 1292400.0 889800.0 ;
      RECT  1282200.0 903600.0 1292400.0 917400.0 ;
      RECT  1282200.0 931200.0 1292400.0 917400.0 ;
      RECT  1282200.0 931200.0 1292400.0 945000.0 ;
      RECT  1282200.0 958800.0 1292400.0 945000.0 ;
      RECT  1282200.0 958800.0 1292400.0 972600.0 ;
      RECT  1282200.0 986400.0 1292400.0 972600.0 ;
      RECT  1282200.0 986400.0 1292400.0 1000200.0 ;
      RECT  1282200.0 1014000.0 1292400.0 1000200.0 ;
      RECT  1282200.0 1014000.0 1292400.0 1027800.0 ;
      RECT  1282200.0 1041600.0 1292400.0 1027800.0 ;
      RECT  1282200.0 1041600.0 1292400.0 1055400.0 ;
      RECT  1282200.0 1069200.0 1292400.0 1055400.0 ;
      RECT  1282200.0 1069200.0 1292400.0 1083000.0 ;
      RECT  1282200.0 1096800.0 1292400.0 1083000.0 ;
      RECT  1282200.0 1096800.0 1292400.0 1110600.0 ;
      RECT  1282200.0 1124400.0 1292400.0 1110600.0 ;
      RECT  1282200.0 1124400.0 1292400.0 1138200.0 ;
      RECT  1282200.0 1152000.0 1292400.0 1138200.0 ;
      RECT  1282200.0 1152000.0 1292400.0 1165800.0 ;
      RECT  1282200.0 1179600.0 1292400.0 1165800.0 ;
      RECT  1282200.0 1179600.0 1292400.0 1193400.0 ;
      RECT  1282200.0 1207200.0 1292400.0 1193400.0 ;
      RECT  1282200.0 1207200.0 1292400.0 1221000.0 ;
      RECT  1282200.0 1234800.0 1292400.0 1221000.0 ;
      RECT  1282200.0 1234800.0 1292400.0 1248600.0 ;
      RECT  1282200.0 1262400.0 1292400.0 1248600.0 ;
      RECT  1282200.0 1262400.0 1292400.0 1276200.0 ;
      RECT  1282200.0 1290000.0 1292400.0 1276200.0 ;
      RECT  1282200.0 1290000.0 1292400.0 1303800.0 ;
      RECT  1282200.0 1317600.0 1292400.0 1303800.0 ;
      RECT  1282200.0 1317600.0 1292400.0 1331400.0 ;
      RECT  1282200.0 1345200.0 1292400.0 1331400.0 ;
      RECT  1282200.0 1345200.0 1292400.0 1359000.0 ;
      RECT  1282200.0 1372800.0 1292400.0 1359000.0 ;
      RECT  1282200.0 1372800.0 1292400.0 1386600.0 ;
      RECT  1282200.0 1400400.0 1292400.0 1386600.0 ;
      RECT  1282200.0 1400400.0 1292400.0 1414200.0 ;
      RECT  1282200.0 1428000.0 1292400.0 1414200.0 ;
      RECT  1282200.0 1428000.0 1292400.0 1441800.0 ;
      RECT  1282200.0 1455600.0 1292400.0 1441800.0 ;
      RECT  1282200.0 1455600.0 1292400.0 1469400.0 ;
      RECT  1282200.0 1483200.0 1292400.0 1469400.0 ;
      RECT  1282200.0 1483200.0 1292400.0 1497000.0 ;
      RECT  1282200.0 1510800.0 1292400.0 1497000.0 ;
      RECT  1282200.0 1510800.0 1292400.0 1524600.0 ;
      RECT  1282200.0 1538400.0 1292400.0 1524600.0 ;
      RECT  1282200.0 1538400.0 1292400.0 1552200.0 ;
      RECT  1282200.0 1566000.0 1292400.0 1552200.0 ;
      RECT  1282200.0 1566000.0 1292400.0 1579800.0 ;
      RECT  1282200.0 1593600.0 1292400.0 1579800.0 ;
      RECT  1282200.0 1593600.0 1292400.0 1607400.0 ;
      RECT  1282200.0 1621200.0 1292400.0 1607400.0 ;
      RECT  1282200.0 1621200.0 1292400.0 1635000.0 ;
      RECT  1282200.0 1648800.0 1292400.0 1635000.0 ;
      RECT  1282200.0 1648800.0 1292400.0 1662600.0 ;
      RECT  1282200.0 1676400.0 1292400.0 1662600.0 ;
      RECT  1282200.0 1676400.0 1292400.0 1690200.0 ;
      RECT  1282200.0 1704000.0 1292400.0 1690200.0 ;
      RECT  1282200.0 1704000.0 1292400.0 1717800.0 ;
      RECT  1282200.0 1731600.0 1292400.0 1717800.0 ;
      RECT  1282200.0 1731600.0 1292400.0 1745400.0 ;
      RECT  1282200.0 1759200.0 1292400.0 1745400.0 ;
      RECT  1282200.0 1759200.0 1292400.0 1773000.0 ;
      RECT  1282200.0 1786800.0 1292400.0 1773000.0 ;
      RECT  1282200.0 1786800.0 1292400.0 1800600.0 ;
      RECT  1282200.0 1814400.0 1292400.0 1800600.0 ;
      RECT  1282200.0 1814400.0 1292400.0 1828200.0 ;
      RECT  1282200.0 1842000.0 1292400.0 1828200.0 ;
      RECT  1282200.0 1842000.0 1292400.0 1855800.0 ;
      RECT  1282200.0 1869600.0 1292400.0 1855800.0 ;
      RECT  1282200.0 1869600.0 1292400.0 1883400.0 ;
      RECT  1282200.0 1897200.0 1292400.0 1883400.0 ;
      RECT  1282200.0 1897200.0 1292400.0 1911000.0 ;
      RECT  1282200.0 1924800.0 1292400.0 1911000.0 ;
      RECT  1282200.0 1924800.0 1292400.0 1938600.0 ;
      RECT  1282200.0 1952400.0 1292400.0 1938600.0 ;
      RECT  1282200.0 1952400.0 1292400.0 1966200.0 ;
      RECT  1282200.0 1980000.0 1292400.0 1966200.0 ;
      RECT  1282200.0 1980000.0 1292400.0 1993800.0 ;
      RECT  1282200.0 2007600.0 1292400.0 1993800.0 ;
      RECT  1282200.0 2007600.0 1292400.0 2021400.0 ;
      RECT  1282200.0 2035200.0 1292400.0 2021400.0 ;
      RECT  1282200.0 2035200.0 1292400.0 2049000.0 ;
      RECT  1282200.0 2062800.0 1292400.0 2049000.0 ;
      RECT  1282200.0 2062800.0 1292400.0 2076600.0 ;
      RECT  1282200.0 2090400.0 1292400.0 2076600.0 ;
      RECT  1282200.0 2090400.0 1292400.0 2104200.0 ;
      RECT  1282200.0 2118000.0 1292400.0 2104200.0 ;
      RECT  1282200.0 2118000.0 1292400.0 2131800.0 ;
      RECT  1282200.0 2145600.0 1292400.0 2131800.0 ;
      RECT  1292400.0 379200.0 1302600.0 393000.0 ;
      RECT  1292400.0 406800.0 1302600.0 393000.0 ;
      RECT  1292400.0 406800.0 1302600.0 420600.0 ;
      RECT  1292400.0 434400.0 1302600.0 420600.0 ;
      RECT  1292400.0 434400.0 1302600.0 448200.0 ;
      RECT  1292400.0 462000.0 1302600.0 448200.0 ;
      RECT  1292400.0 462000.0 1302600.0 475800.0 ;
      RECT  1292400.0 489600.0 1302600.0 475800.0 ;
      RECT  1292400.0 489600.0 1302600.0 503400.0 ;
      RECT  1292400.0 517200.0 1302600.0 503400.0 ;
      RECT  1292400.0 517200.0 1302600.0 531000.0 ;
      RECT  1292400.0 544800.0 1302600.0 531000.0 ;
      RECT  1292400.0 544800.0 1302600.0 558600.0 ;
      RECT  1292400.0 572400.0 1302600.0 558600.0 ;
      RECT  1292400.0 572400.0 1302600.0 586200.0 ;
      RECT  1292400.0 600000.0 1302600.0 586200.0 ;
      RECT  1292400.0 600000.0 1302600.0 613800.0 ;
      RECT  1292400.0 627600.0 1302600.0 613800.0 ;
      RECT  1292400.0 627600.0 1302600.0 641400.0 ;
      RECT  1292400.0 655200.0 1302600.0 641400.0 ;
      RECT  1292400.0 655200.0 1302600.0 669000.0 ;
      RECT  1292400.0 682800.0 1302600.0 669000.0 ;
      RECT  1292400.0 682800.0 1302600.0 696600.0 ;
      RECT  1292400.0 710400.0 1302600.0 696600.0 ;
      RECT  1292400.0 710400.0 1302600.0 724200.0 ;
      RECT  1292400.0 738000.0 1302600.0 724200.0 ;
      RECT  1292400.0 738000.0 1302600.0 751800.0 ;
      RECT  1292400.0 765600.0 1302600.0 751800.0 ;
      RECT  1292400.0 765600.0 1302600.0 779400.0 ;
      RECT  1292400.0 793200.0 1302600.0 779400.0 ;
      RECT  1292400.0 793200.0 1302600.0 807000.0 ;
      RECT  1292400.0 820800.0 1302600.0 807000.0 ;
      RECT  1292400.0 820800.0 1302600.0 834600.0 ;
      RECT  1292400.0 848400.0 1302600.0 834600.0 ;
      RECT  1292400.0 848400.0 1302600.0 862200.0 ;
      RECT  1292400.0 876000.0 1302600.0 862200.0 ;
      RECT  1292400.0 876000.0 1302600.0 889800.0 ;
      RECT  1292400.0 903600.0 1302600.0 889800.0 ;
      RECT  1292400.0 903600.0 1302600.0 917400.0 ;
      RECT  1292400.0 931200.0 1302600.0 917400.0 ;
      RECT  1292400.0 931200.0 1302600.0 945000.0 ;
      RECT  1292400.0 958800.0 1302600.0 945000.0 ;
      RECT  1292400.0 958800.0 1302600.0 972600.0 ;
      RECT  1292400.0 986400.0 1302600.0 972600.0 ;
      RECT  1292400.0 986400.0 1302600.0 1000200.0 ;
      RECT  1292400.0 1014000.0 1302600.0 1000200.0 ;
      RECT  1292400.0 1014000.0 1302600.0 1027800.0 ;
      RECT  1292400.0 1041600.0 1302600.0 1027800.0 ;
      RECT  1292400.0 1041600.0 1302600.0 1055400.0 ;
      RECT  1292400.0 1069200.0 1302600.0 1055400.0 ;
      RECT  1292400.0 1069200.0 1302600.0 1083000.0 ;
      RECT  1292400.0 1096800.0 1302600.0 1083000.0 ;
      RECT  1292400.0 1096800.0 1302600.0 1110600.0 ;
      RECT  1292400.0 1124400.0 1302600.0 1110600.0 ;
      RECT  1292400.0 1124400.0 1302600.0 1138200.0 ;
      RECT  1292400.0 1152000.0 1302600.0 1138200.0 ;
      RECT  1292400.0 1152000.0 1302600.0 1165800.0 ;
      RECT  1292400.0 1179600.0 1302600.0 1165800.0 ;
      RECT  1292400.0 1179600.0 1302600.0 1193400.0 ;
      RECT  1292400.0 1207200.0 1302600.0 1193400.0 ;
      RECT  1292400.0 1207200.0 1302600.0 1221000.0 ;
      RECT  1292400.0 1234800.0 1302600.0 1221000.0 ;
      RECT  1292400.0 1234800.0 1302600.0 1248600.0 ;
      RECT  1292400.0 1262400.0 1302600.0 1248600.0 ;
      RECT  1292400.0 1262400.0 1302600.0 1276200.0 ;
      RECT  1292400.0 1290000.0 1302600.0 1276200.0 ;
      RECT  1292400.0 1290000.0 1302600.0 1303800.0 ;
      RECT  1292400.0 1317600.0 1302600.0 1303800.0 ;
      RECT  1292400.0 1317600.0 1302600.0 1331400.0 ;
      RECT  1292400.0 1345200.0 1302600.0 1331400.0 ;
      RECT  1292400.0 1345200.0 1302600.0 1359000.0 ;
      RECT  1292400.0 1372800.0 1302600.0 1359000.0 ;
      RECT  1292400.0 1372800.0 1302600.0 1386600.0 ;
      RECT  1292400.0 1400400.0 1302600.0 1386600.0 ;
      RECT  1292400.0 1400400.0 1302600.0 1414200.0 ;
      RECT  1292400.0 1428000.0 1302600.0 1414200.0 ;
      RECT  1292400.0 1428000.0 1302600.0 1441800.0 ;
      RECT  1292400.0 1455600.0 1302600.0 1441800.0 ;
      RECT  1292400.0 1455600.0 1302600.0 1469400.0 ;
      RECT  1292400.0 1483200.0 1302600.0 1469400.0 ;
      RECT  1292400.0 1483200.0 1302600.0 1497000.0 ;
      RECT  1292400.0 1510800.0 1302600.0 1497000.0 ;
      RECT  1292400.0 1510800.0 1302600.0 1524600.0 ;
      RECT  1292400.0 1538400.0 1302600.0 1524600.0 ;
      RECT  1292400.0 1538400.0 1302600.0 1552200.0 ;
      RECT  1292400.0 1566000.0 1302600.0 1552200.0 ;
      RECT  1292400.0 1566000.0 1302600.0 1579800.0 ;
      RECT  1292400.0 1593600.0 1302600.0 1579800.0 ;
      RECT  1292400.0 1593600.0 1302600.0 1607400.0 ;
      RECT  1292400.0 1621200.0 1302600.0 1607400.0 ;
      RECT  1292400.0 1621200.0 1302600.0 1635000.0 ;
      RECT  1292400.0 1648800.0 1302600.0 1635000.0 ;
      RECT  1292400.0 1648800.0 1302600.0 1662600.0 ;
      RECT  1292400.0 1676400.0 1302600.0 1662600.0 ;
      RECT  1292400.0 1676400.0 1302600.0 1690200.0 ;
      RECT  1292400.0 1704000.0 1302600.0 1690200.0 ;
      RECT  1292400.0 1704000.0 1302600.0 1717800.0 ;
      RECT  1292400.0 1731600.0 1302600.0 1717800.0 ;
      RECT  1292400.0 1731600.0 1302600.0 1745400.0 ;
      RECT  1292400.0 1759200.0 1302600.0 1745400.0 ;
      RECT  1292400.0 1759200.0 1302600.0 1773000.0 ;
      RECT  1292400.0 1786800.0 1302600.0 1773000.0 ;
      RECT  1292400.0 1786800.0 1302600.0 1800600.0 ;
      RECT  1292400.0 1814400.0 1302600.0 1800600.0 ;
      RECT  1292400.0 1814400.0 1302600.0 1828200.0 ;
      RECT  1292400.0 1842000.0 1302600.0 1828200.0 ;
      RECT  1292400.0 1842000.0 1302600.0 1855800.0 ;
      RECT  1292400.0 1869600.0 1302600.0 1855800.0 ;
      RECT  1292400.0 1869600.0 1302600.0 1883400.0 ;
      RECT  1292400.0 1897200.0 1302600.0 1883400.0 ;
      RECT  1292400.0 1897200.0 1302600.0 1911000.0 ;
      RECT  1292400.0 1924800.0 1302600.0 1911000.0 ;
      RECT  1292400.0 1924800.0 1302600.0 1938600.0 ;
      RECT  1292400.0 1952400.0 1302600.0 1938600.0 ;
      RECT  1292400.0 1952400.0 1302600.0 1966200.0 ;
      RECT  1292400.0 1980000.0 1302600.0 1966200.0 ;
      RECT  1292400.0 1980000.0 1302600.0 1993800.0 ;
      RECT  1292400.0 2007600.0 1302600.0 1993800.0 ;
      RECT  1292400.0 2007600.0 1302600.0 2021400.0 ;
      RECT  1292400.0 2035200.0 1302600.0 2021400.0 ;
      RECT  1292400.0 2035200.0 1302600.0 2049000.0 ;
      RECT  1292400.0 2062800.0 1302600.0 2049000.0 ;
      RECT  1292400.0 2062800.0 1302600.0 2076600.0 ;
      RECT  1292400.0 2090400.0 1302600.0 2076600.0 ;
      RECT  1292400.0 2090400.0 1302600.0 2104200.0 ;
      RECT  1292400.0 2118000.0 1302600.0 2104200.0 ;
      RECT  1292400.0 2118000.0 1302600.0 2131800.0 ;
      RECT  1292400.0 2145600.0 1302600.0 2131800.0 ;
      RECT  1302600.0 379200.0 1312800.0 393000.0 ;
      RECT  1302600.0 406800.0 1312800.0 393000.0 ;
      RECT  1302600.0 406800.0 1312800.0 420600.0 ;
      RECT  1302600.0 434400.0 1312800.0 420600.0 ;
      RECT  1302600.0 434400.0 1312800.0 448200.0 ;
      RECT  1302600.0 462000.0 1312800.0 448200.0 ;
      RECT  1302600.0 462000.0 1312800.0 475800.0 ;
      RECT  1302600.0 489600.0 1312800.0 475800.0 ;
      RECT  1302600.0 489600.0 1312800.0 503400.0 ;
      RECT  1302600.0 517200.0 1312800.0 503400.0 ;
      RECT  1302600.0 517200.0 1312800.0 531000.0 ;
      RECT  1302600.0 544800.0 1312800.0 531000.0 ;
      RECT  1302600.0 544800.0 1312800.0 558600.0 ;
      RECT  1302600.0 572400.0 1312800.0 558600.0 ;
      RECT  1302600.0 572400.0 1312800.0 586200.0 ;
      RECT  1302600.0 600000.0 1312800.0 586200.0 ;
      RECT  1302600.0 600000.0 1312800.0 613800.0 ;
      RECT  1302600.0 627600.0 1312800.0 613800.0 ;
      RECT  1302600.0 627600.0 1312800.0 641400.0 ;
      RECT  1302600.0 655200.0 1312800.0 641400.0 ;
      RECT  1302600.0 655200.0 1312800.0 669000.0 ;
      RECT  1302600.0 682800.0 1312800.0 669000.0 ;
      RECT  1302600.0 682800.0 1312800.0 696600.0 ;
      RECT  1302600.0 710400.0 1312800.0 696600.0 ;
      RECT  1302600.0 710400.0 1312800.0 724200.0 ;
      RECT  1302600.0 738000.0 1312800.0 724200.0 ;
      RECT  1302600.0 738000.0 1312800.0 751800.0 ;
      RECT  1302600.0 765600.0 1312800.0 751800.0 ;
      RECT  1302600.0 765600.0 1312800.0 779400.0 ;
      RECT  1302600.0 793200.0 1312800.0 779400.0 ;
      RECT  1302600.0 793200.0 1312800.0 807000.0 ;
      RECT  1302600.0 820800.0 1312800.0 807000.0 ;
      RECT  1302600.0 820800.0 1312800.0 834600.0 ;
      RECT  1302600.0 848400.0 1312800.0 834600.0 ;
      RECT  1302600.0 848400.0 1312800.0 862200.0 ;
      RECT  1302600.0 876000.0 1312800.0 862200.0 ;
      RECT  1302600.0 876000.0 1312800.0 889800.0 ;
      RECT  1302600.0 903600.0 1312800.0 889800.0 ;
      RECT  1302600.0 903600.0 1312800.0 917400.0 ;
      RECT  1302600.0 931200.0 1312800.0 917400.0 ;
      RECT  1302600.0 931200.0 1312800.0 945000.0 ;
      RECT  1302600.0 958800.0 1312800.0 945000.0 ;
      RECT  1302600.0 958800.0 1312800.0 972600.0 ;
      RECT  1302600.0 986400.0 1312800.0 972600.0 ;
      RECT  1302600.0 986400.0 1312800.0 1000200.0 ;
      RECT  1302600.0 1014000.0 1312800.0 1000200.0 ;
      RECT  1302600.0 1014000.0 1312800.0 1027800.0 ;
      RECT  1302600.0 1041600.0 1312800.0 1027800.0 ;
      RECT  1302600.0 1041600.0 1312800.0 1055400.0 ;
      RECT  1302600.0 1069200.0 1312800.0 1055400.0 ;
      RECT  1302600.0 1069200.0 1312800.0 1083000.0 ;
      RECT  1302600.0 1096800.0 1312800.0 1083000.0 ;
      RECT  1302600.0 1096800.0 1312800.0 1110600.0 ;
      RECT  1302600.0 1124400.0 1312800.0 1110600.0 ;
      RECT  1302600.0 1124400.0 1312800.0 1138200.0 ;
      RECT  1302600.0 1152000.0 1312800.0 1138200.0 ;
      RECT  1302600.0 1152000.0 1312800.0 1165800.0 ;
      RECT  1302600.0 1179600.0 1312800.0 1165800.0 ;
      RECT  1302600.0 1179600.0 1312800.0 1193400.0 ;
      RECT  1302600.0 1207200.0 1312800.0 1193400.0 ;
      RECT  1302600.0 1207200.0 1312800.0 1221000.0 ;
      RECT  1302600.0 1234800.0 1312800.0 1221000.0 ;
      RECT  1302600.0 1234800.0 1312800.0 1248600.0 ;
      RECT  1302600.0 1262400.0 1312800.0 1248600.0 ;
      RECT  1302600.0 1262400.0 1312800.0 1276200.0 ;
      RECT  1302600.0 1290000.0 1312800.0 1276200.0 ;
      RECT  1302600.0 1290000.0 1312800.0 1303800.0 ;
      RECT  1302600.0 1317600.0 1312800.0 1303800.0 ;
      RECT  1302600.0 1317600.0 1312800.0 1331400.0 ;
      RECT  1302600.0 1345200.0 1312800.0 1331400.0 ;
      RECT  1302600.0 1345200.0 1312800.0 1359000.0 ;
      RECT  1302600.0 1372800.0 1312800.0 1359000.0 ;
      RECT  1302600.0 1372800.0 1312800.0 1386600.0 ;
      RECT  1302600.0 1400400.0 1312800.0 1386600.0 ;
      RECT  1302600.0 1400400.0 1312800.0 1414200.0 ;
      RECT  1302600.0 1428000.0 1312800.0 1414200.0 ;
      RECT  1302600.0 1428000.0 1312800.0 1441800.0 ;
      RECT  1302600.0 1455600.0 1312800.0 1441800.0 ;
      RECT  1302600.0 1455600.0 1312800.0 1469400.0 ;
      RECT  1302600.0 1483200.0 1312800.0 1469400.0 ;
      RECT  1302600.0 1483200.0 1312800.0 1497000.0 ;
      RECT  1302600.0 1510800.0 1312800.0 1497000.0 ;
      RECT  1302600.0 1510800.0 1312800.0 1524600.0 ;
      RECT  1302600.0 1538400.0 1312800.0 1524600.0 ;
      RECT  1302600.0 1538400.0 1312800.0 1552200.0 ;
      RECT  1302600.0 1566000.0 1312800.0 1552200.0 ;
      RECT  1302600.0 1566000.0 1312800.0 1579800.0 ;
      RECT  1302600.0 1593600.0 1312800.0 1579800.0 ;
      RECT  1302600.0 1593600.0 1312800.0 1607400.0 ;
      RECT  1302600.0 1621200.0 1312800.0 1607400.0 ;
      RECT  1302600.0 1621200.0 1312800.0 1635000.0 ;
      RECT  1302600.0 1648800.0 1312800.0 1635000.0 ;
      RECT  1302600.0 1648800.0 1312800.0 1662600.0 ;
      RECT  1302600.0 1676400.0 1312800.0 1662600.0 ;
      RECT  1302600.0 1676400.0 1312800.0 1690200.0 ;
      RECT  1302600.0 1704000.0 1312800.0 1690200.0 ;
      RECT  1302600.0 1704000.0 1312800.0 1717800.0 ;
      RECT  1302600.0 1731600.0 1312800.0 1717800.0 ;
      RECT  1302600.0 1731600.0 1312800.0 1745400.0 ;
      RECT  1302600.0 1759200.0 1312800.0 1745400.0 ;
      RECT  1302600.0 1759200.0 1312800.0 1773000.0 ;
      RECT  1302600.0 1786800.0 1312800.0 1773000.0 ;
      RECT  1302600.0 1786800.0 1312800.0 1800600.0 ;
      RECT  1302600.0 1814400.0 1312800.0 1800600.0 ;
      RECT  1302600.0 1814400.0 1312800.0 1828200.0 ;
      RECT  1302600.0 1842000.0 1312800.0 1828200.0 ;
      RECT  1302600.0 1842000.0 1312800.0 1855800.0 ;
      RECT  1302600.0 1869600.0 1312800.0 1855800.0 ;
      RECT  1302600.0 1869600.0 1312800.0 1883400.0 ;
      RECT  1302600.0 1897200.0 1312800.0 1883400.0 ;
      RECT  1302600.0 1897200.0 1312800.0 1911000.0 ;
      RECT  1302600.0 1924800.0 1312800.0 1911000.0 ;
      RECT  1302600.0 1924800.0 1312800.0 1938600.0 ;
      RECT  1302600.0 1952400.0 1312800.0 1938600.0 ;
      RECT  1302600.0 1952400.0 1312800.0 1966200.0 ;
      RECT  1302600.0 1980000.0 1312800.0 1966200.0 ;
      RECT  1302600.0 1980000.0 1312800.0 1993800.0 ;
      RECT  1302600.0 2007600.0 1312800.0 1993800.0 ;
      RECT  1302600.0 2007600.0 1312800.0 2021400.0 ;
      RECT  1302600.0 2035200.0 1312800.0 2021400.0 ;
      RECT  1302600.0 2035200.0 1312800.0 2049000.0 ;
      RECT  1302600.0 2062800.0 1312800.0 2049000.0 ;
      RECT  1302600.0 2062800.0 1312800.0 2076600.0 ;
      RECT  1302600.0 2090400.0 1312800.0 2076600.0 ;
      RECT  1302600.0 2090400.0 1312800.0 2104200.0 ;
      RECT  1302600.0 2118000.0 1312800.0 2104200.0 ;
      RECT  1302600.0 2118000.0 1312800.0 2131800.0 ;
      RECT  1302600.0 2145600.0 1312800.0 2131800.0 ;
      RECT  1312800.0 379200.0 1323000.0 393000.0 ;
      RECT  1312800.0 406800.0 1323000.0 393000.0 ;
      RECT  1312800.0 406800.0 1323000.0 420600.0 ;
      RECT  1312800.0 434400.0 1323000.0 420600.0 ;
      RECT  1312800.0 434400.0 1323000.0 448200.0 ;
      RECT  1312800.0 462000.0 1323000.0 448200.0 ;
      RECT  1312800.0 462000.0 1323000.0 475800.0 ;
      RECT  1312800.0 489600.0 1323000.0 475800.0 ;
      RECT  1312800.0 489600.0 1323000.0 503400.0 ;
      RECT  1312800.0 517200.0 1323000.0 503400.0 ;
      RECT  1312800.0 517200.0 1323000.0 531000.0 ;
      RECT  1312800.0 544800.0 1323000.0 531000.0 ;
      RECT  1312800.0 544800.0 1323000.0 558600.0 ;
      RECT  1312800.0 572400.0 1323000.0 558600.0 ;
      RECT  1312800.0 572400.0 1323000.0 586200.0 ;
      RECT  1312800.0 600000.0 1323000.0 586200.0 ;
      RECT  1312800.0 600000.0 1323000.0 613800.0 ;
      RECT  1312800.0 627600.0 1323000.0 613800.0 ;
      RECT  1312800.0 627600.0 1323000.0 641400.0 ;
      RECT  1312800.0 655200.0 1323000.0 641400.0 ;
      RECT  1312800.0 655200.0 1323000.0 669000.0 ;
      RECT  1312800.0 682800.0 1323000.0 669000.0 ;
      RECT  1312800.0 682800.0 1323000.0 696600.0 ;
      RECT  1312800.0 710400.0 1323000.0 696600.0 ;
      RECT  1312800.0 710400.0 1323000.0 724200.0 ;
      RECT  1312800.0 738000.0 1323000.0 724200.0 ;
      RECT  1312800.0 738000.0 1323000.0 751800.0 ;
      RECT  1312800.0 765600.0 1323000.0 751800.0 ;
      RECT  1312800.0 765600.0 1323000.0 779400.0 ;
      RECT  1312800.0 793200.0 1323000.0 779400.0 ;
      RECT  1312800.0 793200.0 1323000.0 807000.0 ;
      RECT  1312800.0 820800.0 1323000.0 807000.0 ;
      RECT  1312800.0 820800.0 1323000.0 834600.0 ;
      RECT  1312800.0 848400.0 1323000.0 834600.0 ;
      RECT  1312800.0 848400.0 1323000.0 862200.0 ;
      RECT  1312800.0 876000.0 1323000.0 862200.0 ;
      RECT  1312800.0 876000.0 1323000.0 889800.0 ;
      RECT  1312800.0 903600.0 1323000.0 889800.0 ;
      RECT  1312800.0 903600.0 1323000.0 917400.0 ;
      RECT  1312800.0 931200.0 1323000.0 917400.0 ;
      RECT  1312800.0 931200.0 1323000.0 945000.0 ;
      RECT  1312800.0 958800.0 1323000.0 945000.0 ;
      RECT  1312800.0 958800.0 1323000.0 972600.0 ;
      RECT  1312800.0 986400.0 1323000.0 972600.0 ;
      RECT  1312800.0 986400.0 1323000.0 1000200.0 ;
      RECT  1312800.0 1014000.0 1323000.0 1000200.0 ;
      RECT  1312800.0 1014000.0 1323000.0 1027800.0 ;
      RECT  1312800.0 1041600.0 1323000.0 1027800.0 ;
      RECT  1312800.0 1041600.0 1323000.0 1055400.0 ;
      RECT  1312800.0 1069200.0 1323000.0 1055400.0 ;
      RECT  1312800.0 1069200.0 1323000.0 1083000.0 ;
      RECT  1312800.0 1096800.0 1323000.0 1083000.0 ;
      RECT  1312800.0 1096800.0 1323000.0 1110600.0 ;
      RECT  1312800.0 1124400.0 1323000.0 1110600.0 ;
      RECT  1312800.0 1124400.0 1323000.0 1138200.0 ;
      RECT  1312800.0 1152000.0 1323000.0 1138200.0 ;
      RECT  1312800.0 1152000.0 1323000.0 1165800.0 ;
      RECT  1312800.0 1179600.0 1323000.0 1165800.0 ;
      RECT  1312800.0 1179600.0 1323000.0 1193400.0 ;
      RECT  1312800.0 1207200.0 1323000.0 1193400.0 ;
      RECT  1312800.0 1207200.0 1323000.0 1221000.0 ;
      RECT  1312800.0 1234800.0 1323000.0 1221000.0 ;
      RECT  1312800.0 1234800.0 1323000.0 1248600.0 ;
      RECT  1312800.0 1262400.0 1323000.0 1248600.0 ;
      RECT  1312800.0 1262400.0 1323000.0 1276200.0 ;
      RECT  1312800.0 1290000.0 1323000.0 1276200.0 ;
      RECT  1312800.0 1290000.0 1323000.0 1303800.0 ;
      RECT  1312800.0 1317600.0 1323000.0 1303800.0 ;
      RECT  1312800.0 1317600.0 1323000.0 1331400.0 ;
      RECT  1312800.0 1345200.0 1323000.0 1331400.0 ;
      RECT  1312800.0 1345200.0 1323000.0 1359000.0 ;
      RECT  1312800.0 1372800.0 1323000.0 1359000.0 ;
      RECT  1312800.0 1372800.0 1323000.0 1386600.0 ;
      RECT  1312800.0 1400400.0 1323000.0 1386600.0 ;
      RECT  1312800.0 1400400.0 1323000.0 1414200.0 ;
      RECT  1312800.0 1428000.0 1323000.0 1414200.0 ;
      RECT  1312800.0 1428000.0 1323000.0 1441800.0 ;
      RECT  1312800.0 1455600.0 1323000.0 1441800.0 ;
      RECT  1312800.0 1455600.0 1323000.0 1469400.0 ;
      RECT  1312800.0 1483200.0 1323000.0 1469400.0 ;
      RECT  1312800.0 1483200.0 1323000.0 1497000.0 ;
      RECT  1312800.0 1510800.0 1323000.0 1497000.0 ;
      RECT  1312800.0 1510800.0 1323000.0 1524600.0 ;
      RECT  1312800.0 1538400.0 1323000.0 1524600.0 ;
      RECT  1312800.0 1538400.0 1323000.0 1552200.0 ;
      RECT  1312800.0 1566000.0 1323000.0 1552200.0 ;
      RECT  1312800.0 1566000.0 1323000.0 1579800.0 ;
      RECT  1312800.0 1593600.0 1323000.0 1579800.0 ;
      RECT  1312800.0 1593600.0 1323000.0 1607400.0 ;
      RECT  1312800.0 1621200.0 1323000.0 1607400.0 ;
      RECT  1312800.0 1621200.0 1323000.0 1635000.0 ;
      RECT  1312800.0 1648800.0 1323000.0 1635000.0 ;
      RECT  1312800.0 1648800.0 1323000.0 1662600.0 ;
      RECT  1312800.0 1676400.0 1323000.0 1662600.0 ;
      RECT  1312800.0 1676400.0 1323000.0 1690200.0 ;
      RECT  1312800.0 1704000.0 1323000.0 1690200.0 ;
      RECT  1312800.0 1704000.0 1323000.0 1717800.0 ;
      RECT  1312800.0 1731600.0 1323000.0 1717800.0 ;
      RECT  1312800.0 1731600.0 1323000.0 1745400.0 ;
      RECT  1312800.0 1759200.0 1323000.0 1745400.0 ;
      RECT  1312800.0 1759200.0 1323000.0 1773000.0 ;
      RECT  1312800.0 1786800.0 1323000.0 1773000.0 ;
      RECT  1312800.0 1786800.0 1323000.0 1800600.0 ;
      RECT  1312800.0 1814400.0 1323000.0 1800600.0 ;
      RECT  1312800.0 1814400.0 1323000.0 1828200.0 ;
      RECT  1312800.0 1842000.0 1323000.0 1828200.0 ;
      RECT  1312800.0 1842000.0 1323000.0 1855800.0 ;
      RECT  1312800.0 1869600.0 1323000.0 1855800.0 ;
      RECT  1312800.0 1869600.0 1323000.0 1883400.0 ;
      RECT  1312800.0 1897200.0 1323000.0 1883400.0 ;
      RECT  1312800.0 1897200.0 1323000.0 1911000.0 ;
      RECT  1312800.0 1924800.0 1323000.0 1911000.0 ;
      RECT  1312800.0 1924800.0 1323000.0 1938600.0 ;
      RECT  1312800.0 1952400.0 1323000.0 1938600.0 ;
      RECT  1312800.0 1952400.0 1323000.0 1966200.0 ;
      RECT  1312800.0 1980000.0 1323000.0 1966200.0 ;
      RECT  1312800.0 1980000.0 1323000.0 1993800.0 ;
      RECT  1312800.0 2007600.0 1323000.0 1993800.0 ;
      RECT  1312800.0 2007600.0 1323000.0 2021400.0 ;
      RECT  1312800.0 2035200.0 1323000.0 2021400.0 ;
      RECT  1312800.0 2035200.0 1323000.0 2049000.0 ;
      RECT  1312800.0 2062800.0 1323000.0 2049000.0 ;
      RECT  1312800.0 2062800.0 1323000.0 2076600.0 ;
      RECT  1312800.0 2090400.0 1323000.0 2076600.0 ;
      RECT  1312800.0 2090400.0 1323000.0 2104200.0 ;
      RECT  1312800.0 2118000.0 1323000.0 2104200.0 ;
      RECT  1312800.0 2118000.0 1323000.0 2131800.0 ;
      RECT  1312800.0 2145600.0 1323000.0 2131800.0 ;
      RECT  1323000.0 379200.0 1333200.0 393000.0 ;
      RECT  1323000.0 406800.0 1333200.0 393000.0 ;
      RECT  1323000.0 406800.0 1333200.0 420600.0 ;
      RECT  1323000.0 434400.0 1333200.0 420600.0 ;
      RECT  1323000.0 434400.0 1333200.0 448200.0 ;
      RECT  1323000.0 462000.0 1333200.0 448200.0 ;
      RECT  1323000.0 462000.0 1333200.0 475800.0 ;
      RECT  1323000.0 489600.0 1333200.0 475800.0 ;
      RECT  1323000.0 489600.0 1333200.0 503400.0 ;
      RECT  1323000.0 517200.0 1333200.0 503400.0 ;
      RECT  1323000.0 517200.0 1333200.0 531000.0 ;
      RECT  1323000.0 544800.0 1333200.0 531000.0 ;
      RECT  1323000.0 544800.0 1333200.0 558600.0 ;
      RECT  1323000.0 572400.0 1333200.0 558600.0 ;
      RECT  1323000.0 572400.0 1333200.0 586200.0 ;
      RECT  1323000.0 600000.0 1333200.0 586200.0 ;
      RECT  1323000.0 600000.0 1333200.0 613800.0 ;
      RECT  1323000.0 627600.0 1333200.0 613800.0 ;
      RECT  1323000.0 627600.0 1333200.0 641400.0 ;
      RECT  1323000.0 655200.0 1333200.0 641400.0 ;
      RECT  1323000.0 655200.0 1333200.0 669000.0 ;
      RECT  1323000.0 682800.0 1333200.0 669000.0 ;
      RECT  1323000.0 682800.0 1333200.0 696600.0 ;
      RECT  1323000.0 710400.0 1333200.0 696600.0 ;
      RECT  1323000.0 710400.0 1333200.0 724200.0 ;
      RECT  1323000.0 738000.0 1333200.0 724200.0 ;
      RECT  1323000.0 738000.0 1333200.0 751800.0 ;
      RECT  1323000.0 765600.0 1333200.0 751800.0 ;
      RECT  1323000.0 765600.0 1333200.0 779400.0 ;
      RECT  1323000.0 793200.0 1333200.0 779400.0 ;
      RECT  1323000.0 793200.0 1333200.0 807000.0 ;
      RECT  1323000.0 820800.0 1333200.0 807000.0 ;
      RECT  1323000.0 820800.0 1333200.0 834600.0 ;
      RECT  1323000.0 848400.0 1333200.0 834600.0 ;
      RECT  1323000.0 848400.0 1333200.0 862200.0 ;
      RECT  1323000.0 876000.0 1333200.0 862200.0 ;
      RECT  1323000.0 876000.0 1333200.0 889800.0 ;
      RECT  1323000.0 903600.0 1333200.0 889800.0 ;
      RECT  1323000.0 903600.0 1333200.0 917400.0 ;
      RECT  1323000.0 931200.0 1333200.0 917400.0 ;
      RECT  1323000.0 931200.0 1333200.0 945000.0 ;
      RECT  1323000.0 958800.0 1333200.0 945000.0 ;
      RECT  1323000.0 958800.0 1333200.0 972600.0 ;
      RECT  1323000.0 986400.0 1333200.0 972600.0 ;
      RECT  1323000.0 986400.0 1333200.0 1000200.0 ;
      RECT  1323000.0 1014000.0 1333200.0 1000200.0 ;
      RECT  1323000.0 1014000.0 1333200.0 1027800.0 ;
      RECT  1323000.0 1041600.0 1333200.0 1027800.0 ;
      RECT  1323000.0 1041600.0 1333200.0 1055400.0 ;
      RECT  1323000.0 1069200.0 1333200.0 1055400.0 ;
      RECT  1323000.0 1069200.0 1333200.0 1083000.0 ;
      RECT  1323000.0 1096800.0 1333200.0 1083000.0 ;
      RECT  1323000.0 1096800.0 1333200.0 1110600.0 ;
      RECT  1323000.0 1124400.0 1333200.0 1110600.0 ;
      RECT  1323000.0 1124400.0 1333200.0 1138200.0 ;
      RECT  1323000.0 1152000.0 1333200.0 1138200.0 ;
      RECT  1323000.0 1152000.0 1333200.0 1165800.0 ;
      RECT  1323000.0 1179600.0 1333200.0 1165800.0 ;
      RECT  1323000.0 1179600.0 1333200.0 1193400.0 ;
      RECT  1323000.0 1207200.0 1333200.0 1193400.0 ;
      RECT  1323000.0 1207200.0 1333200.0 1221000.0 ;
      RECT  1323000.0 1234800.0 1333200.0 1221000.0 ;
      RECT  1323000.0 1234800.0 1333200.0 1248600.0 ;
      RECT  1323000.0 1262400.0 1333200.0 1248600.0 ;
      RECT  1323000.0 1262400.0 1333200.0 1276200.0 ;
      RECT  1323000.0 1290000.0 1333200.0 1276200.0 ;
      RECT  1323000.0 1290000.0 1333200.0 1303800.0 ;
      RECT  1323000.0 1317600.0 1333200.0 1303800.0 ;
      RECT  1323000.0 1317600.0 1333200.0 1331400.0 ;
      RECT  1323000.0 1345200.0 1333200.0 1331400.0 ;
      RECT  1323000.0 1345200.0 1333200.0 1359000.0 ;
      RECT  1323000.0 1372800.0 1333200.0 1359000.0 ;
      RECT  1323000.0 1372800.0 1333200.0 1386600.0 ;
      RECT  1323000.0 1400400.0 1333200.0 1386600.0 ;
      RECT  1323000.0 1400400.0 1333200.0 1414200.0 ;
      RECT  1323000.0 1428000.0 1333200.0 1414200.0 ;
      RECT  1323000.0 1428000.0 1333200.0 1441800.0 ;
      RECT  1323000.0 1455600.0 1333200.0 1441800.0 ;
      RECT  1323000.0 1455600.0 1333200.0 1469400.0 ;
      RECT  1323000.0 1483200.0 1333200.0 1469400.0 ;
      RECT  1323000.0 1483200.0 1333200.0 1497000.0 ;
      RECT  1323000.0 1510800.0 1333200.0 1497000.0 ;
      RECT  1323000.0 1510800.0 1333200.0 1524600.0 ;
      RECT  1323000.0 1538400.0 1333200.0 1524600.0 ;
      RECT  1323000.0 1538400.0 1333200.0 1552200.0 ;
      RECT  1323000.0 1566000.0 1333200.0 1552200.0 ;
      RECT  1323000.0 1566000.0 1333200.0 1579800.0 ;
      RECT  1323000.0 1593600.0 1333200.0 1579800.0 ;
      RECT  1323000.0 1593600.0 1333200.0 1607400.0 ;
      RECT  1323000.0 1621200.0 1333200.0 1607400.0 ;
      RECT  1323000.0 1621200.0 1333200.0 1635000.0 ;
      RECT  1323000.0 1648800.0 1333200.0 1635000.0 ;
      RECT  1323000.0 1648800.0 1333200.0 1662600.0 ;
      RECT  1323000.0 1676400.0 1333200.0 1662600.0 ;
      RECT  1323000.0 1676400.0 1333200.0 1690200.0 ;
      RECT  1323000.0 1704000.0 1333200.0 1690200.0 ;
      RECT  1323000.0 1704000.0 1333200.0 1717800.0 ;
      RECT  1323000.0 1731600.0 1333200.0 1717800.0 ;
      RECT  1323000.0 1731600.0 1333200.0 1745400.0 ;
      RECT  1323000.0 1759200.0 1333200.0 1745400.0 ;
      RECT  1323000.0 1759200.0 1333200.0 1773000.0 ;
      RECT  1323000.0 1786800.0 1333200.0 1773000.0 ;
      RECT  1323000.0 1786800.0 1333200.0 1800600.0 ;
      RECT  1323000.0 1814400.0 1333200.0 1800600.0 ;
      RECT  1323000.0 1814400.0 1333200.0 1828200.0 ;
      RECT  1323000.0 1842000.0 1333200.0 1828200.0 ;
      RECT  1323000.0 1842000.0 1333200.0 1855800.0 ;
      RECT  1323000.0 1869600.0 1333200.0 1855800.0 ;
      RECT  1323000.0 1869600.0 1333200.0 1883400.0 ;
      RECT  1323000.0 1897200.0 1333200.0 1883400.0 ;
      RECT  1323000.0 1897200.0 1333200.0 1911000.0 ;
      RECT  1323000.0 1924800.0 1333200.0 1911000.0 ;
      RECT  1323000.0 1924800.0 1333200.0 1938600.0 ;
      RECT  1323000.0 1952400.0 1333200.0 1938600.0 ;
      RECT  1323000.0 1952400.0 1333200.0 1966200.0 ;
      RECT  1323000.0 1980000.0 1333200.0 1966200.0 ;
      RECT  1323000.0 1980000.0 1333200.0 1993800.0 ;
      RECT  1323000.0 2007600.0 1333200.0 1993800.0 ;
      RECT  1323000.0 2007600.0 1333200.0 2021400.0 ;
      RECT  1323000.0 2035200.0 1333200.0 2021400.0 ;
      RECT  1323000.0 2035200.0 1333200.0 2049000.0 ;
      RECT  1323000.0 2062800.0 1333200.0 2049000.0 ;
      RECT  1323000.0 2062800.0 1333200.0 2076600.0 ;
      RECT  1323000.0 2090400.0 1333200.0 2076600.0 ;
      RECT  1323000.0 2090400.0 1333200.0 2104200.0 ;
      RECT  1323000.0 2118000.0 1333200.0 2104200.0 ;
      RECT  1323000.0 2118000.0 1333200.0 2131800.0 ;
      RECT  1323000.0 2145600.0 1333200.0 2131800.0 ;
      RECT  1333200.0 379200.0 1343400.0 393000.0 ;
      RECT  1333200.0 406800.0 1343400.0 393000.0 ;
      RECT  1333200.0 406800.0 1343400.0 420600.0 ;
      RECT  1333200.0 434400.0 1343400.0 420600.0 ;
      RECT  1333200.0 434400.0 1343400.0 448200.0 ;
      RECT  1333200.0 462000.0 1343400.0 448200.0 ;
      RECT  1333200.0 462000.0 1343400.0 475800.0 ;
      RECT  1333200.0 489600.0 1343400.0 475800.0 ;
      RECT  1333200.0 489600.0 1343400.0 503400.0 ;
      RECT  1333200.0 517200.0 1343400.0 503400.0 ;
      RECT  1333200.0 517200.0 1343400.0 531000.0 ;
      RECT  1333200.0 544800.0 1343400.0 531000.0 ;
      RECT  1333200.0 544800.0 1343400.0 558600.0 ;
      RECT  1333200.0 572400.0 1343400.0 558600.0 ;
      RECT  1333200.0 572400.0 1343400.0 586200.0 ;
      RECT  1333200.0 600000.0 1343400.0 586200.0 ;
      RECT  1333200.0 600000.0 1343400.0 613800.0 ;
      RECT  1333200.0 627600.0 1343400.0 613800.0 ;
      RECT  1333200.0 627600.0 1343400.0 641400.0 ;
      RECT  1333200.0 655200.0 1343400.0 641400.0 ;
      RECT  1333200.0 655200.0 1343400.0 669000.0 ;
      RECT  1333200.0 682800.0 1343400.0 669000.0 ;
      RECT  1333200.0 682800.0 1343400.0 696600.0 ;
      RECT  1333200.0 710400.0 1343400.0 696600.0 ;
      RECT  1333200.0 710400.0 1343400.0 724200.0 ;
      RECT  1333200.0 738000.0 1343400.0 724200.0 ;
      RECT  1333200.0 738000.0 1343400.0 751800.0 ;
      RECT  1333200.0 765600.0 1343400.0 751800.0 ;
      RECT  1333200.0 765600.0 1343400.0 779400.0 ;
      RECT  1333200.0 793200.0 1343400.0 779400.0 ;
      RECT  1333200.0 793200.0 1343400.0 807000.0 ;
      RECT  1333200.0 820800.0 1343400.0 807000.0 ;
      RECT  1333200.0 820800.0 1343400.0 834600.0 ;
      RECT  1333200.0 848400.0 1343400.0 834600.0 ;
      RECT  1333200.0 848400.0 1343400.0 862200.0 ;
      RECT  1333200.0 876000.0 1343400.0 862200.0 ;
      RECT  1333200.0 876000.0 1343400.0 889800.0 ;
      RECT  1333200.0 903600.0 1343400.0 889800.0 ;
      RECT  1333200.0 903600.0 1343400.0 917400.0 ;
      RECT  1333200.0 931200.0 1343400.0 917400.0 ;
      RECT  1333200.0 931200.0 1343400.0 945000.0 ;
      RECT  1333200.0 958800.0 1343400.0 945000.0 ;
      RECT  1333200.0 958800.0 1343400.0 972600.0 ;
      RECT  1333200.0 986400.0 1343400.0 972600.0 ;
      RECT  1333200.0 986400.0 1343400.0 1000200.0 ;
      RECT  1333200.0 1014000.0 1343400.0 1000200.0 ;
      RECT  1333200.0 1014000.0 1343400.0 1027800.0 ;
      RECT  1333200.0 1041600.0 1343400.0 1027800.0 ;
      RECT  1333200.0 1041600.0 1343400.0 1055400.0 ;
      RECT  1333200.0 1069200.0 1343400.0 1055400.0 ;
      RECT  1333200.0 1069200.0 1343400.0 1083000.0 ;
      RECT  1333200.0 1096800.0 1343400.0 1083000.0 ;
      RECT  1333200.0 1096800.0 1343400.0 1110600.0 ;
      RECT  1333200.0 1124400.0 1343400.0 1110600.0 ;
      RECT  1333200.0 1124400.0 1343400.0 1138200.0 ;
      RECT  1333200.0 1152000.0 1343400.0 1138200.0 ;
      RECT  1333200.0 1152000.0 1343400.0 1165800.0 ;
      RECT  1333200.0 1179600.0 1343400.0 1165800.0 ;
      RECT  1333200.0 1179600.0 1343400.0 1193400.0 ;
      RECT  1333200.0 1207200.0 1343400.0 1193400.0 ;
      RECT  1333200.0 1207200.0 1343400.0 1221000.0 ;
      RECT  1333200.0 1234800.0 1343400.0 1221000.0 ;
      RECT  1333200.0 1234800.0 1343400.0 1248600.0 ;
      RECT  1333200.0 1262400.0 1343400.0 1248600.0 ;
      RECT  1333200.0 1262400.0 1343400.0 1276200.0 ;
      RECT  1333200.0 1290000.0 1343400.0 1276200.0 ;
      RECT  1333200.0 1290000.0 1343400.0 1303800.0 ;
      RECT  1333200.0 1317600.0 1343400.0 1303800.0 ;
      RECT  1333200.0 1317600.0 1343400.0 1331400.0 ;
      RECT  1333200.0 1345200.0 1343400.0 1331400.0 ;
      RECT  1333200.0 1345200.0 1343400.0 1359000.0 ;
      RECT  1333200.0 1372800.0 1343400.0 1359000.0 ;
      RECT  1333200.0 1372800.0 1343400.0 1386600.0 ;
      RECT  1333200.0 1400400.0 1343400.0 1386600.0 ;
      RECT  1333200.0 1400400.0 1343400.0 1414200.0 ;
      RECT  1333200.0 1428000.0 1343400.0 1414200.0 ;
      RECT  1333200.0 1428000.0 1343400.0 1441800.0 ;
      RECT  1333200.0 1455600.0 1343400.0 1441800.0 ;
      RECT  1333200.0 1455600.0 1343400.0 1469400.0 ;
      RECT  1333200.0 1483200.0 1343400.0 1469400.0 ;
      RECT  1333200.0 1483200.0 1343400.0 1497000.0 ;
      RECT  1333200.0 1510800.0 1343400.0 1497000.0 ;
      RECT  1333200.0 1510800.0 1343400.0 1524600.0 ;
      RECT  1333200.0 1538400.0 1343400.0 1524600.0 ;
      RECT  1333200.0 1538400.0 1343400.0 1552200.0 ;
      RECT  1333200.0 1566000.0 1343400.0 1552200.0 ;
      RECT  1333200.0 1566000.0 1343400.0 1579800.0 ;
      RECT  1333200.0 1593600.0 1343400.0 1579800.0 ;
      RECT  1333200.0 1593600.0 1343400.0 1607400.0 ;
      RECT  1333200.0 1621200.0 1343400.0 1607400.0 ;
      RECT  1333200.0 1621200.0 1343400.0 1635000.0 ;
      RECT  1333200.0 1648800.0 1343400.0 1635000.0 ;
      RECT  1333200.0 1648800.0 1343400.0 1662600.0 ;
      RECT  1333200.0 1676400.0 1343400.0 1662600.0 ;
      RECT  1333200.0 1676400.0 1343400.0 1690200.0 ;
      RECT  1333200.0 1704000.0 1343400.0 1690200.0 ;
      RECT  1333200.0 1704000.0 1343400.0 1717800.0 ;
      RECT  1333200.0 1731600.0 1343400.0 1717800.0 ;
      RECT  1333200.0 1731600.0 1343400.0 1745400.0 ;
      RECT  1333200.0 1759200.0 1343400.0 1745400.0 ;
      RECT  1333200.0 1759200.0 1343400.0 1773000.0 ;
      RECT  1333200.0 1786800.0 1343400.0 1773000.0 ;
      RECT  1333200.0 1786800.0 1343400.0 1800600.0 ;
      RECT  1333200.0 1814400.0 1343400.0 1800600.0 ;
      RECT  1333200.0 1814400.0 1343400.0 1828200.0 ;
      RECT  1333200.0 1842000.0 1343400.0 1828200.0 ;
      RECT  1333200.0 1842000.0 1343400.0 1855800.0 ;
      RECT  1333200.0 1869600.0 1343400.0 1855800.0 ;
      RECT  1333200.0 1869600.0 1343400.0 1883400.0 ;
      RECT  1333200.0 1897200.0 1343400.0 1883400.0 ;
      RECT  1333200.0 1897200.0 1343400.0 1911000.0 ;
      RECT  1333200.0 1924800.0 1343400.0 1911000.0 ;
      RECT  1333200.0 1924800.0 1343400.0 1938600.0 ;
      RECT  1333200.0 1952400.0 1343400.0 1938600.0 ;
      RECT  1333200.0 1952400.0 1343400.0 1966200.0 ;
      RECT  1333200.0 1980000.0 1343400.0 1966200.0 ;
      RECT  1333200.0 1980000.0 1343400.0 1993800.0 ;
      RECT  1333200.0 2007600.0 1343400.0 1993800.0 ;
      RECT  1333200.0 2007600.0 1343400.0 2021400.0 ;
      RECT  1333200.0 2035200.0 1343400.0 2021400.0 ;
      RECT  1333200.0 2035200.0 1343400.0 2049000.0 ;
      RECT  1333200.0 2062800.0 1343400.0 2049000.0 ;
      RECT  1333200.0 2062800.0 1343400.0 2076600.0 ;
      RECT  1333200.0 2090400.0 1343400.0 2076600.0 ;
      RECT  1333200.0 2090400.0 1343400.0 2104200.0 ;
      RECT  1333200.0 2118000.0 1343400.0 2104200.0 ;
      RECT  1333200.0 2118000.0 1343400.0 2131800.0 ;
      RECT  1333200.0 2145600.0 1343400.0 2131800.0 ;
      RECT  1343400.0 379200.0 1353600.0 393000.0 ;
      RECT  1343400.0 406800.0 1353600.0 393000.0 ;
      RECT  1343400.0 406800.0 1353600.0 420600.0 ;
      RECT  1343400.0 434400.0 1353600.0 420600.0 ;
      RECT  1343400.0 434400.0 1353600.0 448200.0 ;
      RECT  1343400.0 462000.0 1353600.0 448200.0 ;
      RECT  1343400.0 462000.0 1353600.0 475800.0 ;
      RECT  1343400.0 489600.0 1353600.0 475800.0 ;
      RECT  1343400.0 489600.0 1353600.0 503400.0 ;
      RECT  1343400.0 517200.0 1353600.0 503400.0 ;
      RECT  1343400.0 517200.0 1353600.0 531000.0 ;
      RECT  1343400.0 544800.0 1353600.0 531000.0 ;
      RECT  1343400.0 544800.0 1353600.0 558600.0 ;
      RECT  1343400.0 572400.0 1353600.0 558600.0 ;
      RECT  1343400.0 572400.0 1353600.0 586200.0 ;
      RECT  1343400.0 600000.0 1353600.0 586200.0 ;
      RECT  1343400.0 600000.0 1353600.0 613800.0 ;
      RECT  1343400.0 627600.0 1353600.0 613800.0 ;
      RECT  1343400.0 627600.0 1353600.0 641400.0 ;
      RECT  1343400.0 655200.0 1353600.0 641400.0 ;
      RECT  1343400.0 655200.0 1353600.0 669000.0 ;
      RECT  1343400.0 682800.0 1353600.0 669000.0 ;
      RECT  1343400.0 682800.0 1353600.0 696600.0 ;
      RECT  1343400.0 710400.0 1353600.0 696600.0 ;
      RECT  1343400.0 710400.0 1353600.0 724200.0 ;
      RECT  1343400.0 738000.0 1353600.0 724200.0 ;
      RECT  1343400.0 738000.0 1353600.0 751800.0 ;
      RECT  1343400.0 765600.0 1353600.0 751800.0 ;
      RECT  1343400.0 765600.0 1353600.0 779400.0 ;
      RECT  1343400.0 793200.0 1353600.0 779400.0 ;
      RECT  1343400.0 793200.0 1353600.0 807000.0 ;
      RECT  1343400.0 820800.0 1353600.0 807000.0 ;
      RECT  1343400.0 820800.0 1353600.0 834600.0 ;
      RECT  1343400.0 848400.0 1353600.0 834600.0 ;
      RECT  1343400.0 848400.0 1353600.0 862200.0 ;
      RECT  1343400.0 876000.0 1353600.0 862200.0 ;
      RECT  1343400.0 876000.0 1353600.0 889800.0 ;
      RECT  1343400.0 903600.0 1353600.0 889800.0 ;
      RECT  1343400.0 903600.0 1353600.0 917400.0 ;
      RECT  1343400.0 931200.0 1353600.0 917400.0 ;
      RECT  1343400.0 931200.0 1353600.0 945000.0 ;
      RECT  1343400.0 958800.0 1353600.0 945000.0 ;
      RECT  1343400.0 958800.0 1353600.0 972600.0 ;
      RECT  1343400.0 986400.0 1353600.0 972600.0 ;
      RECT  1343400.0 986400.0 1353600.0 1000200.0 ;
      RECT  1343400.0 1014000.0 1353600.0 1000200.0 ;
      RECT  1343400.0 1014000.0 1353600.0 1027800.0 ;
      RECT  1343400.0 1041600.0 1353600.0 1027800.0 ;
      RECT  1343400.0 1041600.0 1353600.0 1055400.0 ;
      RECT  1343400.0 1069200.0 1353600.0 1055400.0 ;
      RECT  1343400.0 1069200.0 1353600.0 1083000.0 ;
      RECT  1343400.0 1096800.0 1353600.0 1083000.0 ;
      RECT  1343400.0 1096800.0 1353600.0 1110600.0 ;
      RECT  1343400.0 1124400.0 1353600.0 1110600.0 ;
      RECT  1343400.0 1124400.0 1353600.0 1138200.0 ;
      RECT  1343400.0 1152000.0 1353600.0 1138200.0 ;
      RECT  1343400.0 1152000.0 1353600.0 1165800.0 ;
      RECT  1343400.0 1179600.0 1353600.0 1165800.0 ;
      RECT  1343400.0 1179600.0 1353600.0 1193400.0 ;
      RECT  1343400.0 1207200.0 1353600.0 1193400.0 ;
      RECT  1343400.0 1207200.0 1353600.0 1221000.0 ;
      RECT  1343400.0 1234800.0 1353600.0 1221000.0 ;
      RECT  1343400.0 1234800.0 1353600.0 1248600.0 ;
      RECT  1343400.0 1262400.0 1353600.0 1248600.0 ;
      RECT  1343400.0 1262400.0 1353600.0 1276200.0 ;
      RECT  1343400.0 1290000.0 1353600.0 1276200.0 ;
      RECT  1343400.0 1290000.0 1353600.0 1303800.0 ;
      RECT  1343400.0 1317600.0 1353600.0 1303800.0 ;
      RECT  1343400.0 1317600.0 1353600.0 1331400.0 ;
      RECT  1343400.0 1345200.0 1353600.0 1331400.0 ;
      RECT  1343400.0 1345200.0 1353600.0 1359000.0 ;
      RECT  1343400.0 1372800.0 1353600.0 1359000.0 ;
      RECT  1343400.0 1372800.0 1353600.0 1386600.0 ;
      RECT  1343400.0 1400400.0 1353600.0 1386600.0 ;
      RECT  1343400.0 1400400.0 1353600.0 1414200.0 ;
      RECT  1343400.0 1428000.0 1353600.0 1414200.0 ;
      RECT  1343400.0 1428000.0 1353600.0 1441800.0 ;
      RECT  1343400.0 1455600.0 1353600.0 1441800.0 ;
      RECT  1343400.0 1455600.0 1353600.0 1469400.0 ;
      RECT  1343400.0 1483200.0 1353600.0 1469400.0 ;
      RECT  1343400.0 1483200.0 1353600.0 1497000.0 ;
      RECT  1343400.0 1510800.0 1353600.0 1497000.0 ;
      RECT  1343400.0 1510800.0 1353600.0 1524600.0 ;
      RECT  1343400.0 1538400.0 1353600.0 1524600.0 ;
      RECT  1343400.0 1538400.0 1353600.0 1552200.0 ;
      RECT  1343400.0 1566000.0 1353600.0 1552200.0 ;
      RECT  1343400.0 1566000.0 1353600.0 1579800.0 ;
      RECT  1343400.0 1593600.0 1353600.0 1579800.0 ;
      RECT  1343400.0 1593600.0 1353600.0 1607400.0 ;
      RECT  1343400.0 1621200.0 1353600.0 1607400.0 ;
      RECT  1343400.0 1621200.0 1353600.0 1635000.0 ;
      RECT  1343400.0 1648800.0 1353600.0 1635000.0 ;
      RECT  1343400.0 1648800.0 1353600.0 1662600.0 ;
      RECT  1343400.0 1676400.0 1353600.0 1662600.0 ;
      RECT  1343400.0 1676400.0 1353600.0 1690200.0 ;
      RECT  1343400.0 1704000.0 1353600.0 1690200.0 ;
      RECT  1343400.0 1704000.0 1353600.0 1717800.0 ;
      RECT  1343400.0 1731600.0 1353600.0 1717800.0 ;
      RECT  1343400.0 1731600.0 1353600.0 1745400.0 ;
      RECT  1343400.0 1759200.0 1353600.0 1745400.0 ;
      RECT  1343400.0 1759200.0 1353600.0 1773000.0 ;
      RECT  1343400.0 1786800.0 1353600.0 1773000.0 ;
      RECT  1343400.0 1786800.0 1353600.0 1800600.0 ;
      RECT  1343400.0 1814400.0 1353600.0 1800600.0 ;
      RECT  1343400.0 1814400.0 1353600.0 1828200.0 ;
      RECT  1343400.0 1842000.0 1353600.0 1828200.0 ;
      RECT  1343400.0 1842000.0 1353600.0 1855800.0 ;
      RECT  1343400.0 1869600.0 1353600.0 1855800.0 ;
      RECT  1343400.0 1869600.0 1353600.0 1883400.0 ;
      RECT  1343400.0 1897200.0 1353600.0 1883400.0 ;
      RECT  1343400.0 1897200.0 1353600.0 1911000.0 ;
      RECT  1343400.0 1924800.0 1353600.0 1911000.0 ;
      RECT  1343400.0 1924800.0 1353600.0 1938600.0 ;
      RECT  1343400.0 1952400.0 1353600.0 1938600.0 ;
      RECT  1343400.0 1952400.0 1353600.0 1966200.0 ;
      RECT  1343400.0 1980000.0 1353600.0 1966200.0 ;
      RECT  1343400.0 1980000.0 1353600.0 1993800.0 ;
      RECT  1343400.0 2007600.0 1353600.0 1993800.0 ;
      RECT  1343400.0 2007600.0 1353600.0 2021400.0 ;
      RECT  1343400.0 2035200.0 1353600.0 2021400.0 ;
      RECT  1343400.0 2035200.0 1353600.0 2049000.0 ;
      RECT  1343400.0 2062800.0 1353600.0 2049000.0 ;
      RECT  1343400.0 2062800.0 1353600.0 2076600.0 ;
      RECT  1343400.0 2090400.0 1353600.0 2076600.0 ;
      RECT  1343400.0 2090400.0 1353600.0 2104200.0 ;
      RECT  1343400.0 2118000.0 1353600.0 2104200.0 ;
      RECT  1343400.0 2118000.0 1353600.0 2131800.0 ;
      RECT  1343400.0 2145600.0 1353600.0 2131800.0 ;
      RECT  1353600.0 379200.0 1363800.0 393000.0 ;
      RECT  1353600.0 406800.0 1363800.0 393000.0 ;
      RECT  1353600.0 406800.0 1363800.0 420600.0 ;
      RECT  1353600.0 434400.0 1363800.0 420600.0 ;
      RECT  1353600.0 434400.0 1363800.0 448200.0 ;
      RECT  1353600.0 462000.0 1363800.0 448200.0 ;
      RECT  1353600.0 462000.0 1363800.0 475800.0 ;
      RECT  1353600.0 489600.0 1363800.0 475800.0 ;
      RECT  1353600.0 489600.0 1363800.0 503400.0 ;
      RECT  1353600.0 517200.0 1363800.0 503400.0 ;
      RECT  1353600.0 517200.0 1363800.0 531000.0 ;
      RECT  1353600.0 544800.0 1363800.0 531000.0 ;
      RECT  1353600.0 544800.0 1363800.0 558600.0 ;
      RECT  1353600.0 572400.0 1363800.0 558600.0 ;
      RECT  1353600.0 572400.0 1363800.0 586200.0 ;
      RECT  1353600.0 600000.0 1363800.0 586200.0 ;
      RECT  1353600.0 600000.0 1363800.0 613800.0 ;
      RECT  1353600.0 627600.0 1363800.0 613800.0 ;
      RECT  1353600.0 627600.0 1363800.0 641400.0 ;
      RECT  1353600.0 655200.0 1363800.0 641400.0 ;
      RECT  1353600.0 655200.0 1363800.0 669000.0 ;
      RECT  1353600.0 682800.0 1363800.0 669000.0 ;
      RECT  1353600.0 682800.0 1363800.0 696600.0 ;
      RECT  1353600.0 710400.0 1363800.0 696600.0 ;
      RECT  1353600.0 710400.0 1363800.0 724200.0 ;
      RECT  1353600.0 738000.0 1363800.0 724200.0 ;
      RECT  1353600.0 738000.0 1363800.0 751800.0 ;
      RECT  1353600.0 765600.0 1363800.0 751800.0 ;
      RECT  1353600.0 765600.0 1363800.0 779400.0 ;
      RECT  1353600.0 793200.0 1363800.0 779400.0 ;
      RECT  1353600.0 793200.0 1363800.0 807000.0 ;
      RECT  1353600.0 820800.0 1363800.0 807000.0 ;
      RECT  1353600.0 820800.0 1363800.0 834600.0 ;
      RECT  1353600.0 848400.0 1363800.0 834600.0 ;
      RECT  1353600.0 848400.0 1363800.0 862200.0 ;
      RECT  1353600.0 876000.0 1363800.0 862200.0 ;
      RECT  1353600.0 876000.0 1363800.0 889800.0 ;
      RECT  1353600.0 903600.0 1363800.0 889800.0 ;
      RECT  1353600.0 903600.0 1363800.0 917400.0 ;
      RECT  1353600.0 931200.0 1363800.0 917400.0 ;
      RECT  1353600.0 931200.0 1363800.0 945000.0 ;
      RECT  1353600.0 958800.0 1363800.0 945000.0 ;
      RECT  1353600.0 958800.0 1363800.0 972600.0 ;
      RECT  1353600.0 986400.0 1363800.0 972600.0 ;
      RECT  1353600.0 986400.0 1363800.0 1000200.0 ;
      RECT  1353600.0 1014000.0 1363800.0 1000200.0 ;
      RECT  1353600.0 1014000.0 1363800.0 1027800.0 ;
      RECT  1353600.0 1041600.0 1363800.0 1027800.0 ;
      RECT  1353600.0 1041600.0 1363800.0 1055400.0 ;
      RECT  1353600.0 1069200.0 1363800.0 1055400.0 ;
      RECT  1353600.0 1069200.0 1363800.0 1083000.0 ;
      RECT  1353600.0 1096800.0 1363800.0 1083000.0 ;
      RECT  1353600.0 1096800.0 1363800.0 1110600.0 ;
      RECT  1353600.0 1124400.0 1363800.0 1110600.0 ;
      RECT  1353600.0 1124400.0 1363800.0 1138200.0 ;
      RECT  1353600.0 1152000.0 1363800.0 1138200.0 ;
      RECT  1353600.0 1152000.0 1363800.0 1165800.0 ;
      RECT  1353600.0 1179600.0 1363800.0 1165800.0 ;
      RECT  1353600.0 1179600.0 1363800.0 1193400.0 ;
      RECT  1353600.0 1207200.0 1363800.0 1193400.0 ;
      RECT  1353600.0 1207200.0 1363800.0 1221000.0 ;
      RECT  1353600.0 1234800.0 1363800.0 1221000.0 ;
      RECT  1353600.0 1234800.0 1363800.0 1248600.0 ;
      RECT  1353600.0 1262400.0 1363800.0 1248600.0 ;
      RECT  1353600.0 1262400.0 1363800.0 1276200.0 ;
      RECT  1353600.0 1290000.0 1363800.0 1276200.0 ;
      RECT  1353600.0 1290000.0 1363800.0 1303800.0 ;
      RECT  1353600.0 1317600.0 1363800.0 1303800.0 ;
      RECT  1353600.0 1317600.0 1363800.0 1331400.0 ;
      RECT  1353600.0 1345200.0 1363800.0 1331400.0 ;
      RECT  1353600.0 1345200.0 1363800.0 1359000.0 ;
      RECT  1353600.0 1372800.0 1363800.0 1359000.0 ;
      RECT  1353600.0 1372800.0 1363800.0 1386600.0 ;
      RECT  1353600.0 1400400.0 1363800.0 1386600.0 ;
      RECT  1353600.0 1400400.0 1363800.0 1414200.0 ;
      RECT  1353600.0 1428000.0 1363800.0 1414200.0 ;
      RECT  1353600.0 1428000.0 1363800.0 1441800.0 ;
      RECT  1353600.0 1455600.0 1363800.0 1441800.0 ;
      RECT  1353600.0 1455600.0 1363800.0 1469400.0 ;
      RECT  1353600.0 1483200.0 1363800.0 1469400.0 ;
      RECT  1353600.0 1483200.0 1363800.0 1497000.0 ;
      RECT  1353600.0 1510800.0 1363800.0 1497000.0 ;
      RECT  1353600.0 1510800.0 1363800.0 1524600.0 ;
      RECT  1353600.0 1538400.0 1363800.0 1524600.0 ;
      RECT  1353600.0 1538400.0 1363800.0 1552200.0 ;
      RECT  1353600.0 1566000.0 1363800.0 1552200.0 ;
      RECT  1353600.0 1566000.0 1363800.0 1579800.0 ;
      RECT  1353600.0 1593600.0 1363800.0 1579800.0 ;
      RECT  1353600.0 1593600.0 1363800.0 1607400.0 ;
      RECT  1353600.0 1621200.0 1363800.0 1607400.0 ;
      RECT  1353600.0 1621200.0 1363800.0 1635000.0 ;
      RECT  1353600.0 1648800.0 1363800.0 1635000.0 ;
      RECT  1353600.0 1648800.0 1363800.0 1662600.0 ;
      RECT  1353600.0 1676400.0 1363800.0 1662600.0 ;
      RECT  1353600.0 1676400.0 1363800.0 1690200.0 ;
      RECT  1353600.0 1704000.0 1363800.0 1690200.0 ;
      RECT  1353600.0 1704000.0 1363800.0 1717800.0 ;
      RECT  1353600.0 1731600.0 1363800.0 1717800.0 ;
      RECT  1353600.0 1731600.0 1363800.0 1745400.0 ;
      RECT  1353600.0 1759200.0 1363800.0 1745400.0 ;
      RECT  1353600.0 1759200.0 1363800.0 1773000.0 ;
      RECT  1353600.0 1786800.0 1363800.0 1773000.0 ;
      RECT  1353600.0 1786800.0 1363800.0 1800600.0 ;
      RECT  1353600.0 1814400.0 1363800.0 1800600.0 ;
      RECT  1353600.0 1814400.0 1363800.0 1828200.0 ;
      RECT  1353600.0 1842000.0 1363800.0 1828200.0 ;
      RECT  1353600.0 1842000.0 1363800.0 1855800.0 ;
      RECT  1353600.0 1869600.0 1363800.0 1855800.0 ;
      RECT  1353600.0 1869600.0 1363800.0 1883400.0 ;
      RECT  1353600.0 1897200.0 1363800.0 1883400.0 ;
      RECT  1353600.0 1897200.0 1363800.0 1911000.0 ;
      RECT  1353600.0 1924800.0 1363800.0 1911000.0 ;
      RECT  1353600.0 1924800.0 1363800.0 1938600.0 ;
      RECT  1353600.0 1952400.0 1363800.0 1938600.0 ;
      RECT  1353600.0 1952400.0 1363800.0 1966200.0 ;
      RECT  1353600.0 1980000.0 1363800.0 1966200.0 ;
      RECT  1353600.0 1980000.0 1363800.0 1993800.0 ;
      RECT  1353600.0 2007600.0 1363800.0 1993800.0 ;
      RECT  1353600.0 2007600.0 1363800.0 2021400.0 ;
      RECT  1353600.0 2035200.0 1363800.0 2021400.0 ;
      RECT  1353600.0 2035200.0 1363800.0 2049000.0 ;
      RECT  1353600.0 2062800.0 1363800.0 2049000.0 ;
      RECT  1353600.0 2062800.0 1363800.0 2076600.0 ;
      RECT  1353600.0 2090400.0 1363800.0 2076600.0 ;
      RECT  1353600.0 2090400.0 1363800.0 2104200.0 ;
      RECT  1353600.0 2118000.0 1363800.0 2104200.0 ;
      RECT  1353600.0 2118000.0 1363800.0 2131800.0 ;
      RECT  1353600.0 2145600.0 1363800.0 2131800.0 ;
      RECT  1363800.0 379200.0 1374000.0 393000.0 ;
      RECT  1363800.0 406800.0 1374000.0 393000.0 ;
      RECT  1363800.0 406800.0 1374000.0 420600.0 ;
      RECT  1363800.0 434400.0 1374000.0 420600.0 ;
      RECT  1363800.0 434400.0 1374000.0 448200.0 ;
      RECT  1363800.0 462000.0 1374000.0 448200.0 ;
      RECT  1363800.0 462000.0 1374000.0 475800.0 ;
      RECT  1363800.0 489600.0 1374000.0 475800.0 ;
      RECT  1363800.0 489600.0 1374000.0 503400.0 ;
      RECT  1363800.0 517200.0 1374000.0 503400.0 ;
      RECT  1363800.0 517200.0 1374000.0 531000.0 ;
      RECT  1363800.0 544800.0 1374000.0 531000.0 ;
      RECT  1363800.0 544800.0 1374000.0 558600.0 ;
      RECT  1363800.0 572400.0 1374000.0 558600.0 ;
      RECT  1363800.0 572400.0 1374000.0 586200.0 ;
      RECT  1363800.0 600000.0 1374000.0 586200.0 ;
      RECT  1363800.0 600000.0 1374000.0 613800.0 ;
      RECT  1363800.0 627600.0 1374000.0 613800.0 ;
      RECT  1363800.0 627600.0 1374000.0 641400.0 ;
      RECT  1363800.0 655200.0 1374000.0 641400.0 ;
      RECT  1363800.0 655200.0 1374000.0 669000.0 ;
      RECT  1363800.0 682800.0 1374000.0 669000.0 ;
      RECT  1363800.0 682800.0 1374000.0 696600.0 ;
      RECT  1363800.0 710400.0 1374000.0 696600.0 ;
      RECT  1363800.0 710400.0 1374000.0 724200.0 ;
      RECT  1363800.0 738000.0 1374000.0 724200.0 ;
      RECT  1363800.0 738000.0 1374000.0 751800.0 ;
      RECT  1363800.0 765600.0 1374000.0 751800.0 ;
      RECT  1363800.0 765600.0 1374000.0 779400.0 ;
      RECT  1363800.0 793200.0 1374000.0 779400.0 ;
      RECT  1363800.0 793200.0 1374000.0 807000.0 ;
      RECT  1363800.0 820800.0 1374000.0 807000.0 ;
      RECT  1363800.0 820800.0 1374000.0 834600.0 ;
      RECT  1363800.0 848400.0 1374000.0 834600.0 ;
      RECT  1363800.0 848400.0 1374000.0 862200.0 ;
      RECT  1363800.0 876000.0 1374000.0 862200.0 ;
      RECT  1363800.0 876000.0 1374000.0 889800.0 ;
      RECT  1363800.0 903600.0 1374000.0 889800.0 ;
      RECT  1363800.0 903600.0 1374000.0 917400.0 ;
      RECT  1363800.0 931200.0 1374000.0 917400.0 ;
      RECT  1363800.0 931200.0 1374000.0 945000.0 ;
      RECT  1363800.0 958800.0 1374000.0 945000.0 ;
      RECT  1363800.0 958800.0 1374000.0 972600.0 ;
      RECT  1363800.0 986400.0 1374000.0 972600.0 ;
      RECT  1363800.0 986400.0 1374000.0 1000200.0 ;
      RECT  1363800.0 1014000.0 1374000.0 1000200.0 ;
      RECT  1363800.0 1014000.0 1374000.0 1027800.0 ;
      RECT  1363800.0 1041600.0 1374000.0 1027800.0 ;
      RECT  1363800.0 1041600.0 1374000.0 1055400.0 ;
      RECT  1363800.0 1069200.0 1374000.0 1055400.0 ;
      RECT  1363800.0 1069200.0 1374000.0 1083000.0 ;
      RECT  1363800.0 1096800.0 1374000.0 1083000.0 ;
      RECT  1363800.0 1096800.0 1374000.0 1110600.0 ;
      RECT  1363800.0 1124400.0 1374000.0 1110600.0 ;
      RECT  1363800.0 1124400.0 1374000.0 1138200.0 ;
      RECT  1363800.0 1152000.0 1374000.0 1138200.0 ;
      RECT  1363800.0 1152000.0 1374000.0 1165800.0 ;
      RECT  1363800.0 1179600.0 1374000.0 1165800.0 ;
      RECT  1363800.0 1179600.0 1374000.0 1193400.0 ;
      RECT  1363800.0 1207200.0 1374000.0 1193400.0 ;
      RECT  1363800.0 1207200.0 1374000.0 1221000.0 ;
      RECT  1363800.0 1234800.0 1374000.0 1221000.0 ;
      RECT  1363800.0 1234800.0 1374000.0 1248600.0 ;
      RECT  1363800.0 1262400.0 1374000.0 1248600.0 ;
      RECT  1363800.0 1262400.0 1374000.0 1276200.0 ;
      RECT  1363800.0 1290000.0 1374000.0 1276200.0 ;
      RECT  1363800.0 1290000.0 1374000.0 1303800.0 ;
      RECT  1363800.0 1317600.0 1374000.0 1303800.0 ;
      RECT  1363800.0 1317600.0 1374000.0 1331400.0 ;
      RECT  1363800.0 1345200.0 1374000.0 1331400.0 ;
      RECT  1363800.0 1345200.0 1374000.0 1359000.0 ;
      RECT  1363800.0 1372800.0 1374000.0 1359000.0 ;
      RECT  1363800.0 1372800.0 1374000.0 1386600.0 ;
      RECT  1363800.0 1400400.0 1374000.0 1386600.0 ;
      RECT  1363800.0 1400400.0 1374000.0 1414200.0 ;
      RECT  1363800.0 1428000.0 1374000.0 1414200.0 ;
      RECT  1363800.0 1428000.0 1374000.0 1441800.0 ;
      RECT  1363800.0 1455600.0 1374000.0 1441800.0 ;
      RECT  1363800.0 1455600.0 1374000.0 1469400.0 ;
      RECT  1363800.0 1483200.0 1374000.0 1469400.0 ;
      RECT  1363800.0 1483200.0 1374000.0 1497000.0 ;
      RECT  1363800.0 1510800.0 1374000.0 1497000.0 ;
      RECT  1363800.0 1510800.0 1374000.0 1524600.0 ;
      RECT  1363800.0 1538400.0 1374000.0 1524600.0 ;
      RECT  1363800.0 1538400.0 1374000.0 1552200.0 ;
      RECT  1363800.0 1566000.0 1374000.0 1552200.0 ;
      RECT  1363800.0 1566000.0 1374000.0 1579800.0 ;
      RECT  1363800.0 1593600.0 1374000.0 1579800.0 ;
      RECT  1363800.0 1593600.0 1374000.0 1607400.0 ;
      RECT  1363800.0 1621200.0 1374000.0 1607400.0 ;
      RECT  1363800.0 1621200.0 1374000.0 1635000.0 ;
      RECT  1363800.0 1648800.0 1374000.0 1635000.0 ;
      RECT  1363800.0 1648800.0 1374000.0 1662600.0 ;
      RECT  1363800.0 1676400.0 1374000.0 1662600.0 ;
      RECT  1363800.0 1676400.0 1374000.0 1690200.0 ;
      RECT  1363800.0 1704000.0 1374000.0 1690200.0 ;
      RECT  1363800.0 1704000.0 1374000.0 1717800.0 ;
      RECT  1363800.0 1731600.0 1374000.0 1717800.0 ;
      RECT  1363800.0 1731600.0 1374000.0 1745400.0 ;
      RECT  1363800.0 1759200.0 1374000.0 1745400.0 ;
      RECT  1363800.0 1759200.0 1374000.0 1773000.0 ;
      RECT  1363800.0 1786800.0 1374000.0 1773000.0 ;
      RECT  1363800.0 1786800.0 1374000.0 1800600.0 ;
      RECT  1363800.0 1814400.0 1374000.0 1800600.0 ;
      RECT  1363800.0 1814400.0 1374000.0 1828200.0 ;
      RECT  1363800.0 1842000.0 1374000.0 1828200.0 ;
      RECT  1363800.0 1842000.0 1374000.0 1855800.0 ;
      RECT  1363800.0 1869600.0 1374000.0 1855800.0 ;
      RECT  1363800.0 1869600.0 1374000.0 1883400.0 ;
      RECT  1363800.0 1897200.0 1374000.0 1883400.0 ;
      RECT  1363800.0 1897200.0 1374000.0 1911000.0 ;
      RECT  1363800.0 1924800.0 1374000.0 1911000.0 ;
      RECT  1363800.0 1924800.0 1374000.0 1938600.0 ;
      RECT  1363800.0 1952400.0 1374000.0 1938600.0 ;
      RECT  1363800.0 1952400.0 1374000.0 1966200.0 ;
      RECT  1363800.0 1980000.0 1374000.0 1966200.0 ;
      RECT  1363800.0 1980000.0 1374000.0 1993800.0 ;
      RECT  1363800.0 2007600.0 1374000.0 1993800.0 ;
      RECT  1363800.0 2007600.0 1374000.0 2021400.0 ;
      RECT  1363800.0 2035200.0 1374000.0 2021400.0 ;
      RECT  1363800.0 2035200.0 1374000.0 2049000.0 ;
      RECT  1363800.0 2062800.0 1374000.0 2049000.0 ;
      RECT  1363800.0 2062800.0 1374000.0 2076600.0 ;
      RECT  1363800.0 2090400.0 1374000.0 2076600.0 ;
      RECT  1363800.0 2090400.0 1374000.0 2104200.0 ;
      RECT  1363800.0 2118000.0 1374000.0 2104200.0 ;
      RECT  1363800.0 2118000.0 1374000.0 2131800.0 ;
      RECT  1363800.0 2145600.0 1374000.0 2131800.0 ;
      RECT  1374000.0 379200.0 1384200.0 393000.0 ;
      RECT  1374000.0 406800.0 1384200.0 393000.0 ;
      RECT  1374000.0 406800.0 1384200.0 420600.0 ;
      RECT  1374000.0 434400.0 1384200.0 420600.0 ;
      RECT  1374000.0 434400.0 1384200.0 448200.0 ;
      RECT  1374000.0 462000.0 1384200.0 448200.0 ;
      RECT  1374000.0 462000.0 1384200.0 475800.0 ;
      RECT  1374000.0 489600.0 1384200.0 475800.0 ;
      RECT  1374000.0 489600.0 1384200.0 503400.0 ;
      RECT  1374000.0 517200.0 1384200.0 503400.0 ;
      RECT  1374000.0 517200.0 1384200.0 531000.0 ;
      RECT  1374000.0 544800.0 1384200.0 531000.0 ;
      RECT  1374000.0 544800.0 1384200.0 558600.0 ;
      RECT  1374000.0 572400.0 1384200.0 558600.0 ;
      RECT  1374000.0 572400.0 1384200.0 586200.0 ;
      RECT  1374000.0 600000.0 1384200.0 586200.0 ;
      RECT  1374000.0 600000.0 1384200.0 613800.0 ;
      RECT  1374000.0 627600.0 1384200.0 613800.0 ;
      RECT  1374000.0 627600.0 1384200.0 641400.0 ;
      RECT  1374000.0 655200.0 1384200.0 641400.0 ;
      RECT  1374000.0 655200.0 1384200.0 669000.0 ;
      RECT  1374000.0 682800.0 1384200.0 669000.0 ;
      RECT  1374000.0 682800.0 1384200.0 696600.0 ;
      RECT  1374000.0 710400.0 1384200.0 696600.0 ;
      RECT  1374000.0 710400.0 1384200.0 724200.0 ;
      RECT  1374000.0 738000.0 1384200.0 724200.0 ;
      RECT  1374000.0 738000.0 1384200.0 751800.0 ;
      RECT  1374000.0 765600.0 1384200.0 751800.0 ;
      RECT  1374000.0 765600.0 1384200.0 779400.0 ;
      RECT  1374000.0 793200.0 1384200.0 779400.0 ;
      RECT  1374000.0 793200.0 1384200.0 807000.0 ;
      RECT  1374000.0 820800.0 1384200.0 807000.0 ;
      RECT  1374000.0 820800.0 1384200.0 834600.0 ;
      RECT  1374000.0 848400.0 1384200.0 834600.0 ;
      RECT  1374000.0 848400.0 1384200.0 862200.0 ;
      RECT  1374000.0 876000.0 1384200.0 862200.0 ;
      RECT  1374000.0 876000.0 1384200.0 889800.0 ;
      RECT  1374000.0 903600.0 1384200.0 889800.0 ;
      RECT  1374000.0 903600.0 1384200.0 917400.0 ;
      RECT  1374000.0 931200.0 1384200.0 917400.0 ;
      RECT  1374000.0 931200.0 1384200.0 945000.0 ;
      RECT  1374000.0 958800.0 1384200.0 945000.0 ;
      RECT  1374000.0 958800.0 1384200.0 972600.0 ;
      RECT  1374000.0 986400.0 1384200.0 972600.0 ;
      RECT  1374000.0 986400.0 1384200.0 1000200.0 ;
      RECT  1374000.0 1014000.0 1384200.0 1000200.0 ;
      RECT  1374000.0 1014000.0 1384200.0 1027800.0 ;
      RECT  1374000.0 1041600.0 1384200.0 1027800.0 ;
      RECT  1374000.0 1041600.0 1384200.0 1055400.0 ;
      RECT  1374000.0 1069200.0 1384200.0 1055400.0 ;
      RECT  1374000.0 1069200.0 1384200.0 1083000.0 ;
      RECT  1374000.0 1096800.0 1384200.0 1083000.0 ;
      RECT  1374000.0 1096800.0 1384200.0 1110600.0 ;
      RECT  1374000.0 1124400.0 1384200.0 1110600.0 ;
      RECT  1374000.0 1124400.0 1384200.0 1138200.0 ;
      RECT  1374000.0 1152000.0 1384200.0 1138200.0 ;
      RECT  1374000.0 1152000.0 1384200.0 1165800.0 ;
      RECT  1374000.0 1179600.0 1384200.0 1165800.0 ;
      RECT  1374000.0 1179600.0 1384200.0 1193400.0 ;
      RECT  1374000.0 1207200.0 1384200.0 1193400.0 ;
      RECT  1374000.0 1207200.0 1384200.0 1221000.0 ;
      RECT  1374000.0 1234800.0 1384200.0 1221000.0 ;
      RECT  1374000.0 1234800.0 1384200.0 1248600.0 ;
      RECT  1374000.0 1262400.0 1384200.0 1248600.0 ;
      RECT  1374000.0 1262400.0 1384200.0 1276200.0 ;
      RECT  1374000.0 1290000.0 1384200.0 1276200.0 ;
      RECT  1374000.0 1290000.0 1384200.0 1303800.0 ;
      RECT  1374000.0 1317600.0 1384200.0 1303800.0 ;
      RECT  1374000.0 1317600.0 1384200.0 1331400.0 ;
      RECT  1374000.0 1345200.0 1384200.0 1331400.0 ;
      RECT  1374000.0 1345200.0 1384200.0 1359000.0 ;
      RECT  1374000.0 1372800.0 1384200.0 1359000.0 ;
      RECT  1374000.0 1372800.0 1384200.0 1386600.0 ;
      RECT  1374000.0 1400400.0 1384200.0 1386600.0 ;
      RECT  1374000.0 1400400.0 1384200.0 1414200.0 ;
      RECT  1374000.0 1428000.0 1384200.0 1414200.0 ;
      RECT  1374000.0 1428000.0 1384200.0 1441800.0 ;
      RECT  1374000.0 1455600.0 1384200.0 1441800.0 ;
      RECT  1374000.0 1455600.0 1384200.0 1469400.0 ;
      RECT  1374000.0 1483200.0 1384200.0 1469400.0 ;
      RECT  1374000.0 1483200.0 1384200.0 1497000.0 ;
      RECT  1374000.0 1510800.0 1384200.0 1497000.0 ;
      RECT  1374000.0 1510800.0 1384200.0 1524600.0 ;
      RECT  1374000.0 1538400.0 1384200.0 1524600.0 ;
      RECT  1374000.0 1538400.0 1384200.0 1552200.0 ;
      RECT  1374000.0 1566000.0 1384200.0 1552200.0 ;
      RECT  1374000.0 1566000.0 1384200.0 1579800.0 ;
      RECT  1374000.0 1593600.0 1384200.0 1579800.0 ;
      RECT  1374000.0 1593600.0 1384200.0 1607400.0 ;
      RECT  1374000.0 1621200.0 1384200.0 1607400.0 ;
      RECT  1374000.0 1621200.0 1384200.0 1635000.0 ;
      RECT  1374000.0 1648800.0 1384200.0 1635000.0 ;
      RECT  1374000.0 1648800.0 1384200.0 1662600.0 ;
      RECT  1374000.0 1676400.0 1384200.0 1662600.0 ;
      RECT  1374000.0 1676400.0 1384200.0 1690200.0 ;
      RECT  1374000.0 1704000.0 1384200.0 1690200.0 ;
      RECT  1374000.0 1704000.0 1384200.0 1717800.0 ;
      RECT  1374000.0 1731600.0 1384200.0 1717800.0 ;
      RECT  1374000.0 1731600.0 1384200.0 1745400.0 ;
      RECT  1374000.0 1759200.0 1384200.0 1745400.0 ;
      RECT  1374000.0 1759200.0 1384200.0 1773000.0 ;
      RECT  1374000.0 1786800.0 1384200.0 1773000.0 ;
      RECT  1374000.0 1786800.0 1384200.0 1800600.0 ;
      RECT  1374000.0 1814400.0 1384200.0 1800600.0 ;
      RECT  1374000.0 1814400.0 1384200.0 1828200.0 ;
      RECT  1374000.0 1842000.0 1384200.0 1828200.0 ;
      RECT  1374000.0 1842000.0 1384200.0 1855800.0 ;
      RECT  1374000.0 1869600.0 1384200.0 1855800.0 ;
      RECT  1374000.0 1869600.0 1384200.0 1883400.0 ;
      RECT  1374000.0 1897200.0 1384200.0 1883400.0 ;
      RECT  1374000.0 1897200.0 1384200.0 1911000.0 ;
      RECT  1374000.0 1924800.0 1384200.0 1911000.0 ;
      RECT  1374000.0 1924800.0 1384200.0 1938600.0 ;
      RECT  1374000.0 1952400.0 1384200.0 1938600.0 ;
      RECT  1374000.0 1952400.0 1384200.0 1966200.0 ;
      RECT  1374000.0 1980000.0 1384200.0 1966200.0 ;
      RECT  1374000.0 1980000.0 1384200.0 1993800.0 ;
      RECT  1374000.0 2007600.0 1384200.0 1993800.0 ;
      RECT  1374000.0 2007600.0 1384200.0 2021400.0 ;
      RECT  1374000.0 2035200.0 1384200.0 2021400.0 ;
      RECT  1374000.0 2035200.0 1384200.0 2049000.0 ;
      RECT  1374000.0 2062800.0 1384200.0 2049000.0 ;
      RECT  1374000.0 2062800.0 1384200.0 2076600.0 ;
      RECT  1374000.0 2090400.0 1384200.0 2076600.0 ;
      RECT  1374000.0 2090400.0 1384200.0 2104200.0 ;
      RECT  1374000.0 2118000.0 1384200.0 2104200.0 ;
      RECT  1374000.0 2118000.0 1384200.0 2131800.0 ;
      RECT  1374000.0 2145600.0 1384200.0 2131800.0 ;
      RECT  1384200.0 379200.0 1394400.0 393000.0 ;
      RECT  1384200.0 406800.0 1394400.0 393000.0 ;
      RECT  1384200.0 406800.0 1394400.0 420600.0 ;
      RECT  1384200.0 434400.0 1394400.0 420600.0 ;
      RECT  1384200.0 434400.0 1394400.0 448200.0 ;
      RECT  1384200.0 462000.0 1394400.0 448200.0 ;
      RECT  1384200.0 462000.0 1394400.0 475800.0 ;
      RECT  1384200.0 489600.0 1394400.0 475800.0 ;
      RECT  1384200.0 489600.0 1394400.0 503400.0 ;
      RECT  1384200.0 517200.0 1394400.0 503400.0 ;
      RECT  1384200.0 517200.0 1394400.0 531000.0 ;
      RECT  1384200.0 544800.0 1394400.0 531000.0 ;
      RECT  1384200.0 544800.0 1394400.0 558600.0 ;
      RECT  1384200.0 572400.0 1394400.0 558600.0 ;
      RECT  1384200.0 572400.0 1394400.0 586200.0 ;
      RECT  1384200.0 600000.0 1394400.0 586200.0 ;
      RECT  1384200.0 600000.0 1394400.0 613800.0 ;
      RECT  1384200.0 627600.0 1394400.0 613800.0 ;
      RECT  1384200.0 627600.0 1394400.0 641400.0 ;
      RECT  1384200.0 655200.0 1394400.0 641400.0 ;
      RECT  1384200.0 655200.0 1394400.0 669000.0 ;
      RECT  1384200.0 682800.0 1394400.0 669000.0 ;
      RECT  1384200.0 682800.0 1394400.0 696600.0 ;
      RECT  1384200.0 710400.0 1394400.0 696600.0 ;
      RECT  1384200.0 710400.0 1394400.0 724200.0 ;
      RECT  1384200.0 738000.0 1394400.0 724200.0 ;
      RECT  1384200.0 738000.0 1394400.0 751800.0 ;
      RECT  1384200.0 765600.0 1394400.0 751800.0 ;
      RECT  1384200.0 765600.0 1394400.0 779400.0 ;
      RECT  1384200.0 793200.0 1394400.0 779400.0 ;
      RECT  1384200.0 793200.0 1394400.0 807000.0 ;
      RECT  1384200.0 820800.0 1394400.0 807000.0 ;
      RECT  1384200.0 820800.0 1394400.0 834600.0 ;
      RECT  1384200.0 848400.0 1394400.0 834600.0 ;
      RECT  1384200.0 848400.0 1394400.0 862200.0 ;
      RECT  1384200.0 876000.0 1394400.0 862200.0 ;
      RECT  1384200.0 876000.0 1394400.0 889800.0 ;
      RECT  1384200.0 903600.0 1394400.0 889800.0 ;
      RECT  1384200.0 903600.0 1394400.0 917400.0 ;
      RECT  1384200.0 931200.0 1394400.0 917400.0 ;
      RECT  1384200.0 931200.0 1394400.0 945000.0 ;
      RECT  1384200.0 958800.0 1394400.0 945000.0 ;
      RECT  1384200.0 958800.0 1394400.0 972600.0 ;
      RECT  1384200.0 986400.0 1394400.0 972600.0 ;
      RECT  1384200.0 986400.0 1394400.0 1000200.0 ;
      RECT  1384200.0 1014000.0 1394400.0 1000200.0 ;
      RECT  1384200.0 1014000.0 1394400.0 1027800.0 ;
      RECT  1384200.0 1041600.0 1394400.0 1027800.0 ;
      RECT  1384200.0 1041600.0 1394400.0 1055400.0 ;
      RECT  1384200.0 1069200.0 1394400.0 1055400.0 ;
      RECT  1384200.0 1069200.0 1394400.0 1083000.0 ;
      RECT  1384200.0 1096800.0 1394400.0 1083000.0 ;
      RECT  1384200.0 1096800.0 1394400.0 1110600.0 ;
      RECT  1384200.0 1124400.0 1394400.0 1110600.0 ;
      RECT  1384200.0 1124400.0 1394400.0 1138200.0 ;
      RECT  1384200.0 1152000.0 1394400.0 1138200.0 ;
      RECT  1384200.0 1152000.0 1394400.0 1165800.0 ;
      RECT  1384200.0 1179600.0 1394400.0 1165800.0 ;
      RECT  1384200.0 1179600.0 1394400.0 1193400.0 ;
      RECT  1384200.0 1207200.0 1394400.0 1193400.0 ;
      RECT  1384200.0 1207200.0 1394400.0 1221000.0 ;
      RECT  1384200.0 1234800.0 1394400.0 1221000.0 ;
      RECT  1384200.0 1234800.0 1394400.0 1248600.0 ;
      RECT  1384200.0 1262400.0 1394400.0 1248600.0 ;
      RECT  1384200.0 1262400.0 1394400.0 1276200.0 ;
      RECT  1384200.0 1290000.0 1394400.0 1276200.0 ;
      RECT  1384200.0 1290000.0 1394400.0 1303800.0 ;
      RECT  1384200.0 1317600.0 1394400.0 1303800.0 ;
      RECT  1384200.0 1317600.0 1394400.0 1331400.0 ;
      RECT  1384200.0 1345200.0 1394400.0 1331400.0 ;
      RECT  1384200.0 1345200.0 1394400.0 1359000.0 ;
      RECT  1384200.0 1372800.0 1394400.0 1359000.0 ;
      RECT  1384200.0 1372800.0 1394400.0 1386600.0 ;
      RECT  1384200.0 1400400.0 1394400.0 1386600.0 ;
      RECT  1384200.0 1400400.0 1394400.0 1414200.0 ;
      RECT  1384200.0 1428000.0 1394400.0 1414200.0 ;
      RECT  1384200.0 1428000.0 1394400.0 1441800.0 ;
      RECT  1384200.0 1455600.0 1394400.0 1441800.0 ;
      RECT  1384200.0 1455600.0 1394400.0 1469400.0 ;
      RECT  1384200.0 1483200.0 1394400.0 1469400.0 ;
      RECT  1384200.0 1483200.0 1394400.0 1497000.0 ;
      RECT  1384200.0 1510800.0 1394400.0 1497000.0 ;
      RECT  1384200.0 1510800.0 1394400.0 1524600.0 ;
      RECT  1384200.0 1538400.0 1394400.0 1524600.0 ;
      RECT  1384200.0 1538400.0 1394400.0 1552200.0 ;
      RECT  1384200.0 1566000.0 1394400.0 1552200.0 ;
      RECT  1384200.0 1566000.0 1394400.0 1579800.0 ;
      RECT  1384200.0 1593600.0 1394400.0 1579800.0 ;
      RECT  1384200.0 1593600.0 1394400.0 1607400.0 ;
      RECT  1384200.0 1621200.0 1394400.0 1607400.0 ;
      RECT  1384200.0 1621200.0 1394400.0 1635000.0 ;
      RECT  1384200.0 1648800.0 1394400.0 1635000.0 ;
      RECT  1384200.0 1648800.0 1394400.0 1662600.0 ;
      RECT  1384200.0 1676400.0 1394400.0 1662600.0 ;
      RECT  1384200.0 1676400.0 1394400.0 1690200.0 ;
      RECT  1384200.0 1704000.0 1394400.0 1690200.0 ;
      RECT  1384200.0 1704000.0 1394400.0 1717800.0 ;
      RECT  1384200.0 1731600.0 1394400.0 1717800.0 ;
      RECT  1384200.0 1731600.0 1394400.0 1745400.0 ;
      RECT  1384200.0 1759200.0 1394400.0 1745400.0 ;
      RECT  1384200.0 1759200.0 1394400.0 1773000.0 ;
      RECT  1384200.0 1786800.0 1394400.0 1773000.0 ;
      RECT  1384200.0 1786800.0 1394400.0 1800600.0 ;
      RECT  1384200.0 1814400.0 1394400.0 1800600.0 ;
      RECT  1384200.0 1814400.0 1394400.0 1828200.0 ;
      RECT  1384200.0 1842000.0 1394400.0 1828200.0 ;
      RECT  1384200.0 1842000.0 1394400.0 1855800.0 ;
      RECT  1384200.0 1869600.0 1394400.0 1855800.0 ;
      RECT  1384200.0 1869600.0 1394400.0 1883400.0 ;
      RECT  1384200.0 1897200.0 1394400.0 1883400.0 ;
      RECT  1384200.0 1897200.0 1394400.0 1911000.0 ;
      RECT  1384200.0 1924800.0 1394400.0 1911000.0 ;
      RECT  1384200.0 1924800.0 1394400.0 1938600.0 ;
      RECT  1384200.0 1952400.0 1394400.0 1938600.0 ;
      RECT  1384200.0 1952400.0 1394400.0 1966200.0 ;
      RECT  1384200.0 1980000.0 1394400.0 1966200.0 ;
      RECT  1384200.0 1980000.0 1394400.0 1993800.0 ;
      RECT  1384200.0 2007600.0 1394400.0 1993800.0 ;
      RECT  1384200.0 2007600.0 1394400.0 2021400.0 ;
      RECT  1384200.0 2035200.0 1394400.0 2021400.0 ;
      RECT  1384200.0 2035200.0 1394400.0 2049000.0 ;
      RECT  1384200.0 2062800.0 1394400.0 2049000.0 ;
      RECT  1384200.0 2062800.0 1394400.0 2076600.0 ;
      RECT  1384200.0 2090400.0 1394400.0 2076600.0 ;
      RECT  1384200.0 2090400.0 1394400.0 2104200.0 ;
      RECT  1384200.0 2118000.0 1394400.0 2104200.0 ;
      RECT  1384200.0 2118000.0 1394400.0 2131800.0 ;
      RECT  1384200.0 2145600.0 1394400.0 2131800.0 ;
      RECT  1394400.0 379200.0 1404600.0 393000.0 ;
      RECT  1394400.0 406800.0 1404600.0 393000.0 ;
      RECT  1394400.0 406800.0 1404600.0 420600.0 ;
      RECT  1394400.0 434400.0 1404600.0 420600.0 ;
      RECT  1394400.0 434400.0 1404600.0 448200.0 ;
      RECT  1394400.0 462000.0 1404600.0 448200.0 ;
      RECT  1394400.0 462000.0 1404600.0 475800.0 ;
      RECT  1394400.0 489600.0 1404600.0 475800.0 ;
      RECT  1394400.0 489600.0 1404600.0 503400.0 ;
      RECT  1394400.0 517200.0 1404600.0 503400.0 ;
      RECT  1394400.0 517200.0 1404600.0 531000.0 ;
      RECT  1394400.0 544800.0 1404600.0 531000.0 ;
      RECT  1394400.0 544800.0 1404600.0 558600.0 ;
      RECT  1394400.0 572400.0 1404600.0 558600.0 ;
      RECT  1394400.0 572400.0 1404600.0 586200.0 ;
      RECT  1394400.0 600000.0 1404600.0 586200.0 ;
      RECT  1394400.0 600000.0 1404600.0 613800.0 ;
      RECT  1394400.0 627600.0 1404600.0 613800.0 ;
      RECT  1394400.0 627600.0 1404600.0 641400.0 ;
      RECT  1394400.0 655200.0 1404600.0 641400.0 ;
      RECT  1394400.0 655200.0 1404600.0 669000.0 ;
      RECT  1394400.0 682800.0 1404600.0 669000.0 ;
      RECT  1394400.0 682800.0 1404600.0 696600.0 ;
      RECT  1394400.0 710400.0 1404600.0 696600.0 ;
      RECT  1394400.0 710400.0 1404600.0 724200.0 ;
      RECT  1394400.0 738000.0 1404600.0 724200.0 ;
      RECT  1394400.0 738000.0 1404600.0 751800.0 ;
      RECT  1394400.0 765600.0 1404600.0 751800.0 ;
      RECT  1394400.0 765600.0 1404600.0 779400.0 ;
      RECT  1394400.0 793200.0 1404600.0 779400.0 ;
      RECT  1394400.0 793200.0 1404600.0 807000.0 ;
      RECT  1394400.0 820800.0 1404600.0 807000.0 ;
      RECT  1394400.0 820800.0 1404600.0 834600.0 ;
      RECT  1394400.0 848400.0 1404600.0 834600.0 ;
      RECT  1394400.0 848400.0 1404600.0 862200.0 ;
      RECT  1394400.0 876000.0 1404600.0 862200.0 ;
      RECT  1394400.0 876000.0 1404600.0 889800.0 ;
      RECT  1394400.0 903600.0 1404600.0 889800.0 ;
      RECT  1394400.0 903600.0 1404600.0 917400.0 ;
      RECT  1394400.0 931200.0 1404600.0 917400.0 ;
      RECT  1394400.0 931200.0 1404600.0 945000.0 ;
      RECT  1394400.0 958800.0 1404600.0 945000.0 ;
      RECT  1394400.0 958800.0 1404600.0 972600.0 ;
      RECT  1394400.0 986400.0 1404600.0 972600.0 ;
      RECT  1394400.0 986400.0 1404600.0 1000200.0 ;
      RECT  1394400.0 1014000.0 1404600.0 1000200.0 ;
      RECT  1394400.0 1014000.0 1404600.0 1027800.0 ;
      RECT  1394400.0 1041600.0 1404600.0 1027800.0 ;
      RECT  1394400.0 1041600.0 1404600.0 1055400.0 ;
      RECT  1394400.0 1069200.0 1404600.0 1055400.0 ;
      RECT  1394400.0 1069200.0 1404600.0 1083000.0 ;
      RECT  1394400.0 1096800.0 1404600.0 1083000.0 ;
      RECT  1394400.0 1096800.0 1404600.0 1110600.0 ;
      RECT  1394400.0 1124400.0 1404600.0 1110600.0 ;
      RECT  1394400.0 1124400.0 1404600.0 1138200.0 ;
      RECT  1394400.0 1152000.0 1404600.0 1138200.0 ;
      RECT  1394400.0 1152000.0 1404600.0 1165800.0 ;
      RECT  1394400.0 1179600.0 1404600.0 1165800.0 ;
      RECT  1394400.0 1179600.0 1404600.0 1193400.0 ;
      RECT  1394400.0 1207200.0 1404600.0 1193400.0 ;
      RECT  1394400.0 1207200.0 1404600.0 1221000.0 ;
      RECT  1394400.0 1234800.0 1404600.0 1221000.0 ;
      RECT  1394400.0 1234800.0 1404600.0 1248600.0 ;
      RECT  1394400.0 1262400.0 1404600.0 1248600.0 ;
      RECT  1394400.0 1262400.0 1404600.0 1276200.0 ;
      RECT  1394400.0 1290000.0 1404600.0 1276200.0 ;
      RECT  1394400.0 1290000.0 1404600.0 1303800.0 ;
      RECT  1394400.0 1317600.0 1404600.0 1303800.0 ;
      RECT  1394400.0 1317600.0 1404600.0 1331400.0 ;
      RECT  1394400.0 1345200.0 1404600.0 1331400.0 ;
      RECT  1394400.0 1345200.0 1404600.0 1359000.0 ;
      RECT  1394400.0 1372800.0 1404600.0 1359000.0 ;
      RECT  1394400.0 1372800.0 1404600.0 1386600.0 ;
      RECT  1394400.0 1400400.0 1404600.0 1386600.0 ;
      RECT  1394400.0 1400400.0 1404600.0 1414200.0 ;
      RECT  1394400.0 1428000.0 1404600.0 1414200.0 ;
      RECT  1394400.0 1428000.0 1404600.0 1441800.0 ;
      RECT  1394400.0 1455600.0 1404600.0 1441800.0 ;
      RECT  1394400.0 1455600.0 1404600.0 1469400.0 ;
      RECT  1394400.0 1483200.0 1404600.0 1469400.0 ;
      RECT  1394400.0 1483200.0 1404600.0 1497000.0 ;
      RECT  1394400.0 1510800.0 1404600.0 1497000.0 ;
      RECT  1394400.0 1510800.0 1404600.0 1524600.0 ;
      RECT  1394400.0 1538400.0 1404600.0 1524600.0 ;
      RECT  1394400.0 1538400.0 1404600.0 1552200.0 ;
      RECT  1394400.0 1566000.0 1404600.0 1552200.0 ;
      RECT  1394400.0 1566000.0 1404600.0 1579800.0 ;
      RECT  1394400.0 1593600.0 1404600.0 1579800.0 ;
      RECT  1394400.0 1593600.0 1404600.0 1607400.0 ;
      RECT  1394400.0 1621200.0 1404600.0 1607400.0 ;
      RECT  1394400.0 1621200.0 1404600.0 1635000.0 ;
      RECT  1394400.0 1648800.0 1404600.0 1635000.0 ;
      RECT  1394400.0 1648800.0 1404600.0 1662600.0 ;
      RECT  1394400.0 1676400.0 1404600.0 1662600.0 ;
      RECT  1394400.0 1676400.0 1404600.0 1690200.0 ;
      RECT  1394400.0 1704000.0 1404600.0 1690200.0 ;
      RECT  1394400.0 1704000.0 1404600.0 1717800.0 ;
      RECT  1394400.0 1731600.0 1404600.0 1717800.0 ;
      RECT  1394400.0 1731600.0 1404600.0 1745400.0 ;
      RECT  1394400.0 1759200.0 1404600.0 1745400.0 ;
      RECT  1394400.0 1759200.0 1404600.0 1773000.0 ;
      RECT  1394400.0 1786800.0 1404600.0 1773000.0 ;
      RECT  1394400.0 1786800.0 1404600.0 1800600.0 ;
      RECT  1394400.0 1814400.0 1404600.0 1800600.0 ;
      RECT  1394400.0 1814400.0 1404600.0 1828200.0 ;
      RECT  1394400.0 1842000.0 1404600.0 1828200.0 ;
      RECT  1394400.0 1842000.0 1404600.0 1855800.0 ;
      RECT  1394400.0 1869600.0 1404600.0 1855800.0 ;
      RECT  1394400.0 1869600.0 1404600.0 1883400.0 ;
      RECT  1394400.0 1897200.0 1404600.0 1883400.0 ;
      RECT  1394400.0 1897200.0 1404600.0 1911000.0 ;
      RECT  1394400.0 1924800.0 1404600.0 1911000.0 ;
      RECT  1394400.0 1924800.0 1404600.0 1938600.0 ;
      RECT  1394400.0 1952400.0 1404600.0 1938600.0 ;
      RECT  1394400.0 1952400.0 1404600.0 1966200.0 ;
      RECT  1394400.0 1980000.0 1404600.0 1966200.0 ;
      RECT  1394400.0 1980000.0 1404600.0 1993800.0 ;
      RECT  1394400.0 2007600.0 1404600.0 1993800.0 ;
      RECT  1394400.0 2007600.0 1404600.0 2021400.0 ;
      RECT  1394400.0 2035200.0 1404600.0 2021400.0 ;
      RECT  1394400.0 2035200.0 1404600.0 2049000.0 ;
      RECT  1394400.0 2062800.0 1404600.0 2049000.0 ;
      RECT  1394400.0 2062800.0 1404600.0 2076600.0 ;
      RECT  1394400.0 2090400.0 1404600.0 2076600.0 ;
      RECT  1394400.0 2090400.0 1404600.0 2104200.0 ;
      RECT  1394400.0 2118000.0 1404600.0 2104200.0 ;
      RECT  1394400.0 2118000.0 1404600.0 2131800.0 ;
      RECT  1394400.0 2145600.0 1404600.0 2131800.0 ;
      RECT  1404600.0 379200.0 1414800.0 393000.0 ;
      RECT  1404600.0 406800.0 1414800.0 393000.0 ;
      RECT  1404600.0 406800.0 1414800.0 420600.0 ;
      RECT  1404600.0 434400.0 1414800.0 420600.0 ;
      RECT  1404600.0 434400.0 1414800.0 448200.0 ;
      RECT  1404600.0 462000.0 1414800.0 448200.0 ;
      RECT  1404600.0 462000.0 1414800.0 475800.0 ;
      RECT  1404600.0 489600.0 1414800.0 475800.0 ;
      RECT  1404600.0 489600.0 1414800.0 503400.0 ;
      RECT  1404600.0 517200.0 1414800.0 503400.0 ;
      RECT  1404600.0 517200.0 1414800.0 531000.0 ;
      RECT  1404600.0 544800.0 1414800.0 531000.0 ;
      RECT  1404600.0 544800.0 1414800.0 558600.0 ;
      RECT  1404600.0 572400.0 1414800.0 558600.0 ;
      RECT  1404600.0 572400.0 1414800.0 586200.0 ;
      RECT  1404600.0 600000.0 1414800.0 586200.0 ;
      RECT  1404600.0 600000.0 1414800.0 613800.0 ;
      RECT  1404600.0 627600.0 1414800.0 613800.0 ;
      RECT  1404600.0 627600.0 1414800.0 641400.0 ;
      RECT  1404600.0 655200.0 1414800.0 641400.0 ;
      RECT  1404600.0 655200.0 1414800.0 669000.0 ;
      RECT  1404600.0 682800.0 1414800.0 669000.0 ;
      RECT  1404600.0 682800.0 1414800.0 696600.0 ;
      RECT  1404600.0 710400.0 1414800.0 696600.0 ;
      RECT  1404600.0 710400.0 1414800.0 724200.0 ;
      RECT  1404600.0 738000.0 1414800.0 724200.0 ;
      RECT  1404600.0 738000.0 1414800.0 751800.0 ;
      RECT  1404600.0 765600.0 1414800.0 751800.0 ;
      RECT  1404600.0 765600.0 1414800.0 779400.0 ;
      RECT  1404600.0 793200.0 1414800.0 779400.0 ;
      RECT  1404600.0 793200.0 1414800.0 807000.0 ;
      RECT  1404600.0 820800.0 1414800.0 807000.0 ;
      RECT  1404600.0 820800.0 1414800.0 834600.0 ;
      RECT  1404600.0 848400.0 1414800.0 834600.0 ;
      RECT  1404600.0 848400.0 1414800.0 862200.0 ;
      RECT  1404600.0 876000.0 1414800.0 862200.0 ;
      RECT  1404600.0 876000.0 1414800.0 889800.0 ;
      RECT  1404600.0 903600.0 1414800.0 889800.0 ;
      RECT  1404600.0 903600.0 1414800.0 917400.0 ;
      RECT  1404600.0 931200.0 1414800.0 917400.0 ;
      RECT  1404600.0 931200.0 1414800.0 945000.0 ;
      RECT  1404600.0 958800.0 1414800.0 945000.0 ;
      RECT  1404600.0 958800.0 1414800.0 972600.0 ;
      RECT  1404600.0 986400.0 1414800.0 972600.0 ;
      RECT  1404600.0 986400.0 1414800.0 1000200.0 ;
      RECT  1404600.0 1014000.0 1414800.0 1000200.0 ;
      RECT  1404600.0 1014000.0 1414800.0 1027800.0 ;
      RECT  1404600.0 1041600.0 1414800.0 1027800.0 ;
      RECT  1404600.0 1041600.0 1414800.0 1055400.0 ;
      RECT  1404600.0 1069200.0 1414800.0 1055400.0 ;
      RECT  1404600.0 1069200.0 1414800.0 1083000.0 ;
      RECT  1404600.0 1096800.0 1414800.0 1083000.0 ;
      RECT  1404600.0 1096800.0 1414800.0 1110600.0 ;
      RECT  1404600.0 1124400.0 1414800.0 1110600.0 ;
      RECT  1404600.0 1124400.0 1414800.0 1138200.0 ;
      RECT  1404600.0 1152000.0 1414800.0 1138200.0 ;
      RECT  1404600.0 1152000.0 1414800.0 1165800.0 ;
      RECT  1404600.0 1179600.0 1414800.0 1165800.0 ;
      RECT  1404600.0 1179600.0 1414800.0 1193400.0 ;
      RECT  1404600.0 1207200.0 1414800.0 1193400.0 ;
      RECT  1404600.0 1207200.0 1414800.0 1221000.0 ;
      RECT  1404600.0 1234800.0 1414800.0 1221000.0 ;
      RECT  1404600.0 1234800.0 1414800.0 1248600.0 ;
      RECT  1404600.0 1262400.0 1414800.0 1248600.0 ;
      RECT  1404600.0 1262400.0 1414800.0 1276200.0 ;
      RECT  1404600.0 1290000.0 1414800.0 1276200.0 ;
      RECT  1404600.0 1290000.0 1414800.0 1303800.0 ;
      RECT  1404600.0 1317600.0 1414800.0 1303800.0 ;
      RECT  1404600.0 1317600.0 1414800.0 1331400.0 ;
      RECT  1404600.0 1345200.0 1414800.0 1331400.0 ;
      RECT  1404600.0 1345200.0 1414800.0 1359000.0 ;
      RECT  1404600.0 1372800.0 1414800.0 1359000.0 ;
      RECT  1404600.0 1372800.0 1414800.0 1386600.0 ;
      RECT  1404600.0 1400400.0 1414800.0 1386600.0 ;
      RECT  1404600.0 1400400.0 1414800.0 1414200.0 ;
      RECT  1404600.0 1428000.0 1414800.0 1414200.0 ;
      RECT  1404600.0 1428000.0 1414800.0 1441800.0 ;
      RECT  1404600.0 1455600.0 1414800.0 1441800.0 ;
      RECT  1404600.0 1455600.0 1414800.0 1469400.0 ;
      RECT  1404600.0 1483200.0 1414800.0 1469400.0 ;
      RECT  1404600.0 1483200.0 1414800.0 1497000.0 ;
      RECT  1404600.0 1510800.0 1414800.0 1497000.0 ;
      RECT  1404600.0 1510800.0 1414800.0 1524600.0 ;
      RECT  1404600.0 1538400.0 1414800.0 1524600.0 ;
      RECT  1404600.0 1538400.0 1414800.0 1552200.0 ;
      RECT  1404600.0 1566000.0 1414800.0 1552200.0 ;
      RECT  1404600.0 1566000.0 1414800.0 1579800.0 ;
      RECT  1404600.0 1593600.0 1414800.0 1579800.0 ;
      RECT  1404600.0 1593600.0 1414800.0 1607400.0 ;
      RECT  1404600.0 1621200.0 1414800.0 1607400.0 ;
      RECT  1404600.0 1621200.0 1414800.0 1635000.0 ;
      RECT  1404600.0 1648800.0 1414800.0 1635000.0 ;
      RECT  1404600.0 1648800.0 1414800.0 1662600.0 ;
      RECT  1404600.0 1676400.0 1414800.0 1662600.0 ;
      RECT  1404600.0 1676400.0 1414800.0 1690200.0 ;
      RECT  1404600.0 1704000.0 1414800.0 1690200.0 ;
      RECT  1404600.0 1704000.0 1414800.0 1717800.0 ;
      RECT  1404600.0 1731600.0 1414800.0 1717800.0 ;
      RECT  1404600.0 1731600.0 1414800.0 1745400.0 ;
      RECT  1404600.0 1759200.0 1414800.0 1745400.0 ;
      RECT  1404600.0 1759200.0 1414800.0 1773000.0 ;
      RECT  1404600.0 1786800.0 1414800.0 1773000.0 ;
      RECT  1404600.0 1786800.0 1414800.0 1800600.0 ;
      RECT  1404600.0 1814400.0 1414800.0 1800600.0 ;
      RECT  1404600.0 1814400.0 1414800.0 1828200.0 ;
      RECT  1404600.0 1842000.0 1414800.0 1828200.0 ;
      RECT  1404600.0 1842000.0 1414800.0 1855800.0 ;
      RECT  1404600.0 1869600.0 1414800.0 1855800.0 ;
      RECT  1404600.0 1869600.0 1414800.0 1883400.0 ;
      RECT  1404600.0 1897200.0 1414800.0 1883400.0 ;
      RECT  1404600.0 1897200.0 1414800.0 1911000.0 ;
      RECT  1404600.0 1924800.0 1414800.0 1911000.0 ;
      RECT  1404600.0 1924800.0 1414800.0 1938600.0 ;
      RECT  1404600.0 1952400.0 1414800.0 1938600.0 ;
      RECT  1404600.0 1952400.0 1414800.0 1966200.0 ;
      RECT  1404600.0 1980000.0 1414800.0 1966200.0 ;
      RECT  1404600.0 1980000.0 1414800.0 1993800.0 ;
      RECT  1404600.0 2007600.0 1414800.0 1993800.0 ;
      RECT  1404600.0 2007600.0 1414800.0 2021400.0 ;
      RECT  1404600.0 2035200.0 1414800.0 2021400.0 ;
      RECT  1404600.0 2035200.0 1414800.0 2049000.0 ;
      RECT  1404600.0 2062800.0 1414800.0 2049000.0 ;
      RECT  1404600.0 2062800.0 1414800.0 2076600.0 ;
      RECT  1404600.0 2090400.0 1414800.0 2076600.0 ;
      RECT  1404600.0 2090400.0 1414800.0 2104200.0 ;
      RECT  1404600.0 2118000.0 1414800.0 2104200.0 ;
      RECT  1404600.0 2118000.0 1414800.0 2131800.0 ;
      RECT  1404600.0 2145600.0 1414800.0 2131800.0 ;
      RECT  1414800.0 379200.0 1425000.0 393000.0 ;
      RECT  1414800.0 406800.0 1425000.0 393000.0 ;
      RECT  1414800.0 406800.0 1425000.0 420600.0 ;
      RECT  1414800.0 434400.0 1425000.0 420600.0 ;
      RECT  1414800.0 434400.0 1425000.0 448200.0 ;
      RECT  1414800.0 462000.0 1425000.0 448200.0 ;
      RECT  1414800.0 462000.0 1425000.0 475800.0 ;
      RECT  1414800.0 489600.0 1425000.0 475800.0 ;
      RECT  1414800.0 489600.0 1425000.0 503400.0 ;
      RECT  1414800.0 517200.0 1425000.0 503400.0 ;
      RECT  1414800.0 517200.0 1425000.0 531000.0 ;
      RECT  1414800.0 544800.0 1425000.0 531000.0 ;
      RECT  1414800.0 544800.0 1425000.0 558600.0 ;
      RECT  1414800.0 572400.0 1425000.0 558600.0 ;
      RECT  1414800.0 572400.0 1425000.0 586200.0 ;
      RECT  1414800.0 600000.0 1425000.0 586200.0 ;
      RECT  1414800.0 600000.0 1425000.0 613800.0 ;
      RECT  1414800.0 627600.0 1425000.0 613800.0 ;
      RECT  1414800.0 627600.0 1425000.0 641400.0 ;
      RECT  1414800.0 655200.0 1425000.0 641400.0 ;
      RECT  1414800.0 655200.0 1425000.0 669000.0 ;
      RECT  1414800.0 682800.0 1425000.0 669000.0 ;
      RECT  1414800.0 682800.0 1425000.0 696600.0 ;
      RECT  1414800.0 710400.0 1425000.0 696600.0 ;
      RECT  1414800.0 710400.0 1425000.0 724200.0 ;
      RECT  1414800.0 738000.0 1425000.0 724200.0 ;
      RECT  1414800.0 738000.0 1425000.0 751800.0 ;
      RECT  1414800.0 765600.0 1425000.0 751800.0 ;
      RECT  1414800.0 765600.0 1425000.0 779400.0 ;
      RECT  1414800.0 793200.0 1425000.0 779400.0 ;
      RECT  1414800.0 793200.0 1425000.0 807000.0 ;
      RECT  1414800.0 820800.0 1425000.0 807000.0 ;
      RECT  1414800.0 820800.0 1425000.0 834600.0 ;
      RECT  1414800.0 848400.0 1425000.0 834600.0 ;
      RECT  1414800.0 848400.0 1425000.0 862200.0 ;
      RECT  1414800.0 876000.0 1425000.0 862200.0 ;
      RECT  1414800.0 876000.0 1425000.0 889800.0 ;
      RECT  1414800.0 903600.0 1425000.0 889800.0 ;
      RECT  1414800.0 903600.0 1425000.0 917400.0 ;
      RECT  1414800.0 931200.0 1425000.0 917400.0 ;
      RECT  1414800.0 931200.0 1425000.0 945000.0 ;
      RECT  1414800.0 958800.0 1425000.0 945000.0 ;
      RECT  1414800.0 958800.0 1425000.0 972600.0 ;
      RECT  1414800.0 986400.0 1425000.0 972600.0 ;
      RECT  1414800.0 986400.0 1425000.0 1000200.0 ;
      RECT  1414800.0 1014000.0 1425000.0 1000200.0 ;
      RECT  1414800.0 1014000.0 1425000.0 1027800.0 ;
      RECT  1414800.0 1041600.0 1425000.0 1027800.0 ;
      RECT  1414800.0 1041600.0 1425000.0 1055400.0 ;
      RECT  1414800.0 1069200.0 1425000.0 1055400.0 ;
      RECT  1414800.0 1069200.0 1425000.0 1083000.0 ;
      RECT  1414800.0 1096800.0 1425000.0 1083000.0 ;
      RECT  1414800.0 1096800.0 1425000.0 1110600.0 ;
      RECT  1414800.0 1124400.0 1425000.0 1110600.0 ;
      RECT  1414800.0 1124400.0 1425000.0 1138200.0 ;
      RECT  1414800.0 1152000.0 1425000.0 1138200.0 ;
      RECT  1414800.0 1152000.0 1425000.0 1165800.0 ;
      RECT  1414800.0 1179600.0 1425000.0 1165800.0 ;
      RECT  1414800.0 1179600.0 1425000.0 1193400.0 ;
      RECT  1414800.0 1207200.0 1425000.0 1193400.0 ;
      RECT  1414800.0 1207200.0 1425000.0 1221000.0 ;
      RECT  1414800.0 1234800.0 1425000.0 1221000.0 ;
      RECT  1414800.0 1234800.0 1425000.0 1248600.0 ;
      RECT  1414800.0 1262400.0 1425000.0 1248600.0 ;
      RECT  1414800.0 1262400.0 1425000.0 1276200.0 ;
      RECT  1414800.0 1290000.0 1425000.0 1276200.0 ;
      RECT  1414800.0 1290000.0 1425000.0 1303800.0 ;
      RECT  1414800.0 1317600.0 1425000.0 1303800.0 ;
      RECT  1414800.0 1317600.0 1425000.0 1331400.0 ;
      RECT  1414800.0 1345200.0 1425000.0 1331400.0 ;
      RECT  1414800.0 1345200.0 1425000.0 1359000.0 ;
      RECT  1414800.0 1372800.0 1425000.0 1359000.0 ;
      RECT  1414800.0 1372800.0 1425000.0 1386600.0 ;
      RECT  1414800.0 1400400.0 1425000.0 1386600.0 ;
      RECT  1414800.0 1400400.0 1425000.0 1414200.0 ;
      RECT  1414800.0 1428000.0 1425000.0 1414200.0 ;
      RECT  1414800.0 1428000.0 1425000.0 1441800.0 ;
      RECT  1414800.0 1455600.0 1425000.0 1441800.0 ;
      RECT  1414800.0 1455600.0 1425000.0 1469400.0 ;
      RECT  1414800.0 1483200.0 1425000.0 1469400.0 ;
      RECT  1414800.0 1483200.0 1425000.0 1497000.0 ;
      RECT  1414800.0 1510800.0 1425000.0 1497000.0 ;
      RECT  1414800.0 1510800.0 1425000.0 1524600.0 ;
      RECT  1414800.0 1538400.0 1425000.0 1524600.0 ;
      RECT  1414800.0 1538400.0 1425000.0 1552200.0 ;
      RECT  1414800.0 1566000.0 1425000.0 1552200.0 ;
      RECT  1414800.0 1566000.0 1425000.0 1579800.0 ;
      RECT  1414800.0 1593600.0 1425000.0 1579800.0 ;
      RECT  1414800.0 1593600.0 1425000.0 1607400.0 ;
      RECT  1414800.0 1621200.0 1425000.0 1607400.0 ;
      RECT  1414800.0 1621200.0 1425000.0 1635000.0 ;
      RECT  1414800.0 1648800.0 1425000.0 1635000.0 ;
      RECT  1414800.0 1648800.0 1425000.0 1662600.0 ;
      RECT  1414800.0 1676400.0 1425000.0 1662600.0 ;
      RECT  1414800.0 1676400.0 1425000.0 1690200.0 ;
      RECT  1414800.0 1704000.0 1425000.0 1690200.0 ;
      RECT  1414800.0 1704000.0 1425000.0 1717800.0 ;
      RECT  1414800.0 1731600.0 1425000.0 1717800.0 ;
      RECT  1414800.0 1731600.0 1425000.0 1745400.0 ;
      RECT  1414800.0 1759200.0 1425000.0 1745400.0 ;
      RECT  1414800.0 1759200.0 1425000.0 1773000.0 ;
      RECT  1414800.0 1786800.0 1425000.0 1773000.0 ;
      RECT  1414800.0 1786800.0 1425000.0 1800600.0 ;
      RECT  1414800.0 1814400.0 1425000.0 1800600.0 ;
      RECT  1414800.0 1814400.0 1425000.0 1828200.0 ;
      RECT  1414800.0 1842000.0 1425000.0 1828200.0 ;
      RECT  1414800.0 1842000.0 1425000.0 1855800.0 ;
      RECT  1414800.0 1869600.0 1425000.0 1855800.0 ;
      RECT  1414800.0 1869600.0 1425000.0 1883400.0 ;
      RECT  1414800.0 1897200.0 1425000.0 1883400.0 ;
      RECT  1414800.0 1897200.0 1425000.0 1911000.0 ;
      RECT  1414800.0 1924800.0 1425000.0 1911000.0 ;
      RECT  1414800.0 1924800.0 1425000.0 1938600.0 ;
      RECT  1414800.0 1952400.0 1425000.0 1938600.0 ;
      RECT  1414800.0 1952400.0 1425000.0 1966200.0 ;
      RECT  1414800.0 1980000.0 1425000.0 1966200.0 ;
      RECT  1414800.0 1980000.0 1425000.0 1993800.0 ;
      RECT  1414800.0 2007600.0 1425000.0 1993800.0 ;
      RECT  1414800.0 2007600.0 1425000.0 2021400.0 ;
      RECT  1414800.0 2035200.0 1425000.0 2021400.0 ;
      RECT  1414800.0 2035200.0 1425000.0 2049000.0 ;
      RECT  1414800.0 2062800.0 1425000.0 2049000.0 ;
      RECT  1414800.0 2062800.0 1425000.0 2076600.0 ;
      RECT  1414800.0 2090400.0 1425000.0 2076600.0 ;
      RECT  1414800.0 2090400.0 1425000.0 2104200.0 ;
      RECT  1414800.0 2118000.0 1425000.0 2104200.0 ;
      RECT  1414800.0 2118000.0 1425000.0 2131800.0 ;
      RECT  1414800.0 2145600.0 1425000.0 2131800.0 ;
      RECT  1425000.0 379200.0 1435200.0 393000.0 ;
      RECT  1425000.0 406800.0 1435200.0 393000.0 ;
      RECT  1425000.0 406800.0 1435200.0 420600.0 ;
      RECT  1425000.0 434400.0 1435200.0 420600.0 ;
      RECT  1425000.0 434400.0 1435200.0 448200.0 ;
      RECT  1425000.0 462000.0 1435200.0 448200.0 ;
      RECT  1425000.0 462000.0 1435200.0 475800.0 ;
      RECT  1425000.0 489600.0 1435200.0 475800.0 ;
      RECT  1425000.0 489600.0 1435200.0 503400.0 ;
      RECT  1425000.0 517200.0 1435200.0 503400.0 ;
      RECT  1425000.0 517200.0 1435200.0 531000.0 ;
      RECT  1425000.0 544800.0 1435200.0 531000.0 ;
      RECT  1425000.0 544800.0 1435200.0 558600.0 ;
      RECT  1425000.0 572400.0 1435200.0 558600.0 ;
      RECT  1425000.0 572400.0 1435200.0 586200.0 ;
      RECT  1425000.0 600000.0 1435200.0 586200.0 ;
      RECT  1425000.0 600000.0 1435200.0 613800.0 ;
      RECT  1425000.0 627600.0 1435200.0 613800.0 ;
      RECT  1425000.0 627600.0 1435200.0 641400.0 ;
      RECT  1425000.0 655200.0 1435200.0 641400.0 ;
      RECT  1425000.0 655200.0 1435200.0 669000.0 ;
      RECT  1425000.0 682800.0 1435200.0 669000.0 ;
      RECT  1425000.0 682800.0 1435200.0 696600.0 ;
      RECT  1425000.0 710400.0 1435200.0 696600.0 ;
      RECT  1425000.0 710400.0 1435200.0 724200.0 ;
      RECT  1425000.0 738000.0 1435200.0 724200.0 ;
      RECT  1425000.0 738000.0 1435200.0 751800.0 ;
      RECT  1425000.0 765600.0 1435200.0 751800.0 ;
      RECT  1425000.0 765600.0 1435200.0 779400.0 ;
      RECT  1425000.0 793200.0 1435200.0 779400.0 ;
      RECT  1425000.0 793200.0 1435200.0 807000.0 ;
      RECT  1425000.0 820800.0 1435200.0 807000.0 ;
      RECT  1425000.0 820800.0 1435200.0 834600.0 ;
      RECT  1425000.0 848400.0 1435200.0 834600.0 ;
      RECT  1425000.0 848400.0 1435200.0 862200.0 ;
      RECT  1425000.0 876000.0 1435200.0 862200.0 ;
      RECT  1425000.0 876000.0 1435200.0 889800.0 ;
      RECT  1425000.0 903600.0 1435200.0 889800.0 ;
      RECT  1425000.0 903600.0 1435200.0 917400.0 ;
      RECT  1425000.0 931200.0 1435200.0 917400.0 ;
      RECT  1425000.0 931200.0 1435200.0 945000.0 ;
      RECT  1425000.0 958800.0 1435200.0 945000.0 ;
      RECT  1425000.0 958800.0 1435200.0 972600.0 ;
      RECT  1425000.0 986400.0 1435200.0 972600.0 ;
      RECT  1425000.0 986400.0 1435200.0 1000200.0 ;
      RECT  1425000.0 1014000.0 1435200.0 1000200.0 ;
      RECT  1425000.0 1014000.0 1435200.0 1027800.0 ;
      RECT  1425000.0 1041600.0 1435200.0 1027800.0 ;
      RECT  1425000.0 1041600.0 1435200.0 1055400.0 ;
      RECT  1425000.0 1069200.0 1435200.0 1055400.0 ;
      RECT  1425000.0 1069200.0 1435200.0 1083000.0 ;
      RECT  1425000.0 1096800.0 1435200.0 1083000.0 ;
      RECT  1425000.0 1096800.0 1435200.0 1110600.0 ;
      RECT  1425000.0 1124400.0 1435200.0 1110600.0 ;
      RECT  1425000.0 1124400.0 1435200.0 1138200.0 ;
      RECT  1425000.0 1152000.0 1435200.0 1138200.0 ;
      RECT  1425000.0 1152000.0 1435200.0 1165800.0 ;
      RECT  1425000.0 1179600.0 1435200.0 1165800.0 ;
      RECT  1425000.0 1179600.0 1435200.0 1193400.0 ;
      RECT  1425000.0 1207200.0 1435200.0 1193400.0 ;
      RECT  1425000.0 1207200.0 1435200.0 1221000.0 ;
      RECT  1425000.0 1234800.0 1435200.0 1221000.0 ;
      RECT  1425000.0 1234800.0 1435200.0 1248600.0 ;
      RECT  1425000.0 1262400.0 1435200.0 1248600.0 ;
      RECT  1425000.0 1262400.0 1435200.0 1276200.0 ;
      RECT  1425000.0 1290000.0 1435200.0 1276200.0 ;
      RECT  1425000.0 1290000.0 1435200.0 1303800.0 ;
      RECT  1425000.0 1317600.0 1435200.0 1303800.0 ;
      RECT  1425000.0 1317600.0 1435200.0 1331400.0 ;
      RECT  1425000.0 1345200.0 1435200.0 1331400.0 ;
      RECT  1425000.0 1345200.0 1435200.0 1359000.0 ;
      RECT  1425000.0 1372800.0 1435200.0 1359000.0 ;
      RECT  1425000.0 1372800.0 1435200.0 1386600.0 ;
      RECT  1425000.0 1400400.0 1435200.0 1386600.0 ;
      RECT  1425000.0 1400400.0 1435200.0 1414200.0 ;
      RECT  1425000.0 1428000.0 1435200.0 1414200.0 ;
      RECT  1425000.0 1428000.0 1435200.0 1441800.0 ;
      RECT  1425000.0 1455600.0 1435200.0 1441800.0 ;
      RECT  1425000.0 1455600.0 1435200.0 1469400.0 ;
      RECT  1425000.0 1483200.0 1435200.0 1469400.0 ;
      RECT  1425000.0 1483200.0 1435200.0 1497000.0 ;
      RECT  1425000.0 1510800.0 1435200.0 1497000.0 ;
      RECT  1425000.0 1510800.0 1435200.0 1524600.0 ;
      RECT  1425000.0 1538400.0 1435200.0 1524600.0 ;
      RECT  1425000.0 1538400.0 1435200.0 1552200.0 ;
      RECT  1425000.0 1566000.0 1435200.0 1552200.0 ;
      RECT  1425000.0 1566000.0 1435200.0 1579800.0 ;
      RECT  1425000.0 1593600.0 1435200.0 1579800.0 ;
      RECT  1425000.0 1593600.0 1435200.0 1607400.0 ;
      RECT  1425000.0 1621200.0 1435200.0 1607400.0 ;
      RECT  1425000.0 1621200.0 1435200.0 1635000.0 ;
      RECT  1425000.0 1648800.0 1435200.0 1635000.0 ;
      RECT  1425000.0 1648800.0 1435200.0 1662600.0 ;
      RECT  1425000.0 1676400.0 1435200.0 1662600.0 ;
      RECT  1425000.0 1676400.0 1435200.0 1690200.0 ;
      RECT  1425000.0 1704000.0 1435200.0 1690200.0 ;
      RECT  1425000.0 1704000.0 1435200.0 1717800.0 ;
      RECT  1425000.0 1731600.0 1435200.0 1717800.0 ;
      RECT  1425000.0 1731600.0 1435200.0 1745400.0 ;
      RECT  1425000.0 1759200.0 1435200.0 1745400.0 ;
      RECT  1425000.0 1759200.0 1435200.0 1773000.0 ;
      RECT  1425000.0 1786800.0 1435200.0 1773000.0 ;
      RECT  1425000.0 1786800.0 1435200.0 1800600.0 ;
      RECT  1425000.0 1814400.0 1435200.0 1800600.0 ;
      RECT  1425000.0 1814400.0 1435200.0 1828200.0 ;
      RECT  1425000.0 1842000.0 1435200.0 1828200.0 ;
      RECT  1425000.0 1842000.0 1435200.0 1855800.0 ;
      RECT  1425000.0 1869600.0 1435200.0 1855800.0 ;
      RECT  1425000.0 1869600.0 1435200.0 1883400.0 ;
      RECT  1425000.0 1897200.0 1435200.0 1883400.0 ;
      RECT  1425000.0 1897200.0 1435200.0 1911000.0 ;
      RECT  1425000.0 1924800.0 1435200.0 1911000.0 ;
      RECT  1425000.0 1924800.0 1435200.0 1938600.0 ;
      RECT  1425000.0 1952400.0 1435200.0 1938600.0 ;
      RECT  1425000.0 1952400.0 1435200.0 1966200.0 ;
      RECT  1425000.0 1980000.0 1435200.0 1966200.0 ;
      RECT  1425000.0 1980000.0 1435200.0 1993800.0 ;
      RECT  1425000.0 2007600.0 1435200.0 1993800.0 ;
      RECT  1425000.0 2007600.0 1435200.0 2021400.0 ;
      RECT  1425000.0 2035200.0 1435200.0 2021400.0 ;
      RECT  1425000.0 2035200.0 1435200.0 2049000.0 ;
      RECT  1425000.0 2062800.0 1435200.0 2049000.0 ;
      RECT  1425000.0 2062800.0 1435200.0 2076600.0 ;
      RECT  1425000.0 2090400.0 1435200.0 2076600.0 ;
      RECT  1425000.0 2090400.0 1435200.0 2104200.0 ;
      RECT  1425000.0 2118000.0 1435200.0 2104200.0 ;
      RECT  1425000.0 2118000.0 1435200.0 2131800.0 ;
      RECT  1425000.0 2145600.0 1435200.0 2131800.0 ;
      RECT  1435200.0 379200.0 1445400.0 393000.0 ;
      RECT  1435200.0 406800.0 1445400.0 393000.0 ;
      RECT  1435200.0 406800.0 1445400.0 420600.0 ;
      RECT  1435200.0 434400.0 1445400.0 420600.0 ;
      RECT  1435200.0 434400.0 1445400.0 448200.0 ;
      RECT  1435200.0 462000.0 1445400.0 448200.0 ;
      RECT  1435200.0 462000.0 1445400.0 475800.0 ;
      RECT  1435200.0 489600.0 1445400.0 475800.0 ;
      RECT  1435200.0 489600.0 1445400.0 503400.0 ;
      RECT  1435200.0 517200.0 1445400.0 503400.0 ;
      RECT  1435200.0 517200.0 1445400.0 531000.0 ;
      RECT  1435200.0 544800.0 1445400.0 531000.0 ;
      RECT  1435200.0 544800.0 1445400.0 558600.0 ;
      RECT  1435200.0 572400.0 1445400.0 558600.0 ;
      RECT  1435200.0 572400.0 1445400.0 586200.0 ;
      RECT  1435200.0 600000.0 1445400.0 586200.0 ;
      RECT  1435200.0 600000.0 1445400.0 613800.0 ;
      RECT  1435200.0 627600.0 1445400.0 613800.0 ;
      RECT  1435200.0 627600.0 1445400.0 641400.0 ;
      RECT  1435200.0 655200.0 1445400.0 641400.0 ;
      RECT  1435200.0 655200.0 1445400.0 669000.0 ;
      RECT  1435200.0 682800.0 1445400.0 669000.0 ;
      RECT  1435200.0 682800.0 1445400.0 696600.0 ;
      RECT  1435200.0 710400.0 1445400.0 696600.0 ;
      RECT  1435200.0 710400.0 1445400.0 724200.0 ;
      RECT  1435200.0 738000.0 1445400.0 724200.0 ;
      RECT  1435200.0 738000.0 1445400.0 751800.0 ;
      RECT  1435200.0 765600.0 1445400.0 751800.0 ;
      RECT  1435200.0 765600.0 1445400.0 779400.0 ;
      RECT  1435200.0 793200.0 1445400.0 779400.0 ;
      RECT  1435200.0 793200.0 1445400.0 807000.0 ;
      RECT  1435200.0 820800.0 1445400.0 807000.0 ;
      RECT  1435200.0 820800.0 1445400.0 834600.0 ;
      RECT  1435200.0 848400.0 1445400.0 834600.0 ;
      RECT  1435200.0 848400.0 1445400.0 862200.0 ;
      RECT  1435200.0 876000.0 1445400.0 862200.0 ;
      RECT  1435200.0 876000.0 1445400.0 889800.0 ;
      RECT  1435200.0 903600.0 1445400.0 889800.0 ;
      RECT  1435200.0 903600.0 1445400.0 917400.0 ;
      RECT  1435200.0 931200.0 1445400.0 917400.0 ;
      RECT  1435200.0 931200.0 1445400.0 945000.0 ;
      RECT  1435200.0 958800.0 1445400.0 945000.0 ;
      RECT  1435200.0 958800.0 1445400.0 972600.0 ;
      RECT  1435200.0 986400.0 1445400.0 972600.0 ;
      RECT  1435200.0 986400.0 1445400.0 1000200.0 ;
      RECT  1435200.0 1014000.0 1445400.0 1000200.0 ;
      RECT  1435200.0 1014000.0 1445400.0 1027800.0 ;
      RECT  1435200.0 1041600.0 1445400.0 1027800.0 ;
      RECT  1435200.0 1041600.0 1445400.0 1055400.0 ;
      RECT  1435200.0 1069200.0 1445400.0 1055400.0 ;
      RECT  1435200.0 1069200.0 1445400.0 1083000.0 ;
      RECT  1435200.0 1096800.0 1445400.0 1083000.0 ;
      RECT  1435200.0 1096800.0 1445400.0 1110600.0 ;
      RECT  1435200.0 1124400.0 1445400.0 1110600.0 ;
      RECT  1435200.0 1124400.0 1445400.0 1138200.0 ;
      RECT  1435200.0 1152000.0 1445400.0 1138200.0 ;
      RECT  1435200.0 1152000.0 1445400.0 1165800.0 ;
      RECT  1435200.0 1179600.0 1445400.0 1165800.0 ;
      RECT  1435200.0 1179600.0 1445400.0 1193400.0 ;
      RECT  1435200.0 1207200.0 1445400.0 1193400.0 ;
      RECT  1435200.0 1207200.0 1445400.0 1221000.0 ;
      RECT  1435200.0 1234800.0 1445400.0 1221000.0 ;
      RECT  1435200.0 1234800.0 1445400.0 1248600.0 ;
      RECT  1435200.0 1262400.0 1445400.0 1248600.0 ;
      RECT  1435200.0 1262400.0 1445400.0 1276200.0 ;
      RECT  1435200.0 1290000.0 1445400.0 1276200.0 ;
      RECT  1435200.0 1290000.0 1445400.0 1303800.0 ;
      RECT  1435200.0 1317600.0 1445400.0 1303800.0 ;
      RECT  1435200.0 1317600.0 1445400.0 1331400.0 ;
      RECT  1435200.0 1345200.0 1445400.0 1331400.0 ;
      RECT  1435200.0 1345200.0 1445400.0 1359000.0 ;
      RECT  1435200.0 1372800.0 1445400.0 1359000.0 ;
      RECT  1435200.0 1372800.0 1445400.0 1386600.0 ;
      RECT  1435200.0 1400400.0 1445400.0 1386600.0 ;
      RECT  1435200.0 1400400.0 1445400.0 1414200.0 ;
      RECT  1435200.0 1428000.0 1445400.0 1414200.0 ;
      RECT  1435200.0 1428000.0 1445400.0 1441800.0 ;
      RECT  1435200.0 1455600.0 1445400.0 1441800.0 ;
      RECT  1435200.0 1455600.0 1445400.0 1469400.0 ;
      RECT  1435200.0 1483200.0 1445400.0 1469400.0 ;
      RECT  1435200.0 1483200.0 1445400.0 1497000.0 ;
      RECT  1435200.0 1510800.0 1445400.0 1497000.0 ;
      RECT  1435200.0 1510800.0 1445400.0 1524600.0 ;
      RECT  1435200.0 1538400.0 1445400.0 1524600.0 ;
      RECT  1435200.0 1538400.0 1445400.0 1552200.0 ;
      RECT  1435200.0 1566000.0 1445400.0 1552200.0 ;
      RECT  1435200.0 1566000.0 1445400.0 1579800.0 ;
      RECT  1435200.0 1593600.0 1445400.0 1579800.0 ;
      RECT  1435200.0 1593600.0 1445400.0 1607400.0 ;
      RECT  1435200.0 1621200.0 1445400.0 1607400.0 ;
      RECT  1435200.0 1621200.0 1445400.0 1635000.0 ;
      RECT  1435200.0 1648800.0 1445400.0 1635000.0 ;
      RECT  1435200.0 1648800.0 1445400.0 1662600.0 ;
      RECT  1435200.0 1676400.0 1445400.0 1662600.0 ;
      RECT  1435200.0 1676400.0 1445400.0 1690200.0 ;
      RECT  1435200.0 1704000.0 1445400.0 1690200.0 ;
      RECT  1435200.0 1704000.0 1445400.0 1717800.0 ;
      RECT  1435200.0 1731600.0 1445400.0 1717800.0 ;
      RECT  1435200.0 1731600.0 1445400.0 1745400.0 ;
      RECT  1435200.0 1759200.0 1445400.0 1745400.0 ;
      RECT  1435200.0 1759200.0 1445400.0 1773000.0 ;
      RECT  1435200.0 1786800.0 1445400.0 1773000.0 ;
      RECT  1435200.0 1786800.0 1445400.0 1800600.0 ;
      RECT  1435200.0 1814400.0 1445400.0 1800600.0 ;
      RECT  1435200.0 1814400.0 1445400.0 1828200.0 ;
      RECT  1435200.0 1842000.0 1445400.0 1828200.0 ;
      RECT  1435200.0 1842000.0 1445400.0 1855800.0 ;
      RECT  1435200.0 1869600.0 1445400.0 1855800.0 ;
      RECT  1435200.0 1869600.0 1445400.0 1883400.0 ;
      RECT  1435200.0 1897200.0 1445400.0 1883400.0 ;
      RECT  1435200.0 1897200.0 1445400.0 1911000.0 ;
      RECT  1435200.0 1924800.0 1445400.0 1911000.0 ;
      RECT  1435200.0 1924800.0 1445400.0 1938600.0 ;
      RECT  1435200.0 1952400.0 1445400.0 1938600.0 ;
      RECT  1435200.0 1952400.0 1445400.0 1966200.0 ;
      RECT  1435200.0 1980000.0 1445400.0 1966200.0 ;
      RECT  1435200.0 1980000.0 1445400.0 1993800.0 ;
      RECT  1435200.0 2007600.0 1445400.0 1993800.0 ;
      RECT  1435200.0 2007600.0 1445400.0 2021400.0 ;
      RECT  1435200.0 2035200.0 1445400.0 2021400.0 ;
      RECT  1435200.0 2035200.0 1445400.0 2049000.0 ;
      RECT  1435200.0 2062800.0 1445400.0 2049000.0 ;
      RECT  1435200.0 2062800.0 1445400.0 2076600.0 ;
      RECT  1435200.0 2090400.0 1445400.0 2076600.0 ;
      RECT  1435200.0 2090400.0 1445400.0 2104200.0 ;
      RECT  1435200.0 2118000.0 1445400.0 2104200.0 ;
      RECT  1435200.0 2118000.0 1445400.0 2131800.0 ;
      RECT  1435200.0 2145600.0 1445400.0 2131800.0 ;
      RECT  1445400.0 379200.0 1455600.0 393000.0 ;
      RECT  1445400.0 406800.0 1455600.0 393000.0 ;
      RECT  1445400.0 406800.0 1455600.0 420600.0 ;
      RECT  1445400.0 434400.0 1455600.0 420600.0 ;
      RECT  1445400.0 434400.0 1455600.0 448200.0 ;
      RECT  1445400.0 462000.0 1455600.0 448200.0 ;
      RECT  1445400.0 462000.0 1455600.0 475800.0 ;
      RECT  1445400.0 489600.0 1455600.0 475800.0 ;
      RECT  1445400.0 489600.0 1455600.0 503400.0 ;
      RECT  1445400.0 517200.0 1455600.0 503400.0 ;
      RECT  1445400.0 517200.0 1455600.0 531000.0 ;
      RECT  1445400.0 544800.0 1455600.0 531000.0 ;
      RECT  1445400.0 544800.0 1455600.0 558600.0 ;
      RECT  1445400.0 572400.0 1455600.0 558600.0 ;
      RECT  1445400.0 572400.0 1455600.0 586200.0 ;
      RECT  1445400.0 600000.0 1455600.0 586200.0 ;
      RECT  1445400.0 600000.0 1455600.0 613800.0 ;
      RECT  1445400.0 627600.0 1455600.0 613800.0 ;
      RECT  1445400.0 627600.0 1455600.0 641400.0 ;
      RECT  1445400.0 655200.0 1455600.0 641400.0 ;
      RECT  1445400.0 655200.0 1455600.0 669000.0 ;
      RECT  1445400.0 682800.0 1455600.0 669000.0 ;
      RECT  1445400.0 682800.0 1455600.0 696600.0 ;
      RECT  1445400.0 710400.0 1455600.0 696600.0 ;
      RECT  1445400.0 710400.0 1455600.0 724200.0 ;
      RECT  1445400.0 738000.0 1455600.0 724200.0 ;
      RECT  1445400.0 738000.0 1455600.0 751800.0 ;
      RECT  1445400.0 765600.0 1455600.0 751800.0 ;
      RECT  1445400.0 765600.0 1455600.0 779400.0 ;
      RECT  1445400.0 793200.0 1455600.0 779400.0 ;
      RECT  1445400.0 793200.0 1455600.0 807000.0 ;
      RECT  1445400.0 820800.0 1455600.0 807000.0 ;
      RECT  1445400.0 820800.0 1455600.0 834600.0 ;
      RECT  1445400.0 848400.0 1455600.0 834600.0 ;
      RECT  1445400.0 848400.0 1455600.0 862200.0 ;
      RECT  1445400.0 876000.0 1455600.0 862200.0 ;
      RECT  1445400.0 876000.0 1455600.0 889800.0 ;
      RECT  1445400.0 903600.0 1455600.0 889800.0 ;
      RECT  1445400.0 903600.0 1455600.0 917400.0 ;
      RECT  1445400.0 931200.0 1455600.0 917400.0 ;
      RECT  1445400.0 931200.0 1455600.0 945000.0 ;
      RECT  1445400.0 958800.0 1455600.0 945000.0 ;
      RECT  1445400.0 958800.0 1455600.0 972600.0 ;
      RECT  1445400.0 986400.0 1455600.0 972600.0 ;
      RECT  1445400.0 986400.0 1455600.0 1000200.0 ;
      RECT  1445400.0 1014000.0 1455600.0 1000200.0 ;
      RECT  1445400.0 1014000.0 1455600.0 1027800.0 ;
      RECT  1445400.0 1041600.0 1455600.0 1027800.0 ;
      RECT  1445400.0 1041600.0 1455600.0 1055400.0 ;
      RECT  1445400.0 1069200.0 1455600.0 1055400.0 ;
      RECT  1445400.0 1069200.0 1455600.0 1083000.0 ;
      RECT  1445400.0 1096800.0 1455600.0 1083000.0 ;
      RECT  1445400.0 1096800.0 1455600.0 1110600.0 ;
      RECT  1445400.0 1124400.0 1455600.0 1110600.0 ;
      RECT  1445400.0 1124400.0 1455600.0 1138200.0 ;
      RECT  1445400.0 1152000.0 1455600.0 1138200.0 ;
      RECT  1445400.0 1152000.0 1455600.0 1165800.0 ;
      RECT  1445400.0 1179600.0 1455600.0 1165800.0 ;
      RECT  1445400.0 1179600.0 1455600.0 1193400.0 ;
      RECT  1445400.0 1207200.0 1455600.0 1193400.0 ;
      RECT  1445400.0 1207200.0 1455600.0 1221000.0 ;
      RECT  1445400.0 1234800.0 1455600.0 1221000.0 ;
      RECT  1445400.0 1234800.0 1455600.0 1248600.0 ;
      RECT  1445400.0 1262400.0 1455600.0 1248600.0 ;
      RECT  1445400.0 1262400.0 1455600.0 1276200.0 ;
      RECT  1445400.0 1290000.0 1455600.0 1276200.0 ;
      RECT  1445400.0 1290000.0 1455600.0 1303800.0 ;
      RECT  1445400.0 1317600.0 1455600.0 1303800.0 ;
      RECT  1445400.0 1317600.0 1455600.0 1331400.0 ;
      RECT  1445400.0 1345200.0 1455600.0 1331400.0 ;
      RECT  1445400.0 1345200.0 1455600.0 1359000.0 ;
      RECT  1445400.0 1372800.0 1455600.0 1359000.0 ;
      RECT  1445400.0 1372800.0 1455600.0 1386600.0 ;
      RECT  1445400.0 1400400.0 1455600.0 1386600.0 ;
      RECT  1445400.0 1400400.0 1455600.0 1414200.0 ;
      RECT  1445400.0 1428000.0 1455600.0 1414200.0 ;
      RECT  1445400.0 1428000.0 1455600.0 1441800.0 ;
      RECT  1445400.0 1455600.0 1455600.0 1441800.0 ;
      RECT  1445400.0 1455600.0 1455600.0 1469400.0 ;
      RECT  1445400.0 1483200.0 1455600.0 1469400.0 ;
      RECT  1445400.0 1483200.0 1455600.0 1497000.0 ;
      RECT  1445400.0 1510800.0 1455600.0 1497000.0 ;
      RECT  1445400.0 1510800.0 1455600.0 1524600.0 ;
      RECT  1445400.0 1538400.0 1455600.0 1524600.0 ;
      RECT  1445400.0 1538400.0 1455600.0 1552200.0 ;
      RECT  1445400.0 1566000.0 1455600.0 1552200.0 ;
      RECT  1445400.0 1566000.0 1455600.0 1579800.0 ;
      RECT  1445400.0 1593600.0 1455600.0 1579800.0 ;
      RECT  1445400.0 1593600.0 1455600.0 1607400.0 ;
      RECT  1445400.0 1621200.0 1455600.0 1607400.0 ;
      RECT  1445400.0 1621200.0 1455600.0 1635000.0 ;
      RECT  1445400.0 1648800.0 1455600.0 1635000.0 ;
      RECT  1445400.0 1648800.0 1455600.0 1662600.0 ;
      RECT  1445400.0 1676400.0 1455600.0 1662600.0 ;
      RECT  1445400.0 1676400.0 1455600.0 1690200.0 ;
      RECT  1445400.0 1704000.0 1455600.0 1690200.0 ;
      RECT  1445400.0 1704000.0 1455600.0 1717800.0 ;
      RECT  1445400.0 1731600.0 1455600.0 1717800.0 ;
      RECT  1445400.0 1731600.0 1455600.0 1745400.0 ;
      RECT  1445400.0 1759200.0 1455600.0 1745400.0 ;
      RECT  1445400.0 1759200.0 1455600.0 1773000.0 ;
      RECT  1445400.0 1786800.0 1455600.0 1773000.0 ;
      RECT  1445400.0 1786800.0 1455600.0 1800600.0 ;
      RECT  1445400.0 1814400.0 1455600.0 1800600.0 ;
      RECT  1445400.0 1814400.0 1455600.0 1828200.0 ;
      RECT  1445400.0 1842000.0 1455600.0 1828200.0 ;
      RECT  1445400.0 1842000.0 1455600.0 1855800.0 ;
      RECT  1445400.0 1869600.0 1455600.0 1855800.0 ;
      RECT  1445400.0 1869600.0 1455600.0 1883400.0 ;
      RECT  1445400.0 1897200.0 1455600.0 1883400.0 ;
      RECT  1445400.0 1897200.0 1455600.0 1911000.0 ;
      RECT  1445400.0 1924800.0 1455600.0 1911000.0 ;
      RECT  1445400.0 1924800.0 1455600.0 1938600.0 ;
      RECT  1445400.0 1952400.0 1455600.0 1938600.0 ;
      RECT  1445400.0 1952400.0 1455600.0 1966200.0 ;
      RECT  1445400.0 1980000.0 1455600.0 1966200.0 ;
      RECT  1445400.0 1980000.0 1455600.0 1993800.0 ;
      RECT  1445400.0 2007600.0 1455600.0 1993800.0 ;
      RECT  1445400.0 2007600.0 1455600.0 2021400.0 ;
      RECT  1445400.0 2035200.0 1455600.0 2021400.0 ;
      RECT  1445400.0 2035200.0 1455600.0 2049000.0 ;
      RECT  1445400.0 2062800.0 1455600.0 2049000.0 ;
      RECT  1445400.0 2062800.0 1455600.0 2076600.0 ;
      RECT  1445400.0 2090400.0 1455600.0 2076600.0 ;
      RECT  1445400.0 2090400.0 1455600.0 2104200.0 ;
      RECT  1445400.0 2118000.0 1455600.0 2104200.0 ;
      RECT  1445400.0 2118000.0 1455600.0 2131800.0 ;
      RECT  1445400.0 2145600.0 1455600.0 2131800.0 ;
      RECT  1455600.0 379200.0 1465800.0 393000.0 ;
      RECT  1455600.0 406800.0 1465800.0 393000.0 ;
      RECT  1455600.0 406800.0 1465800.0 420600.0 ;
      RECT  1455600.0 434400.0 1465800.0 420600.0 ;
      RECT  1455600.0 434400.0 1465800.0 448200.0 ;
      RECT  1455600.0 462000.0 1465800.0 448200.0 ;
      RECT  1455600.0 462000.0 1465800.0 475800.0 ;
      RECT  1455600.0 489600.0 1465800.0 475800.0 ;
      RECT  1455600.0 489600.0 1465800.0 503400.0 ;
      RECT  1455600.0 517200.0 1465800.0 503400.0 ;
      RECT  1455600.0 517200.0 1465800.0 531000.0 ;
      RECT  1455600.0 544800.0 1465800.0 531000.0 ;
      RECT  1455600.0 544800.0 1465800.0 558600.0 ;
      RECT  1455600.0 572400.0 1465800.0 558600.0 ;
      RECT  1455600.0 572400.0 1465800.0 586200.0 ;
      RECT  1455600.0 600000.0 1465800.0 586200.0 ;
      RECT  1455600.0 600000.0 1465800.0 613800.0 ;
      RECT  1455600.0 627600.0 1465800.0 613800.0 ;
      RECT  1455600.0 627600.0 1465800.0 641400.0 ;
      RECT  1455600.0 655200.0 1465800.0 641400.0 ;
      RECT  1455600.0 655200.0 1465800.0 669000.0 ;
      RECT  1455600.0 682800.0 1465800.0 669000.0 ;
      RECT  1455600.0 682800.0 1465800.0 696600.0 ;
      RECT  1455600.0 710400.0 1465800.0 696600.0 ;
      RECT  1455600.0 710400.0 1465800.0 724200.0 ;
      RECT  1455600.0 738000.0 1465800.0 724200.0 ;
      RECT  1455600.0 738000.0 1465800.0 751800.0 ;
      RECT  1455600.0 765600.0 1465800.0 751800.0 ;
      RECT  1455600.0 765600.0 1465800.0 779400.0 ;
      RECT  1455600.0 793200.0 1465800.0 779400.0 ;
      RECT  1455600.0 793200.0 1465800.0 807000.0 ;
      RECT  1455600.0 820800.0 1465800.0 807000.0 ;
      RECT  1455600.0 820800.0 1465800.0 834600.0 ;
      RECT  1455600.0 848400.0 1465800.0 834600.0 ;
      RECT  1455600.0 848400.0 1465800.0 862200.0 ;
      RECT  1455600.0 876000.0 1465800.0 862200.0 ;
      RECT  1455600.0 876000.0 1465800.0 889800.0 ;
      RECT  1455600.0 903600.0 1465800.0 889800.0 ;
      RECT  1455600.0 903600.0 1465800.0 917400.0 ;
      RECT  1455600.0 931200.0 1465800.0 917400.0 ;
      RECT  1455600.0 931200.0 1465800.0 945000.0 ;
      RECT  1455600.0 958800.0 1465800.0 945000.0 ;
      RECT  1455600.0 958800.0 1465800.0 972600.0 ;
      RECT  1455600.0 986400.0 1465800.0 972600.0 ;
      RECT  1455600.0 986400.0 1465800.0 1000200.0 ;
      RECT  1455600.0 1014000.0 1465800.0 1000200.0 ;
      RECT  1455600.0 1014000.0 1465800.0 1027800.0 ;
      RECT  1455600.0 1041600.0 1465800.0 1027800.0 ;
      RECT  1455600.0 1041600.0 1465800.0 1055400.0 ;
      RECT  1455600.0 1069200.0 1465800.0 1055400.0 ;
      RECT  1455600.0 1069200.0 1465800.0 1083000.0 ;
      RECT  1455600.0 1096800.0 1465800.0 1083000.0 ;
      RECT  1455600.0 1096800.0 1465800.0 1110600.0 ;
      RECT  1455600.0 1124400.0 1465800.0 1110600.0 ;
      RECT  1455600.0 1124400.0 1465800.0 1138200.0 ;
      RECT  1455600.0 1152000.0 1465800.0 1138200.0 ;
      RECT  1455600.0 1152000.0 1465800.0 1165800.0 ;
      RECT  1455600.0 1179600.0 1465800.0 1165800.0 ;
      RECT  1455600.0 1179600.0 1465800.0 1193400.0 ;
      RECT  1455600.0 1207200.0 1465800.0 1193400.0 ;
      RECT  1455600.0 1207200.0 1465800.0 1221000.0 ;
      RECT  1455600.0 1234800.0 1465800.0 1221000.0 ;
      RECT  1455600.0 1234800.0 1465800.0 1248600.0 ;
      RECT  1455600.0 1262400.0 1465800.0 1248600.0 ;
      RECT  1455600.0 1262400.0 1465800.0 1276200.0 ;
      RECT  1455600.0 1290000.0 1465800.0 1276200.0 ;
      RECT  1455600.0 1290000.0 1465800.0 1303800.0 ;
      RECT  1455600.0 1317600.0 1465800.0 1303800.0 ;
      RECT  1455600.0 1317600.0 1465800.0 1331400.0 ;
      RECT  1455600.0 1345200.0 1465800.0 1331400.0 ;
      RECT  1455600.0 1345200.0 1465800.0 1359000.0 ;
      RECT  1455600.0 1372800.0 1465800.0 1359000.0 ;
      RECT  1455600.0 1372800.0 1465800.0 1386600.0 ;
      RECT  1455600.0 1400400.0 1465800.0 1386600.0 ;
      RECT  1455600.0 1400400.0 1465800.0 1414200.0 ;
      RECT  1455600.0 1428000.0 1465800.0 1414200.0 ;
      RECT  1455600.0 1428000.0 1465800.0 1441800.0 ;
      RECT  1455600.0 1455600.0 1465800.0 1441800.0 ;
      RECT  1455600.0 1455600.0 1465800.0 1469400.0 ;
      RECT  1455600.0 1483200.0 1465800.0 1469400.0 ;
      RECT  1455600.0 1483200.0 1465800.0 1497000.0 ;
      RECT  1455600.0 1510800.0 1465800.0 1497000.0 ;
      RECT  1455600.0 1510800.0 1465800.0 1524600.0 ;
      RECT  1455600.0 1538400.0 1465800.0 1524600.0 ;
      RECT  1455600.0 1538400.0 1465800.0 1552200.0 ;
      RECT  1455600.0 1566000.0 1465800.0 1552200.0 ;
      RECT  1455600.0 1566000.0 1465800.0 1579800.0 ;
      RECT  1455600.0 1593600.0 1465800.0 1579800.0 ;
      RECT  1455600.0 1593600.0 1465800.0 1607400.0 ;
      RECT  1455600.0 1621200.0 1465800.0 1607400.0 ;
      RECT  1455600.0 1621200.0 1465800.0 1635000.0 ;
      RECT  1455600.0 1648800.0 1465800.0 1635000.0 ;
      RECT  1455600.0 1648800.0 1465800.0 1662600.0 ;
      RECT  1455600.0 1676400.0 1465800.0 1662600.0 ;
      RECT  1455600.0 1676400.0 1465800.0 1690200.0 ;
      RECT  1455600.0 1704000.0 1465800.0 1690200.0 ;
      RECT  1455600.0 1704000.0 1465800.0 1717800.0 ;
      RECT  1455600.0 1731600.0 1465800.0 1717800.0 ;
      RECT  1455600.0 1731600.0 1465800.0 1745400.0 ;
      RECT  1455600.0 1759200.0 1465800.0 1745400.0 ;
      RECT  1455600.0 1759200.0 1465800.0 1773000.0 ;
      RECT  1455600.0 1786800.0 1465800.0 1773000.0 ;
      RECT  1455600.0 1786800.0 1465800.0 1800600.0 ;
      RECT  1455600.0 1814400.0 1465800.0 1800600.0 ;
      RECT  1455600.0 1814400.0 1465800.0 1828200.0 ;
      RECT  1455600.0 1842000.0 1465800.0 1828200.0 ;
      RECT  1455600.0 1842000.0 1465800.0 1855800.0 ;
      RECT  1455600.0 1869600.0 1465800.0 1855800.0 ;
      RECT  1455600.0 1869600.0 1465800.0 1883400.0 ;
      RECT  1455600.0 1897200.0 1465800.0 1883400.0 ;
      RECT  1455600.0 1897200.0 1465800.0 1911000.0 ;
      RECT  1455600.0 1924800.0 1465800.0 1911000.0 ;
      RECT  1455600.0 1924800.0 1465800.0 1938600.0 ;
      RECT  1455600.0 1952400.0 1465800.0 1938600.0 ;
      RECT  1455600.0 1952400.0 1465800.0 1966200.0 ;
      RECT  1455600.0 1980000.0 1465800.0 1966200.0 ;
      RECT  1455600.0 1980000.0 1465800.0 1993800.0 ;
      RECT  1455600.0 2007600.0 1465800.0 1993800.0 ;
      RECT  1455600.0 2007600.0 1465800.0 2021400.0 ;
      RECT  1455600.0 2035200.0 1465800.0 2021400.0 ;
      RECT  1455600.0 2035200.0 1465800.0 2049000.0 ;
      RECT  1455600.0 2062800.0 1465800.0 2049000.0 ;
      RECT  1455600.0 2062800.0 1465800.0 2076600.0 ;
      RECT  1455600.0 2090400.0 1465800.0 2076600.0 ;
      RECT  1455600.0 2090400.0 1465800.0 2104200.0 ;
      RECT  1455600.0 2118000.0 1465800.0 2104200.0 ;
      RECT  1455600.0 2118000.0 1465800.0 2131800.0 ;
      RECT  1455600.0 2145600.0 1465800.0 2131800.0 ;
      RECT  1465800.0 379200.0 1476000.0 393000.0 ;
      RECT  1465800.0 406800.0 1476000.0 393000.0 ;
      RECT  1465800.0 406800.0 1476000.0 420600.0 ;
      RECT  1465800.0 434400.0 1476000.0 420600.0 ;
      RECT  1465800.0 434400.0 1476000.0 448200.0 ;
      RECT  1465800.0 462000.0 1476000.0 448200.0 ;
      RECT  1465800.0 462000.0 1476000.0 475800.0 ;
      RECT  1465800.0 489600.0 1476000.0 475800.0 ;
      RECT  1465800.0 489600.0 1476000.0 503400.0 ;
      RECT  1465800.0 517200.0 1476000.0 503400.0 ;
      RECT  1465800.0 517200.0 1476000.0 531000.0 ;
      RECT  1465800.0 544800.0 1476000.0 531000.0 ;
      RECT  1465800.0 544800.0 1476000.0 558600.0 ;
      RECT  1465800.0 572400.0 1476000.0 558600.0 ;
      RECT  1465800.0 572400.0 1476000.0 586200.0 ;
      RECT  1465800.0 600000.0 1476000.0 586200.0 ;
      RECT  1465800.0 600000.0 1476000.0 613800.0 ;
      RECT  1465800.0 627600.0 1476000.0 613800.0 ;
      RECT  1465800.0 627600.0 1476000.0 641400.0 ;
      RECT  1465800.0 655200.0 1476000.0 641400.0 ;
      RECT  1465800.0 655200.0 1476000.0 669000.0 ;
      RECT  1465800.0 682800.0 1476000.0 669000.0 ;
      RECT  1465800.0 682800.0 1476000.0 696600.0 ;
      RECT  1465800.0 710400.0 1476000.0 696600.0 ;
      RECT  1465800.0 710400.0 1476000.0 724200.0 ;
      RECT  1465800.0 738000.0 1476000.0 724200.0 ;
      RECT  1465800.0 738000.0 1476000.0 751800.0 ;
      RECT  1465800.0 765600.0 1476000.0 751800.0 ;
      RECT  1465800.0 765600.0 1476000.0 779400.0 ;
      RECT  1465800.0 793200.0 1476000.0 779400.0 ;
      RECT  1465800.0 793200.0 1476000.0 807000.0 ;
      RECT  1465800.0 820800.0 1476000.0 807000.0 ;
      RECT  1465800.0 820800.0 1476000.0 834600.0 ;
      RECT  1465800.0 848400.0 1476000.0 834600.0 ;
      RECT  1465800.0 848400.0 1476000.0 862200.0 ;
      RECT  1465800.0 876000.0 1476000.0 862200.0 ;
      RECT  1465800.0 876000.0 1476000.0 889800.0 ;
      RECT  1465800.0 903600.0 1476000.0 889800.0 ;
      RECT  1465800.0 903600.0 1476000.0 917400.0 ;
      RECT  1465800.0 931200.0 1476000.0 917400.0 ;
      RECT  1465800.0 931200.0 1476000.0 945000.0 ;
      RECT  1465800.0 958800.0 1476000.0 945000.0 ;
      RECT  1465800.0 958800.0 1476000.0 972600.0 ;
      RECT  1465800.0 986400.0 1476000.0 972600.0 ;
      RECT  1465800.0 986400.0 1476000.0 1000200.0 ;
      RECT  1465800.0 1014000.0 1476000.0 1000200.0 ;
      RECT  1465800.0 1014000.0 1476000.0 1027800.0 ;
      RECT  1465800.0 1041600.0 1476000.0 1027800.0 ;
      RECT  1465800.0 1041600.0 1476000.0 1055400.0 ;
      RECT  1465800.0 1069200.0 1476000.0 1055400.0 ;
      RECT  1465800.0 1069200.0 1476000.0 1083000.0 ;
      RECT  1465800.0 1096800.0 1476000.0 1083000.0 ;
      RECT  1465800.0 1096800.0 1476000.0 1110600.0 ;
      RECT  1465800.0 1124400.0 1476000.0 1110600.0 ;
      RECT  1465800.0 1124400.0 1476000.0 1138200.0 ;
      RECT  1465800.0 1152000.0 1476000.0 1138200.0 ;
      RECT  1465800.0 1152000.0 1476000.0 1165800.0 ;
      RECT  1465800.0 1179600.0 1476000.0 1165800.0 ;
      RECT  1465800.0 1179600.0 1476000.0 1193400.0 ;
      RECT  1465800.0 1207200.0 1476000.0 1193400.0 ;
      RECT  1465800.0 1207200.0 1476000.0 1221000.0 ;
      RECT  1465800.0 1234800.0 1476000.0 1221000.0 ;
      RECT  1465800.0 1234800.0 1476000.0 1248600.0 ;
      RECT  1465800.0 1262400.0 1476000.0 1248600.0 ;
      RECT  1465800.0 1262400.0 1476000.0 1276200.0 ;
      RECT  1465800.0 1290000.0 1476000.0 1276200.0 ;
      RECT  1465800.0 1290000.0 1476000.0 1303800.0 ;
      RECT  1465800.0 1317600.0 1476000.0 1303800.0 ;
      RECT  1465800.0 1317600.0 1476000.0 1331400.0 ;
      RECT  1465800.0 1345200.0 1476000.0 1331400.0 ;
      RECT  1465800.0 1345200.0 1476000.0 1359000.0 ;
      RECT  1465800.0 1372800.0 1476000.0 1359000.0 ;
      RECT  1465800.0 1372800.0 1476000.0 1386600.0 ;
      RECT  1465800.0 1400400.0 1476000.0 1386600.0 ;
      RECT  1465800.0 1400400.0 1476000.0 1414200.0 ;
      RECT  1465800.0 1428000.0 1476000.0 1414200.0 ;
      RECT  1465800.0 1428000.0 1476000.0 1441800.0 ;
      RECT  1465800.0 1455600.0 1476000.0 1441800.0 ;
      RECT  1465800.0 1455600.0 1476000.0 1469400.0 ;
      RECT  1465800.0 1483200.0 1476000.0 1469400.0 ;
      RECT  1465800.0 1483200.0 1476000.0 1497000.0 ;
      RECT  1465800.0 1510800.0 1476000.0 1497000.0 ;
      RECT  1465800.0 1510800.0 1476000.0 1524600.0 ;
      RECT  1465800.0 1538400.0 1476000.0 1524600.0 ;
      RECT  1465800.0 1538400.0 1476000.0 1552200.0 ;
      RECT  1465800.0 1566000.0 1476000.0 1552200.0 ;
      RECT  1465800.0 1566000.0 1476000.0 1579800.0 ;
      RECT  1465800.0 1593600.0 1476000.0 1579800.0 ;
      RECT  1465800.0 1593600.0 1476000.0 1607400.0 ;
      RECT  1465800.0 1621200.0 1476000.0 1607400.0 ;
      RECT  1465800.0 1621200.0 1476000.0 1635000.0 ;
      RECT  1465800.0 1648800.0 1476000.0 1635000.0 ;
      RECT  1465800.0 1648800.0 1476000.0 1662600.0 ;
      RECT  1465800.0 1676400.0 1476000.0 1662600.0 ;
      RECT  1465800.0 1676400.0 1476000.0 1690200.0 ;
      RECT  1465800.0 1704000.0 1476000.0 1690200.0 ;
      RECT  1465800.0 1704000.0 1476000.0 1717800.0 ;
      RECT  1465800.0 1731600.0 1476000.0 1717800.0 ;
      RECT  1465800.0 1731600.0 1476000.0 1745400.0 ;
      RECT  1465800.0 1759200.0 1476000.0 1745400.0 ;
      RECT  1465800.0 1759200.0 1476000.0 1773000.0 ;
      RECT  1465800.0 1786800.0 1476000.0 1773000.0 ;
      RECT  1465800.0 1786800.0 1476000.0 1800600.0 ;
      RECT  1465800.0 1814400.0 1476000.0 1800600.0 ;
      RECT  1465800.0 1814400.0 1476000.0 1828200.0 ;
      RECT  1465800.0 1842000.0 1476000.0 1828200.0 ;
      RECT  1465800.0 1842000.0 1476000.0 1855800.0 ;
      RECT  1465800.0 1869600.0 1476000.0 1855800.0 ;
      RECT  1465800.0 1869600.0 1476000.0 1883400.0 ;
      RECT  1465800.0 1897200.0 1476000.0 1883400.0 ;
      RECT  1465800.0 1897200.0 1476000.0 1911000.0 ;
      RECT  1465800.0 1924800.0 1476000.0 1911000.0 ;
      RECT  1465800.0 1924800.0 1476000.0 1938600.0 ;
      RECT  1465800.0 1952400.0 1476000.0 1938600.0 ;
      RECT  1465800.0 1952400.0 1476000.0 1966200.0 ;
      RECT  1465800.0 1980000.0 1476000.0 1966200.0 ;
      RECT  1465800.0 1980000.0 1476000.0 1993800.0 ;
      RECT  1465800.0 2007600.0 1476000.0 1993800.0 ;
      RECT  1465800.0 2007600.0 1476000.0 2021400.0 ;
      RECT  1465800.0 2035200.0 1476000.0 2021400.0 ;
      RECT  1465800.0 2035200.0 1476000.0 2049000.0 ;
      RECT  1465800.0 2062800.0 1476000.0 2049000.0 ;
      RECT  1465800.0 2062800.0 1476000.0 2076600.0 ;
      RECT  1465800.0 2090400.0 1476000.0 2076600.0 ;
      RECT  1465800.0 2090400.0 1476000.0 2104200.0 ;
      RECT  1465800.0 2118000.0 1476000.0 2104200.0 ;
      RECT  1465800.0 2118000.0 1476000.0 2131800.0 ;
      RECT  1465800.0 2145600.0 1476000.0 2131800.0 ;
      RECT  1476000.0 379200.0 1486200.0 393000.0 ;
      RECT  1476000.0 406800.0 1486200.0 393000.0 ;
      RECT  1476000.0 406800.0 1486200.0 420600.0 ;
      RECT  1476000.0 434400.0 1486200.0 420600.0 ;
      RECT  1476000.0 434400.0 1486200.0 448200.0 ;
      RECT  1476000.0 462000.0 1486200.0 448200.0 ;
      RECT  1476000.0 462000.0 1486200.0 475800.0 ;
      RECT  1476000.0 489600.0 1486200.0 475800.0 ;
      RECT  1476000.0 489600.0 1486200.0 503400.0 ;
      RECT  1476000.0 517200.0 1486200.0 503400.0 ;
      RECT  1476000.0 517200.0 1486200.0 531000.0 ;
      RECT  1476000.0 544800.0 1486200.0 531000.0 ;
      RECT  1476000.0 544800.0 1486200.0 558600.0 ;
      RECT  1476000.0 572400.0 1486200.0 558600.0 ;
      RECT  1476000.0 572400.0 1486200.0 586200.0 ;
      RECT  1476000.0 600000.0 1486200.0 586200.0 ;
      RECT  1476000.0 600000.0 1486200.0 613800.0 ;
      RECT  1476000.0 627600.0 1486200.0 613800.0 ;
      RECT  1476000.0 627600.0 1486200.0 641400.0 ;
      RECT  1476000.0 655200.0 1486200.0 641400.0 ;
      RECT  1476000.0 655200.0 1486200.0 669000.0 ;
      RECT  1476000.0 682800.0 1486200.0 669000.0 ;
      RECT  1476000.0 682800.0 1486200.0 696600.0 ;
      RECT  1476000.0 710400.0 1486200.0 696600.0 ;
      RECT  1476000.0 710400.0 1486200.0 724200.0 ;
      RECT  1476000.0 738000.0 1486200.0 724200.0 ;
      RECT  1476000.0 738000.0 1486200.0 751800.0 ;
      RECT  1476000.0 765600.0 1486200.0 751800.0 ;
      RECT  1476000.0 765600.0 1486200.0 779400.0 ;
      RECT  1476000.0 793200.0 1486200.0 779400.0 ;
      RECT  1476000.0 793200.0 1486200.0 807000.0 ;
      RECT  1476000.0 820800.0 1486200.0 807000.0 ;
      RECT  1476000.0 820800.0 1486200.0 834600.0 ;
      RECT  1476000.0 848400.0 1486200.0 834600.0 ;
      RECT  1476000.0 848400.0 1486200.0 862200.0 ;
      RECT  1476000.0 876000.0 1486200.0 862200.0 ;
      RECT  1476000.0 876000.0 1486200.0 889800.0 ;
      RECT  1476000.0 903600.0 1486200.0 889800.0 ;
      RECT  1476000.0 903600.0 1486200.0 917400.0 ;
      RECT  1476000.0 931200.0 1486200.0 917400.0 ;
      RECT  1476000.0 931200.0 1486200.0 945000.0 ;
      RECT  1476000.0 958800.0 1486200.0 945000.0 ;
      RECT  1476000.0 958800.0 1486200.0 972600.0 ;
      RECT  1476000.0 986400.0 1486200.0 972600.0 ;
      RECT  1476000.0 986400.0 1486200.0 1000200.0 ;
      RECT  1476000.0 1014000.0 1486200.0 1000200.0 ;
      RECT  1476000.0 1014000.0 1486200.0 1027800.0 ;
      RECT  1476000.0 1041600.0 1486200.0 1027800.0 ;
      RECT  1476000.0 1041600.0 1486200.0 1055400.0 ;
      RECT  1476000.0 1069200.0 1486200.0 1055400.0 ;
      RECT  1476000.0 1069200.0 1486200.0 1083000.0 ;
      RECT  1476000.0 1096800.0 1486200.0 1083000.0 ;
      RECT  1476000.0 1096800.0 1486200.0 1110600.0 ;
      RECT  1476000.0 1124400.0 1486200.0 1110600.0 ;
      RECT  1476000.0 1124400.0 1486200.0 1138200.0 ;
      RECT  1476000.0 1152000.0 1486200.0 1138200.0 ;
      RECT  1476000.0 1152000.0 1486200.0 1165800.0 ;
      RECT  1476000.0 1179600.0 1486200.0 1165800.0 ;
      RECT  1476000.0 1179600.0 1486200.0 1193400.0 ;
      RECT  1476000.0 1207200.0 1486200.0 1193400.0 ;
      RECT  1476000.0 1207200.0 1486200.0 1221000.0 ;
      RECT  1476000.0 1234800.0 1486200.0 1221000.0 ;
      RECT  1476000.0 1234800.0 1486200.0 1248600.0 ;
      RECT  1476000.0 1262400.0 1486200.0 1248600.0 ;
      RECT  1476000.0 1262400.0 1486200.0 1276200.0 ;
      RECT  1476000.0 1290000.0 1486200.0 1276200.0 ;
      RECT  1476000.0 1290000.0 1486200.0 1303800.0 ;
      RECT  1476000.0 1317600.0 1486200.0 1303800.0 ;
      RECT  1476000.0 1317600.0 1486200.0 1331400.0 ;
      RECT  1476000.0 1345200.0 1486200.0 1331400.0 ;
      RECT  1476000.0 1345200.0 1486200.0 1359000.0 ;
      RECT  1476000.0 1372800.0 1486200.0 1359000.0 ;
      RECT  1476000.0 1372800.0 1486200.0 1386600.0 ;
      RECT  1476000.0 1400400.0 1486200.0 1386600.0 ;
      RECT  1476000.0 1400400.0 1486200.0 1414200.0 ;
      RECT  1476000.0 1428000.0 1486200.0 1414200.0 ;
      RECT  1476000.0 1428000.0 1486200.0 1441800.0 ;
      RECT  1476000.0 1455600.0 1486200.0 1441800.0 ;
      RECT  1476000.0 1455600.0 1486200.0 1469400.0 ;
      RECT  1476000.0 1483200.0 1486200.0 1469400.0 ;
      RECT  1476000.0 1483200.0 1486200.0 1497000.0 ;
      RECT  1476000.0 1510800.0 1486200.0 1497000.0 ;
      RECT  1476000.0 1510800.0 1486200.0 1524600.0 ;
      RECT  1476000.0 1538400.0 1486200.0 1524600.0 ;
      RECT  1476000.0 1538400.0 1486200.0 1552200.0 ;
      RECT  1476000.0 1566000.0 1486200.0 1552200.0 ;
      RECT  1476000.0 1566000.0 1486200.0 1579800.0 ;
      RECT  1476000.0 1593600.0 1486200.0 1579800.0 ;
      RECT  1476000.0 1593600.0 1486200.0 1607400.0 ;
      RECT  1476000.0 1621200.0 1486200.0 1607400.0 ;
      RECT  1476000.0 1621200.0 1486200.0 1635000.0 ;
      RECT  1476000.0 1648800.0 1486200.0 1635000.0 ;
      RECT  1476000.0 1648800.0 1486200.0 1662600.0 ;
      RECT  1476000.0 1676400.0 1486200.0 1662600.0 ;
      RECT  1476000.0 1676400.0 1486200.0 1690200.0 ;
      RECT  1476000.0 1704000.0 1486200.0 1690200.0 ;
      RECT  1476000.0 1704000.0 1486200.0 1717800.0 ;
      RECT  1476000.0 1731600.0 1486200.0 1717800.0 ;
      RECT  1476000.0 1731600.0 1486200.0 1745400.0 ;
      RECT  1476000.0 1759200.0 1486200.0 1745400.0 ;
      RECT  1476000.0 1759200.0 1486200.0 1773000.0 ;
      RECT  1476000.0 1786800.0 1486200.0 1773000.0 ;
      RECT  1476000.0 1786800.0 1486200.0 1800600.0 ;
      RECT  1476000.0 1814400.0 1486200.0 1800600.0 ;
      RECT  1476000.0 1814400.0 1486200.0 1828200.0 ;
      RECT  1476000.0 1842000.0 1486200.0 1828200.0 ;
      RECT  1476000.0 1842000.0 1486200.0 1855800.0 ;
      RECT  1476000.0 1869600.0 1486200.0 1855800.0 ;
      RECT  1476000.0 1869600.0 1486200.0 1883400.0 ;
      RECT  1476000.0 1897200.0 1486200.0 1883400.0 ;
      RECT  1476000.0 1897200.0 1486200.0 1911000.0 ;
      RECT  1476000.0 1924800.0 1486200.0 1911000.0 ;
      RECT  1476000.0 1924800.0 1486200.0 1938600.0 ;
      RECT  1476000.0 1952400.0 1486200.0 1938600.0 ;
      RECT  1476000.0 1952400.0 1486200.0 1966200.0 ;
      RECT  1476000.0 1980000.0 1486200.0 1966200.0 ;
      RECT  1476000.0 1980000.0 1486200.0 1993800.0 ;
      RECT  1476000.0 2007600.0 1486200.0 1993800.0 ;
      RECT  1476000.0 2007600.0 1486200.0 2021400.0 ;
      RECT  1476000.0 2035200.0 1486200.0 2021400.0 ;
      RECT  1476000.0 2035200.0 1486200.0 2049000.0 ;
      RECT  1476000.0 2062800.0 1486200.0 2049000.0 ;
      RECT  1476000.0 2062800.0 1486200.0 2076600.0 ;
      RECT  1476000.0 2090400.0 1486200.0 2076600.0 ;
      RECT  1476000.0 2090400.0 1486200.0 2104200.0 ;
      RECT  1476000.0 2118000.0 1486200.0 2104200.0 ;
      RECT  1476000.0 2118000.0 1486200.0 2131800.0 ;
      RECT  1476000.0 2145600.0 1486200.0 2131800.0 ;
      RECT  1486200.0 379200.0 1496400.0 393000.0 ;
      RECT  1486200.0 406800.0 1496400.0 393000.0 ;
      RECT  1486200.0 406800.0 1496400.0 420600.0 ;
      RECT  1486200.0 434400.0 1496400.0 420600.0 ;
      RECT  1486200.0 434400.0 1496400.0 448200.0 ;
      RECT  1486200.0 462000.0 1496400.0 448200.0 ;
      RECT  1486200.0 462000.0 1496400.0 475800.0 ;
      RECT  1486200.0 489600.0 1496400.0 475800.0 ;
      RECT  1486200.0 489600.0 1496400.0 503400.0 ;
      RECT  1486200.0 517200.0 1496400.0 503400.0 ;
      RECT  1486200.0 517200.0 1496400.0 531000.0 ;
      RECT  1486200.0 544800.0 1496400.0 531000.0 ;
      RECT  1486200.0 544800.0 1496400.0 558600.0 ;
      RECT  1486200.0 572400.0 1496400.0 558600.0 ;
      RECT  1486200.0 572400.0 1496400.0 586200.0 ;
      RECT  1486200.0 600000.0 1496400.0 586200.0 ;
      RECT  1486200.0 600000.0 1496400.0 613800.0 ;
      RECT  1486200.0 627600.0 1496400.0 613800.0 ;
      RECT  1486200.0 627600.0 1496400.0 641400.0 ;
      RECT  1486200.0 655200.0 1496400.0 641400.0 ;
      RECT  1486200.0 655200.0 1496400.0 669000.0 ;
      RECT  1486200.0 682800.0 1496400.0 669000.0 ;
      RECT  1486200.0 682800.0 1496400.0 696600.0 ;
      RECT  1486200.0 710400.0 1496400.0 696600.0 ;
      RECT  1486200.0 710400.0 1496400.0 724200.0 ;
      RECT  1486200.0 738000.0 1496400.0 724200.0 ;
      RECT  1486200.0 738000.0 1496400.0 751800.0 ;
      RECT  1486200.0 765600.0 1496400.0 751800.0 ;
      RECT  1486200.0 765600.0 1496400.0 779400.0 ;
      RECT  1486200.0 793200.0 1496400.0 779400.0 ;
      RECT  1486200.0 793200.0 1496400.0 807000.0 ;
      RECT  1486200.0 820800.0 1496400.0 807000.0 ;
      RECT  1486200.0 820800.0 1496400.0 834600.0 ;
      RECT  1486200.0 848400.0 1496400.0 834600.0 ;
      RECT  1486200.0 848400.0 1496400.0 862200.0 ;
      RECT  1486200.0 876000.0 1496400.0 862200.0 ;
      RECT  1486200.0 876000.0 1496400.0 889800.0 ;
      RECT  1486200.0 903600.0 1496400.0 889800.0 ;
      RECT  1486200.0 903600.0 1496400.0 917400.0 ;
      RECT  1486200.0 931200.0 1496400.0 917400.0 ;
      RECT  1486200.0 931200.0 1496400.0 945000.0 ;
      RECT  1486200.0 958800.0 1496400.0 945000.0 ;
      RECT  1486200.0 958800.0 1496400.0 972600.0 ;
      RECT  1486200.0 986400.0 1496400.0 972600.0 ;
      RECT  1486200.0 986400.0 1496400.0 1000200.0 ;
      RECT  1486200.0 1014000.0 1496400.0 1000200.0 ;
      RECT  1486200.0 1014000.0 1496400.0 1027800.0 ;
      RECT  1486200.0 1041600.0 1496400.0 1027800.0 ;
      RECT  1486200.0 1041600.0 1496400.0 1055400.0 ;
      RECT  1486200.0 1069200.0 1496400.0 1055400.0 ;
      RECT  1486200.0 1069200.0 1496400.0 1083000.0 ;
      RECT  1486200.0 1096800.0 1496400.0 1083000.0 ;
      RECT  1486200.0 1096800.0 1496400.0 1110600.0 ;
      RECT  1486200.0 1124400.0 1496400.0 1110600.0 ;
      RECT  1486200.0 1124400.0 1496400.0 1138200.0 ;
      RECT  1486200.0 1152000.0 1496400.0 1138200.0 ;
      RECT  1486200.0 1152000.0 1496400.0 1165800.0 ;
      RECT  1486200.0 1179600.0 1496400.0 1165800.0 ;
      RECT  1486200.0 1179600.0 1496400.0 1193400.0 ;
      RECT  1486200.0 1207200.0 1496400.0 1193400.0 ;
      RECT  1486200.0 1207200.0 1496400.0 1221000.0 ;
      RECT  1486200.0 1234800.0 1496400.0 1221000.0 ;
      RECT  1486200.0 1234800.0 1496400.0 1248600.0 ;
      RECT  1486200.0 1262400.0 1496400.0 1248600.0 ;
      RECT  1486200.0 1262400.0 1496400.0 1276200.0 ;
      RECT  1486200.0 1290000.0 1496400.0 1276200.0 ;
      RECT  1486200.0 1290000.0 1496400.0 1303800.0 ;
      RECT  1486200.0 1317600.0 1496400.0 1303800.0 ;
      RECT  1486200.0 1317600.0 1496400.0 1331400.0 ;
      RECT  1486200.0 1345200.0 1496400.0 1331400.0 ;
      RECT  1486200.0 1345200.0 1496400.0 1359000.0 ;
      RECT  1486200.0 1372800.0 1496400.0 1359000.0 ;
      RECT  1486200.0 1372800.0 1496400.0 1386600.0 ;
      RECT  1486200.0 1400400.0 1496400.0 1386600.0 ;
      RECT  1486200.0 1400400.0 1496400.0 1414200.0 ;
      RECT  1486200.0 1428000.0 1496400.0 1414200.0 ;
      RECT  1486200.0 1428000.0 1496400.0 1441800.0 ;
      RECT  1486200.0 1455600.0 1496400.0 1441800.0 ;
      RECT  1486200.0 1455600.0 1496400.0 1469400.0 ;
      RECT  1486200.0 1483200.0 1496400.0 1469400.0 ;
      RECT  1486200.0 1483200.0 1496400.0 1497000.0 ;
      RECT  1486200.0 1510800.0 1496400.0 1497000.0 ;
      RECT  1486200.0 1510800.0 1496400.0 1524600.0 ;
      RECT  1486200.0 1538400.0 1496400.0 1524600.0 ;
      RECT  1486200.0 1538400.0 1496400.0 1552200.0 ;
      RECT  1486200.0 1566000.0 1496400.0 1552200.0 ;
      RECT  1486200.0 1566000.0 1496400.0 1579800.0 ;
      RECT  1486200.0 1593600.0 1496400.0 1579800.0 ;
      RECT  1486200.0 1593600.0 1496400.0 1607400.0 ;
      RECT  1486200.0 1621200.0 1496400.0 1607400.0 ;
      RECT  1486200.0 1621200.0 1496400.0 1635000.0 ;
      RECT  1486200.0 1648800.0 1496400.0 1635000.0 ;
      RECT  1486200.0 1648800.0 1496400.0 1662600.0 ;
      RECT  1486200.0 1676400.0 1496400.0 1662600.0 ;
      RECT  1486200.0 1676400.0 1496400.0 1690200.0 ;
      RECT  1486200.0 1704000.0 1496400.0 1690200.0 ;
      RECT  1486200.0 1704000.0 1496400.0 1717800.0 ;
      RECT  1486200.0 1731600.0 1496400.0 1717800.0 ;
      RECT  1486200.0 1731600.0 1496400.0 1745400.0 ;
      RECT  1486200.0 1759200.0 1496400.0 1745400.0 ;
      RECT  1486200.0 1759200.0 1496400.0 1773000.0 ;
      RECT  1486200.0 1786800.0 1496400.0 1773000.0 ;
      RECT  1486200.0 1786800.0 1496400.0 1800600.0 ;
      RECT  1486200.0 1814400.0 1496400.0 1800600.0 ;
      RECT  1486200.0 1814400.0 1496400.0 1828200.0 ;
      RECT  1486200.0 1842000.0 1496400.0 1828200.0 ;
      RECT  1486200.0 1842000.0 1496400.0 1855800.0 ;
      RECT  1486200.0 1869600.0 1496400.0 1855800.0 ;
      RECT  1486200.0 1869600.0 1496400.0 1883400.0 ;
      RECT  1486200.0 1897200.0 1496400.0 1883400.0 ;
      RECT  1486200.0 1897200.0 1496400.0 1911000.0 ;
      RECT  1486200.0 1924800.0 1496400.0 1911000.0 ;
      RECT  1486200.0 1924800.0 1496400.0 1938600.0 ;
      RECT  1486200.0 1952400.0 1496400.0 1938600.0 ;
      RECT  1486200.0 1952400.0 1496400.0 1966200.0 ;
      RECT  1486200.0 1980000.0 1496400.0 1966200.0 ;
      RECT  1486200.0 1980000.0 1496400.0 1993800.0 ;
      RECT  1486200.0 2007600.0 1496400.0 1993800.0 ;
      RECT  1486200.0 2007600.0 1496400.0 2021400.0 ;
      RECT  1486200.0 2035200.0 1496400.0 2021400.0 ;
      RECT  1486200.0 2035200.0 1496400.0 2049000.0 ;
      RECT  1486200.0 2062800.0 1496400.0 2049000.0 ;
      RECT  1486200.0 2062800.0 1496400.0 2076600.0 ;
      RECT  1486200.0 2090400.0 1496400.0 2076600.0 ;
      RECT  1486200.0 2090400.0 1496400.0 2104200.0 ;
      RECT  1486200.0 2118000.0 1496400.0 2104200.0 ;
      RECT  1486200.0 2118000.0 1496400.0 2131800.0 ;
      RECT  1486200.0 2145600.0 1496400.0 2131800.0 ;
      RECT  1496400.0 379200.0 1506600.0 393000.0 ;
      RECT  1496400.0 406800.0 1506600.0 393000.0 ;
      RECT  1496400.0 406800.0 1506600.0 420600.0 ;
      RECT  1496400.0 434400.0 1506600.0 420600.0 ;
      RECT  1496400.0 434400.0 1506600.0 448200.0 ;
      RECT  1496400.0 462000.0 1506600.0 448200.0 ;
      RECT  1496400.0 462000.0 1506600.0 475800.0 ;
      RECT  1496400.0 489600.0 1506600.0 475800.0 ;
      RECT  1496400.0 489600.0 1506600.0 503400.0 ;
      RECT  1496400.0 517200.0 1506600.0 503400.0 ;
      RECT  1496400.0 517200.0 1506600.0 531000.0 ;
      RECT  1496400.0 544800.0 1506600.0 531000.0 ;
      RECT  1496400.0 544800.0 1506600.0 558600.0 ;
      RECT  1496400.0 572400.0 1506600.0 558600.0 ;
      RECT  1496400.0 572400.0 1506600.0 586200.0 ;
      RECT  1496400.0 600000.0 1506600.0 586200.0 ;
      RECT  1496400.0 600000.0 1506600.0 613800.0 ;
      RECT  1496400.0 627600.0 1506600.0 613800.0 ;
      RECT  1496400.0 627600.0 1506600.0 641400.0 ;
      RECT  1496400.0 655200.0 1506600.0 641400.0 ;
      RECT  1496400.0 655200.0 1506600.0 669000.0 ;
      RECT  1496400.0 682800.0 1506600.0 669000.0 ;
      RECT  1496400.0 682800.0 1506600.0 696600.0 ;
      RECT  1496400.0 710400.0 1506600.0 696600.0 ;
      RECT  1496400.0 710400.0 1506600.0 724200.0 ;
      RECT  1496400.0 738000.0 1506600.0 724200.0 ;
      RECT  1496400.0 738000.0 1506600.0 751800.0 ;
      RECT  1496400.0 765600.0 1506600.0 751800.0 ;
      RECT  1496400.0 765600.0 1506600.0 779400.0 ;
      RECT  1496400.0 793200.0 1506600.0 779400.0 ;
      RECT  1496400.0 793200.0 1506600.0 807000.0 ;
      RECT  1496400.0 820800.0 1506600.0 807000.0 ;
      RECT  1496400.0 820800.0 1506600.0 834600.0 ;
      RECT  1496400.0 848400.0 1506600.0 834600.0 ;
      RECT  1496400.0 848400.0 1506600.0 862200.0 ;
      RECT  1496400.0 876000.0 1506600.0 862200.0 ;
      RECT  1496400.0 876000.0 1506600.0 889800.0 ;
      RECT  1496400.0 903600.0 1506600.0 889800.0 ;
      RECT  1496400.0 903600.0 1506600.0 917400.0 ;
      RECT  1496400.0 931200.0 1506600.0 917400.0 ;
      RECT  1496400.0 931200.0 1506600.0 945000.0 ;
      RECT  1496400.0 958800.0 1506600.0 945000.0 ;
      RECT  1496400.0 958800.0 1506600.0 972600.0 ;
      RECT  1496400.0 986400.0 1506600.0 972600.0 ;
      RECT  1496400.0 986400.0 1506600.0 1000200.0 ;
      RECT  1496400.0 1014000.0 1506600.0 1000200.0 ;
      RECT  1496400.0 1014000.0 1506600.0 1027800.0 ;
      RECT  1496400.0 1041600.0 1506600.0 1027800.0 ;
      RECT  1496400.0 1041600.0 1506600.0 1055400.0 ;
      RECT  1496400.0 1069200.0 1506600.0 1055400.0 ;
      RECT  1496400.0 1069200.0 1506600.0 1083000.0 ;
      RECT  1496400.0 1096800.0 1506600.0 1083000.0 ;
      RECT  1496400.0 1096800.0 1506600.0 1110600.0 ;
      RECT  1496400.0 1124400.0 1506600.0 1110600.0 ;
      RECT  1496400.0 1124400.0 1506600.0 1138200.0 ;
      RECT  1496400.0 1152000.0 1506600.0 1138200.0 ;
      RECT  1496400.0 1152000.0 1506600.0 1165800.0 ;
      RECT  1496400.0 1179600.0 1506600.0 1165800.0 ;
      RECT  1496400.0 1179600.0 1506600.0 1193400.0 ;
      RECT  1496400.0 1207200.0 1506600.0 1193400.0 ;
      RECT  1496400.0 1207200.0 1506600.0 1221000.0 ;
      RECT  1496400.0 1234800.0 1506600.0 1221000.0 ;
      RECT  1496400.0 1234800.0 1506600.0 1248600.0 ;
      RECT  1496400.0 1262400.0 1506600.0 1248600.0 ;
      RECT  1496400.0 1262400.0 1506600.0 1276200.0 ;
      RECT  1496400.0 1290000.0 1506600.0 1276200.0 ;
      RECT  1496400.0 1290000.0 1506600.0 1303800.0 ;
      RECT  1496400.0 1317600.0 1506600.0 1303800.0 ;
      RECT  1496400.0 1317600.0 1506600.0 1331400.0 ;
      RECT  1496400.0 1345200.0 1506600.0 1331400.0 ;
      RECT  1496400.0 1345200.0 1506600.0 1359000.0 ;
      RECT  1496400.0 1372800.0 1506600.0 1359000.0 ;
      RECT  1496400.0 1372800.0 1506600.0 1386600.0 ;
      RECT  1496400.0 1400400.0 1506600.0 1386600.0 ;
      RECT  1496400.0 1400400.0 1506600.0 1414200.0 ;
      RECT  1496400.0 1428000.0 1506600.0 1414200.0 ;
      RECT  1496400.0 1428000.0 1506600.0 1441800.0 ;
      RECT  1496400.0 1455600.0 1506600.0 1441800.0 ;
      RECT  1496400.0 1455600.0 1506600.0 1469400.0 ;
      RECT  1496400.0 1483200.0 1506600.0 1469400.0 ;
      RECT  1496400.0 1483200.0 1506600.0 1497000.0 ;
      RECT  1496400.0 1510800.0 1506600.0 1497000.0 ;
      RECT  1496400.0 1510800.0 1506600.0 1524600.0 ;
      RECT  1496400.0 1538400.0 1506600.0 1524600.0 ;
      RECT  1496400.0 1538400.0 1506600.0 1552200.0 ;
      RECT  1496400.0 1566000.0 1506600.0 1552200.0 ;
      RECT  1496400.0 1566000.0 1506600.0 1579800.0 ;
      RECT  1496400.0 1593600.0 1506600.0 1579800.0 ;
      RECT  1496400.0 1593600.0 1506600.0 1607400.0 ;
      RECT  1496400.0 1621200.0 1506600.0 1607400.0 ;
      RECT  1496400.0 1621200.0 1506600.0 1635000.0 ;
      RECT  1496400.0 1648800.0 1506600.0 1635000.0 ;
      RECT  1496400.0 1648800.0 1506600.0 1662600.0 ;
      RECT  1496400.0 1676400.0 1506600.0 1662600.0 ;
      RECT  1496400.0 1676400.0 1506600.0 1690200.0 ;
      RECT  1496400.0 1704000.0 1506600.0 1690200.0 ;
      RECT  1496400.0 1704000.0 1506600.0 1717800.0 ;
      RECT  1496400.0 1731600.0 1506600.0 1717800.0 ;
      RECT  1496400.0 1731600.0 1506600.0 1745400.0 ;
      RECT  1496400.0 1759200.0 1506600.0 1745400.0 ;
      RECT  1496400.0 1759200.0 1506600.0 1773000.0 ;
      RECT  1496400.0 1786800.0 1506600.0 1773000.0 ;
      RECT  1496400.0 1786800.0 1506600.0 1800600.0 ;
      RECT  1496400.0 1814400.0 1506600.0 1800600.0 ;
      RECT  1496400.0 1814400.0 1506600.0 1828200.0 ;
      RECT  1496400.0 1842000.0 1506600.0 1828200.0 ;
      RECT  1496400.0 1842000.0 1506600.0 1855800.0 ;
      RECT  1496400.0 1869600.0 1506600.0 1855800.0 ;
      RECT  1496400.0 1869600.0 1506600.0 1883400.0 ;
      RECT  1496400.0 1897200.0 1506600.0 1883400.0 ;
      RECT  1496400.0 1897200.0 1506600.0 1911000.0 ;
      RECT  1496400.0 1924800.0 1506600.0 1911000.0 ;
      RECT  1496400.0 1924800.0 1506600.0 1938600.0 ;
      RECT  1496400.0 1952400.0 1506600.0 1938600.0 ;
      RECT  1496400.0 1952400.0 1506600.0 1966200.0 ;
      RECT  1496400.0 1980000.0 1506600.0 1966200.0 ;
      RECT  1496400.0 1980000.0 1506600.0 1993800.0 ;
      RECT  1496400.0 2007600.0 1506600.0 1993800.0 ;
      RECT  1496400.0 2007600.0 1506600.0 2021400.0 ;
      RECT  1496400.0 2035200.0 1506600.0 2021400.0 ;
      RECT  1496400.0 2035200.0 1506600.0 2049000.0 ;
      RECT  1496400.0 2062800.0 1506600.0 2049000.0 ;
      RECT  1496400.0 2062800.0 1506600.0 2076600.0 ;
      RECT  1496400.0 2090400.0 1506600.0 2076600.0 ;
      RECT  1496400.0 2090400.0 1506600.0 2104200.0 ;
      RECT  1496400.0 2118000.0 1506600.0 2104200.0 ;
      RECT  1496400.0 2118000.0 1506600.0 2131800.0 ;
      RECT  1496400.0 2145600.0 1506600.0 2131800.0 ;
      RECT  1506600.0 379200.0 1516800.0 393000.0 ;
      RECT  1506600.0 406800.0 1516800.0 393000.0 ;
      RECT  1506600.0 406800.0 1516800.0 420600.0 ;
      RECT  1506600.0 434400.0 1516800.0 420600.0 ;
      RECT  1506600.0 434400.0 1516800.0 448200.0 ;
      RECT  1506600.0 462000.0 1516800.0 448200.0 ;
      RECT  1506600.0 462000.0 1516800.0 475800.0 ;
      RECT  1506600.0 489600.0 1516800.0 475800.0 ;
      RECT  1506600.0 489600.0 1516800.0 503400.0 ;
      RECT  1506600.0 517200.0 1516800.0 503400.0 ;
      RECT  1506600.0 517200.0 1516800.0 531000.0 ;
      RECT  1506600.0 544800.0 1516800.0 531000.0 ;
      RECT  1506600.0 544800.0 1516800.0 558600.0 ;
      RECT  1506600.0 572400.0 1516800.0 558600.0 ;
      RECT  1506600.0 572400.0 1516800.0 586200.0 ;
      RECT  1506600.0 600000.0 1516800.0 586200.0 ;
      RECT  1506600.0 600000.0 1516800.0 613800.0 ;
      RECT  1506600.0 627600.0 1516800.0 613800.0 ;
      RECT  1506600.0 627600.0 1516800.0 641400.0 ;
      RECT  1506600.0 655200.0 1516800.0 641400.0 ;
      RECT  1506600.0 655200.0 1516800.0 669000.0 ;
      RECT  1506600.0 682800.0 1516800.0 669000.0 ;
      RECT  1506600.0 682800.0 1516800.0 696600.0 ;
      RECT  1506600.0 710400.0 1516800.0 696600.0 ;
      RECT  1506600.0 710400.0 1516800.0 724200.0 ;
      RECT  1506600.0 738000.0 1516800.0 724200.0 ;
      RECT  1506600.0 738000.0 1516800.0 751800.0 ;
      RECT  1506600.0 765600.0 1516800.0 751800.0 ;
      RECT  1506600.0 765600.0 1516800.0 779400.0 ;
      RECT  1506600.0 793200.0 1516800.0 779400.0 ;
      RECT  1506600.0 793200.0 1516800.0 807000.0 ;
      RECT  1506600.0 820800.0 1516800.0 807000.0 ;
      RECT  1506600.0 820800.0 1516800.0 834600.0 ;
      RECT  1506600.0 848400.0 1516800.0 834600.0 ;
      RECT  1506600.0 848400.0 1516800.0 862200.0 ;
      RECT  1506600.0 876000.0 1516800.0 862200.0 ;
      RECT  1506600.0 876000.0 1516800.0 889800.0 ;
      RECT  1506600.0 903600.0 1516800.0 889800.0 ;
      RECT  1506600.0 903600.0 1516800.0 917400.0 ;
      RECT  1506600.0 931200.0 1516800.0 917400.0 ;
      RECT  1506600.0 931200.0 1516800.0 945000.0 ;
      RECT  1506600.0 958800.0 1516800.0 945000.0 ;
      RECT  1506600.0 958800.0 1516800.0 972600.0 ;
      RECT  1506600.0 986400.0 1516800.0 972600.0 ;
      RECT  1506600.0 986400.0 1516800.0 1000200.0 ;
      RECT  1506600.0 1014000.0 1516800.0 1000200.0 ;
      RECT  1506600.0 1014000.0 1516800.0 1027800.0 ;
      RECT  1506600.0 1041600.0 1516800.0 1027800.0 ;
      RECT  1506600.0 1041600.0 1516800.0 1055400.0 ;
      RECT  1506600.0 1069200.0 1516800.0 1055400.0 ;
      RECT  1506600.0 1069200.0 1516800.0 1083000.0 ;
      RECT  1506600.0 1096800.0 1516800.0 1083000.0 ;
      RECT  1506600.0 1096800.0 1516800.0 1110600.0 ;
      RECT  1506600.0 1124400.0 1516800.0 1110600.0 ;
      RECT  1506600.0 1124400.0 1516800.0 1138200.0 ;
      RECT  1506600.0 1152000.0 1516800.0 1138200.0 ;
      RECT  1506600.0 1152000.0 1516800.0 1165800.0 ;
      RECT  1506600.0 1179600.0 1516800.0 1165800.0 ;
      RECT  1506600.0 1179600.0 1516800.0 1193400.0 ;
      RECT  1506600.0 1207200.0 1516800.0 1193400.0 ;
      RECT  1506600.0 1207200.0 1516800.0 1221000.0 ;
      RECT  1506600.0 1234800.0 1516800.0 1221000.0 ;
      RECT  1506600.0 1234800.0 1516800.0 1248600.0 ;
      RECT  1506600.0 1262400.0 1516800.0 1248600.0 ;
      RECT  1506600.0 1262400.0 1516800.0 1276200.0 ;
      RECT  1506600.0 1290000.0 1516800.0 1276200.0 ;
      RECT  1506600.0 1290000.0 1516800.0 1303800.0 ;
      RECT  1506600.0 1317600.0 1516800.0 1303800.0 ;
      RECT  1506600.0 1317600.0 1516800.0 1331400.0 ;
      RECT  1506600.0 1345200.0 1516800.0 1331400.0 ;
      RECT  1506600.0 1345200.0 1516800.0 1359000.0 ;
      RECT  1506600.0 1372800.0 1516800.0 1359000.0 ;
      RECT  1506600.0 1372800.0 1516800.0 1386600.0 ;
      RECT  1506600.0 1400400.0 1516800.0 1386600.0 ;
      RECT  1506600.0 1400400.0 1516800.0 1414200.0 ;
      RECT  1506600.0 1428000.0 1516800.0 1414200.0 ;
      RECT  1506600.0 1428000.0 1516800.0 1441800.0 ;
      RECT  1506600.0 1455600.0 1516800.0 1441800.0 ;
      RECT  1506600.0 1455600.0 1516800.0 1469400.0 ;
      RECT  1506600.0 1483200.0 1516800.0 1469400.0 ;
      RECT  1506600.0 1483200.0 1516800.0 1497000.0 ;
      RECT  1506600.0 1510800.0 1516800.0 1497000.0 ;
      RECT  1506600.0 1510800.0 1516800.0 1524600.0 ;
      RECT  1506600.0 1538400.0 1516800.0 1524600.0 ;
      RECT  1506600.0 1538400.0 1516800.0 1552200.0 ;
      RECT  1506600.0 1566000.0 1516800.0 1552200.0 ;
      RECT  1506600.0 1566000.0 1516800.0 1579800.0 ;
      RECT  1506600.0 1593600.0 1516800.0 1579800.0 ;
      RECT  1506600.0 1593600.0 1516800.0 1607400.0 ;
      RECT  1506600.0 1621200.0 1516800.0 1607400.0 ;
      RECT  1506600.0 1621200.0 1516800.0 1635000.0 ;
      RECT  1506600.0 1648800.0 1516800.0 1635000.0 ;
      RECT  1506600.0 1648800.0 1516800.0 1662600.0 ;
      RECT  1506600.0 1676400.0 1516800.0 1662600.0 ;
      RECT  1506600.0 1676400.0 1516800.0 1690200.0 ;
      RECT  1506600.0 1704000.0 1516800.0 1690200.0 ;
      RECT  1506600.0 1704000.0 1516800.0 1717800.0 ;
      RECT  1506600.0 1731600.0 1516800.0 1717800.0 ;
      RECT  1506600.0 1731600.0 1516800.0 1745400.0 ;
      RECT  1506600.0 1759200.0 1516800.0 1745400.0 ;
      RECT  1506600.0 1759200.0 1516800.0 1773000.0 ;
      RECT  1506600.0 1786800.0 1516800.0 1773000.0 ;
      RECT  1506600.0 1786800.0 1516800.0 1800600.0 ;
      RECT  1506600.0 1814400.0 1516800.0 1800600.0 ;
      RECT  1506600.0 1814400.0 1516800.0 1828200.0 ;
      RECT  1506600.0 1842000.0 1516800.0 1828200.0 ;
      RECT  1506600.0 1842000.0 1516800.0 1855800.0 ;
      RECT  1506600.0 1869600.0 1516800.0 1855800.0 ;
      RECT  1506600.0 1869600.0 1516800.0 1883400.0 ;
      RECT  1506600.0 1897200.0 1516800.0 1883400.0 ;
      RECT  1506600.0 1897200.0 1516800.0 1911000.0 ;
      RECT  1506600.0 1924800.0 1516800.0 1911000.0 ;
      RECT  1506600.0 1924800.0 1516800.0 1938600.0 ;
      RECT  1506600.0 1952400.0 1516800.0 1938600.0 ;
      RECT  1506600.0 1952400.0 1516800.0 1966200.0 ;
      RECT  1506600.0 1980000.0 1516800.0 1966200.0 ;
      RECT  1506600.0 1980000.0 1516800.0 1993800.0 ;
      RECT  1506600.0 2007600.0 1516800.0 1993800.0 ;
      RECT  1506600.0 2007600.0 1516800.0 2021400.0 ;
      RECT  1506600.0 2035200.0 1516800.0 2021400.0 ;
      RECT  1506600.0 2035200.0 1516800.0 2049000.0 ;
      RECT  1506600.0 2062800.0 1516800.0 2049000.0 ;
      RECT  1506600.0 2062800.0 1516800.0 2076600.0 ;
      RECT  1506600.0 2090400.0 1516800.0 2076600.0 ;
      RECT  1506600.0 2090400.0 1516800.0 2104200.0 ;
      RECT  1506600.0 2118000.0 1516800.0 2104200.0 ;
      RECT  1506600.0 2118000.0 1516800.0 2131800.0 ;
      RECT  1506600.0 2145600.0 1516800.0 2131800.0 ;
      RECT  1516800.0 379200.0 1527000.0 393000.0 ;
      RECT  1516800.0 406800.0 1527000.0 393000.0 ;
      RECT  1516800.0 406800.0 1527000.0 420600.0 ;
      RECT  1516800.0 434400.0 1527000.0 420600.0 ;
      RECT  1516800.0 434400.0 1527000.0 448200.0 ;
      RECT  1516800.0 462000.0 1527000.0 448200.0 ;
      RECT  1516800.0 462000.0 1527000.0 475800.0 ;
      RECT  1516800.0 489600.0 1527000.0 475800.0 ;
      RECT  1516800.0 489600.0 1527000.0 503400.0 ;
      RECT  1516800.0 517200.0 1527000.0 503400.0 ;
      RECT  1516800.0 517200.0 1527000.0 531000.0 ;
      RECT  1516800.0 544800.0 1527000.0 531000.0 ;
      RECT  1516800.0 544800.0 1527000.0 558600.0 ;
      RECT  1516800.0 572400.0 1527000.0 558600.0 ;
      RECT  1516800.0 572400.0 1527000.0 586200.0 ;
      RECT  1516800.0 600000.0 1527000.0 586200.0 ;
      RECT  1516800.0 600000.0 1527000.0 613800.0 ;
      RECT  1516800.0 627600.0 1527000.0 613800.0 ;
      RECT  1516800.0 627600.0 1527000.0 641400.0 ;
      RECT  1516800.0 655200.0 1527000.0 641400.0 ;
      RECT  1516800.0 655200.0 1527000.0 669000.0 ;
      RECT  1516800.0 682800.0 1527000.0 669000.0 ;
      RECT  1516800.0 682800.0 1527000.0 696600.0 ;
      RECT  1516800.0 710400.0 1527000.0 696600.0 ;
      RECT  1516800.0 710400.0 1527000.0 724200.0 ;
      RECT  1516800.0 738000.0 1527000.0 724200.0 ;
      RECT  1516800.0 738000.0 1527000.0 751800.0 ;
      RECT  1516800.0 765600.0 1527000.0 751800.0 ;
      RECT  1516800.0 765600.0 1527000.0 779400.0 ;
      RECT  1516800.0 793200.0 1527000.0 779400.0 ;
      RECT  1516800.0 793200.0 1527000.0 807000.0 ;
      RECT  1516800.0 820800.0 1527000.0 807000.0 ;
      RECT  1516800.0 820800.0 1527000.0 834600.0 ;
      RECT  1516800.0 848400.0 1527000.0 834600.0 ;
      RECT  1516800.0 848400.0 1527000.0 862200.0 ;
      RECT  1516800.0 876000.0 1527000.0 862200.0 ;
      RECT  1516800.0 876000.0 1527000.0 889800.0 ;
      RECT  1516800.0 903600.0 1527000.0 889800.0 ;
      RECT  1516800.0 903600.0 1527000.0 917400.0 ;
      RECT  1516800.0 931200.0 1527000.0 917400.0 ;
      RECT  1516800.0 931200.0 1527000.0 945000.0 ;
      RECT  1516800.0 958800.0 1527000.0 945000.0 ;
      RECT  1516800.0 958800.0 1527000.0 972600.0 ;
      RECT  1516800.0 986400.0 1527000.0 972600.0 ;
      RECT  1516800.0 986400.0 1527000.0 1000200.0 ;
      RECT  1516800.0 1014000.0 1527000.0 1000200.0 ;
      RECT  1516800.0 1014000.0 1527000.0 1027800.0 ;
      RECT  1516800.0 1041600.0 1527000.0 1027800.0 ;
      RECT  1516800.0 1041600.0 1527000.0 1055400.0 ;
      RECT  1516800.0 1069200.0 1527000.0 1055400.0 ;
      RECT  1516800.0 1069200.0 1527000.0 1083000.0 ;
      RECT  1516800.0 1096800.0 1527000.0 1083000.0 ;
      RECT  1516800.0 1096800.0 1527000.0 1110600.0 ;
      RECT  1516800.0 1124400.0 1527000.0 1110600.0 ;
      RECT  1516800.0 1124400.0 1527000.0 1138200.0 ;
      RECT  1516800.0 1152000.0 1527000.0 1138200.0 ;
      RECT  1516800.0 1152000.0 1527000.0 1165800.0 ;
      RECT  1516800.0 1179600.0 1527000.0 1165800.0 ;
      RECT  1516800.0 1179600.0 1527000.0 1193400.0 ;
      RECT  1516800.0 1207200.0 1527000.0 1193400.0 ;
      RECT  1516800.0 1207200.0 1527000.0 1221000.0 ;
      RECT  1516800.0 1234800.0 1527000.0 1221000.0 ;
      RECT  1516800.0 1234800.0 1527000.0 1248600.0 ;
      RECT  1516800.0 1262400.0 1527000.0 1248600.0 ;
      RECT  1516800.0 1262400.0 1527000.0 1276200.0 ;
      RECT  1516800.0 1290000.0 1527000.0 1276200.0 ;
      RECT  1516800.0 1290000.0 1527000.0 1303800.0 ;
      RECT  1516800.0 1317600.0 1527000.0 1303800.0 ;
      RECT  1516800.0 1317600.0 1527000.0 1331400.0 ;
      RECT  1516800.0 1345200.0 1527000.0 1331400.0 ;
      RECT  1516800.0 1345200.0 1527000.0 1359000.0 ;
      RECT  1516800.0 1372800.0 1527000.0 1359000.0 ;
      RECT  1516800.0 1372800.0 1527000.0 1386600.0 ;
      RECT  1516800.0 1400400.0 1527000.0 1386600.0 ;
      RECT  1516800.0 1400400.0 1527000.0 1414200.0 ;
      RECT  1516800.0 1428000.0 1527000.0 1414200.0 ;
      RECT  1516800.0 1428000.0 1527000.0 1441800.0 ;
      RECT  1516800.0 1455600.0 1527000.0 1441800.0 ;
      RECT  1516800.0 1455600.0 1527000.0 1469400.0 ;
      RECT  1516800.0 1483200.0 1527000.0 1469400.0 ;
      RECT  1516800.0 1483200.0 1527000.0 1497000.0 ;
      RECT  1516800.0 1510800.0 1527000.0 1497000.0 ;
      RECT  1516800.0 1510800.0 1527000.0 1524600.0 ;
      RECT  1516800.0 1538400.0 1527000.0 1524600.0 ;
      RECT  1516800.0 1538400.0 1527000.0 1552200.0 ;
      RECT  1516800.0 1566000.0 1527000.0 1552200.0 ;
      RECT  1516800.0 1566000.0 1527000.0 1579800.0 ;
      RECT  1516800.0 1593600.0 1527000.0 1579800.0 ;
      RECT  1516800.0 1593600.0 1527000.0 1607400.0 ;
      RECT  1516800.0 1621200.0 1527000.0 1607400.0 ;
      RECT  1516800.0 1621200.0 1527000.0 1635000.0 ;
      RECT  1516800.0 1648800.0 1527000.0 1635000.0 ;
      RECT  1516800.0 1648800.0 1527000.0 1662600.0 ;
      RECT  1516800.0 1676400.0 1527000.0 1662600.0 ;
      RECT  1516800.0 1676400.0 1527000.0 1690200.0 ;
      RECT  1516800.0 1704000.0 1527000.0 1690200.0 ;
      RECT  1516800.0 1704000.0 1527000.0 1717800.0 ;
      RECT  1516800.0 1731600.0 1527000.0 1717800.0 ;
      RECT  1516800.0 1731600.0 1527000.0 1745400.0 ;
      RECT  1516800.0 1759200.0 1527000.0 1745400.0 ;
      RECT  1516800.0 1759200.0 1527000.0 1773000.0 ;
      RECT  1516800.0 1786800.0 1527000.0 1773000.0 ;
      RECT  1516800.0 1786800.0 1527000.0 1800600.0 ;
      RECT  1516800.0 1814400.0 1527000.0 1800600.0 ;
      RECT  1516800.0 1814400.0 1527000.0 1828200.0 ;
      RECT  1516800.0 1842000.0 1527000.0 1828200.0 ;
      RECT  1516800.0 1842000.0 1527000.0 1855800.0 ;
      RECT  1516800.0 1869600.0 1527000.0 1855800.0 ;
      RECT  1516800.0 1869600.0 1527000.0 1883400.0 ;
      RECT  1516800.0 1897200.0 1527000.0 1883400.0 ;
      RECT  1516800.0 1897200.0 1527000.0 1911000.0 ;
      RECT  1516800.0 1924800.0 1527000.0 1911000.0 ;
      RECT  1516800.0 1924800.0 1527000.0 1938600.0 ;
      RECT  1516800.0 1952400.0 1527000.0 1938600.0 ;
      RECT  1516800.0 1952400.0 1527000.0 1966200.0 ;
      RECT  1516800.0 1980000.0 1527000.0 1966200.0 ;
      RECT  1516800.0 1980000.0 1527000.0 1993800.0 ;
      RECT  1516800.0 2007600.0 1527000.0 1993800.0 ;
      RECT  1516800.0 2007600.0 1527000.0 2021400.0 ;
      RECT  1516800.0 2035200.0 1527000.0 2021400.0 ;
      RECT  1516800.0 2035200.0 1527000.0 2049000.0 ;
      RECT  1516800.0 2062800.0 1527000.0 2049000.0 ;
      RECT  1516800.0 2062800.0 1527000.0 2076600.0 ;
      RECT  1516800.0 2090400.0 1527000.0 2076600.0 ;
      RECT  1516800.0 2090400.0 1527000.0 2104200.0 ;
      RECT  1516800.0 2118000.0 1527000.0 2104200.0 ;
      RECT  1516800.0 2118000.0 1527000.0 2131800.0 ;
      RECT  1516800.0 2145600.0 1527000.0 2131800.0 ;
      RECT  220800.0 380700.0 1527600.0 381900.0 ;
      RECT  220800.0 404100.0 1527600.0 405300.0 ;
      RECT  220800.0 408300.0 1527600.0 409500.0 ;
      RECT  220800.0 431700.0 1527600.0 432900.0 ;
      RECT  220800.0 435900.0 1527600.0 437100.0 ;
      RECT  220800.0 459300.0 1527600.0 460500.0 ;
      RECT  220800.0 463500.0 1527600.0 464700.0 ;
      RECT  220800.0 486900.0 1527600.0 488100.0 ;
      RECT  220800.0 491100.0 1527600.0 492300.0 ;
      RECT  220800.0 514500.0 1527600.0 515700.0 ;
      RECT  220800.0 518700.0 1527600.0 519900.0 ;
      RECT  220800.0 542100.0 1527600.0 543300.0 ;
      RECT  220800.0 546300.0 1527600.0 547500.0 ;
      RECT  220800.0 569700.0 1527600.0 570900.0 ;
      RECT  220800.0 573900.0 1527600.0 575100.0 ;
      RECT  220800.0 597300.0 1527600.0 598500.0 ;
      RECT  220800.0 601500.0 1527600.0 602700.0 ;
      RECT  220800.0 624900.0 1527600.0 626100.0 ;
      RECT  220800.0 629100.0 1527600.0 630300.0 ;
      RECT  220800.0 652500.0 1527600.0 653700.0 ;
      RECT  220800.0 656700.0 1527600.0 657900.0 ;
      RECT  220800.0 680100.0 1527600.0 681300.0 ;
      RECT  220800.0 684300.0 1527600.0 685500.0 ;
      RECT  220800.0 707700.0 1527600.0 708900.0 ;
      RECT  220800.0 711900.0 1527600.0 713100.0 ;
      RECT  220800.0 735300.0 1527600.0 736500.0 ;
      RECT  220800.0 739500.0 1527600.0 740700.0 ;
      RECT  220800.0 762900.0 1527600.0 764100.0 ;
      RECT  220800.0 767100.0 1527600.0 768300.0 ;
      RECT  220800.0 790500.0 1527600.0 791700.0 ;
      RECT  220800.0 794700.0 1527600.0 795900.0 ;
      RECT  220800.0 818100.0 1527600.0 819300.0 ;
      RECT  220800.0 822300.0 1527600.0 823500.0 ;
      RECT  220800.0 845700.0 1527600.0 846900.0 ;
      RECT  220800.0 849900.0 1527600.0 851100.0 ;
      RECT  220800.0 873300.0 1527600.0 874500.0 ;
      RECT  220800.0 877500.0 1527600.0 878700.0 ;
      RECT  220800.0 900900.0 1527600.0 902100.0 ;
      RECT  220800.0 905100.0 1527600.0 906300.0 ;
      RECT  220800.0 928500.0 1527600.0 929700.0 ;
      RECT  220800.0 932700.0 1527600.0 933900.0 ;
      RECT  220800.0 956100.0 1527600.0 957300.0 ;
      RECT  220800.0 960300.0 1527600.0 961500.0 ;
      RECT  220800.0 983700.0 1527600.0 984900.0 ;
      RECT  220800.0 987900.0 1527600.0 989100.0 ;
      RECT  220800.0 1011300.0 1527600.0 1012500.0 ;
      RECT  220800.0 1015500.0 1527600.0 1016700.0 ;
      RECT  220800.0 1038900.0 1527600.0 1040100.0 ;
      RECT  220800.0 1043100.0 1527600.0 1044300.0 ;
      RECT  220800.0 1066500.0 1527600.0 1067700.0 ;
      RECT  220800.0 1070700.0 1527600.0 1071900.0 ;
      RECT  220800.0 1094100.0 1527600.0 1095300.0 ;
      RECT  220800.0 1098300.0 1527600.0 1099500.0 ;
      RECT  220800.0 1121700.0 1527600.0 1122900.0 ;
      RECT  220800.0 1125900.0 1527600.0 1127100.0 ;
      RECT  220800.0 1149300.0 1527600.0 1150500.0 ;
      RECT  220800.0 1153500.0 1527600.0 1154700.0 ;
      RECT  220800.0 1176900.0 1527600.0 1178100.0 ;
      RECT  220800.0 1181100.0 1527600.0 1182300.0 ;
      RECT  220800.0 1204500.0 1527600.0 1205700.0 ;
      RECT  220800.0 1208700.0 1527600.0 1209900.0 ;
      RECT  220800.0 1232100.0 1527600.0 1233300.0 ;
      RECT  220800.0 1236300.0 1527600.0 1237500.0 ;
      RECT  220800.0 1259700.0 1527600.0 1260900.0 ;
      RECT  220800.0 1263900.0 1527600.0 1265100.0 ;
      RECT  220800.0 1287300.0 1527600.0 1288500.0 ;
      RECT  220800.0 1291500.0 1527600.0 1292700.0 ;
      RECT  220800.0 1314900.0 1527600.0 1316100.0 ;
      RECT  220800.0 1319100.0 1527600.0 1320300.0 ;
      RECT  220800.0 1342500.0 1527600.0 1343700.0 ;
      RECT  220800.0 1346700.0 1527600.0 1347900.0 ;
      RECT  220800.0 1370100.0 1527600.0 1371300.0 ;
      RECT  220800.0 1374300.0 1527600.0 1375500.0 ;
      RECT  220800.0 1397700.0 1527600.0 1398900.0 ;
      RECT  220800.0 1401900.0 1527600.0 1403100.0 ;
      RECT  220800.0 1425300.0 1527600.0 1426500.0 ;
      RECT  220800.0 1429500.0 1527600.0 1430700.0 ;
      RECT  220800.0 1452900.0 1527600.0 1454100.0 ;
      RECT  220800.0 1457100.0 1527600.0 1458300.0 ;
      RECT  220800.0 1480500.0 1527600.0 1481700.0 ;
      RECT  220800.0 1484700.0 1527600.0 1485900.0 ;
      RECT  220800.0 1508100.0 1527600.0 1509300.0 ;
      RECT  220800.0 1512300.0 1527600.0 1513500.0 ;
      RECT  220800.0 1535700.0 1527600.0 1536900.0 ;
      RECT  220800.0 1539900.0 1527600.0 1541100.0 ;
      RECT  220800.0 1563300.0 1527600.0 1564500.0 ;
      RECT  220800.0 1567500.0 1527600.0 1568700.0 ;
      RECT  220800.0 1590900.0 1527600.0 1592100.0 ;
      RECT  220800.0 1595100.0 1527600.0 1596300.0 ;
      RECT  220800.0 1618500.0 1527600.0 1619700.0 ;
      RECT  220800.0 1622700.0 1527600.0 1623900.0 ;
      RECT  220800.0 1646100.0 1527600.0 1647300.0 ;
      RECT  220800.0 1650300.0 1527600.0 1651500.0 ;
      RECT  220800.0 1673700.0 1527600.0 1674900.0 ;
      RECT  220800.0 1677900.0 1527600.0 1679100.0 ;
      RECT  220800.0 1701300.0 1527600.0 1702500.0 ;
      RECT  220800.0 1705500.0 1527600.0 1706700.0 ;
      RECT  220800.0 1728900.0 1527600.0 1730100.0 ;
      RECT  220800.0 1733100.0 1527600.0 1734300.0 ;
      RECT  220800.0 1756500.0 1527600.0 1757700.0 ;
      RECT  220800.0 1760700.0 1527600.0 1761900.0 ;
      RECT  220800.0 1784100.0 1527600.0 1785300.0 ;
      RECT  220800.0 1788300.0 1527600.0 1789500.0 ;
      RECT  220800.0 1811700.0 1527600.0 1812900.0 ;
      RECT  220800.0 1815900.0 1527600.0 1817100.0 ;
      RECT  220800.0 1839300.0 1527600.0 1840500.0 ;
      RECT  220800.0 1843500.0 1527600.0 1844700.0 ;
      RECT  220800.0 1866900.0 1527600.0 1868100.0 ;
      RECT  220800.0 1871100.0 1527600.0 1872300.0 ;
      RECT  220800.0 1894500.0 1527600.0 1895700.0 ;
      RECT  220800.0 1898700.0 1527600.0 1899900.0 ;
      RECT  220800.0 1922100.0 1527600.0 1923300.0 ;
      RECT  220800.0 1926300.0 1527600.0 1927500.0 ;
      RECT  220800.0 1949700.0 1527600.0 1950900.0 ;
      RECT  220800.0 1953900.0 1527600.0 1955100.0 ;
      RECT  220800.0 1977300.0 1527600.0 1978500.0 ;
      RECT  220800.0 1981500.0 1527600.0 1982700.0 ;
      RECT  220800.0 2004900.0 1527600.0 2006100.0 ;
      RECT  220800.0 2009100.0 1527600.0 2010300.0 ;
      RECT  220800.0 2032500.0 1527600.0 2033700.0 ;
      RECT  220800.0 2036700.0 1527600.0 2037900.0 ;
      RECT  220800.0 2060100.0 1527600.0 2061300.0 ;
      RECT  220800.0 2064300.0 1527600.0 2065500.0 ;
      RECT  220800.0 2087700.0 1527600.0 2088900.0 ;
      RECT  220800.0 2091900.0 1527600.0 2093100.0 ;
      RECT  220800.0 2115300.0 1527600.0 2116500.0 ;
      RECT  220800.0 2119500.0 1527600.0 2120700.0 ;
      RECT  220800.0 2142900.0 1527600.0 2144100.0 ;
      RECT  220800.0 392400.0 1527600.0 393300.0 ;
      RECT  220800.0 420000.0 1527600.0 420900.0 ;
      RECT  220800.0 447600.0 1527600.0 448500.0 ;
      RECT  220800.0 475200.0 1527600.0 476100.0 ;
      RECT  220800.0 502800.0 1527600.0 503700.0 ;
      RECT  220800.0 530400.0 1527600.0 531300.0 ;
      RECT  220800.0 558000.0 1527600.0 558900.0 ;
      RECT  220800.0 585600.0 1527600.0 586500.0 ;
      RECT  220800.0 613200.0 1527600.0 614100.0 ;
      RECT  220800.0 640800.0 1527600.0 641700.0 ;
      RECT  220800.0 668400.0 1527600.0 669300.0 ;
      RECT  220800.0 696000.0 1527600.0 696900.0 ;
      RECT  220800.0 723600.0 1527600.0 724500.0 ;
      RECT  220800.0 751200.0 1527600.0 752100.0 ;
      RECT  220800.0 778800.0 1527600.0 779700.0 ;
      RECT  220800.0 806400.0 1527600.0 807300.0 ;
      RECT  220800.0 834000.0 1527600.0 834900.0 ;
      RECT  220800.0 861600.0 1527600.0 862500.0 ;
      RECT  220800.0 889200.0 1527600.0 890100.0 ;
      RECT  220800.0 916800.0 1527600.0 917700.0 ;
      RECT  220800.0 944400.0 1527600.0 945300.0 ;
      RECT  220800.0 972000.0 1527600.0 972900.0 ;
      RECT  220800.0 999600.0 1527600.0 1000500.0 ;
      RECT  220800.0 1027200.0 1527600.0 1028100.0 ;
      RECT  220800.0 1054800.0 1527600.0 1055700.0 ;
      RECT  220800.0 1082400.0 1527600.0 1083300.0 ;
      RECT  220800.0 1110000.0 1527600.0 1110900.0 ;
      RECT  220800.0 1137600.0 1527600.0 1138500.0 ;
      RECT  220800.0 1165200.0 1527600.0 1166100.0 ;
      RECT  220800.0 1192800.0 1527600.0 1193700.0 ;
      RECT  220800.0 1220400.0 1527600.0 1221300.0 ;
      RECT  220800.0 1248000.0 1527600.0 1248900.0 ;
      RECT  220800.0 1275600.0 1527600.0 1276500.0 ;
      RECT  220800.0 1303200.0 1527600.0 1304100.0 ;
      RECT  220800.0 1330800.0 1527600.0 1331700.0 ;
      RECT  220800.0 1358400.0 1527600.0 1359300.0 ;
      RECT  220800.0 1386000.0 1527600.0 1386900.0 ;
      RECT  220800.0 1413600.0 1527600.0 1414500.0 ;
      RECT  220800.0 1441200.0 1527600.0 1442100.0 ;
      RECT  220800.0 1468800.0 1527600.0 1469700.0 ;
      RECT  220800.0 1496400.0 1527600.0 1497300.0 ;
      RECT  220800.0 1524000.0 1527600.0 1524900.0 ;
      RECT  220800.0 1551600.0 1527600.0 1552500.0 ;
      RECT  220800.0 1579200.0 1527600.0 1580100.0 ;
      RECT  220800.0 1606800.0 1527600.0 1607700.0 ;
      RECT  220800.0 1634400.0 1527600.0 1635300.0 ;
      RECT  220800.0 1662000.0 1527600.0 1662900.0 ;
      RECT  220800.0 1689600.0 1527600.0 1690500.0 ;
      RECT  220800.0 1717200.0 1527600.0 1718100.0 ;
      RECT  220800.0 1744800.0 1527600.0 1745700.0 ;
      RECT  220800.0 1772400.0 1527600.0 1773300.0 ;
      RECT  220800.0 1800000.0 1527600.0 1800900.0 ;
      RECT  220800.0 1827600.0 1527600.0 1828500.0 ;
      RECT  220800.0 1855200.0 1527600.0 1856100.0 ;
      RECT  220800.0 1882800.0 1527600.0 1883700.0 ;
      RECT  220800.0 1910400.0 1527600.0 1911300.0 ;
      RECT  220800.0 1938000.0 1527600.0 1938900.0 ;
      RECT  220800.0 1965600.0 1527600.0 1966500.0 ;
      RECT  220800.0 1993200.0 1527600.0 1994100.0 ;
      RECT  220800.0 2020800.0 1527600.0 2021700.0 ;
      RECT  220800.0 2048400.0 1527600.0 2049300.0 ;
      RECT  220800.0 2076000.0 1527600.0 2076900.0 ;
      RECT  220800.0 2103600.0 1527600.0 2104500.0 ;
      RECT  220800.0 2131200.0 1527600.0 2132100.0 ;
      RECT  226800.0 2158800.0 228000.0 2166000.0 ;
      RECT  224400.0 2151600.0 225600.0 2152800.0 ;
      RECT  226800.0 2151600.0 228000.0 2152800.0 ;
      RECT  226800.0 2151600.0 228000.0 2152800.0 ;
      RECT  224400.0 2151600.0 225600.0 2152800.0 ;
      RECT  224400.0 2158800.0 225600.0 2160000.0 ;
      RECT  226800.0 2158800.0 228000.0 2160000.0 ;
      RECT  226800.0 2158800.0 228000.0 2160000.0 ;
      RECT  224400.0 2158800.0 225600.0 2160000.0 ;
      RECT  226800.0 2158800.0 228000.0 2160000.0 ;
      RECT  229200.0 2158800.0 230400.0 2160000.0 ;
      RECT  229200.0 2158800.0 230400.0 2160000.0 ;
      RECT  226800.0 2158800.0 228000.0 2160000.0 ;
      RECT  226500.0 2153850.0 225300.0 2155050.0 ;
      RECT  226800.0 2164200.0 228000.0 2165400.0 ;
      RECT  224400.0 2151600.0 225600.0 2152800.0 ;
      RECT  226800.0 2151600.0 228000.0 2152800.0 ;
      RECT  224400.0 2158800.0 225600.0 2160000.0 ;
      RECT  229200.0 2158800.0 230400.0 2160000.0 ;
      RECT  221400.0 2154000.0 231600.0 2154900.0 ;
      RECT  221400.0 2165100.0 231600.0 2166000.0 ;
      RECT  237000.0 2158800.0 238200.0 2166000.0 ;
      RECT  234600.0 2151600.0 235800.0 2152800.0 ;
      RECT  237000.0 2151600.0 238200.0 2152800.0 ;
      RECT  237000.0 2151600.0 238200.0 2152800.0 ;
      RECT  234600.0 2151600.0 235800.0 2152800.0 ;
      RECT  234600.0 2158800.0 235800.0 2160000.0 ;
      RECT  237000.0 2158800.0 238200.0 2160000.0 ;
      RECT  237000.0 2158800.0 238200.0 2160000.0 ;
      RECT  234600.0 2158800.0 235800.0 2160000.0 ;
      RECT  237000.0 2158800.0 238200.0 2160000.0 ;
      RECT  239400.0 2158800.0 240600.0 2160000.0 ;
      RECT  239400.0 2158800.0 240600.0 2160000.0 ;
      RECT  237000.0 2158800.0 238200.0 2160000.0 ;
      RECT  236700.0 2153850.0 235500.0 2155050.0 ;
      RECT  237000.0 2164200.0 238200.0 2165400.0 ;
      RECT  234600.0 2151600.0 235800.0 2152800.0 ;
      RECT  237000.0 2151600.0 238200.0 2152800.0 ;
      RECT  234600.0 2158800.0 235800.0 2160000.0 ;
      RECT  239400.0 2158800.0 240600.0 2160000.0 ;
      RECT  231600.0 2154000.0 241800.0 2154900.0 ;
      RECT  231600.0 2165100.0 241800.0 2166000.0 ;
      RECT  247200.0 2158800.0 248400.0 2166000.0 ;
      RECT  244800.0 2151600.0 246000.0 2152800.0 ;
      RECT  247200.0 2151600.0 248400.0 2152800.0 ;
      RECT  247200.0 2151600.0 248400.0 2152800.0 ;
      RECT  244800.0 2151600.0 246000.0 2152800.0 ;
      RECT  244800.0 2158800.0 246000.0 2160000.0 ;
      RECT  247200.0 2158800.0 248400.0 2160000.0 ;
      RECT  247200.0 2158800.0 248400.0 2160000.0 ;
      RECT  244800.0 2158800.0 246000.0 2160000.0 ;
      RECT  247200.0 2158800.0 248400.0 2160000.0 ;
      RECT  249600.0 2158800.0 250800.0 2160000.0 ;
      RECT  249600.0 2158800.0 250800.0 2160000.0 ;
      RECT  247200.0 2158800.0 248400.0 2160000.0 ;
      RECT  246900.0 2153850.0 245700.0 2155050.0 ;
      RECT  247200.0 2164200.0 248400.0 2165400.0 ;
      RECT  244800.0 2151600.0 246000.0 2152800.0 ;
      RECT  247200.0 2151600.0 248400.0 2152800.0 ;
      RECT  244800.0 2158800.0 246000.0 2160000.0 ;
      RECT  249600.0 2158800.0 250800.0 2160000.0 ;
      RECT  241800.0 2154000.0 252000.0 2154900.0 ;
      RECT  241800.0 2165100.0 252000.0 2166000.0 ;
      RECT  257400.0 2158800.0 258600.0 2166000.0 ;
      RECT  255000.0 2151600.0 256200.0 2152800.0 ;
      RECT  257400.0 2151600.0 258600.0 2152800.0 ;
      RECT  257400.0 2151600.0 258600.0 2152800.0 ;
      RECT  255000.0 2151600.0 256200.0 2152800.0 ;
      RECT  255000.0 2158800.0 256200.0 2160000.0 ;
      RECT  257400.0 2158800.0 258600.0 2160000.0 ;
      RECT  257400.0 2158800.0 258600.0 2160000.0 ;
      RECT  255000.0 2158800.0 256200.0 2160000.0 ;
      RECT  257400.0 2158800.0 258600.0 2160000.0 ;
      RECT  259800.0 2158800.0 261000.0 2160000.0 ;
      RECT  259800.0 2158800.0 261000.0 2160000.0 ;
      RECT  257400.0 2158800.0 258600.0 2160000.0 ;
      RECT  257100.0 2153850.0 255900.0 2155050.0 ;
      RECT  257400.0 2164200.0 258600.0 2165400.0 ;
      RECT  255000.0 2151600.0 256200.0 2152800.0 ;
      RECT  257400.0 2151600.0 258600.0 2152800.0 ;
      RECT  255000.0 2158800.0 256200.0 2160000.0 ;
      RECT  259800.0 2158800.0 261000.0 2160000.0 ;
      RECT  252000.0 2154000.0 262200.0 2154900.0 ;
      RECT  252000.0 2165100.0 262200.0 2166000.0 ;
      RECT  267600.0 2158800.0 268800.0 2166000.0 ;
      RECT  265200.0 2151600.0 266400.0 2152800.0 ;
      RECT  267600.0 2151600.0 268800.0 2152800.0 ;
      RECT  267600.0 2151600.0 268800.0 2152800.0 ;
      RECT  265200.0 2151600.0 266400.0 2152800.0 ;
      RECT  265200.0 2158800.0 266400.0 2160000.0 ;
      RECT  267600.0 2158800.0 268800.0 2160000.0 ;
      RECT  267600.0 2158800.0 268800.0 2160000.0 ;
      RECT  265200.0 2158800.0 266400.0 2160000.0 ;
      RECT  267600.0 2158800.0 268800.0 2160000.0 ;
      RECT  270000.0 2158800.0 271200.0 2160000.0 ;
      RECT  270000.0 2158800.0 271200.0 2160000.0 ;
      RECT  267600.0 2158800.0 268800.0 2160000.0 ;
      RECT  267300.0 2153850.0 266100.0 2155050.0 ;
      RECT  267600.0 2164200.0 268800.0 2165400.0 ;
      RECT  265200.0 2151600.0 266400.0 2152800.0 ;
      RECT  267600.0 2151600.0 268800.0 2152800.0 ;
      RECT  265200.0 2158800.0 266400.0 2160000.0 ;
      RECT  270000.0 2158800.0 271200.0 2160000.0 ;
      RECT  262200.0 2154000.0 272400.0 2154900.0 ;
      RECT  262200.0 2165100.0 272400.0 2166000.0 ;
      RECT  277800.0 2158800.0 279000.0 2166000.0 ;
      RECT  275400.0 2151600.0 276600.0 2152800.0 ;
      RECT  277800.0 2151600.0 279000.0 2152800.0 ;
      RECT  277800.0 2151600.0 279000.0 2152800.0 ;
      RECT  275400.0 2151600.0 276600.0 2152800.0 ;
      RECT  275400.0 2158800.0 276600.0 2160000.0 ;
      RECT  277800.0 2158800.0 279000.0 2160000.0 ;
      RECT  277800.0 2158800.0 279000.0 2160000.0 ;
      RECT  275400.0 2158800.0 276600.0 2160000.0 ;
      RECT  277800.0 2158800.0 279000.0 2160000.0 ;
      RECT  280200.0 2158800.0 281400.0 2160000.0 ;
      RECT  280200.0 2158800.0 281400.0 2160000.0 ;
      RECT  277800.0 2158800.0 279000.0 2160000.0 ;
      RECT  277500.0 2153850.0 276300.0 2155050.0 ;
      RECT  277800.0 2164200.0 279000.0 2165400.0 ;
      RECT  275400.0 2151600.0 276600.0 2152800.0 ;
      RECT  277800.0 2151600.0 279000.0 2152800.0 ;
      RECT  275400.0 2158800.0 276600.0 2160000.0 ;
      RECT  280200.0 2158800.0 281400.0 2160000.0 ;
      RECT  272400.0 2154000.0 282600.0 2154900.0 ;
      RECT  272400.0 2165100.0 282600.0 2166000.0 ;
      RECT  288000.0 2158800.0 289200.0 2166000.0 ;
      RECT  285600.0 2151600.0 286800.0 2152800.0 ;
      RECT  288000.0 2151600.0 289200.0 2152800.0 ;
      RECT  288000.0 2151600.0 289200.0 2152800.0 ;
      RECT  285600.0 2151600.0 286800.0 2152800.0 ;
      RECT  285600.0 2158800.0 286800.0 2160000.0 ;
      RECT  288000.0 2158800.0 289200.0 2160000.0 ;
      RECT  288000.0 2158800.0 289200.0 2160000.0 ;
      RECT  285600.0 2158800.0 286800.0 2160000.0 ;
      RECT  288000.0 2158800.0 289200.0 2160000.0 ;
      RECT  290400.0 2158800.0 291600.0 2160000.0 ;
      RECT  290400.0 2158800.0 291600.0 2160000.0 ;
      RECT  288000.0 2158800.0 289200.0 2160000.0 ;
      RECT  287700.0 2153850.0 286500.0 2155050.0 ;
      RECT  288000.0 2164200.0 289200.0 2165400.0 ;
      RECT  285600.0 2151600.0 286800.0 2152800.0 ;
      RECT  288000.0 2151600.0 289200.0 2152800.0 ;
      RECT  285600.0 2158800.0 286800.0 2160000.0 ;
      RECT  290400.0 2158800.0 291600.0 2160000.0 ;
      RECT  282600.0 2154000.0 292800.0 2154900.0 ;
      RECT  282600.0 2165100.0 292800.0 2166000.0 ;
      RECT  298200.0 2158800.0 299400.0 2166000.0 ;
      RECT  295800.0 2151600.0 297000.0 2152800.0 ;
      RECT  298200.0 2151600.0 299400.0 2152800.0 ;
      RECT  298200.0 2151600.0 299400.0 2152800.0 ;
      RECT  295800.0 2151600.0 297000.0 2152800.0 ;
      RECT  295800.0 2158800.0 297000.0 2160000.0 ;
      RECT  298200.0 2158800.0 299400.0 2160000.0 ;
      RECT  298200.0 2158800.0 299400.0 2160000.0 ;
      RECT  295800.0 2158800.0 297000.0 2160000.0 ;
      RECT  298200.0 2158800.0 299400.0 2160000.0 ;
      RECT  300600.0 2158800.0 301800.0 2160000.0 ;
      RECT  300600.0 2158800.0 301800.0 2160000.0 ;
      RECT  298200.0 2158800.0 299400.0 2160000.0 ;
      RECT  297900.0 2153850.0 296700.0 2155050.0 ;
      RECT  298200.0 2164200.0 299400.0 2165400.0 ;
      RECT  295800.0 2151600.0 297000.0 2152800.0 ;
      RECT  298200.0 2151600.0 299400.0 2152800.0 ;
      RECT  295800.0 2158800.0 297000.0 2160000.0 ;
      RECT  300600.0 2158800.0 301800.0 2160000.0 ;
      RECT  292800.0 2154000.0 303000.0 2154900.0 ;
      RECT  292800.0 2165100.0 303000.0 2166000.0 ;
      RECT  308400.0 2158800.0 309600.0 2166000.0 ;
      RECT  306000.0 2151600.0 307200.0 2152800.0 ;
      RECT  308400.0 2151600.0 309600.0 2152800.0 ;
      RECT  308400.0 2151600.0 309600.0 2152800.0 ;
      RECT  306000.0 2151600.0 307200.0 2152800.0 ;
      RECT  306000.0 2158800.0 307200.0 2160000.0 ;
      RECT  308400.0 2158800.0 309600.0 2160000.0 ;
      RECT  308400.0 2158800.0 309600.0 2160000.0 ;
      RECT  306000.0 2158800.0 307200.0 2160000.0 ;
      RECT  308400.0 2158800.0 309600.0 2160000.0 ;
      RECT  310800.0 2158800.0 312000.0 2160000.0 ;
      RECT  310800.0 2158800.0 312000.0 2160000.0 ;
      RECT  308400.0 2158800.0 309600.0 2160000.0 ;
      RECT  308100.0 2153850.0 306900.0 2155050.0 ;
      RECT  308400.0 2164200.0 309600.0 2165400.0 ;
      RECT  306000.0 2151600.0 307200.0 2152800.0 ;
      RECT  308400.0 2151600.0 309600.0 2152800.0 ;
      RECT  306000.0 2158800.0 307200.0 2160000.0 ;
      RECT  310800.0 2158800.0 312000.0 2160000.0 ;
      RECT  303000.0 2154000.0 313200.0 2154900.0 ;
      RECT  303000.0 2165100.0 313200.0 2166000.0 ;
      RECT  318600.0 2158800.0 319800.0 2166000.0 ;
      RECT  316200.0 2151600.0 317400.0 2152800.0 ;
      RECT  318600.0 2151600.0 319800.0 2152800.0 ;
      RECT  318600.0 2151600.0 319800.0 2152800.0 ;
      RECT  316200.0 2151600.0 317400.0 2152800.0 ;
      RECT  316200.0 2158800.0 317400.0 2160000.0 ;
      RECT  318600.0 2158800.0 319800.0 2160000.0 ;
      RECT  318600.0 2158800.0 319800.0 2160000.0 ;
      RECT  316200.0 2158800.0 317400.0 2160000.0 ;
      RECT  318600.0 2158800.0 319800.0 2160000.0 ;
      RECT  321000.0 2158800.0 322200.0 2160000.0 ;
      RECT  321000.0 2158800.0 322200.0 2160000.0 ;
      RECT  318600.0 2158800.0 319800.0 2160000.0 ;
      RECT  318300.0 2153850.0 317100.0 2155050.0 ;
      RECT  318600.0 2164200.0 319800.0 2165400.0 ;
      RECT  316200.0 2151600.0 317400.0 2152800.0 ;
      RECT  318600.0 2151600.0 319800.0 2152800.0 ;
      RECT  316200.0 2158800.0 317400.0 2160000.0 ;
      RECT  321000.0 2158800.0 322200.0 2160000.0 ;
      RECT  313200.0 2154000.0 323400.0 2154900.0 ;
      RECT  313200.0 2165100.0 323400.0 2166000.0 ;
      RECT  328800.0 2158800.0 330000.0 2166000.0 ;
      RECT  326400.0 2151600.0 327600.0 2152800.0 ;
      RECT  328800.0 2151600.0 330000.0 2152800.0 ;
      RECT  328800.0 2151600.0 330000.0 2152800.0 ;
      RECT  326400.0 2151600.0 327600.0 2152800.0 ;
      RECT  326400.0 2158800.0 327600.0 2160000.0 ;
      RECT  328800.0 2158800.0 330000.0 2160000.0 ;
      RECT  328800.0 2158800.0 330000.0 2160000.0 ;
      RECT  326400.0 2158800.0 327600.0 2160000.0 ;
      RECT  328800.0 2158800.0 330000.0 2160000.0 ;
      RECT  331200.0 2158800.0 332400.0 2160000.0 ;
      RECT  331200.0 2158800.0 332400.0 2160000.0 ;
      RECT  328800.0 2158800.0 330000.0 2160000.0 ;
      RECT  328500.0 2153850.0 327300.0 2155050.0 ;
      RECT  328800.0 2164200.0 330000.0 2165400.0 ;
      RECT  326400.0 2151600.0 327600.0 2152800.0 ;
      RECT  328800.0 2151600.0 330000.0 2152800.0 ;
      RECT  326400.0 2158800.0 327600.0 2160000.0 ;
      RECT  331200.0 2158800.0 332400.0 2160000.0 ;
      RECT  323400.0 2154000.0 333600.0 2154900.0 ;
      RECT  323400.0 2165100.0 333600.0 2166000.0 ;
      RECT  339000.0 2158800.0 340200.0 2166000.0 ;
      RECT  336600.0 2151600.0 337800.0 2152800.0 ;
      RECT  339000.0 2151600.0 340200.0 2152800.0 ;
      RECT  339000.0 2151600.0 340200.0 2152800.0 ;
      RECT  336600.0 2151600.0 337800.0 2152800.0 ;
      RECT  336600.0 2158800.0 337800.0 2160000.0 ;
      RECT  339000.0 2158800.0 340200.0 2160000.0 ;
      RECT  339000.0 2158800.0 340200.0 2160000.0 ;
      RECT  336600.0 2158800.0 337800.0 2160000.0 ;
      RECT  339000.0 2158800.0 340200.0 2160000.0 ;
      RECT  341400.0 2158800.0 342600.0 2160000.0 ;
      RECT  341400.0 2158800.0 342600.0 2160000.0 ;
      RECT  339000.0 2158800.0 340200.0 2160000.0 ;
      RECT  338700.0 2153850.0 337500.0 2155050.0 ;
      RECT  339000.0 2164200.0 340200.0 2165400.0 ;
      RECT  336600.0 2151600.0 337800.0 2152800.0 ;
      RECT  339000.0 2151600.0 340200.0 2152800.0 ;
      RECT  336600.0 2158800.0 337800.0 2160000.0 ;
      RECT  341400.0 2158800.0 342600.0 2160000.0 ;
      RECT  333600.0 2154000.0 343800.0 2154900.0 ;
      RECT  333600.0 2165100.0 343800.0 2166000.0 ;
      RECT  349200.0 2158800.0 350400.0 2166000.0 ;
      RECT  346800.0 2151600.0 348000.0 2152800.0 ;
      RECT  349200.0 2151600.0 350400.0 2152800.0 ;
      RECT  349200.0 2151600.0 350400.0 2152800.0 ;
      RECT  346800.0 2151600.0 348000.0 2152800.0 ;
      RECT  346800.0 2158800.0 348000.0 2160000.0 ;
      RECT  349200.0 2158800.0 350400.0 2160000.0 ;
      RECT  349200.0 2158800.0 350400.0 2160000.0 ;
      RECT  346800.0 2158800.0 348000.0 2160000.0 ;
      RECT  349200.0 2158800.0 350400.0 2160000.0 ;
      RECT  351600.0 2158800.0 352800.0 2160000.0 ;
      RECT  351600.0 2158800.0 352800.0 2160000.0 ;
      RECT  349200.0 2158800.0 350400.0 2160000.0 ;
      RECT  348900.0 2153850.0 347700.0 2155050.0 ;
      RECT  349200.0 2164200.0 350400.0 2165400.0 ;
      RECT  346800.0 2151600.0 348000.0 2152800.0 ;
      RECT  349200.0 2151600.0 350400.0 2152800.0 ;
      RECT  346800.0 2158800.0 348000.0 2160000.0 ;
      RECT  351600.0 2158800.0 352800.0 2160000.0 ;
      RECT  343800.0 2154000.0 354000.0 2154900.0 ;
      RECT  343800.0 2165100.0 354000.0 2166000.0 ;
      RECT  359400.0 2158800.0 360600.0 2166000.0 ;
      RECT  357000.0 2151600.0 358200.0 2152800.0 ;
      RECT  359400.0 2151600.0 360600.0 2152800.0 ;
      RECT  359400.0 2151600.0 360600.0 2152800.0 ;
      RECT  357000.0 2151600.0 358200.0 2152800.0 ;
      RECT  357000.0 2158800.0 358200.0 2160000.0 ;
      RECT  359400.0 2158800.0 360600.0 2160000.0 ;
      RECT  359400.0 2158800.0 360600.0 2160000.0 ;
      RECT  357000.0 2158800.0 358200.0 2160000.0 ;
      RECT  359400.0 2158800.0 360600.0 2160000.0 ;
      RECT  361800.0 2158800.0 363000.0 2160000.0 ;
      RECT  361800.0 2158800.0 363000.0 2160000.0 ;
      RECT  359400.0 2158800.0 360600.0 2160000.0 ;
      RECT  359100.0 2153850.0 357900.0 2155050.0 ;
      RECT  359400.0 2164200.0 360600.0 2165400.0 ;
      RECT  357000.0 2151600.0 358200.0 2152800.0 ;
      RECT  359400.0 2151600.0 360600.0 2152800.0 ;
      RECT  357000.0 2158800.0 358200.0 2160000.0 ;
      RECT  361800.0 2158800.0 363000.0 2160000.0 ;
      RECT  354000.0 2154000.0 364200.0 2154900.0 ;
      RECT  354000.0 2165100.0 364200.0 2166000.0 ;
      RECT  369600.0 2158800.0 370800.0 2166000.0 ;
      RECT  367200.0 2151600.0 368400.0 2152800.0 ;
      RECT  369600.0 2151600.0 370800.0 2152800.0 ;
      RECT  369600.0 2151600.0 370800.0 2152800.0 ;
      RECT  367200.0 2151600.0 368400.0 2152800.0 ;
      RECT  367200.0 2158800.0 368400.0 2160000.0 ;
      RECT  369600.0 2158800.0 370800.0 2160000.0 ;
      RECT  369600.0 2158800.0 370800.0 2160000.0 ;
      RECT  367200.0 2158800.0 368400.0 2160000.0 ;
      RECT  369600.0 2158800.0 370800.0 2160000.0 ;
      RECT  372000.0 2158800.0 373200.0 2160000.0 ;
      RECT  372000.0 2158800.0 373200.0 2160000.0 ;
      RECT  369600.0 2158800.0 370800.0 2160000.0 ;
      RECT  369300.0 2153850.0 368100.0 2155050.0 ;
      RECT  369600.0 2164200.0 370800.0 2165400.0 ;
      RECT  367200.0 2151600.0 368400.0 2152800.0 ;
      RECT  369600.0 2151600.0 370800.0 2152800.0 ;
      RECT  367200.0 2158800.0 368400.0 2160000.0 ;
      RECT  372000.0 2158800.0 373200.0 2160000.0 ;
      RECT  364200.0 2154000.0 374400.0 2154900.0 ;
      RECT  364200.0 2165100.0 374400.0 2166000.0 ;
      RECT  379800.0 2158800.0 381000.0 2166000.0 ;
      RECT  377400.0 2151600.0 378600.0 2152800.0 ;
      RECT  379800.0 2151600.0 381000.0 2152800.0 ;
      RECT  379800.0 2151600.0 381000.0 2152800.0 ;
      RECT  377400.0 2151600.0 378600.0 2152800.0 ;
      RECT  377400.0 2158800.0 378600.0 2160000.0 ;
      RECT  379800.0 2158800.0 381000.0 2160000.0 ;
      RECT  379800.0 2158800.0 381000.0 2160000.0 ;
      RECT  377400.0 2158800.0 378600.0 2160000.0 ;
      RECT  379800.0 2158800.0 381000.0 2160000.0 ;
      RECT  382200.0 2158800.0 383400.0 2160000.0 ;
      RECT  382200.0 2158800.0 383400.0 2160000.0 ;
      RECT  379800.0 2158800.0 381000.0 2160000.0 ;
      RECT  379500.0 2153850.0 378300.0 2155050.0 ;
      RECT  379800.0 2164200.0 381000.0 2165400.0 ;
      RECT  377400.0 2151600.0 378600.0 2152800.0 ;
      RECT  379800.0 2151600.0 381000.0 2152800.0 ;
      RECT  377400.0 2158800.0 378600.0 2160000.0 ;
      RECT  382200.0 2158800.0 383400.0 2160000.0 ;
      RECT  374400.0 2154000.0 384600.0 2154900.0 ;
      RECT  374400.0 2165100.0 384600.0 2166000.0 ;
      RECT  390000.0 2158800.0 391200.0 2166000.0 ;
      RECT  387600.0 2151600.0 388800.0 2152800.0 ;
      RECT  390000.0 2151600.0 391200.0 2152800.0 ;
      RECT  390000.0 2151600.0 391200.0 2152800.0 ;
      RECT  387600.0 2151600.0 388800.0 2152800.0 ;
      RECT  387600.0 2158800.0 388800.0 2160000.0 ;
      RECT  390000.0 2158800.0 391200.0 2160000.0 ;
      RECT  390000.0 2158800.0 391200.0 2160000.0 ;
      RECT  387600.0 2158800.0 388800.0 2160000.0 ;
      RECT  390000.0 2158800.0 391200.0 2160000.0 ;
      RECT  392400.0 2158800.0 393600.0 2160000.0 ;
      RECT  392400.0 2158800.0 393600.0 2160000.0 ;
      RECT  390000.0 2158800.0 391200.0 2160000.0 ;
      RECT  389700.0 2153850.0 388500.0 2155050.0 ;
      RECT  390000.0 2164200.0 391200.0 2165400.0 ;
      RECT  387600.0 2151600.0 388800.0 2152800.0 ;
      RECT  390000.0 2151600.0 391200.0 2152800.0 ;
      RECT  387600.0 2158800.0 388800.0 2160000.0 ;
      RECT  392400.0 2158800.0 393600.0 2160000.0 ;
      RECT  384600.0 2154000.0 394800.0 2154900.0 ;
      RECT  384600.0 2165100.0 394800.0 2166000.0 ;
      RECT  400200.0 2158800.0 401400.0 2166000.0 ;
      RECT  397800.0 2151600.0 399000.0 2152800.0 ;
      RECT  400200.0 2151600.0 401400.0 2152800.0 ;
      RECT  400200.0 2151600.0 401400.0 2152800.0 ;
      RECT  397800.0 2151600.0 399000.0 2152800.0 ;
      RECT  397800.0 2158800.0 399000.0 2160000.0 ;
      RECT  400200.0 2158800.0 401400.0 2160000.0 ;
      RECT  400200.0 2158800.0 401400.0 2160000.0 ;
      RECT  397800.0 2158800.0 399000.0 2160000.0 ;
      RECT  400200.0 2158800.0 401400.0 2160000.0 ;
      RECT  402600.0 2158800.0 403800.0 2160000.0 ;
      RECT  402600.0 2158800.0 403800.0 2160000.0 ;
      RECT  400200.0 2158800.0 401400.0 2160000.0 ;
      RECT  399900.0 2153850.0 398700.0 2155050.0 ;
      RECT  400200.0 2164200.0 401400.0 2165400.0 ;
      RECT  397800.0 2151600.0 399000.0 2152800.0 ;
      RECT  400200.0 2151600.0 401400.0 2152800.0 ;
      RECT  397800.0 2158800.0 399000.0 2160000.0 ;
      RECT  402600.0 2158800.0 403800.0 2160000.0 ;
      RECT  394800.0 2154000.0 405000.0 2154900.0 ;
      RECT  394800.0 2165100.0 405000.0 2166000.0 ;
      RECT  410400.0 2158800.0 411600.0 2166000.0 ;
      RECT  408000.0 2151600.0 409200.0 2152800.0 ;
      RECT  410400.0 2151600.0 411600.0 2152800.0 ;
      RECT  410400.0 2151600.0 411600.0 2152800.0 ;
      RECT  408000.0 2151600.0 409200.0 2152800.0 ;
      RECT  408000.0 2158800.0 409200.0 2160000.0 ;
      RECT  410400.0 2158800.0 411600.0 2160000.0 ;
      RECT  410400.0 2158800.0 411600.0 2160000.0 ;
      RECT  408000.0 2158800.0 409200.0 2160000.0 ;
      RECT  410400.0 2158800.0 411600.0 2160000.0 ;
      RECT  412800.0 2158800.0 414000.0 2160000.0 ;
      RECT  412800.0 2158800.0 414000.0 2160000.0 ;
      RECT  410400.0 2158800.0 411600.0 2160000.0 ;
      RECT  410100.0 2153850.0 408900.0 2155050.0 ;
      RECT  410400.0 2164200.0 411600.0 2165400.0 ;
      RECT  408000.0 2151600.0 409200.0 2152800.0 ;
      RECT  410400.0 2151600.0 411600.0 2152800.0 ;
      RECT  408000.0 2158800.0 409200.0 2160000.0 ;
      RECT  412800.0 2158800.0 414000.0 2160000.0 ;
      RECT  405000.0 2154000.0 415200.0 2154900.0 ;
      RECT  405000.0 2165100.0 415200.0 2166000.0 ;
      RECT  420600.0 2158800.0 421800.0 2166000.0 ;
      RECT  418200.0 2151600.0 419400.0 2152800.0 ;
      RECT  420600.0 2151600.0 421800.0 2152800.0 ;
      RECT  420600.0 2151600.0 421800.0 2152800.0 ;
      RECT  418200.0 2151600.0 419400.0 2152800.0 ;
      RECT  418200.0 2158800.0 419400.0 2160000.0 ;
      RECT  420600.0 2158800.0 421800.0 2160000.0 ;
      RECT  420600.0 2158800.0 421800.0 2160000.0 ;
      RECT  418200.0 2158800.0 419400.0 2160000.0 ;
      RECT  420600.0 2158800.0 421800.0 2160000.0 ;
      RECT  423000.0 2158800.0 424200.0 2160000.0 ;
      RECT  423000.0 2158800.0 424200.0 2160000.0 ;
      RECT  420600.0 2158800.0 421800.0 2160000.0 ;
      RECT  420300.0 2153850.0 419100.0 2155050.0 ;
      RECT  420600.0 2164200.0 421800.0 2165400.0 ;
      RECT  418200.0 2151600.0 419400.0 2152800.0 ;
      RECT  420600.0 2151600.0 421800.0 2152800.0 ;
      RECT  418200.0 2158800.0 419400.0 2160000.0 ;
      RECT  423000.0 2158800.0 424200.0 2160000.0 ;
      RECT  415200.0 2154000.0 425400.0 2154900.0 ;
      RECT  415200.0 2165100.0 425400.0 2166000.0 ;
      RECT  430800.0 2158800.0 432000.0 2166000.0 ;
      RECT  428400.0 2151600.0 429600.0 2152800.0 ;
      RECT  430800.0 2151600.0 432000.0 2152800.0 ;
      RECT  430800.0 2151600.0 432000.0 2152800.0 ;
      RECT  428400.0 2151600.0 429600.0 2152800.0 ;
      RECT  428400.0 2158800.0 429600.0 2160000.0 ;
      RECT  430800.0 2158800.0 432000.0 2160000.0 ;
      RECT  430800.0 2158800.0 432000.0 2160000.0 ;
      RECT  428400.0 2158800.0 429600.0 2160000.0 ;
      RECT  430800.0 2158800.0 432000.0 2160000.0 ;
      RECT  433200.0 2158800.0 434400.0 2160000.0 ;
      RECT  433200.0 2158800.0 434400.0 2160000.0 ;
      RECT  430800.0 2158800.0 432000.0 2160000.0 ;
      RECT  430500.0 2153850.0 429300.0 2155050.0 ;
      RECT  430800.0 2164200.0 432000.0 2165400.0 ;
      RECT  428400.0 2151600.0 429600.0 2152800.0 ;
      RECT  430800.0 2151600.0 432000.0 2152800.0 ;
      RECT  428400.0 2158800.0 429600.0 2160000.0 ;
      RECT  433200.0 2158800.0 434400.0 2160000.0 ;
      RECT  425400.0 2154000.0 435600.0 2154900.0 ;
      RECT  425400.0 2165100.0 435600.0 2166000.0 ;
      RECT  441000.0 2158800.0 442200.0 2166000.0 ;
      RECT  438600.0 2151600.0 439800.0 2152800.0 ;
      RECT  441000.0 2151600.0 442200.0 2152800.0 ;
      RECT  441000.0 2151600.0 442200.0 2152800.0 ;
      RECT  438600.0 2151600.0 439800.0 2152800.0 ;
      RECT  438600.0 2158800.0 439800.0 2160000.0 ;
      RECT  441000.0 2158800.0 442200.0 2160000.0 ;
      RECT  441000.0 2158800.0 442200.0 2160000.0 ;
      RECT  438600.0 2158800.0 439800.0 2160000.0 ;
      RECT  441000.0 2158800.0 442200.0 2160000.0 ;
      RECT  443400.0 2158800.0 444600.0 2160000.0 ;
      RECT  443400.0 2158800.0 444600.0 2160000.0 ;
      RECT  441000.0 2158800.0 442200.0 2160000.0 ;
      RECT  440700.0 2153850.0 439500.0 2155050.0 ;
      RECT  441000.0 2164200.0 442200.0 2165400.0 ;
      RECT  438600.0 2151600.0 439800.0 2152800.0 ;
      RECT  441000.0 2151600.0 442200.0 2152800.0 ;
      RECT  438600.0 2158800.0 439800.0 2160000.0 ;
      RECT  443400.0 2158800.0 444600.0 2160000.0 ;
      RECT  435600.0 2154000.0 445800.0 2154900.0 ;
      RECT  435600.0 2165100.0 445800.0 2166000.0 ;
      RECT  451200.0 2158800.0 452400.0 2166000.0 ;
      RECT  448800.0 2151600.0 450000.0 2152800.0 ;
      RECT  451200.0 2151600.0 452400.0 2152800.0 ;
      RECT  451200.0 2151600.0 452400.0 2152800.0 ;
      RECT  448800.0 2151600.0 450000.0 2152800.0 ;
      RECT  448800.0 2158800.0 450000.0 2160000.0 ;
      RECT  451200.0 2158800.0 452400.0 2160000.0 ;
      RECT  451200.0 2158800.0 452400.0 2160000.0 ;
      RECT  448800.0 2158800.0 450000.0 2160000.0 ;
      RECT  451200.0 2158800.0 452400.0 2160000.0 ;
      RECT  453600.0 2158800.0 454800.0 2160000.0 ;
      RECT  453600.0 2158800.0 454800.0 2160000.0 ;
      RECT  451200.0 2158800.0 452400.0 2160000.0 ;
      RECT  450900.0 2153850.0 449700.0 2155050.0 ;
      RECT  451200.0 2164200.0 452400.0 2165400.0 ;
      RECT  448800.0 2151600.0 450000.0 2152800.0 ;
      RECT  451200.0 2151600.0 452400.0 2152800.0 ;
      RECT  448800.0 2158800.0 450000.0 2160000.0 ;
      RECT  453600.0 2158800.0 454800.0 2160000.0 ;
      RECT  445800.0 2154000.0 456000.0 2154900.0 ;
      RECT  445800.0 2165100.0 456000.0 2166000.0 ;
      RECT  461400.0 2158800.0 462600.0 2166000.0 ;
      RECT  459000.0 2151600.0 460200.0 2152800.0 ;
      RECT  461400.0 2151600.0 462600.0 2152800.0 ;
      RECT  461400.0 2151600.0 462600.0 2152800.0 ;
      RECT  459000.0 2151600.0 460200.0 2152800.0 ;
      RECT  459000.0 2158800.0 460200.0 2160000.0 ;
      RECT  461400.0 2158800.0 462600.0 2160000.0 ;
      RECT  461400.0 2158800.0 462600.0 2160000.0 ;
      RECT  459000.0 2158800.0 460200.0 2160000.0 ;
      RECT  461400.0 2158800.0 462600.0 2160000.0 ;
      RECT  463800.0 2158800.0 465000.0 2160000.0 ;
      RECT  463800.0 2158800.0 465000.0 2160000.0 ;
      RECT  461400.0 2158800.0 462600.0 2160000.0 ;
      RECT  461100.0 2153850.0 459900.0 2155050.0 ;
      RECT  461400.0 2164200.0 462600.0 2165400.0 ;
      RECT  459000.0 2151600.0 460200.0 2152800.0 ;
      RECT  461400.0 2151600.0 462600.0 2152800.0 ;
      RECT  459000.0 2158800.0 460200.0 2160000.0 ;
      RECT  463800.0 2158800.0 465000.0 2160000.0 ;
      RECT  456000.0 2154000.0 466200.0 2154900.0 ;
      RECT  456000.0 2165100.0 466200.0 2166000.0 ;
      RECT  471600.0 2158800.0 472800.0 2166000.0 ;
      RECT  469200.0 2151600.0 470400.0 2152800.0 ;
      RECT  471600.0 2151600.0 472800.0 2152800.0 ;
      RECT  471600.0 2151600.0 472800.0 2152800.0 ;
      RECT  469200.0 2151600.0 470400.0 2152800.0 ;
      RECT  469200.0 2158800.0 470400.0 2160000.0 ;
      RECT  471600.0 2158800.0 472800.0 2160000.0 ;
      RECT  471600.0 2158800.0 472800.0 2160000.0 ;
      RECT  469200.0 2158800.0 470400.0 2160000.0 ;
      RECT  471600.0 2158800.0 472800.0 2160000.0 ;
      RECT  474000.0 2158800.0 475200.0 2160000.0 ;
      RECT  474000.0 2158800.0 475200.0 2160000.0 ;
      RECT  471600.0 2158800.0 472800.0 2160000.0 ;
      RECT  471300.0 2153850.0 470100.0 2155050.0 ;
      RECT  471600.0 2164200.0 472800.0 2165400.0 ;
      RECT  469200.0 2151600.0 470400.0 2152800.0 ;
      RECT  471600.0 2151600.0 472800.0 2152800.0 ;
      RECT  469200.0 2158800.0 470400.0 2160000.0 ;
      RECT  474000.0 2158800.0 475200.0 2160000.0 ;
      RECT  466200.0 2154000.0 476400.0 2154900.0 ;
      RECT  466200.0 2165100.0 476400.0 2166000.0 ;
      RECT  481800.0 2158800.0 483000.0 2166000.0 ;
      RECT  479400.0 2151600.0 480600.0 2152800.0 ;
      RECT  481800.0 2151600.0 483000.0 2152800.0 ;
      RECT  481800.0 2151600.0 483000.0 2152800.0 ;
      RECT  479400.0 2151600.0 480600.0 2152800.0 ;
      RECT  479400.0 2158800.0 480600.0 2160000.0 ;
      RECT  481800.0 2158800.0 483000.0 2160000.0 ;
      RECT  481800.0 2158800.0 483000.0 2160000.0 ;
      RECT  479400.0 2158800.0 480600.0 2160000.0 ;
      RECT  481800.0 2158800.0 483000.0 2160000.0 ;
      RECT  484200.0 2158800.0 485400.0 2160000.0 ;
      RECT  484200.0 2158800.0 485400.0 2160000.0 ;
      RECT  481800.0 2158800.0 483000.0 2160000.0 ;
      RECT  481500.0 2153850.0 480300.0 2155050.0 ;
      RECT  481800.0 2164200.0 483000.0 2165400.0 ;
      RECT  479400.0 2151600.0 480600.0 2152800.0 ;
      RECT  481800.0 2151600.0 483000.0 2152800.0 ;
      RECT  479400.0 2158800.0 480600.0 2160000.0 ;
      RECT  484200.0 2158800.0 485400.0 2160000.0 ;
      RECT  476400.0 2154000.0 486600.0 2154900.0 ;
      RECT  476400.0 2165100.0 486600.0 2166000.0 ;
      RECT  492000.0 2158800.0 493200.0 2166000.0 ;
      RECT  489600.0 2151600.0 490800.0 2152800.0 ;
      RECT  492000.0 2151600.0 493200.0 2152800.0 ;
      RECT  492000.0 2151600.0 493200.0 2152800.0 ;
      RECT  489600.0 2151600.0 490800.0 2152800.0 ;
      RECT  489600.0 2158800.0 490800.0 2160000.0 ;
      RECT  492000.0 2158800.0 493200.0 2160000.0 ;
      RECT  492000.0 2158800.0 493200.0 2160000.0 ;
      RECT  489600.0 2158800.0 490800.0 2160000.0 ;
      RECT  492000.0 2158800.0 493200.0 2160000.0 ;
      RECT  494400.0 2158800.0 495600.0 2160000.0 ;
      RECT  494400.0 2158800.0 495600.0 2160000.0 ;
      RECT  492000.0 2158800.0 493200.0 2160000.0 ;
      RECT  491700.0 2153850.0 490500.0 2155050.0 ;
      RECT  492000.0 2164200.0 493200.0 2165400.0 ;
      RECT  489600.0 2151600.0 490800.0 2152800.0 ;
      RECT  492000.0 2151600.0 493200.0 2152800.0 ;
      RECT  489600.0 2158800.0 490800.0 2160000.0 ;
      RECT  494400.0 2158800.0 495600.0 2160000.0 ;
      RECT  486600.0 2154000.0 496800.0 2154900.0 ;
      RECT  486600.0 2165100.0 496800.0 2166000.0 ;
      RECT  502200.0 2158800.0 503400.0 2166000.0 ;
      RECT  499800.0 2151600.0 501000.0 2152800.0 ;
      RECT  502200.0 2151600.0 503400.0 2152800.0 ;
      RECT  502200.0 2151600.0 503400.0 2152800.0 ;
      RECT  499800.0 2151600.0 501000.0 2152800.0 ;
      RECT  499800.0 2158800.0 501000.0 2160000.0 ;
      RECT  502200.0 2158800.0 503400.0 2160000.0 ;
      RECT  502200.0 2158800.0 503400.0 2160000.0 ;
      RECT  499800.0 2158800.0 501000.0 2160000.0 ;
      RECT  502200.0 2158800.0 503400.0 2160000.0 ;
      RECT  504600.0 2158800.0 505800.0 2160000.0 ;
      RECT  504600.0 2158800.0 505800.0 2160000.0 ;
      RECT  502200.0 2158800.0 503400.0 2160000.0 ;
      RECT  501900.0 2153850.0 500700.0 2155050.0 ;
      RECT  502200.0 2164200.0 503400.0 2165400.0 ;
      RECT  499800.0 2151600.0 501000.0 2152800.0 ;
      RECT  502200.0 2151600.0 503400.0 2152800.0 ;
      RECT  499800.0 2158800.0 501000.0 2160000.0 ;
      RECT  504600.0 2158800.0 505800.0 2160000.0 ;
      RECT  496800.0 2154000.0 507000.0 2154900.0 ;
      RECT  496800.0 2165100.0 507000.0 2166000.0 ;
      RECT  512400.0 2158800.0 513600.0 2166000.0 ;
      RECT  510000.0 2151600.0 511200.0 2152800.0 ;
      RECT  512400.0 2151600.0 513600.0 2152800.0 ;
      RECT  512400.0 2151600.0 513600.0 2152800.0 ;
      RECT  510000.0 2151600.0 511200.0 2152800.0 ;
      RECT  510000.0 2158800.0 511200.0 2160000.0 ;
      RECT  512400.0 2158800.0 513600.0 2160000.0 ;
      RECT  512400.0 2158800.0 513600.0 2160000.0 ;
      RECT  510000.0 2158800.0 511200.0 2160000.0 ;
      RECT  512400.0 2158800.0 513600.0 2160000.0 ;
      RECT  514800.0 2158800.0 516000.0 2160000.0 ;
      RECT  514800.0 2158800.0 516000.0 2160000.0 ;
      RECT  512400.0 2158800.0 513600.0 2160000.0 ;
      RECT  512100.0 2153850.0 510900.0 2155050.0 ;
      RECT  512400.0 2164200.0 513600.0 2165400.0 ;
      RECT  510000.0 2151600.0 511200.0 2152800.0 ;
      RECT  512400.0 2151600.0 513600.0 2152800.0 ;
      RECT  510000.0 2158800.0 511200.0 2160000.0 ;
      RECT  514800.0 2158800.0 516000.0 2160000.0 ;
      RECT  507000.0 2154000.0 517200.0 2154900.0 ;
      RECT  507000.0 2165100.0 517200.0 2166000.0 ;
      RECT  522600.0 2158800.0 523800.0 2166000.0 ;
      RECT  520200.0 2151600.0 521400.0 2152800.0 ;
      RECT  522600.0 2151600.0 523800.0 2152800.0 ;
      RECT  522600.0 2151600.0 523800.0 2152800.0 ;
      RECT  520200.0 2151600.0 521400.0 2152800.0 ;
      RECT  520200.0 2158800.0 521400.0 2160000.0 ;
      RECT  522600.0 2158800.0 523800.0 2160000.0 ;
      RECT  522600.0 2158800.0 523800.0 2160000.0 ;
      RECT  520200.0 2158800.0 521400.0 2160000.0 ;
      RECT  522600.0 2158800.0 523800.0 2160000.0 ;
      RECT  525000.0 2158800.0 526200.0 2160000.0 ;
      RECT  525000.0 2158800.0 526200.0 2160000.0 ;
      RECT  522600.0 2158800.0 523800.0 2160000.0 ;
      RECT  522300.0 2153850.0 521100.0 2155050.0 ;
      RECT  522600.0 2164200.0 523800.0 2165400.0 ;
      RECT  520200.0 2151600.0 521400.0 2152800.0 ;
      RECT  522600.0 2151600.0 523800.0 2152800.0 ;
      RECT  520200.0 2158800.0 521400.0 2160000.0 ;
      RECT  525000.0 2158800.0 526200.0 2160000.0 ;
      RECT  517200.0 2154000.0 527400.0 2154900.0 ;
      RECT  517200.0 2165100.0 527400.0 2166000.0 ;
      RECT  532800.0 2158800.0 534000.0 2166000.0 ;
      RECT  530400.0 2151600.0 531600.0 2152800.0 ;
      RECT  532800.0 2151600.0 534000.0 2152800.0 ;
      RECT  532800.0 2151600.0 534000.0 2152800.0 ;
      RECT  530400.0 2151600.0 531600.0 2152800.0 ;
      RECT  530400.0 2158800.0 531600.0 2160000.0 ;
      RECT  532800.0 2158800.0 534000.0 2160000.0 ;
      RECT  532800.0 2158800.0 534000.0 2160000.0 ;
      RECT  530400.0 2158800.0 531600.0 2160000.0 ;
      RECT  532800.0 2158800.0 534000.0 2160000.0 ;
      RECT  535200.0 2158800.0 536400.0 2160000.0 ;
      RECT  535200.0 2158800.0 536400.0 2160000.0 ;
      RECT  532800.0 2158800.0 534000.0 2160000.0 ;
      RECT  532500.0 2153850.0 531300.0 2155050.0 ;
      RECT  532800.0 2164200.0 534000.0 2165400.0 ;
      RECT  530400.0 2151600.0 531600.0 2152800.0 ;
      RECT  532800.0 2151600.0 534000.0 2152800.0 ;
      RECT  530400.0 2158800.0 531600.0 2160000.0 ;
      RECT  535200.0 2158800.0 536400.0 2160000.0 ;
      RECT  527400.0 2154000.0 537600.0 2154900.0 ;
      RECT  527400.0 2165100.0 537600.0 2166000.0 ;
      RECT  543000.0 2158800.0 544200.0 2166000.0 ;
      RECT  540600.0 2151600.0 541800.0 2152800.0 ;
      RECT  543000.0 2151600.0 544200.0 2152800.0 ;
      RECT  543000.0 2151600.0 544200.0 2152800.0 ;
      RECT  540600.0 2151600.0 541800.0 2152800.0 ;
      RECT  540600.0 2158800.0 541800.0 2160000.0 ;
      RECT  543000.0 2158800.0 544200.0 2160000.0 ;
      RECT  543000.0 2158800.0 544200.0 2160000.0 ;
      RECT  540600.0 2158800.0 541800.0 2160000.0 ;
      RECT  543000.0 2158800.0 544200.0 2160000.0 ;
      RECT  545400.0 2158800.0 546600.0 2160000.0 ;
      RECT  545400.0 2158800.0 546600.0 2160000.0 ;
      RECT  543000.0 2158800.0 544200.0 2160000.0 ;
      RECT  542700.0 2153850.0 541500.0 2155050.0 ;
      RECT  543000.0 2164200.0 544200.0 2165400.0 ;
      RECT  540600.0 2151600.0 541800.0 2152800.0 ;
      RECT  543000.0 2151600.0 544200.0 2152800.0 ;
      RECT  540600.0 2158800.0 541800.0 2160000.0 ;
      RECT  545400.0 2158800.0 546600.0 2160000.0 ;
      RECT  537600.0 2154000.0 547800.0 2154900.0 ;
      RECT  537600.0 2165100.0 547800.0 2166000.0 ;
      RECT  553200.0 2158800.0 554400.0 2166000.0 ;
      RECT  550800.0 2151600.0 552000.0 2152800.0 ;
      RECT  553200.0 2151600.0 554400.0 2152800.0 ;
      RECT  553200.0 2151600.0 554400.0 2152800.0 ;
      RECT  550800.0 2151600.0 552000.0 2152800.0 ;
      RECT  550800.0 2158800.0 552000.0 2160000.0 ;
      RECT  553200.0 2158800.0 554400.0 2160000.0 ;
      RECT  553200.0 2158800.0 554400.0 2160000.0 ;
      RECT  550800.0 2158800.0 552000.0 2160000.0 ;
      RECT  553200.0 2158800.0 554400.0 2160000.0 ;
      RECT  555600.0 2158800.0 556800.0 2160000.0 ;
      RECT  555600.0 2158800.0 556800.0 2160000.0 ;
      RECT  553200.0 2158800.0 554400.0 2160000.0 ;
      RECT  552900.0 2153850.0 551700.0 2155050.0 ;
      RECT  553200.0 2164200.0 554400.0 2165400.0 ;
      RECT  550800.0 2151600.0 552000.0 2152800.0 ;
      RECT  553200.0 2151600.0 554400.0 2152800.0 ;
      RECT  550800.0 2158800.0 552000.0 2160000.0 ;
      RECT  555600.0 2158800.0 556800.0 2160000.0 ;
      RECT  547800.0 2154000.0 558000.0 2154900.0 ;
      RECT  547800.0 2165100.0 558000.0 2166000.0 ;
      RECT  563400.0 2158800.0 564600.0 2166000.0 ;
      RECT  561000.0 2151600.0 562200.0 2152800.0 ;
      RECT  563400.0 2151600.0 564600.0 2152800.0 ;
      RECT  563400.0 2151600.0 564600.0 2152800.0 ;
      RECT  561000.0 2151600.0 562200.0 2152800.0 ;
      RECT  561000.0 2158800.0 562200.0 2160000.0 ;
      RECT  563400.0 2158800.0 564600.0 2160000.0 ;
      RECT  563400.0 2158800.0 564600.0 2160000.0 ;
      RECT  561000.0 2158800.0 562200.0 2160000.0 ;
      RECT  563400.0 2158800.0 564600.0 2160000.0 ;
      RECT  565800.0 2158800.0 567000.0 2160000.0 ;
      RECT  565800.0 2158800.0 567000.0 2160000.0 ;
      RECT  563400.0 2158800.0 564600.0 2160000.0 ;
      RECT  563100.0 2153850.0 561900.0 2155050.0 ;
      RECT  563400.0 2164200.0 564600.0 2165400.0 ;
      RECT  561000.0 2151600.0 562200.0 2152800.0 ;
      RECT  563400.0 2151600.0 564600.0 2152800.0 ;
      RECT  561000.0 2158800.0 562200.0 2160000.0 ;
      RECT  565800.0 2158800.0 567000.0 2160000.0 ;
      RECT  558000.0 2154000.0 568200.0 2154900.0 ;
      RECT  558000.0 2165100.0 568200.0 2166000.0 ;
      RECT  573600.0 2158800.0 574800.0 2166000.0 ;
      RECT  571200.0 2151600.0 572400.0 2152800.0 ;
      RECT  573600.0 2151600.0 574800.0 2152800.0 ;
      RECT  573600.0 2151600.0 574800.0 2152800.0 ;
      RECT  571200.0 2151600.0 572400.0 2152800.0 ;
      RECT  571200.0 2158800.0 572400.0 2160000.0 ;
      RECT  573600.0 2158800.0 574800.0 2160000.0 ;
      RECT  573600.0 2158800.0 574800.0 2160000.0 ;
      RECT  571200.0 2158800.0 572400.0 2160000.0 ;
      RECT  573600.0 2158800.0 574800.0 2160000.0 ;
      RECT  576000.0 2158800.0 577200.0 2160000.0 ;
      RECT  576000.0 2158800.0 577200.0 2160000.0 ;
      RECT  573600.0 2158800.0 574800.0 2160000.0 ;
      RECT  573300.0 2153850.0 572100.0 2155050.0 ;
      RECT  573600.0 2164200.0 574800.0 2165400.0 ;
      RECT  571200.0 2151600.0 572400.0 2152800.0 ;
      RECT  573600.0 2151600.0 574800.0 2152800.0 ;
      RECT  571200.0 2158800.0 572400.0 2160000.0 ;
      RECT  576000.0 2158800.0 577200.0 2160000.0 ;
      RECT  568200.0 2154000.0 578400.0 2154900.0 ;
      RECT  568200.0 2165100.0 578400.0 2166000.0 ;
      RECT  583800.0 2158800.0 585000.0 2166000.0 ;
      RECT  581400.0 2151600.0 582600.0 2152800.0 ;
      RECT  583800.0 2151600.0 585000.0 2152800.0 ;
      RECT  583800.0 2151600.0 585000.0 2152800.0 ;
      RECT  581400.0 2151600.0 582600.0 2152800.0 ;
      RECT  581400.0 2158800.0 582600.0 2160000.0 ;
      RECT  583800.0 2158800.0 585000.0 2160000.0 ;
      RECT  583800.0 2158800.0 585000.0 2160000.0 ;
      RECT  581400.0 2158800.0 582600.0 2160000.0 ;
      RECT  583800.0 2158800.0 585000.0 2160000.0 ;
      RECT  586200.0 2158800.0 587400.0 2160000.0 ;
      RECT  586200.0 2158800.0 587400.0 2160000.0 ;
      RECT  583800.0 2158800.0 585000.0 2160000.0 ;
      RECT  583500.0 2153850.0 582300.0 2155050.0 ;
      RECT  583800.0 2164200.0 585000.0 2165400.0 ;
      RECT  581400.0 2151600.0 582600.0 2152800.0 ;
      RECT  583800.0 2151600.0 585000.0 2152800.0 ;
      RECT  581400.0 2158800.0 582600.0 2160000.0 ;
      RECT  586200.0 2158800.0 587400.0 2160000.0 ;
      RECT  578400.0 2154000.0 588600.0 2154900.0 ;
      RECT  578400.0 2165100.0 588600.0 2166000.0 ;
      RECT  594000.0 2158800.0 595200.0 2166000.0 ;
      RECT  591600.0 2151600.0 592800.0 2152800.0 ;
      RECT  594000.0 2151600.0 595200.0 2152800.0 ;
      RECT  594000.0 2151600.0 595200.0 2152800.0 ;
      RECT  591600.0 2151600.0 592800.0 2152800.0 ;
      RECT  591600.0 2158800.0 592800.0 2160000.0 ;
      RECT  594000.0 2158800.0 595200.0 2160000.0 ;
      RECT  594000.0 2158800.0 595200.0 2160000.0 ;
      RECT  591600.0 2158800.0 592800.0 2160000.0 ;
      RECT  594000.0 2158800.0 595200.0 2160000.0 ;
      RECT  596400.0 2158800.0 597600.0 2160000.0 ;
      RECT  596400.0 2158800.0 597600.0 2160000.0 ;
      RECT  594000.0 2158800.0 595200.0 2160000.0 ;
      RECT  593700.0 2153850.0 592500.0 2155050.0 ;
      RECT  594000.0 2164200.0 595200.0 2165400.0 ;
      RECT  591600.0 2151600.0 592800.0 2152800.0 ;
      RECT  594000.0 2151600.0 595200.0 2152800.0 ;
      RECT  591600.0 2158800.0 592800.0 2160000.0 ;
      RECT  596400.0 2158800.0 597600.0 2160000.0 ;
      RECT  588600.0 2154000.0 598800.0 2154900.0 ;
      RECT  588600.0 2165100.0 598800.0 2166000.0 ;
      RECT  604200.0 2158800.0 605400.0 2166000.0 ;
      RECT  601800.0 2151600.0 603000.0 2152800.0 ;
      RECT  604200.0 2151600.0 605400.0 2152800.0 ;
      RECT  604200.0 2151600.0 605400.0 2152800.0 ;
      RECT  601800.0 2151600.0 603000.0 2152800.0 ;
      RECT  601800.0 2158800.0 603000.0 2160000.0 ;
      RECT  604200.0 2158800.0 605400.0 2160000.0 ;
      RECT  604200.0 2158800.0 605400.0 2160000.0 ;
      RECT  601800.0 2158800.0 603000.0 2160000.0 ;
      RECT  604200.0 2158800.0 605400.0 2160000.0 ;
      RECT  606600.0 2158800.0 607800.0 2160000.0 ;
      RECT  606600.0 2158800.0 607800.0 2160000.0 ;
      RECT  604200.0 2158800.0 605400.0 2160000.0 ;
      RECT  603900.0 2153850.0 602700.0 2155050.0 ;
      RECT  604200.0 2164200.0 605400.0 2165400.0 ;
      RECT  601800.0 2151600.0 603000.0 2152800.0 ;
      RECT  604200.0 2151600.0 605400.0 2152800.0 ;
      RECT  601800.0 2158800.0 603000.0 2160000.0 ;
      RECT  606600.0 2158800.0 607800.0 2160000.0 ;
      RECT  598800.0 2154000.0 609000.0 2154900.0 ;
      RECT  598800.0 2165100.0 609000.0 2166000.0 ;
      RECT  614400.0 2158800.0 615600.0 2166000.0 ;
      RECT  612000.0 2151600.0 613200.0 2152800.0 ;
      RECT  614400.0 2151600.0 615600.0 2152800.0 ;
      RECT  614400.0 2151600.0 615600.0 2152800.0 ;
      RECT  612000.0 2151600.0 613200.0 2152800.0 ;
      RECT  612000.0 2158800.0 613200.0 2160000.0 ;
      RECT  614400.0 2158800.0 615600.0 2160000.0 ;
      RECT  614400.0 2158800.0 615600.0 2160000.0 ;
      RECT  612000.0 2158800.0 613200.0 2160000.0 ;
      RECT  614400.0 2158800.0 615600.0 2160000.0 ;
      RECT  616800.0 2158800.0 618000.0 2160000.0 ;
      RECT  616800.0 2158800.0 618000.0 2160000.0 ;
      RECT  614400.0 2158800.0 615600.0 2160000.0 ;
      RECT  614100.0 2153850.0 612900.0 2155050.0 ;
      RECT  614400.0 2164200.0 615600.0 2165400.0 ;
      RECT  612000.0 2151600.0 613200.0 2152800.0 ;
      RECT  614400.0 2151600.0 615600.0 2152800.0 ;
      RECT  612000.0 2158800.0 613200.0 2160000.0 ;
      RECT  616800.0 2158800.0 618000.0 2160000.0 ;
      RECT  609000.0 2154000.0 619200.0 2154900.0 ;
      RECT  609000.0 2165100.0 619200.0 2166000.0 ;
      RECT  624600.0 2158800.0 625800.0 2166000.0 ;
      RECT  622200.0 2151600.0 623400.0 2152800.0 ;
      RECT  624600.0 2151600.0 625800.0 2152800.0 ;
      RECT  624600.0 2151600.0 625800.0 2152800.0 ;
      RECT  622200.0 2151600.0 623400.0 2152800.0 ;
      RECT  622200.0 2158800.0 623400.0 2160000.0 ;
      RECT  624600.0 2158800.0 625800.0 2160000.0 ;
      RECT  624600.0 2158800.0 625800.0 2160000.0 ;
      RECT  622200.0 2158800.0 623400.0 2160000.0 ;
      RECT  624600.0 2158800.0 625800.0 2160000.0 ;
      RECT  627000.0 2158800.0 628200.0 2160000.0 ;
      RECT  627000.0 2158800.0 628200.0 2160000.0 ;
      RECT  624600.0 2158800.0 625800.0 2160000.0 ;
      RECT  624300.0 2153850.0 623100.0 2155050.0 ;
      RECT  624600.0 2164200.0 625800.0 2165400.0 ;
      RECT  622200.0 2151600.0 623400.0 2152800.0 ;
      RECT  624600.0 2151600.0 625800.0 2152800.0 ;
      RECT  622200.0 2158800.0 623400.0 2160000.0 ;
      RECT  627000.0 2158800.0 628200.0 2160000.0 ;
      RECT  619200.0 2154000.0 629400.0 2154900.0 ;
      RECT  619200.0 2165100.0 629400.0 2166000.0 ;
      RECT  634800.0 2158800.0 636000.0 2166000.0 ;
      RECT  632400.0 2151600.0 633600.0 2152800.0 ;
      RECT  634800.0 2151600.0 636000.0 2152800.0 ;
      RECT  634800.0 2151600.0 636000.0 2152800.0 ;
      RECT  632400.0 2151600.0 633600.0 2152800.0 ;
      RECT  632400.0 2158800.0 633600.0 2160000.0 ;
      RECT  634800.0 2158800.0 636000.0 2160000.0 ;
      RECT  634800.0 2158800.0 636000.0 2160000.0 ;
      RECT  632400.0 2158800.0 633600.0 2160000.0 ;
      RECT  634800.0 2158800.0 636000.0 2160000.0 ;
      RECT  637200.0 2158800.0 638400.0 2160000.0 ;
      RECT  637200.0 2158800.0 638400.0 2160000.0 ;
      RECT  634800.0 2158800.0 636000.0 2160000.0 ;
      RECT  634500.0 2153850.0 633300.0 2155050.0 ;
      RECT  634800.0 2164200.0 636000.0 2165400.0 ;
      RECT  632400.0 2151600.0 633600.0 2152800.0 ;
      RECT  634800.0 2151600.0 636000.0 2152800.0 ;
      RECT  632400.0 2158800.0 633600.0 2160000.0 ;
      RECT  637200.0 2158800.0 638400.0 2160000.0 ;
      RECT  629400.0 2154000.0 639600.0 2154900.0 ;
      RECT  629400.0 2165100.0 639600.0 2166000.0 ;
      RECT  645000.0 2158800.0 646200.0 2166000.0 ;
      RECT  642600.0 2151600.0 643800.0 2152800.0 ;
      RECT  645000.0 2151600.0 646200.0 2152800.0 ;
      RECT  645000.0 2151600.0 646200.0 2152800.0 ;
      RECT  642600.0 2151600.0 643800.0 2152800.0 ;
      RECT  642600.0 2158800.0 643800.0 2160000.0 ;
      RECT  645000.0 2158800.0 646200.0 2160000.0 ;
      RECT  645000.0 2158800.0 646200.0 2160000.0 ;
      RECT  642600.0 2158800.0 643800.0 2160000.0 ;
      RECT  645000.0 2158800.0 646200.0 2160000.0 ;
      RECT  647400.0 2158800.0 648600.0 2160000.0 ;
      RECT  647400.0 2158800.0 648600.0 2160000.0 ;
      RECT  645000.0 2158800.0 646200.0 2160000.0 ;
      RECT  644700.0 2153850.0 643500.0 2155050.0 ;
      RECT  645000.0 2164200.0 646200.0 2165400.0 ;
      RECT  642600.0 2151600.0 643800.0 2152800.0 ;
      RECT  645000.0 2151600.0 646200.0 2152800.0 ;
      RECT  642600.0 2158800.0 643800.0 2160000.0 ;
      RECT  647400.0 2158800.0 648600.0 2160000.0 ;
      RECT  639600.0 2154000.0 649800.0 2154900.0 ;
      RECT  639600.0 2165100.0 649800.0 2166000.0 ;
      RECT  655200.0 2158800.0 656400.0 2166000.0 ;
      RECT  652800.0 2151600.0 654000.0 2152800.0 ;
      RECT  655200.0 2151600.0 656400.0 2152800.0 ;
      RECT  655200.0 2151600.0 656400.0 2152800.0 ;
      RECT  652800.0 2151600.0 654000.0 2152800.0 ;
      RECT  652800.0 2158800.0 654000.0 2160000.0 ;
      RECT  655200.0 2158800.0 656400.0 2160000.0 ;
      RECT  655200.0 2158800.0 656400.0 2160000.0 ;
      RECT  652800.0 2158800.0 654000.0 2160000.0 ;
      RECT  655200.0 2158800.0 656400.0 2160000.0 ;
      RECT  657600.0 2158800.0 658800.0 2160000.0 ;
      RECT  657600.0 2158800.0 658800.0 2160000.0 ;
      RECT  655200.0 2158800.0 656400.0 2160000.0 ;
      RECT  654900.0 2153850.0 653700.0 2155050.0 ;
      RECT  655200.0 2164200.0 656400.0 2165400.0 ;
      RECT  652800.0 2151600.0 654000.0 2152800.0 ;
      RECT  655200.0 2151600.0 656400.0 2152800.0 ;
      RECT  652800.0 2158800.0 654000.0 2160000.0 ;
      RECT  657600.0 2158800.0 658800.0 2160000.0 ;
      RECT  649800.0 2154000.0 660000.0 2154900.0 ;
      RECT  649800.0 2165100.0 660000.0 2166000.0 ;
      RECT  665400.0 2158800.0 666600.0 2166000.0 ;
      RECT  663000.0 2151600.0 664200.0 2152800.0 ;
      RECT  665400.0 2151600.0 666600.0 2152800.0 ;
      RECT  665400.0 2151600.0 666600.0 2152800.0 ;
      RECT  663000.0 2151600.0 664200.0 2152800.0 ;
      RECT  663000.0 2158800.0 664200.0 2160000.0 ;
      RECT  665400.0 2158800.0 666600.0 2160000.0 ;
      RECT  665400.0 2158800.0 666600.0 2160000.0 ;
      RECT  663000.0 2158800.0 664200.0 2160000.0 ;
      RECT  665400.0 2158800.0 666600.0 2160000.0 ;
      RECT  667800.0 2158800.0 669000.0 2160000.0 ;
      RECT  667800.0 2158800.0 669000.0 2160000.0 ;
      RECT  665400.0 2158800.0 666600.0 2160000.0 ;
      RECT  665100.0 2153850.0 663900.0 2155050.0 ;
      RECT  665400.0 2164200.0 666600.0 2165400.0 ;
      RECT  663000.0 2151600.0 664200.0 2152800.0 ;
      RECT  665400.0 2151600.0 666600.0 2152800.0 ;
      RECT  663000.0 2158800.0 664200.0 2160000.0 ;
      RECT  667800.0 2158800.0 669000.0 2160000.0 ;
      RECT  660000.0 2154000.0 670200.0 2154900.0 ;
      RECT  660000.0 2165100.0 670200.0 2166000.0 ;
      RECT  675600.0 2158800.0 676800.0 2166000.0 ;
      RECT  673200.0 2151600.0 674400.0 2152800.0 ;
      RECT  675600.0 2151600.0 676800.0 2152800.0 ;
      RECT  675600.0 2151600.0 676800.0 2152800.0 ;
      RECT  673200.0 2151600.0 674400.0 2152800.0 ;
      RECT  673200.0 2158800.0 674400.0 2160000.0 ;
      RECT  675600.0 2158800.0 676800.0 2160000.0 ;
      RECT  675600.0 2158800.0 676800.0 2160000.0 ;
      RECT  673200.0 2158800.0 674400.0 2160000.0 ;
      RECT  675600.0 2158800.0 676800.0 2160000.0 ;
      RECT  678000.0 2158800.0 679200.0 2160000.0 ;
      RECT  678000.0 2158800.0 679200.0 2160000.0 ;
      RECT  675600.0 2158800.0 676800.0 2160000.0 ;
      RECT  675300.0 2153850.0 674100.0 2155050.0 ;
      RECT  675600.0 2164200.0 676800.0 2165400.0 ;
      RECT  673200.0 2151600.0 674400.0 2152800.0 ;
      RECT  675600.0 2151600.0 676800.0 2152800.0 ;
      RECT  673200.0 2158800.0 674400.0 2160000.0 ;
      RECT  678000.0 2158800.0 679200.0 2160000.0 ;
      RECT  670200.0 2154000.0 680400.0 2154900.0 ;
      RECT  670200.0 2165100.0 680400.0 2166000.0 ;
      RECT  685800.0 2158800.0 687000.0 2166000.0 ;
      RECT  683400.0 2151600.0 684600.0 2152800.0 ;
      RECT  685800.0 2151600.0 687000.0 2152800.0 ;
      RECT  685800.0 2151600.0 687000.0 2152800.0 ;
      RECT  683400.0 2151600.0 684600.0 2152800.0 ;
      RECT  683400.0 2158800.0 684600.0 2160000.0 ;
      RECT  685800.0 2158800.0 687000.0 2160000.0 ;
      RECT  685800.0 2158800.0 687000.0 2160000.0 ;
      RECT  683400.0 2158800.0 684600.0 2160000.0 ;
      RECT  685800.0 2158800.0 687000.0 2160000.0 ;
      RECT  688200.0 2158800.0 689400.0 2160000.0 ;
      RECT  688200.0 2158800.0 689400.0 2160000.0 ;
      RECT  685800.0 2158800.0 687000.0 2160000.0 ;
      RECT  685500.0 2153850.0 684300.0 2155050.0 ;
      RECT  685800.0 2164200.0 687000.0 2165400.0 ;
      RECT  683400.0 2151600.0 684600.0 2152800.0 ;
      RECT  685800.0 2151600.0 687000.0 2152800.0 ;
      RECT  683400.0 2158800.0 684600.0 2160000.0 ;
      RECT  688200.0 2158800.0 689400.0 2160000.0 ;
      RECT  680400.0 2154000.0 690600.0 2154900.0 ;
      RECT  680400.0 2165100.0 690600.0 2166000.0 ;
      RECT  696000.0 2158800.0 697200.0 2166000.0 ;
      RECT  693600.0 2151600.0 694800.0 2152800.0 ;
      RECT  696000.0 2151600.0 697200.0 2152800.0 ;
      RECT  696000.0 2151600.0 697200.0 2152800.0 ;
      RECT  693600.0 2151600.0 694800.0 2152800.0 ;
      RECT  693600.0 2158800.0 694800.0 2160000.0 ;
      RECT  696000.0 2158800.0 697200.0 2160000.0 ;
      RECT  696000.0 2158800.0 697200.0 2160000.0 ;
      RECT  693600.0 2158800.0 694800.0 2160000.0 ;
      RECT  696000.0 2158800.0 697200.0 2160000.0 ;
      RECT  698400.0 2158800.0 699600.0 2160000.0 ;
      RECT  698400.0 2158800.0 699600.0 2160000.0 ;
      RECT  696000.0 2158800.0 697200.0 2160000.0 ;
      RECT  695700.0 2153850.0 694500.0 2155050.0 ;
      RECT  696000.0 2164200.0 697200.0 2165400.0 ;
      RECT  693600.0 2151600.0 694800.0 2152800.0 ;
      RECT  696000.0 2151600.0 697200.0 2152800.0 ;
      RECT  693600.0 2158800.0 694800.0 2160000.0 ;
      RECT  698400.0 2158800.0 699600.0 2160000.0 ;
      RECT  690600.0 2154000.0 700800.0 2154900.0 ;
      RECT  690600.0 2165100.0 700800.0 2166000.0 ;
      RECT  706200.0 2158800.0 707400.0 2166000.0 ;
      RECT  703800.0 2151600.0 705000.0 2152800.0 ;
      RECT  706200.0 2151600.0 707400.0 2152800.0 ;
      RECT  706200.0 2151600.0 707400.0 2152800.0 ;
      RECT  703800.0 2151600.0 705000.0 2152800.0 ;
      RECT  703800.0 2158800.0 705000.0 2160000.0 ;
      RECT  706200.0 2158800.0 707400.0 2160000.0 ;
      RECT  706200.0 2158800.0 707400.0 2160000.0 ;
      RECT  703800.0 2158800.0 705000.0 2160000.0 ;
      RECT  706200.0 2158800.0 707400.0 2160000.0 ;
      RECT  708600.0 2158800.0 709800.0 2160000.0 ;
      RECT  708600.0 2158800.0 709800.0 2160000.0 ;
      RECT  706200.0 2158800.0 707400.0 2160000.0 ;
      RECT  705900.0 2153850.0 704700.0 2155050.0 ;
      RECT  706200.0 2164200.0 707400.0 2165400.0 ;
      RECT  703800.0 2151600.0 705000.0 2152800.0 ;
      RECT  706200.0 2151600.0 707400.0 2152800.0 ;
      RECT  703800.0 2158800.0 705000.0 2160000.0 ;
      RECT  708600.0 2158800.0 709800.0 2160000.0 ;
      RECT  700800.0 2154000.0 711000.0 2154900.0 ;
      RECT  700800.0 2165100.0 711000.0 2166000.0 ;
      RECT  716400.0 2158800.0 717600.0 2166000.0 ;
      RECT  714000.0 2151600.0 715200.0 2152800.0 ;
      RECT  716400.0 2151600.0 717600.0 2152800.0 ;
      RECT  716400.0 2151600.0 717600.0 2152800.0 ;
      RECT  714000.0 2151600.0 715200.0 2152800.0 ;
      RECT  714000.0 2158800.0 715200.0 2160000.0 ;
      RECT  716400.0 2158800.0 717600.0 2160000.0 ;
      RECT  716400.0 2158800.0 717600.0 2160000.0 ;
      RECT  714000.0 2158800.0 715200.0 2160000.0 ;
      RECT  716400.0 2158800.0 717600.0 2160000.0 ;
      RECT  718800.0 2158800.0 720000.0 2160000.0 ;
      RECT  718800.0 2158800.0 720000.0 2160000.0 ;
      RECT  716400.0 2158800.0 717600.0 2160000.0 ;
      RECT  716100.0 2153850.0 714900.0 2155050.0 ;
      RECT  716400.0 2164200.0 717600.0 2165400.0 ;
      RECT  714000.0 2151600.0 715200.0 2152800.0 ;
      RECT  716400.0 2151600.0 717600.0 2152800.0 ;
      RECT  714000.0 2158800.0 715200.0 2160000.0 ;
      RECT  718800.0 2158800.0 720000.0 2160000.0 ;
      RECT  711000.0 2154000.0 721200.0 2154900.0 ;
      RECT  711000.0 2165100.0 721200.0 2166000.0 ;
      RECT  726600.0 2158800.0 727800.0 2166000.0 ;
      RECT  724200.0 2151600.0 725400.0 2152800.0 ;
      RECT  726600.0 2151600.0 727800.0 2152800.0 ;
      RECT  726600.0 2151600.0 727800.0 2152800.0 ;
      RECT  724200.0 2151600.0 725400.0 2152800.0 ;
      RECT  724200.0 2158800.0 725400.0 2160000.0 ;
      RECT  726600.0 2158800.0 727800.0 2160000.0 ;
      RECT  726600.0 2158800.0 727800.0 2160000.0 ;
      RECT  724200.0 2158800.0 725400.0 2160000.0 ;
      RECT  726600.0 2158800.0 727800.0 2160000.0 ;
      RECT  729000.0 2158800.0 730200.0 2160000.0 ;
      RECT  729000.0 2158800.0 730200.0 2160000.0 ;
      RECT  726600.0 2158800.0 727800.0 2160000.0 ;
      RECT  726300.0 2153850.0 725100.0 2155050.0 ;
      RECT  726600.0 2164200.0 727800.0 2165400.0 ;
      RECT  724200.0 2151600.0 725400.0 2152800.0 ;
      RECT  726600.0 2151600.0 727800.0 2152800.0 ;
      RECT  724200.0 2158800.0 725400.0 2160000.0 ;
      RECT  729000.0 2158800.0 730200.0 2160000.0 ;
      RECT  721200.0 2154000.0 731400.0 2154900.0 ;
      RECT  721200.0 2165100.0 731400.0 2166000.0 ;
      RECT  736800.0 2158800.0 738000.0 2166000.0 ;
      RECT  734400.0 2151600.0 735600.0 2152800.0 ;
      RECT  736800.0 2151600.0 738000.0 2152800.0 ;
      RECT  736800.0 2151600.0 738000.0 2152800.0 ;
      RECT  734400.0 2151600.0 735600.0 2152800.0 ;
      RECT  734400.0 2158800.0 735600.0 2160000.0 ;
      RECT  736800.0 2158800.0 738000.0 2160000.0 ;
      RECT  736800.0 2158800.0 738000.0 2160000.0 ;
      RECT  734400.0 2158800.0 735600.0 2160000.0 ;
      RECT  736800.0 2158800.0 738000.0 2160000.0 ;
      RECT  739200.0 2158800.0 740400.0 2160000.0 ;
      RECT  739200.0 2158800.0 740400.0 2160000.0 ;
      RECT  736800.0 2158800.0 738000.0 2160000.0 ;
      RECT  736500.0 2153850.0 735300.0 2155050.0 ;
      RECT  736800.0 2164200.0 738000.0 2165400.0 ;
      RECT  734400.0 2151600.0 735600.0 2152800.0 ;
      RECT  736800.0 2151600.0 738000.0 2152800.0 ;
      RECT  734400.0 2158800.0 735600.0 2160000.0 ;
      RECT  739200.0 2158800.0 740400.0 2160000.0 ;
      RECT  731400.0 2154000.0 741600.0 2154900.0 ;
      RECT  731400.0 2165100.0 741600.0 2166000.0 ;
      RECT  747000.0 2158800.0 748200.0 2166000.0 ;
      RECT  744600.0 2151600.0 745800.0 2152800.0 ;
      RECT  747000.0 2151600.0 748200.0 2152800.0 ;
      RECT  747000.0 2151600.0 748200.0 2152800.0 ;
      RECT  744600.0 2151600.0 745800.0 2152800.0 ;
      RECT  744600.0 2158800.0 745800.0 2160000.0 ;
      RECT  747000.0 2158800.0 748200.0 2160000.0 ;
      RECT  747000.0 2158800.0 748200.0 2160000.0 ;
      RECT  744600.0 2158800.0 745800.0 2160000.0 ;
      RECT  747000.0 2158800.0 748200.0 2160000.0 ;
      RECT  749400.0 2158800.0 750600.0 2160000.0 ;
      RECT  749400.0 2158800.0 750600.0 2160000.0 ;
      RECT  747000.0 2158800.0 748200.0 2160000.0 ;
      RECT  746700.0 2153850.0 745500.0 2155050.0 ;
      RECT  747000.0 2164200.0 748200.0 2165400.0 ;
      RECT  744600.0 2151600.0 745800.0 2152800.0 ;
      RECT  747000.0 2151600.0 748200.0 2152800.0 ;
      RECT  744600.0 2158800.0 745800.0 2160000.0 ;
      RECT  749400.0 2158800.0 750600.0 2160000.0 ;
      RECT  741600.0 2154000.0 751800.0 2154900.0 ;
      RECT  741600.0 2165100.0 751800.0 2166000.0 ;
      RECT  757200.0 2158800.0 758400.0 2166000.0 ;
      RECT  754800.0 2151600.0 756000.0 2152800.0 ;
      RECT  757200.0 2151600.0 758400.0 2152800.0 ;
      RECT  757200.0 2151600.0 758400.0 2152800.0 ;
      RECT  754800.0 2151600.0 756000.0 2152800.0 ;
      RECT  754800.0 2158800.0 756000.0 2160000.0 ;
      RECT  757200.0 2158800.0 758400.0 2160000.0 ;
      RECT  757200.0 2158800.0 758400.0 2160000.0 ;
      RECT  754800.0 2158800.0 756000.0 2160000.0 ;
      RECT  757200.0 2158800.0 758400.0 2160000.0 ;
      RECT  759600.0 2158800.0 760800.0 2160000.0 ;
      RECT  759600.0 2158800.0 760800.0 2160000.0 ;
      RECT  757200.0 2158800.0 758400.0 2160000.0 ;
      RECT  756900.0 2153850.0 755700.0 2155050.0 ;
      RECT  757200.0 2164200.0 758400.0 2165400.0 ;
      RECT  754800.0 2151600.0 756000.0 2152800.0 ;
      RECT  757200.0 2151600.0 758400.0 2152800.0 ;
      RECT  754800.0 2158800.0 756000.0 2160000.0 ;
      RECT  759600.0 2158800.0 760800.0 2160000.0 ;
      RECT  751800.0 2154000.0 762000.0 2154900.0 ;
      RECT  751800.0 2165100.0 762000.0 2166000.0 ;
      RECT  767400.0 2158800.0 768600.0 2166000.0 ;
      RECT  765000.0 2151600.0 766200.0 2152800.0 ;
      RECT  767400.0 2151600.0 768600.0 2152800.0 ;
      RECT  767400.0 2151600.0 768600.0 2152800.0 ;
      RECT  765000.0 2151600.0 766200.0 2152800.0 ;
      RECT  765000.0 2158800.0 766200.0 2160000.0 ;
      RECT  767400.0 2158800.0 768600.0 2160000.0 ;
      RECT  767400.0 2158800.0 768600.0 2160000.0 ;
      RECT  765000.0 2158800.0 766200.0 2160000.0 ;
      RECT  767400.0 2158800.0 768600.0 2160000.0 ;
      RECT  769800.0 2158800.0 771000.0 2160000.0 ;
      RECT  769800.0 2158800.0 771000.0 2160000.0 ;
      RECT  767400.0 2158800.0 768600.0 2160000.0 ;
      RECT  767100.0 2153850.0 765900.0 2155050.0 ;
      RECT  767400.0 2164200.0 768600.0 2165400.0 ;
      RECT  765000.0 2151600.0 766200.0 2152800.0 ;
      RECT  767400.0 2151600.0 768600.0 2152800.0 ;
      RECT  765000.0 2158800.0 766200.0 2160000.0 ;
      RECT  769800.0 2158800.0 771000.0 2160000.0 ;
      RECT  762000.0 2154000.0 772200.0 2154900.0 ;
      RECT  762000.0 2165100.0 772200.0 2166000.0 ;
      RECT  777600.0 2158800.0 778800.0 2166000.0 ;
      RECT  775200.0 2151600.0 776400.0 2152800.0 ;
      RECT  777600.0 2151600.0 778800.0 2152800.0 ;
      RECT  777600.0 2151600.0 778800.0 2152800.0 ;
      RECT  775200.0 2151600.0 776400.0 2152800.0 ;
      RECT  775200.0 2158800.0 776400.0 2160000.0 ;
      RECT  777600.0 2158800.0 778800.0 2160000.0 ;
      RECT  777600.0 2158800.0 778800.0 2160000.0 ;
      RECT  775200.0 2158800.0 776400.0 2160000.0 ;
      RECT  777600.0 2158800.0 778800.0 2160000.0 ;
      RECT  780000.0 2158800.0 781200.0 2160000.0 ;
      RECT  780000.0 2158800.0 781200.0 2160000.0 ;
      RECT  777600.0 2158800.0 778800.0 2160000.0 ;
      RECT  777300.0 2153850.0 776100.0 2155050.0 ;
      RECT  777600.0 2164200.0 778800.0 2165400.0 ;
      RECT  775200.0 2151600.0 776400.0 2152800.0 ;
      RECT  777600.0 2151600.0 778800.0 2152800.0 ;
      RECT  775200.0 2158800.0 776400.0 2160000.0 ;
      RECT  780000.0 2158800.0 781200.0 2160000.0 ;
      RECT  772200.0 2154000.0 782400.0 2154900.0 ;
      RECT  772200.0 2165100.0 782400.0 2166000.0 ;
      RECT  787800.0 2158800.0 789000.0 2166000.0 ;
      RECT  785400.0 2151600.0 786600.0 2152800.0 ;
      RECT  787800.0 2151600.0 789000.0 2152800.0 ;
      RECT  787800.0 2151600.0 789000.0 2152800.0 ;
      RECT  785400.0 2151600.0 786600.0 2152800.0 ;
      RECT  785400.0 2158800.0 786600.0 2160000.0 ;
      RECT  787800.0 2158800.0 789000.0 2160000.0 ;
      RECT  787800.0 2158800.0 789000.0 2160000.0 ;
      RECT  785400.0 2158800.0 786600.0 2160000.0 ;
      RECT  787800.0 2158800.0 789000.0 2160000.0 ;
      RECT  790200.0 2158800.0 791400.0 2160000.0 ;
      RECT  790200.0 2158800.0 791400.0 2160000.0 ;
      RECT  787800.0 2158800.0 789000.0 2160000.0 ;
      RECT  787500.0 2153850.0 786300.0 2155050.0 ;
      RECT  787800.0 2164200.0 789000.0 2165400.0 ;
      RECT  785400.0 2151600.0 786600.0 2152800.0 ;
      RECT  787800.0 2151600.0 789000.0 2152800.0 ;
      RECT  785400.0 2158800.0 786600.0 2160000.0 ;
      RECT  790200.0 2158800.0 791400.0 2160000.0 ;
      RECT  782400.0 2154000.0 792600.0 2154900.0 ;
      RECT  782400.0 2165100.0 792600.0 2166000.0 ;
      RECT  798000.0 2158800.0 799200.0 2166000.0 ;
      RECT  795600.0 2151600.0 796800.0 2152800.0 ;
      RECT  798000.0 2151600.0 799200.0 2152800.0 ;
      RECT  798000.0 2151600.0 799200.0 2152800.0 ;
      RECT  795600.0 2151600.0 796800.0 2152800.0 ;
      RECT  795600.0 2158800.0 796800.0 2160000.0 ;
      RECT  798000.0 2158800.0 799200.0 2160000.0 ;
      RECT  798000.0 2158800.0 799200.0 2160000.0 ;
      RECT  795600.0 2158800.0 796800.0 2160000.0 ;
      RECT  798000.0 2158800.0 799200.0 2160000.0 ;
      RECT  800400.0 2158800.0 801600.0 2160000.0 ;
      RECT  800400.0 2158800.0 801600.0 2160000.0 ;
      RECT  798000.0 2158800.0 799200.0 2160000.0 ;
      RECT  797700.0 2153850.0 796500.0 2155050.0 ;
      RECT  798000.0 2164200.0 799200.0 2165400.0 ;
      RECT  795600.0 2151600.0 796800.0 2152800.0 ;
      RECT  798000.0 2151600.0 799200.0 2152800.0 ;
      RECT  795600.0 2158800.0 796800.0 2160000.0 ;
      RECT  800400.0 2158800.0 801600.0 2160000.0 ;
      RECT  792600.0 2154000.0 802800.0 2154900.0 ;
      RECT  792600.0 2165100.0 802800.0 2166000.0 ;
      RECT  808200.0 2158800.0 809400.0 2166000.0 ;
      RECT  805800.0 2151600.0 807000.0 2152800.0 ;
      RECT  808200.0 2151600.0 809400.0 2152800.0 ;
      RECT  808200.0 2151600.0 809400.0 2152800.0 ;
      RECT  805800.0 2151600.0 807000.0 2152800.0 ;
      RECT  805800.0 2158800.0 807000.0 2160000.0 ;
      RECT  808200.0 2158800.0 809400.0 2160000.0 ;
      RECT  808200.0 2158800.0 809400.0 2160000.0 ;
      RECT  805800.0 2158800.0 807000.0 2160000.0 ;
      RECT  808200.0 2158800.0 809400.0 2160000.0 ;
      RECT  810600.0 2158800.0 811800.0 2160000.0 ;
      RECT  810600.0 2158800.0 811800.0 2160000.0 ;
      RECT  808200.0 2158800.0 809400.0 2160000.0 ;
      RECT  807900.0 2153850.0 806700.0 2155050.0 ;
      RECT  808200.0 2164200.0 809400.0 2165400.0 ;
      RECT  805800.0 2151600.0 807000.0 2152800.0 ;
      RECT  808200.0 2151600.0 809400.0 2152800.0 ;
      RECT  805800.0 2158800.0 807000.0 2160000.0 ;
      RECT  810600.0 2158800.0 811800.0 2160000.0 ;
      RECT  802800.0 2154000.0 813000.0 2154900.0 ;
      RECT  802800.0 2165100.0 813000.0 2166000.0 ;
      RECT  818400.0 2158800.0 819600.0 2166000.0 ;
      RECT  816000.0 2151600.0 817200.0 2152800.0 ;
      RECT  818400.0 2151600.0 819600.0 2152800.0 ;
      RECT  818400.0 2151600.0 819600.0 2152800.0 ;
      RECT  816000.0 2151600.0 817200.0 2152800.0 ;
      RECT  816000.0 2158800.0 817200.0 2160000.0 ;
      RECT  818400.0 2158800.0 819600.0 2160000.0 ;
      RECT  818400.0 2158800.0 819600.0 2160000.0 ;
      RECT  816000.0 2158800.0 817200.0 2160000.0 ;
      RECT  818400.0 2158800.0 819600.0 2160000.0 ;
      RECT  820800.0 2158800.0 822000.0 2160000.0 ;
      RECT  820800.0 2158800.0 822000.0 2160000.0 ;
      RECT  818400.0 2158800.0 819600.0 2160000.0 ;
      RECT  818100.0 2153850.0 816900.0 2155050.0 ;
      RECT  818400.0 2164200.0 819600.0 2165400.0 ;
      RECT  816000.0 2151600.0 817200.0 2152800.0 ;
      RECT  818400.0 2151600.0 819600.0 2152800.0 ;
      RECT  816000.0 2158800.0 817200.0 2160000.0 ;
      RECT  820800.0 2158800.0 822000.0 2160000.0 ;
      RECT  813000.0 2154000.0 823200.0 2154900.0 ;
      RECT  813000.0 2165100.0 823200.0 2166000.0 ;
      RECT  828600.0 2158800.0 829800.0 2166000.0 ;
      RECT  826200.0 2151600.0 827400.0 2152800.0 ;
      RECT  828600.0 2151600.0 829800.0 2152800.0 ;
      RECT  828600.0 2151600.0 829800.0 2152800.0 ;
      RECT  826200.0 2151600.0 827400.0 2152800.0 ;
      RECT  826200.0 2158800.0 827400.0 2160000.0 ;
      RECT  828600.0 2158800.0 829800.0 2160000.0 ;
      RECT  828600.0 2158800.0 829800.0 2160000.0 ;
      RECT  826200.0 2158800.0 827400.0 2160000.0 ;
      RECT  828600.0 2158800.0 829800.0 2160000.0 ;
      RECT  831000.0 2158800.0 832200.0 2160000.0 ;
      RECT  831000.0 2158800.0 832200.0 2160000.0 ;
      RECT  828600.0 2158800.0 829800.0 2160000.0 ;
      RECT  828300.0 2153850.0 827100.0 2155050.0 ;
      RECT  828600.0 2164200.0 829800.0 2165400.0 ;
      RECT  826200.0 2151600.0 827400.0 2152800.0 ;
      RECT  828600.0 2151600.0 829800.0 2152800.0 ;
      RECT  826200.0 2158800.0 827400.0 2160000.0 ;
      RECT  831000.0 2158800.0 832200.0 2160000.0 ;
      RECT  823200.0 2154000.0 833400.0 2154900.0 ;
      RECT  823200.0 2165100.0 833400.0 2166000.0 ;
      RECT  838800.0 2158800.0 840000.0 2166000.0 ;
      RECT  836400.0 2151600.0 837600.0 2152800.0 ;
      RECT  838800.0 2151600.0 840000.0 2152800.0 ;
      RECT  838800.0 2151600.0 840000.0 2152800.0 ;
      RECT  836400.0 2151600.0 837600.0 2152800.0 ;
      RECT  836400.0 2158800.0 837600.0 2160000.0 ;
      RECT  838800.0 2158800.0 840000.0 2160000.0 ;
      RECT  838800.0 2158800.0 840000.0 2160000.0 ;
      RECT  836400.0 2158800.0 837600.0 2160000.0 ;
      RECT  838800.0 2158800.0 840000.0 2160000.0 ;
      RECT  841200.0 2158800.0 842400.0 2160000.0 ;
      RECT  841200.0 2158800.0 842400.0 2160000.0 ;
      RECT  838800.0 2158800.0 840000.0 2160000.0 ;
      RECT  838500.0 2153850.0 837300.0 2155050.0 ;
      RECT  838800.0 2164200.0 840000.0 2165400.0 ;
      RECT  836400.0 2151600.0 837600.0 2152800.0 ;
      RECT  838800.0 2151600.0 840000.0 2152800.0 ;
      RECT  836400.0 2158800.0 837600.0 2160000.0 ;
      RECT  841200.0 2158800.0 842400.0 2160000.0 ;
      RECT  833400.0 2154000.0 843600.0 2154900.0 ;
      RECT  833400.0 2165100.0 843600.0 2166000.0 ;
      RECT  849000.0 2158800.0 850200.0 2166000.0 ;
      RECT  846600.0 2151600.0 847800.0 2152800.0 ;
      RECT  849000.0 2151600.0 850200.0 2152800.0 ;
      RECT  849000.0 2151600.0 850200.0 2152800.0 ;
      RECT  846600.0 2151600.0 847800.0 2152800.0 ;
      RECT  846600.0 2158800.0 847800.0 2160000.0 ;
      RECT  849000.0 2158800.0 850200.0 2160000.0 ;
      RECT  849000.0 2158800.0 850200.0 2160000.0 ;
      RECT  846600.0 2158800.0 847800.0 2160000.0 ;
      RECT  849000.0 2158800.0 850200.0 2160000.0 ;
      RECT  851400.0 2158800.0 852600.0 2160000.0 ;
      RECT  851400.0 2158800.0 852600.0 2160000.0 ;
      RECT  849000.0 2158800.0 850200.0 2160000.0 ;
      RECT  848700.0 2153850.0 847500.0 2155050.0 ;
      RECT  849000.0 2164200.0 850200.0 2165400.0 ;
      RECT  846600.0 2151600.0 847800.0 2152800.0 ;
      RECT  849000.0 2151600.0 850200.0 2152800.0 ;
      RECT  846600.0 2158800.0 847800.0 2160000.0 ;
      RECT  851400.0 2158800.0 852600.0 2160000.0 ;
      RECT  843600.0 2154000.0 853800.0 2154900.0 ;
      RECT  843600.0 2165100.0 853800.0 2166000.0 ;
      RECT  859200.0 2158800.0 860400.0 2166000.0 ;
      RECT  856800.0 2151600.0 858000.0 2152800.0 ;
      RECT  859200.0 2151600.0 860400.0 2152800.0 ;
      RECT  859200.0 2151600.0 860400.0 2152800.0 ;
      RECT  856800.0 2151600.0 858000.0 2152800.0 ;
      RECT  856800.0 2158800.0 858000.0 2160000.0 ;
      RECT  859200.0 2158800.0 860400.0 2160000.0 ;
      RECT  859200.0 2158800.0 860400.0 2160000.0 ;
      RECT  856800.0 2158800.0 858000.0 2160000.0 ;
      RECT  859200.0 2158800.0 860400.0 2160000.0 ;
      RECT  861600.0 2158800.0 862800.0 2160000.0 ;
      RECT  861600.0 2158800.0 862800.0 2160000.0 ;
      RECT  859200.0 2158800.0 860400.0 2160000.0 ;
      RECT  858900.0 2153850.0 857700.0 2155050.0 ;
      RECT  859200.0 2164200.0 860400.0 2165400.0 ;
      RECT  856800.0 2151600.0 858000.0 2152800.0 ;
      RECT  859200.0 2151600.0 860400.0 2152800.0 ;
      RECT  856800.0 2158800.0 858000.0 2160000.0 ;
      RECT  861600.0 2158800.0 862800.0 2160000.0 ;
      RECT  853800.0 2154000.0 864000.0 2154900.0 ;
      RECT  853800.0 2165100.0 864000.0 2166000.0 ;
      RECT  869400.0 2158800.0 870600.0 2166000.0 ;
      RECT  867000.0 2151600.0 868200.0 2152800.0 ;
      RECT  869400.0 2151600.0 870600.0 2152800.0 ;
      RECT  869400.0 2151600.0 870600.0 2152800.0 ;
      RECT  867000.0 2151600.0 868200.0 2152800.0 ;
      RECT  867000.0 2158800.0 868200.0 2160000.0 ;
      RECT  869400.0 2158800.0 870600.0 2160000.0 ;
      RECT  869400.0 2158800.0 870600.0 2160000.0 ;
      RECT  867000.0 2158800.0 868200.0 2160000.0 ;
      RECT  869400.0 2158800.0 870600.0 2160000.0 ;
      RECT  871800.0 2158800.0 873000.0 2160000.0 ;
      RECT  871800.0 2158800.0 873000.0 2160000.0 ;
      RECT  869400.0 2158800.0 870600.0 2160000.0 ;
      RECT  869100.0 2153850.0 867900.0 2155050.0 ;
      RECT  869400.0 2164200.0 870600.0 2165400.0 ;
      RECT  867000.0 2151600.0 868200.0 2152800.0 ;
      RECT  869400.0 2151600.0 870600.0 2152800.0 ;
      RECT  867000.0 2158800.0 868200.0 2160000.0 ;
      RECT  871800.0 2158800.0 873000.0 2160000.0 ;
      RECT  864000.0 2154000.0 874200.0 2154900.0 ;
      RECT  864000.0 2165100.0 874200.0 2166000.0 ;
      RECT  879600.0 2158800.0 880800.0 2166000.0 ;
      RECT  877200.0 2151600.0 878400.0 2152800.0 ;
      RECT  879600.0 2151600.0 880800.0 2152800.0 ;
      RECT  879600.0 2151600.0 880800.0 2152800.0 ;
      RECT  877200.0 2151600.0 878400.0 2152800.0 ;
      RECT  877200.0 2158800.0 878400.0 2160000.0 ;
      RECT  879600.0 2158800.0 880800.0 2160000.0 ;
      RECT  879600.0 2158800.0 880800.0 2160000.0 ;
      RECT  877200.0 2158800.0 878400.0 2160000.0 ;
      RECT  879600.0 2158800.0 880800.0 2160000.0 ;
      RECT  882000.0 2158800.0 883200.0 2160000.0 ;
      RECT  882000.0 2158800.0 883200.0 2160000.0 ;
      RECT  879600.0 2158800.0 880800.0 2160000.0 ;
      RECT  879300.0 2153850.0 878100.0 2155050.0 ;
      RECT  879600.0 2164200.0 880800.0 2165400.0 ;
      RECT  877200.0 2151600.0 878400.0 2152800.0 ;
      RECT  879600.0 2151600.0 880800.0 2152800.0 ;
      RECT  877200.0 2158800.0 878400.0 2160000.0 ;
      RECT  882000.0 2158800.0 883200.0 2160000.0 ;
      RECT  874200.0 2154000.0 884400.0 2154900.0 ;
      RECT  874200.0 2165100.0 884400.0 2166000.0 ;
      RECT  889800.0 2158800.0 891000.0 2166000.0 ;
      RECT  887400.0 2151600.0 888600.0 2152800.0 ;
      RECT  889800.0 2151600.0 891000.0 2152800.0 ;
      RECT  889800.0 2151600.0 891000.0 2152800.0 ;
      RECT  887400.0 2151600.0 888600.0 2152800.0 ;
      RECT  887400.0 2158800.0 888600.0 2160000.0 ;
      RECT  889800.0 2158800.0 891000.0 2160000.0 ;
      RECT  889800.0 2158800.0 891000.0 2160000.0 ;
      RECT  887400.0 2158800.0 888600.0 2160000.0 ;
      RECT  889800.0 2158800.0 891000.0 2160000.0 ;
      RECT  892200.0 2158800.0 893400.0 2160000.0 ;
      RECT  892200.0 2158800.0 893400.0 2160000.0 ;
      RECT  889800.0 2158800.0 891000.0 2160000.0 ;
      RECT  889500.0 2153850.0 888300.0 2155050.0 ;
      RECT  889800.0 2164200.0 891000.0 2165400.0 ;
      RECT  887400.0 2151600.0 888600.0 2152800.0 ;
      RECT  889800.0 2151600.0 891000.0 2152800.0 ;
      RECT  887400.0 2158800.0 888600.0 2160000.0 ;
      RECT  892200.0 2158800.0 893400.0 2160000.0 ;
      RECT  884400.0 2154000.0 894600.0 2154900.0 ;
      RECT  884400.0 2165100.0 894600.0 2166000.0 ;
      RECT  900000.0 2158800.0 901200.0 2166000.0 ;
      RECT  897600.0 2151600.0 898800.0 2152800.0 ;
      RECT  900000.0 2151600.0 901200.0 2152800.0 ;
      RECT  900000.0 2151600.0 901200.0 2152800.0 ;
      RECT  897600.0 2151600.0 898800.0 2152800.0 ;
      RECT  897600.0 2158800.0 898800.0 2160000.0 ;
      RECT  900000.0 2158800.0 901200.0 2160000.0 ;
      RECT  900000.0 2158800.0 901200.0 2160000.0 ;
      RECT  897600.0 2158800.0 898800.0 2160000.0 ;
      RECT  900000.0 2158800.0 901200.0 2160000.0 ;
      RECT  902400.0 2158800.0 903600.0 2160000.0 ;
      RECT  902400.0 2158800.0 903600.0 2160000.0 ;
      RECT  900000.0 2158800.0 901200.0 2160000.0 ;
      RECT  899700.0 2153850.0 898500.0 2155050.0 ;
      RECT  900000.0 2164200.0 901200.0 2165400.0 ;
      RECT  897600.0 2151600.0 898800.0 2152800.0 ;
      RECT  900000.0 2151600.0 901200.0 2152800.0 ;
      RECT  897600.0 2158800.0 898800.0 2160000.0 ;
      RECT  902400.0 2158800.0 903600.0 2160000.0 ;
      RECT  894600.0 2154000.0 904800.0 2154900.0 ;
      RECT  894600.0 2165100.0 904800.0 2166000.0 ;
      RECT  910200.0 2158800.0 911400.0 2166000.0 ;
      RECT  907800.0 2151600.0 909000.0 2152800.0 ;
      RECT  910200.0 2151600.0 911400.0 2152800.0 ;
      RECT  910200.0 2151600.0 911400.0 2152800.0 ;
      RECT  907800.0 2151600.0 909000.0 2152800.0 ;
      RECT  907800.0 2158800.0 909000.0 2160000.0 ;
      RECT  910200.0 2158800.0 911400.0 2160000.0 ;
      RECT  910200.0 2158800.0 911400.0 2160000.0 ;
      RECT  907800.0 2158800.0 909000.0 2160000.0 ;
      RECT  910200.0 2158800.0 911400.0 2160000.0 ;
      RECT  912600.0 2158800.0 913800.0 2160000.0 ;
      RECT  912600.0 2158800.0 913800.0 2160000.0 ;
      RECT  910200.0 2158800.0 911400.0 2160000.0 ;
      RECT  909900.0 2153850.0 908700.0 2155050.0 ;
      RECT  910200.0 2164200.0 911400.0 2165400.0 ;
      RECT  907800.0 2151600.0 909000.0 2152800.0 ;
      RECT  910200.0 2151600.0 911400.0 2152800.0 ;
      RECT  907800.0 2158800.0 909000.0 2160000.0 ;
      RECT  912600.0 2158800.0 913800.0 2160000.0 ;
      RECT  904800.0 2154000.0 915000.0 2154900.0 ;
      RECT  904800.0 2165100.0 915000.0 2166000.0 ;
      RECT  920400.0 2158800.0 921600.0 2166000.0 ;
      RECT  918000.0 2151600.0 919200.0 2152800.0 ;
      RECT  920400.0 2151600.0 921600.0 2152800.0 ;
      RECT  920400.0 2151600.0 921600.0 2152800.0 ;
      RECT  918000.0 2151600.0 919200.0 2152800.0 ;
      RECT  918000.0 2158800.0 919200.0 2160000.0 ;
      RECT  920400.0 2158800.0 921600.0 2160000.0 ;
      RECT  920400.0 2158800.0 921600.0 2160000.0 ;
      RECT  918000.0 2158800.0 919200.0 2160000.0 ;
      RECT  920400.0 2158800.0 921600.0 2160000.0 ;
      RECT  922800.0 2158800.0 924000.0 2160000.0 ;
      RECT  922800.0 2158800.0 924000.0 2160000.0 ;
      RECT  920400.0 2158800.0 921600.0 2160000.0 ;
      RECT  920100.0 2153850.0 918900.0 2155050.0 ;
      RECT  920400.0 2164200.0 921600.0 2165400.0 ;
      RECT  918000.0 2151600.0 919200.0 2152800.0 ;
      RECT  920400.0 2151600.0 921600.0 2152800.0 ;
      RECT  918000.0 2158800.0 919200.0 2160000.0 ;
      RECT  922800.0 2158800.0 924000.0 2160000.0 ;
      RECT  915000.0 2154000.0 925200.0 2154900.0 ;
      RECT  915000.0 2165100.0 925200.0 2166000.0 ;
      RECT  930600.0 2158800.0 931800.0 2166000.0 ;
      RECT  928200.0 2151600.0 929400.0 2152800.0 ;
      RECT  930600.0 2151600.0 931800.0 2152800.0 ;
      RECT  930600.0 2151600.0 931800.0 2152800.0 ;
      RECT  928200.0 2151600.0 929400.0 2152800.0 ;
      RECT  928200.0 2158800.0 929400.0 2160000.0 ;
      RECT  930600.0 2158800.0 931800.0 2160000.0 ;
      RECT  930600.0 2158800.0 931800.0 2160000.0 ;
      RECT  928200.0 2158800.0 929400.0 2160000.0 ;
      RECT  930600.0 2158800.0 931800.0 2160000.0 ;
      RECT  933000.0 2158800.0 934200.0 2160000.0 ;
      RECT  933000.0 2158800.0 934200.0 2160000.0 ;
      RECT  930600.0 2158800.0 931800.0 2160000.0 ;
      RECT  930300.0 2153850.0 929100.0 2155050.0 ;
      RECT  930600.0 2164200.0 931800.0 2165400.0 ;
      RECT  928200.0 2151600.0 929400.0 2152800.0 ;
      RECT  930600.0 2151600.0 931800.0 2152800.0 ;
      RECT  928200.0 2158800.0 929400.0 2160000.0 ;
      RECT  933000.0 2158800.0 934200.0 2160000.0 ;
      RECT  925200.0 2154000.0 935400.0 2154900.0 ;
      RECT  925200.0 2165100.0 935400.0 2166000.0 ;
      RECT  940800.0 2158800.0 942000.0 2166000.0 ;
      RECT  938400.0 2151600.0 939600.0 2152800.0 ;
      RECT  940800.0 2151600.0 942000.0 2152800.0 ;
      RECT  940800.0 2151600.0 942000.0 2152800.0 ;
      RECT  938400.0 2151600.0 939600.0 2152800.0 ;
      RECT  938400.0 2158800.0 939600.0 2160000.0 ;
      RECT  940800.0 2158800.0 942000.0 2160000.0 ;
      RECT  940800.0 2158800.0 942000.0 2160000.0 ;
      RECT  938400.0 2158800.0 939600.0 2160000.0 ;
      RECT  940800.0 2158800.0 942000.0 2160000.0 ;
      RECT  943200.0 2158800.0 944400.0 2160000.0 ;
      RECT  943200.0 2158800.0 944400.0 2160000.0 ;
      RECT  940800.0 2158800.0 942000.0 2160000.0 ;
      RECT  940500.0 2153850.0 939300.0 2155050.0 ;
      RECT  940800.0 2164200.0 942000.0 2165400.0 ;
      RECT  938400.0 2151600.0 939600.0 2152800.0 ;
      RECT  940800.0 2151600.0 942000.0 2152800.0 ;
      RECT  938400.0 2158800.0 939600.0 2160000.0 ;
      RECT  943200.0 2158800.0 944400.0 2160000.0 ;
      RECT  935400.0 2154000.0 945600.0 2154900.0 ;
      RECT  935400.0 2165100.0 945600.0 2166000.0 ;
      RECT  951000.0 2158800.0 952200.0 2166000.0 ;
      RECT  948600.0 2151600.0 949800.0 2152800.0 ;
      RECT  951000.0 2151600.0 952200.0 2152800.0 ;
      RECT  951000.0 2151600.0 952200.0 2152800.0 ;
      RECT  948600.0 2151600.0 949800.0 2152800.0 ;
      RECT  948600.0 2158800.0 949800.0 2160000.0 ;
      RECT  951000.0 2158800.0 952200.0 2160000.0 ;
      RECT  951000.0 2158800.0 952200.0 2160000.0 ;
      RECT  948600.0 2158800.0 949800.0 2160000.0 ;
      RECT  951000.0 2158800.0 952200.0 2160000.0 ;
      RECT  953400.0 2158800.0 954600.0 2160000.0 ;
      RECT  953400.0 2158800.0 954600.0 2160000.0 ;
      RECT  951000.0 2158800.0 952200.0 2160000.0 ;
      RECT  950700.0 2153850.0 949500.0 2155050.0 ;
      RECT  951000.0 2164200.0 952200.0 2165400.0 ;
      RECT  948600.0 2151600.0 949800.0 2152800.0 ;
      RECT  951000.0 2151600.0 952200.0 2152800.0 ;
      RECT  948600.0 2158800.0 949800.0 2160000.0 ;
      RECT  953400.0 2158800.0 954600.0 2160000.0 ;
      RECT  945600.0 2154000.0 955800.0 2154900.0 ;
      RECT  945600.0 2165100.0 955800.0 2166000.0 ;
      RECT  961200.0 2158800.0 962400.0 2166000.0 ;
      RECT  958800.0 2151600.0 960000.0 2152800.0 ;
      RECT  961200.0 2151600.0 962400.0 2152800.0 ;
      RECT  961200.0 2151600.0 962400.0 2152800.0 ;
      RECT  958800.0 2151600.0 960000.0 2152800.0 ;
      RECT  958800.0 2158800.0 960000.0 2160000.0 ;
      RECT  961200.0 2158800.0 962400.0 2160000.0 ;
      RECT  961200.0 2158800.0 962400.0 2160000.0 ;
      RECT  958800.0 2158800.0 960000.0 2160000.0 ;
      RECT  961200.0 2158800.0 962400.0 2160000.0 ;
      RECT  963600.0 2158800.0 964800.0 2160000.0 ;
      RECT  963600.0 2158800.0 964800.0 2160000.0 ;
      RECT  961200.0 2158800.0 962400.0 2160000.0 ;
      RECT  960900.0 2153850.0 959700.0 2155050.0 ;
      RECT  961200.0 2164200.0 962400.0 2165400.0 ;
      RECT  958800.0 2151600.0 960000.0 2152800.0 ;
      RECT  961200.0 2151600.0 962400.0 2152800.0 ;
      RECT  958800.0 2158800.0 960000.0 2160000.0 ;
      RECT  963600.0 2158800.0 964800.0 2160000.0 ;
      RECT  955800.0 2154000.0 966000.0 2154900.0 ;
      RECT  955800.0 2165100.0 966000.0 2166000.0 ;
      RECT  971400.0 2158800.0 972600.0 2166000.0 ;
      RECT  969000.0 2151600.0 970200.0 2152800.0 ;
      RECT  971400.0 2151600.0 972600.0 2152800.0 ;
      RECT  971400.0 2151600.0 972600.0 2152800.0 ;
      RECT  969000.0 2151600.0 970200.0 2152800.0 ;
      RECT  969000.0 2158800.0 970200.0 2160000.0 ;
      RECT  971400.0 2158800.0 972600.0 2160000.0 ;
      RECT  971400.0 2158800.0 972600.0 2160000.0 ;
      RECT  969000.0 2158800.0 970200.0 2160000.0 ;
      RECT  971400.0 2158800.0 972600.0 2160000.0 ;
      RECT  973800.0 2158800.0 975000.0 2160000.0 ;
      RECT  973800.0 2158800.0 975000.0 2160000.0 ;
      RECT  971400.0 2158800.0 972600.0 2160000.0 ;
      RECT  971100.0 2153850.0 969900.0 2155050.0 ;
      RECT  971400.0 2164200.0 972600.0 2165400.0 ;
      RECT  969000.0 2151600.0 970200.0 2152800.0 ;
      RECT  971400.0 2151600.0 972600.0 2152800.0 ;
      RECT  969000.0 2158800.0 970200.0 2160000.0 ;
      RECT  973800.0 2158800.0 975000.0 2160000.0 ;
      RECT  966000.0 2154000.0 976200.0 2154900.0 ;
      RECT  966000.0 2165100.0 976200.0 2166000.0 ;
      RECT  981600.0 2158800.0 982800.0 2166000.0 ;
      RECT  979200.0 2151600.0 980400.0 2152800.0 ;
      RECT  981600.0 2151600.0 982800.0 2152800.0 ;
      RECT  981600.0 2151600.0 982800.0 2152800.0 ;
      RECT  979200.0 2151600.0 980400.0 2152800.0 ;
      RECT  979200.0 2158800.0 980400.0 2160000.0 ;
      RECT  981600.0 2158800.0 982800.0 2160000.0 ;
      RECT  981600.0 2158800.0 982800.0 2160000.0 ;
      RECT  979200.0 2158800.0 980400.0 2160000.0 ;
      RECT  981600.0 2158800.0 982800.0 2160000.0 ;
      RECT  984000.0 2158800.0 985200.0 2160000.0 ;
      RECT  984000.0 2158800.0 985200.0 2160000.0 ;
      RECT  981600.0 2158800.0 982800.0 2160000.0 ;
      RECT  981300.0 2153850.0 980100.0 2155050.0 ;
      RECT  981600.0 2164200.0 982800.0 2165400.0 ;
      RECT  979200.0 2151600.0 980400.0 2152800.0 ;
      RECT  981600.0 2151600.0 982800.0 2152800.0 ;
      RECT  979200.0 2158800.0 980400.0 2160000.0 ;
      RECT  984000.0 2158800.0 985200.0 2160000.0 ;
      RECT  976200.0 2154000.0 986400.0 2154900.0 ;
      RECT  976200.0 2165100.0 986400.0 2166000.0 ;
      RECT  991800.0 2158800.0 993000.0 2166000.0 ;
      RECT  989400.0 2151600.0 990600.0 2152800.0 ;
      RECT  991800.0 2151600.0 993000.0 2152800.0 ;
      RECT  991800.0 2151600.0 993000.0 2152800.0 ;
      RECT  989400.0 2151600.0 990600.0 2152800.0 ;
      RECT  989400.0 2158800.0 990600.0 2160000.0 ;
      RECT  991800.0 2158800.0 993000.0 2160000.0 ;
      RECT  991800.0 2158800.0 993000.0 2160000.0 ;
      RECT  989400.0 2158800.0 990600.0 2160000.0 ;
      RECT  991800.0 2158800.0 993000.0 2160000.0 ;
      RECT  994200.0 2158800.0 995400.0 2160000.0 ;
      RECT  994200.0 2158800.0 995400.0 2160000.0 ;
      RECT  991800.0 2158800.0 993000.0 2160000.0 ;
      RECT  991500.0 2153850.0 990300.0 2155050.0 ;
      RECT  991800.0 2164200.0 993000.0 2165400.0 ;
      RECT  989400.0 2151600.0 990600.0 2152800.0 ;
      RECT  991800.0 2151600.0 993000.0 2152800.0 ;
      RECT  989400.0 2158800.0 990600.0 2160000.0 ;
      RECT  994200.0 2158800.0 995400.0 2160000.0 ;
      RECT  986400.0 2154000.0 996600.0 2154900.0 ;
      RECT  986400.0 2165100.0 996600.0 2166000.0 ;
      RECT  1002000.0 2158800.0 1003200.0 2166000.0 ;
      RECT  999600.0 2151600.0 1000800.0 2152800.0 ;
      RECT  1002000.0 2151600.0 1003200.0 2152800.0 ;
      RECT  1002000.0 2151600.0 1003200.0 2152800.0 ;
      RECT  999600.0 2151600.0 1000800.0 2152800.0 ;
      RECT  999600.0 2158800.0 1000800.0 2160000.0 ;
      RECT  1002000.0 2158800.0 1003200.0 2160000.0 ;
      RECT  1002000.0 2158800.0 1003200.0 2160000.0 ;
      RECT  999600.0 2158800.0 1000800.0 2160000.0 ;
      RECT  1002000.0 2158800.0 1003200.0 2160000.0 ;
      RECT  1004400.0 2158800.0 1005600.0 2160000.0 ;
      RECT  1004400.0 2158800.0 1005600.0 2160000.0 ;
      RECT  1002000.0 2158800.0 1003200.0 2160000.0 ;
      RECT  1001700.0 2153850.0 1000500.0 2155050.0 ;
      RECT  1002000.0 2164200.0 1003200.0 2165400.0 ;
      RECT  999600.0 2151600.0 1000800.0 2152800.0 ;
      RECT  1002000.0 2151600.0 1003200.0 2152800.0 ;
      RECT  999600.0 2158800.0 1000800.0 2160000.0 ;
      RECT  1004400.0 2158800.0 1005600.0 2160000.0 ;
      RECT  996600.0 2154000.0 1006800.0 2154900.0 ;
      RECT  996600.0 2165100.0 1006800.0 2166000.0 ;
      RECT  1012200.0 2158800.0 1013400.0 2166000.0 ;
      RECT  1009800.0 2151600.0 1011000.0 2152800.0 ;
      RECT  1012200.0 2151600.0 1013400.0 2152800.0 ;
      RECT  1012200.0 2151600.0 1013400.0 2152800.0 ;
      RECT  1009800.0 2151600.0 1011000.0 2152800.0 ;
      RECT  1009800.0 2158800.0 1011000.0 2160000.0 ;
      RECT  1012200.0 2158800.0 1013400.0 2160000.0 ;
      RECT  1012200.0 2158800.0 1013400.0 2160000.0 ;
      RECT  1009800.0 2158800.0 1011000.0 2160000.0 ;
      RECT  1012200.0 2158800.0 1013400.0 2160000.0 ;
      RECT  1014600.0 2158800.0 1015800.0 2160000.0 ;
      RECT  1014600.0 2158800.0 1015800.0 2160000.0 ;
      RECT  1012200.0 2158800.0 1013400.0 2160000.0 ;
      RECT  1011900.0 2153850.0 1010700.0 2155050.0 ;
      RECT  1012200.0 2164200.0 1013400.0 2165400.0 ;
      RECT  1009800.0 2151600.0 1011000.0 2152800.0 ;
      RECT  1012200.0 2151600.0 1013400.0 2152800.0 ;
      RECT  1009800.0 2158800.0 1011000.0 2160000.0 ;
      RECT  1014600.0 2158800.0 1015800.0 2160000.0 ;
      RECT  1006800.0 2154000.0 1017000.0 2154900.0 ;
      RECT  1006800.0 2165100.0 1017000.0 2166000.0 ;
      RECT  1022400.0 2158800.0 1023600.0 2166000.0 ;
      RECT  1020000.0 2151600.0 1021200.0 2152800.0 ;
      RECT  1022400.0 2151600.0 1023600.0 2152800.0 ;
      RECT  1022400.0 2151600.0 1023600.0 2152800.0 ;
      RECT  1020000.0 2151600.0 1021200.0 2152800.0 ;
      RECT  1020000.0 2158800.0 1021200.0 2160000.0 ;
      RECT  1022400.0 2158800.0 1023600.0 2160000.0 ;
      RECT  1022400.0 2158800.0 1023600.0 2160000.0 ;
      RECT  1020000.0 2158800.0 1021200.0 2160000.0 ;
      RECT  1022400.0 2158800.0 1023600.0 2160000.0 ;
      RECT  1024800.0 2158800.0 1026000.0 2160000.0 ;
      RECT  1024800.0 2158800.0 1026000.0 2160000.0 ;
      RECT  1022400.0 2158800.0 1023600.0 2160000.0 ;
      RECT  1022100.0 2153850.0 1020900.0 2155050.0 ;
      RECT  1022400.0 2164200.0 1023600.0 2165400.0 ;
      RECT  1020000.0 2151600.0 1021200.0 2152800.0 ;
      RECT  1022400.0 2151600.0 1023600.0 2152800.0 ;
      RECT  1020000.0 2158800.0 1021200.0 2160000.0 ;
      RECT  1024800.0 2158800.0 1026000.0 2160000.0 ;
      RECT  1017000.0 2154000.0 1027200.0 2154900.0 ;
      RECT  1017000.0 2165100.0 1027200.0 2166000.0 ;
      RECT  1032600.0 2158800.0 1033800.0 2166000.0 ;
      RECT  1030200.0 2151600.0 1031400.0 2152800.0 ;
      RECT  1032600.0 2151600.0 1033800.0 2152800.0 ;
      RECT  1032600.0 2151600.0 1033800.0 2152800.0 ;
      RECT  1030200.0 2151600.0 1031400.0 2152800.0 ;
      RECT  1030200.0 2158800.0 1031400.0 2160000.0 ;
      RECT  1032600.0 2158800.0 1033800.0 2160000.0 ;
      RECT  1032600.0 2158800.0 1033800.0 2160000.0 ;
      RECT  1030200.0 2158800.0 1031400.0 2160000.0 ;
      RECT  1032600.0 2158800.0 1033800.0 2160000.0 ;
      RECT  1035000.0 2158800.0 1036200.0 2160000.0 ;
      RECT  1035000.0 2158800.0 1036200.0 2160000.0 ;
      RECT  1032600.0 2158800.0 1033800.0 2160000.0 ;
      RECT  1032300.0 2153850.0 1031100.0 2155050.0 ;
      RECT  1032600.0 2164200.0 1033800.0 2165400.0 ;
      RECT  1030200.0 2151600.0 1031400.0 2152800.0 ;
      RECT  1032600.0 2151600.0 1033800.0 2152800.0 ;
      RECT  1030200.0 2158800.0 1031400.0 2160000.0 ;
      RECT  1035000.0 2158800.0 1036200.0 2160000.0 ;
      RECT  1027200.0 2154000.0 1037400.0 2154900.0 ;
      RECT  1027200.0 2165100.0 1037400.0 2166000.0 ;
      RECT  1042800.0 2158800.0 1044000.0 2166000.0 ;
      RECT  1040400.0 2151600.0 1041600.0 2152800.0 ;
      RECT  1042800.0 2151600.0 1044000.0 2152800.0 ;
      RECT  1042800.0 2151600.0 1044000.0 2152800.0 ;
      RECT  1040400.0 2151600.0 1041600.0 2152800.0 ;
      RECT  1040400.0 2158800.0 1041600.0 2160000.0 ;
      RECT  1042800.0 2158800.0 1044000.0 2160000.0 ;
      RECT  1042800.0 2158800.0 1044000.0 2160000.0 ;
      RECT  1040400.0 2158800.0 1041600.0 2160000.0 ;
      RECT  1042800.0 2158800.0 1044000.0 2160000.0 ;
      RECT  1045200.0 2158800.0 1046400.0 2160000.0 ;
      RECT  1045200.0 2158800.0 1046400.0 2160000.0 ;
      RECT  1042800.0 2158800.0 1044000.0 2160000.0 ;
      RECT  1042500.0 2153850.0 1041300.0 2155050.0 ;
      RECT  1042800.0 2164200.0 1044000.0 2165400.0 ;
      RECT  1040400.0 2151600.0 1041600.0 2152800.0 ;
      RECT  1042800.0 2151600.0 1044000.0 2152800.0 ;
      RECT  1040400.0 2158800.0 1041600.0 2160000.0 ;
      RECT  1045200.0 2158800.0 1046400.0 2160000.0 ;
      RECT  1037400.0 2154000.0 1047600.0 2154900.0 ;
      RECT  1037400.0 2165100.0 1047600.0 2166000.0 ;
      RECT  1053000.0 2158800.0 1054200.0 2166000.0 ;
      RECT  1050600.0 2151600.0 1051800.0 2152800.0 ;
      RECT  1053000.0 2151600.0 1054200.0 2152800.0 ;
      RECT  1053000.0 2151600.0 1054200.0 2152800.0 ;
      RECT  1050600.0 2151600.0 1051800.0 2152800.0 ;
      RECT  1050600.0 2158800.0 1051800.0 2160000.0 ;
      RECT  1053000.0 2158800.0 1054200.0 2160000.0 ;
      RECT  1053000.0 2158800.0 1054200.0 2160000.0 ;
      RECT  1050600.0 2158800.0 1051800.0 2160000.0 ;
      RECT  1053000.0 2158800.0 1054200.0 2160000.0 ;
      RECT  1055400.0 2158800.0 1056600.0 2160000.0 ;
      RECT  1055400.0 2158800.0 1056600.0 2160000.0 ;
      RECT  1053000.0 2158800.0 1054200.0 2160000.0 ;
      RECT  1052700.0 2153850.0 1051500.0 2155050.0 ;
      RECT  1053000.0 2164200.0 1054200.0 2165400.0 ;
      RECT  1050600.0 2151600.0 1051800.0 2152800.0 ;
      RECT  1053000.0 2151600.0 1054200.0 2152800.0 ;
      RECT  1050600.0 2158800.0 1051800.0 2160000.0 ;
      RECT  1055400.0 2158800.0 1056600.0 2160000.0 ;
      RECT  1047600.0 2154000.0 1057800.0 2154900.0 ;
      RECT  1047600.0 2165100.0 1057800.0 2166000.0 ;
      RECT  1063200.0 2158800.0 1064400.0 2166000.0 ;
      RECT  1060800.0 2151600.0 1062000.0 2152800.0 ;
      RECT  1063200.0 2151600.0 1064400.0 2152800.0 ;
      RECT  1063200.0 2151600.0 1064400.0 2152800.0 ;
      RECT  1060800.0 2151600.0 1062000.0 2152800.0 ;
      RECT  1060800.0 2158800.0 1062000.0 2160000.0 ;
      RECT  1063200.0 2158800.0 1064400.0 2160000.0 ;
      RECT  1063200.0 2158800.0 1064400.0 2160000.0 ;
      RECT  1060800.0 2158800.0 1062000.0 2160000.0 ;
      RECT  1063200.0 2158800.0 1064400.0 2160000.0 ;
      RECT  1065600.0 2158800.0 1066800.0 2160000.0 ;
      RECT  1065600.0 2158800.0 1066800.0 2160000.0 ;
      RECT  1063200.0 2158800.0 1064400.0 2160000.0 ;
      RECT  1062900.0 2153850.0 1061700.0 2155050.0 ;
      RECT  1063200.0 2164200.0 1064400.0 2165400.0 ;
      RECT  1060800.0 2151600.0 1062000.0 2152800.0 ;
      RECT  1063200.0 2151600.0 1064400.0 2152800.0 ;
      RECT  1060800.0 2158800.0 1062000.0 2160000.0 ;
      RECT  1065600.0 2158800.0 1066800.0 2160000.0 ;
      RECT  1057800.0 2154000.0 1068000.0 2154900.0 ;
      RECT  1057800.0 2165100.0 1068000.0 2166000.0 ;
      RECT  1073400.0 2158800.0 1074600.0 2166000.0 ;
      RECT  1071000.0 2151600.0 1072200.0 2152800.0 ;
      RECT  1073400.0 2151600.0 1074600.0 2152800.0 ;
      RECT  1073400.0 2151600.0 1074600.0 2152800.0 ;
      RECT  1071000.0 2151600.0 1072200.0 2152800.0 ;
      RECT  1071000.0 2158800.0 1072200.0 2160000.0 ;
      RECT  1073400.0 2158800.0 1074600.0 2160000.0 ;
      RECT  1073400.0 2158800.0 1074600.0 2160000.0 ;
      RECT  1071000.0 2158800.0 1072200.0 2160000.0 ;
      RECT  1073400.0 2158800.0 1074600.0 2160000.0 ;
      RECT  1075800.0 2158800.0 1077000.0 2160000.0 ;
      RECT  1075800.0 2158800.0 1077000.0 2160000.0 ;
      RECT  1073400.0 2158800.0 1074600.0 2160000.0 ;
      RECT  1073100.0 2153850.0 1071900.0 2155050.0 ;
      RECT  1073400.0 2164200.0 1074600.0 2165400.0 ;
      RECT  1071000.0 2151600.0 1072200.0 2152800.0 ;
      RECT  1073400.0 2151600.0 1074600.0 2152800.0 ;
      RECT  1071000.0 2158800.0 1072200.0 2160000.0 ;
      RECT  1075800.0 2158800.0 1077000.0 2160000.0 ;
      RECT  1068000.0 2154000.0 1078200.0 2154900.0 ;
      RECT  1068000.0 2165100.0 1078200.0 2166000.0 ;
      RECT  1083600.0 2158800.0 1084800.0 2166000.0 ;
      RECT  1081200.0 2151600.0 1082400.0 2152800.0 ;
      RECT  1083600.0 2151600.0 1084800.0 2152800.0 ;
      RECT  1083600.0 2151600.0 1084800.0 2152800.0 ;
      RECT  1081200.0 2151600.0 1082400.0 2152800.0 ;
      RECT  1081200.0 2158800.0 1082400.0 2160000.0 ;
      RECT  1083600.0 2158800.0 1084800.0 2160000.0 ;
      RECT  1083600.0 2158800.0 1084800.0 2160000.0 ;
      RECT  1081200.0 2158800.0 1082400.0 2160000.0 ;
      RECT  1083600.0 2158800.0 1084800.0 2160000.0 ;
      RECT  1086000.0 2158800.0 1087200.0 2160000.0 ;
      RECT  1086000.0 2158800.0 1087200.0 2160000.0 ;
      RECT  1083600.0 2158800.0 1084800.0 2160000.0 ;
      RECT  1083300.0 2153850.0 1082100.0 2155050.0 ;
      RECT  1083600.0 2164200.0 1084800.0 2165400.0 ;
      RECT  1081200.0 2151600.0 1082400.0 2152800.0 ;
      RECT  1083600.0 2151600.0 1084800.0 2152800.0 ;
      RECT  1081200.0 2158800.0 1082400.0 2160000.0 ;
      RECT  1086000.0 2158800.0 1087200.0 2160000.0 ;
      RECT  1078200.0 2154000.0 1088400.0 2154900.0 ;
      RECT  1078200.0 2165100.0 1088400.0 2166000.0 ;
      RECT  1093800.0 2158800.0 1095000.0 2166000.0 ;
      RECT  1091400.0 2151600.0 1092600.0 2152800.0 ;
      RECT  1093800.0 2151600.0 1095000.0 2152800.0 ;
      RECT  1093800.0 2151600.0 1095000.0 2152800.0 ;
      RECT  1091400.0 2151600.0 1092600.0 2152800.0 ;
      RECT  1091400.0 2158800.0 1092600.0 2160000.0 ;
      RECT  1093800.0 2158800.0 1095000.0 2160000.0 ;
      RECT  1093800.0 2158800.0 1095000.0 2160000.0 ;
      RECT  1091400.0 2158800.0 1092600.0 2160000.0 ;
      RECT  1093800.0 2158800.0 1095000.0 2160000.0 ;
      RECT  1096200.0 2158800.0 1097400.0 2160000.0 ;
      RECT  1096200.0 2158800.0 1097400.0 2160000.0 ;
      RECT  1093800.0 2158800.0 1095000.0 2160000.0 ;
      RECT  1093500.0 2153850.0 1092300.0 2155050.0 ;
      RECT  1093800.0 2164200.0 1095000.0 2165400.0 ;
      RECT  1091400.0 2151600.0 1092600.0 2152800.0 ;
      RECT  1093800.0 2151600.0 1095000.0 2152800.0 ;
      RECT  1091400.0 2158800.0 1092600.0 2160000.0 ;
      RECT  1096200.0 2158800.0 1097400.0 2160000.0 ;
      RECT  1088400.0 2154000.0 1098600.0 2154900.0 ;
      RECT  1088400.0 2165100.0 1098600.0 2166000.0 ;
      RECT  1104000.0 2158800.0 1105200.0 2166000.0 ;
      RECT  1101600.0 2151600.0 1102800.0 2152800.0 ;
      RECT  1104000.0 2151600.0 1105200.0 2152800.0 ;
      RECT  1104000.0 2151600.0 1105200.0 2152800.0 ;
      RECT  1101600.0 2151600.0 1102800.0 2152800.0 ;
      RECT  1101600.0 2158800.0 1102800.0 2160000.0 ;
      RECT  1104000.0 2158800.0 1105200.0 2160000.0 ;
      RECT  1104000.0 2158800.0 1105200.0 2160000.0 ;
      RECT  1101600.0 2158800.0 1102800.0 2160000.0 ;
      RECT  1104000.0 2158800.0 1105200.0 2160000.0 ;
      RECT  1106400.0 2158800.0 1107600.0 2160000.0 ;
      RECT  1106400.0 2158800.0 1107600.0 2160000.0 ;
      RECT  1104000.0 2158800.0 1105200.0 2160000.0 ;
      RECT  1103700.0 2153850.0 1102500.0 2155050.0 ;
      RECT  1104000.0 2164200.0 1105200.0 2165400.0 ;
      RECT  1101600.0 2151600.0 1102800.0 2152800.0 ;
      RECT  1104000.0 2151600.0 1105200.0 2152800.0 ;
      RECT  1101600.0 2158800.0 1102800.0 2160000.0 ;
      RECT  1106400.0 2158800.0 1107600.0 2160000.0 ;
      RECT  1098600.0 2154000.0 1108800.0 2154900.0 ;
      RECT  1098600.0 2165100.0 1108800.0 2166000.0 ;
      RECT  1114200.0 2158800.0 1115400.0 2166000.0 ;
      RECT  1111800.0 2151600.0 1113000.0 2152800.0 ;
      RECT  1114200.0 2151600.0 1115400.0 2152800.0 ;
      RECT  1114200.0 2151600.0 1115400.0 2152800.0 ;
      RECT  1111800.0 2151600.0 1113000.0 2152800.0 ;
      RECT  1111800.0 2158800.0 1113000.0 2160000.0 ;
      RECT  1114200.0 2158800.0 1115400.0 2160000.0 ;
      RECT  1114200.0 2158800.0 1115400.0 2160000.0 ;
      RECT  1111800.0 2158800.0 1113000.0 2160000.0 ;
      RECT  1114200.0 2158800.0 1115400.0 2160000.0 ;
      RECT  1116600.0 2158800.0 1117800.0 2160000.0 ;
      RECT  1116600.0 2158800.0 1117800.0 2160000.0 ;
      RECT  1114200.0 2158800.0 1115400.0 2160000.0 ;
      RECT  1113900.0 2153850.0 1112700.0 2155050.0 ;
      RECT  1114200.0 2164200.0 1115400.0 2165400.0 ;
      RECT  1111800.0 2151600.0 1113000.0 2152800.0 ;
      RECT  1114200.0 2151600.0 1115400.0 2152800.0 ;
      RECT  1111800.0 2158800.0 1113000.0 2160000.0 ;
      RECT  1116600.0 2158800.0 1117800.0 2160000.0 ;
      RECT  1108800.0 2154000.0 1119000.0 2154900.0 ;
      RECT  1108800.0 2165100.0 1119000.0 2166000.0 ;
      RECT  1124400.0 2158800.0 1125600.0 2166000.0 ;
      RECT  1122000.0 2151600.0 1123200.0 2152800.0 ;
      RECT  1124400.0 2151600.0 1125600.0 2152800.0 ;
      RECT  1124400.0 2151600.0 1125600.0 2152800.0 ;
      RECT  1122000.0 2151600.0 1123200.0 2152800.0 ;
      RECT  1122000.0 2158800.0 1123200.0 2160000.0 ;
      RECT  1124400.0 2158800.0 1125600.0 2160000.0 ;
      RECT  1124400.0 2158800.0 1125600.0 2160000.0 ;
      RECT  1122000.0 2158800.0 1123200.0 2160000.0 ;
      RECT  1124400.0 2158800.0 1125600.0 2160000.0 ;
      RECT  1126800.0 2158800.0 1128000.0 2160000.0 ;
      RECT  1126800.0 2158800.0 1128000.0 2160000.0 ;
      RECT  1124400.0 2158800.0 1125600.0 2160000.0 ;
      RECT  1124100.0 2153850.0 1122900.0 2155050.0 ;
      RECT  1124400.0 2164200.0 1125600.0 2165400.0 ;
      RECT  1122000.0 2151600.0 1123200.0 2152800.0 ;
      RECT  1124400.0 2151600.0 1125600.0 2152800.0 ;
      RECT  1122000.0 2158800.0 1123200.0 2160000.0 ;
      RECT  1126800.0 2158800.0 1128000.0 2160000.0 ;
      RECT  1119000.0 2154000.0 1129200.0 2154900.0 ;
      RECT  1119000.0 2165100.0 1129200.0 2166000.0 ;
      RECT  1134600.0 2158800.0 1135800.0 2166000.0 ;
      RECT  1132200.0 2151600.0 1133400.0 2152800.0 ;
      RECT  1134600.0 2151600.0 1135800.0 2152800.0 ;
      RECT  1134600.0 2151600.0 1135800.0 2152800.0 ;
      RECT  1132200.0 2151600.0 1133400.0 2152800.0 ;
      RECT  1132200.0 2158800.0 1133400.0 2160000.0 ;
      RECT  1134600.0 2158800.0 1135800.0 2160000.0 ;
      RECT  1134600.0 2158800.0 1135800.0 2160000.0 ;
      RECT  1132200.0 2158800.0 1133400.0 2160000.0 ;
      RECT  1134600.0 2158800.0 1135800.0 2160000.0 ;
      RECT  1137000.0 2158800.0 1138200.0 2160000.0 ;
      RECT  1137000.0 2158800.0 1138200.0 2160000.0 ;
      RECT  1134600.0 2158800.0 1135800.0 2160000.0 ;
      RECT  1134300.0 2153850.0 1133100.0 2155050.0 ;
      RECT  1134600.0 2164200.0 1135800.0 2165400.0 ;
      RECT  1132200.0 2151600.0 1133400.0 2152800.0 ;
      RECT  1134600.0 2151600.0 1135800.0 2152800.0 ;
      RECT  1132200.0 2158800.0 1133400.0 2160000.0 ;
      RECT  1137000.0 2158800.0 1138200.0 2160000.0 ;
      RECT  1129200.0 2154000.0 1139400.0 2154900.0 ;
      RECT  1129200.0 2165100.0 1139400.0 2166000.0 ;
      RECT  1144800.0 2158800.0 1146000.0 2166000.0 ;
      RECT  1142400.0 2151600.0 1143600.0 2152800.0 ;
      RECT  1144800.0 2151600.0 1146000.0 2152800.0 ;
      RECT  1144800.0 2151600.0 1146000.0 2152800.0 ;
      RECT  1142400.0 2151600.0 1143600.0 2152800.0 ;
      RECT  1142400.0 2158800.0 1143600.0 2160000.0 ;
      RECT  1144800.0 2158800.0 1146000.0 2160000.0 ;
      RECT  1144800.0 2158800.0 1146000.0 2160000.0 ;
      RECT  1142400.0 2158800.0 1143600.0 2160000.0 ;
      RECT  1144800.0 2158800.0 1146000.0 2160000.0 ;
      RECT  1147200.0 2158800.0 1148400.0 2160000.0 ;
      RECT  1147200.0 2158800.0 1148400.0 2160000.0 ;
      RECT  1144800.0 2158800.0 1146000.0 2160000.0 ;
      RECT  1144500.0 2153850.0 1143300.0 2155050.0 ;
      RECT  1144800.0 2164200.0 1146000.0 2165400.0 ;
      RECT  1142400.0 2151600.0 1143600.0 2152800.0 ;
      RECT  1144800.0 2151600.0 1146000.0 2152800.0 ;
      RECT  1142400.0 2158800.0 1143600.0 2160000.0 ;
      RECT  1147200.0 2158800.0 1148400.0 2160000.0 ;
      RECT  1139400.0 2154000.0 1149600.0 2154900.0 ;
      RECT  1139400.0 2165100.0 1149600.0 2166000.0 ;
      RECT  1155000.0 2158800.0 1156200.0 2166000.0 ;
      RECT  1152600.0 2151600.0 1153800.0 2152800.0 ;
      RECT  1155000.0 2151600.0 1156200.0 2152800.0 ;
      RECT  1155000.0 2151600.0 1156200.0 2152800.0 ;
      RECT  1152600.0 2151600.0 1153800.0 2152800.0 ;
      RECT  1152600.0 2158800.0 1153800.0 2160000.0 ;
      RECT  1155000.0 2158800.0 1156200.0 2160000.0 ;
      RECT  1155000.0 2158800.0 1156200.0 2160000.0 ;
      RECT  1152600.0 2158800.0 1153800.0 2160000.0 ;
      RECT  1155000.0 2158800.0 1156200.0 2160000.0 ;
      RECT  1157400.0 2158800.0 1158600.0 2160000.0 ;
      RECT  1157400.0 2158800.0 1158600.0 2160000.0 ;
      RECT  1155000.0 2158800.0 1156200.0 2160000.0 ;
      RECT  1154700.0 2153850.0 1153500.0 2155050.0 ;
      RECT  1155000.0 2164200.0 1156200.0 2165400.0 ;
      RECT  1152600.0 2151600.0 1153800.0 2152800.0 ;
      RECT  1155000.0 2151600.0 1156200.0 2152800.0 ;
      RECT  1152600.0 2158800.0 1153800.0 2160000.0 ;
      RECT  1157400.0 2158800.0 1158600.0 2160000.0 ;
      RECT  1149600.0 2154000.0 1159800.0 2154900.0 ;
      RECT  1149600.0 2165100.0 1159800.0 2166000.0 ;
      RECT  1165200.0 2158800.0 1166400.0 2166000.0 ;
      RECT  1162800.0 2151600.0 1164000.0 2152800.0 ;
      RECT  1165200.0 2151600.0 1166400.0 2152800.0 ;
      RECT  1165200.0 2151600.0 1166400.0 2152800.0 ;
      RECT  1162800.0 2151600.0 1164000.0 2152800.0 ;
      RECT  1162800.0 2158800.0 1164000.0 2160000.0 ;
      RECT  1165200.0 2158800.0 1166400.0 2160000.0 ;
      RECT  1165200.0 2158800.0 1166400.0 2160000.0 ;
      RECT  1162800.0 2158800.0 1164000.0 2160000.0 ;
      RECT  1165200.0 2158800.0 1166400.0 2160000.0 ;
      RECT  1167600.0 2158800.0 1168800.0 2160000.0 ;
      RECT  1167600.0 2158800.0 1168800.0 2160000.0 ;
      RECT  1165200.0 2158800.0 1166400.0 2160000.0 ;
      RECT  1164900.0 2153850.0 1163700.0 2155050.0 ;
      RECT  1165200.0 2164200.0 1166400.0 2165400.0 ;
      RECT  1162800.0 2151600.0 1164000.0 2152800.0 ;
      RECT  1165200.0 2151600.0 1166400.0 2152800.0 ;
      RECT  1162800.0 2158800.0 1164000.0 2160000.0 ;
      RECT  1167600.0 2158800.0 1168800.0 2160000.0 ;
      RECT  1159800.0 2154000.0 1170000.0 2154900.0 ;
      RECT  1159800.0 2165100.0 1170000.0 2166000.0 ;
      RECT  1175400.0 2158800.0 1176600.0 2166000.0 ;
      RECT  1173000.0 2151600.0 1174200.0 2152800.0 ;
      RECT  1175400.0 2151600.0 1176600.0 2152800.0 ;
      RECT  1175400.0 2151600.0 1176600.0 2152800.0 ;
      RECT  1173000.0 2151600.0 1174200.0 2152800.0 ;
      RECT  1173000.0 2158800.0 1174200.0 2160000.0 ;
      RECT  1175400.0 2158800.0 1176600.0 2160000.0 ;
      RECT  1175400.0 2158800.0 1176600.0 2160000.0 ;
      RECT  1173000.0 2158800.0 1174200.0 2160000.0 ;
      RECT  1175400.0 2158800.0 1176600.0 2160000.0 ;
      RECT  1177800.0 2158800.0 1179000.0 2160000.0 ;
      RECT  1177800.0 2158800.0 1179000.0 2160000.0 ;
      RECT  1175400.0 2158800.0 1176600.0 2160000.0 ;
      RECT  1175100.0 2153850.0 1173900.0 2155050.0 ;
      RECT  1175400.0 2164200.0 1176600.0 2165400.0 ;
      RECT  1173000.0 2151600.0 1174200.0 2152800.0 ;
      RECT  1175400.0 2151600.0 1176600.0 2152800.0 ;
      RECT  1173000.0 2158800.0 1174200.0 2160000.0 ;
      RECT  1177800.0 2158800.0 1179000.0 2160000.0 ;
      RECT  1170000.0 2154000.0 1180200.0 2154900.0 ;
      RECT  1170000.0 2165100.0 1180200.0 2166000.0 ;
      RECT  1185600.0 2158800.0 1186800.0 2166000.0 ;
      RECT  1183200.0 2151600.0 1184400.0 2152800.0 ;
      RECT  1185600.0 2151600.0 1186800.0 2152800.0 ;
      RECT  1185600.0 2151600.0 1186800.0 2152800.0 ;
      RECT  1183200.0 2151600.0 1184400.0 2152800.0 ;
      RECT  1183200.0 2158800.0 1184400.0 2160000.0 ;
      RECT  1185600.0 2158800.0 1186800.0 2160000.0 ;
      RECT  1185600.0 2158800.0 1186800.0 2160000.0 ;
      RECT  1183200.0 2158800.0 1184400.0 2160000.0 ;
      RECT  1185600.0 2158800.0 1186800.0 2160000.0 ;
      RECT  1188000.0 2158800.0 1189200.0 2160000.0 ;
      RECT  1188000.0 2158800.0 1189200.0 2160000.0 ;
      RECT  1185600.0 2158800.0 1186800.0 2160000.0 ;
      RECT  1185300.0 2153850.0 1184100.0 2155050.0 ;
      RECT  1185600.0 2164200.0 1186800.0 2165400.0 ;
      RECT  1183200.0 2151600.0 1184400.0 2152800.0 ;
      RECT  1185600.0 2151600.0 1186800.0 2152800.0 ;
      RECT  1183200.0 2158800.0 1184400.0 2160000.0 ;
      RECT  1188000.0 2158800.0 1189200.0 2160000.0 ;
      RECT  1180200.0 2154000.0 1190400.0 2154900.0 ;
      RECT  1180200.0 2165100.0 1190400.0 2166000.0 ;
      RECT  1195800.0 2158800.0 1197000.0 2166000.0 ;
      RECT  1193400.0 2151600.0 1194600.0 2152800.0 ;
      RECT  1195800.0 2151600.0 1197000.0 2152800.0 ;
      RECT  1195800.0 2151600.0 1197000.0 2152800.0 ;
      RECT  1193400.0 2151600.0 1194600.0 2152800.0 ;
      RECT  1193400.0 2158800.0 1194600.0 2160000.0 ;
      RECT  1195800.0 2158800.0 1197000.0 2160000.0 ;
      RECT  1195800.0 2158800.0 1197000.0 2160000.0 ;
      RECT  1193400.0 2158800.0 1194600.0 2160000.0 ;
      RECT  1195800.0 2158800.0 1197000.0 2160000.0 ;
      RECT  1198200.0 2158800.0 1199400.0 2160000.0 ;
      RECT  1198200.0 2158800.0 1199400.0 2160000.0 ;
      RECT  1195800.0 2158800.0 1197000.0 2160000.0 ;
      RECT  1195500.0 2153850.0 1194300.0 2155050.0 ;
      RECT  1195800.0 2164200.0 1197000.0 2165400.0 ;
      RECT  1193400.0 2151600.0 1194600.0 2152800.0 ;
      RECT  1195800.0 2151600.0 1197000.0 2152800.0 ;
      RECT  1193400.0 2158800.0 1194600.0 2160000.0 ;
      RECT  1198200.0 2158800.0 1199400.0 2160000.0 ;
      RECT  1190400.0 2154000.0 1200600.0 2154900.0 ;
      RECT  1190400.0 2165100.0 1200600.0 2166000.0 ;
      RECT  1206000.0 2158800.0 1207200.0 2166000.0 ;
      RECT  1203600.0 2151600.0 1204800.0 2152800.0 ;
      RECT  1206000.0 2151600.0 1207200.0 2152800.0 ;
      RECT  1206000.0 2151600.0 1207200.0 2152800.0 ;
      RECT  1203600.0 2151600.0 1204800.0 2152800.0 ;
      RECT  1203600.0 2158800.0 1204800.0 2160000.0 ;
      RECT  1206000.0 2158800.0 1207200.0 2160000.0 ;
      RECT  1206000.0 2158800.0 1207200.0 2160000.0 ;
      RECT  1203600.0 2158800.0 1204800.0 2160000.0 ;
      RECT  1206000.0 2158800.0 1207200.0 2160000.0 ;
      RECT  1208400.0 2158800.0 1209600.0 2160000.0 ;
      RECT  1208400.0 2158800.0 1209600.0 2160000.0 ;
      RECT  1206000.0 2158800.0 1207200.0 2160000.0 ;
      RECT  1205700.0 2153850.0 1204500.0 2155050.0 ;
      RECT  1206000.0 2164200.0 1207200.0 2165400.0 ;
      RECT  1203600.0 2151600.0 1204800.0 2152800.0 ;
      RECT  1206000.0 2151600.0 1207200.0 2152800.0 ;
      RECT  1203600.0 2158800.0 1204800.0 2160000.0 ;
      RECT  1208400.0 2158800.0 1209600.0 2160000.0 ;
      RECT  1200600.0 2154000.0 1210800.0 2154900.0 ;
      RECT  1200600.0 2165100.0 1210800.0 2166000.0 ;
      RECT  1216200.0 2158800.0 1217400.0 2166000.0 ;
      RECT  1213800.0 2151600.0 1215000.0 2152800.0 ;
      RECT  1216200.0 2151600.0 1217400.0 2152800.0 ;
      RECT  1216200.0 2151600.0 1217400.0 2152800.0 ;
      RECT  1213800.0 2151600.0 1215000.0 2152800.0 ;
      RECT  1213800.0 2158800.0 1215000.0 2160000.0 ;
      RECT  1216200.0 2158800.0 1217400.0 2160000.0 ;
      RECT  1216200.0 2158800.0 1217400.0 2160000.0 ;
      RECT  1213800.0 2158800.0 1215000.0 2160000.0 ;
      RECT  1216200.0 2158800.0 1217400.0 2160000.0 ;
      RECT  1218600.0 2158800.0 1219800.0 2160000.0 ;
      RECT  1218600.0 2158800.0 1219800.0 2160000.0 ;
      RECT  1216200.0 2158800.0 1217400.0 2160000.0 ;
      RECT  1215900.0 2153850.0 1214700.0 2155050.0 ;
      RECT  1216200.0 2164200.0 1217400.0 2165400.0 ;
      RECT  1213800.0 2151600.0 1215000.0 2152800.0 ;
      RECT  1216200.0 2151600.0 1217400.0 2152800.0 ;
      RECT  1213800.0 2158800.0 1215000.0 2160000.0 ;
      RECT  1218600.0 2158800.0 1219800.0 2160000.0 ;
      RECT  1210800.0 2154000.0 1221000.0 2154900.0 ;
      RECT  1210800.0 2165100.0 1221000.0 2166000.0 ;
      RECT  1226400.0 2158800.0 1227600.0 2166000.0 ;
      RECT  1224000.0 2151600.0 1225200.0 2152800.0 ;
      RECT  1226400.0 2151600.0 1227600.0 2152800.0 ;
      RECT  1226400.0 2151600.0 1227600.0 2152800.0 ;
      RECT  1224000.0 2151600.0 1225200.0 2152800.0 ;
      RECT  1224000.0 2158800.0 1225200.0 2160000.0 ;
      RECT  1226400.0 2158800.0 1227600.0 2160000.0 ;
      RECT  1226400.0 2158800.0 1227600.0 2160000.0 ;
      RECT  1224000.0 2158800.0 1225200.0 2160000.0 ;
      RECT  1226400.0 2158800.0 1227600.0 2160000.0 ;
      RECT  1228800.0 2158800.0 1230000.0 2160000.0 ;
      RECT  1228800.0 2158800.0 1230000.0 2160000.0 ;
      RECT  1226400.0 2158800.0 1227600.0 2160000.0 ;
      RECT  1226100.0 2153850.0 1224900.0 2155050.0 ;
      RECT  1226400.0 2164200.0 1227600.0 2165400.0 ;
      RECT  1224000.0 2151600.0 1225200.0 2152800.0 ;
      RECT  1226400.0 2151600.0 1227600.0 2152800.0 ;
      RECT  1224000.0 2158800.0 1225200.0 2160000.0 ;
      RECT  1228800.0 2158800.0 1230000.0 2160000.0 ;
      RECT  1221000.0 2154000.0 1231200.0 2154900.0 ;
      RECT  1221000.0 2165100.0 1231200.0 2166000.0 ;
      RECT  1236600.0 2158800.0 1237800.0 2166000.0 ;
      RECT  1234200.0 2151600.0 1235400.0 2152800.0 ;
      RECT  1236600.0 2151600.0 1237800.0 2152800.0 ;
      RECT  1236600.0 2151600.0 1237800.0 2152800.0 ;
      RECT  1234200.0 2151600.0 1235400.0 2152800.0 ;
      RECT  1234200.0 2158800.0 1235400.0 2160000.0 ;
      RECT  1236600.0 2158800.0 1237800.0 2160000.0 ;
      RECT  1236600.0 2158800.0 1237800.0 2160000.0 ;
      RECT  1234200.0 2158800.0 1235400.0 2160000.0 ;
      RECT  1236600.0 2158800.0 1237800.0 2160000.0 ;
      RECT  1239000.0 2158800.0 1240200.0 2160000.0 ;
      RECT  1239000.0 2158800.0 1240200.0 2160000.0 ;
      RECT  1236600.0 2158800.0 1237800.0 2160000.0 ;
      RECT  1236300.0 2153850.0 1235100.0 2155050.0 ;
      RECT  1236600.0 2164200.0 1237800.0 2165400.0 ;
      RECT  1234200.0 2151600.0 1235400.0 2152800.0 ;
      RECT  1236600.0 2151600.0 1237800.0 2152800.0 ;
      RECT  1234200.0 2158800.0 1235400.0 2160000.0 ;
      RECT  1239000.0 2158800.0 1240200.0 2160000.0 ;
      RECT  1231200.0 2154000.0 1241400.0 2154900.0 ;
      RECT  1231200.0 2165100.0 1241400.0 2166000.0 ;
      RECT  1246800.0 2158800.0 1248000.0 2166000.0 ;
      RECT  1244400.0 2151600.0 1245600.0 2152800.0 ;
      RECT  1246800.0 2151600.0 1248000.0 2152800.0 ;
      RECT  1246800.0 2151600.0 1248000.0 2152800.0 ;
      RECT  1244400.0 2151600.0 1245600.0 2152800.0 ;
      RECT  1244400.0 2158800.0 1245600.0 2160000.0 ;
      RECT  1246800.0 2158800.0 1248000.0 2160000.0 ;
      RECT  1246800.0 2158800.0 1248000.0 2160000.0 ;
      RECT  1244400.0 2158800.0 1245600.0 2160000.0 ;
      RECT  1246800.0 2158800.0 1248000.0 2160000.0 ;
      RECT  1249200.0 2158800.0 1250400.0 2160000.0 ;
      RECT  1249200.0 2158800.0 1250400.0 2160000.0 ;
      RECT  1246800.0 2158800.0 1248000.0 2160000.0 ;
      RECT  1246500.0 2153850.0 1245300.0 2155050.0 ;
      RECT  1246800.0 2164200.0 1248000.0 2165400.0 ;
      RECT  1244400.0 2151600.0 1245600.0 2152800.0 ;
      RECT  1246800.0 2151600.0 1248000.0 2152800.0 ;
      RECT  1244400.0 2158800.0 1245600.0 2160000.0 ;
      RECT  1249200.0 2158800.0 1250400.0 2160000.0 ;
      RECT  1241400.0 2154000.0 1251600.0 2154900.0 ;
      RECT  1241400.0 2165100.0 1251600.0 2166000.0 ;
      RECT  1257000.0 2158800.0 1258200.0 2166000.0 ;
      RECT  1254600.0 2151600.0 1255800.0 2152800.0 ;
      RECT  1257000.0 2151600.0 1258200.0 2152800.0 ;
      RECT  1257000.0 2151600.0 1258200.0 2152800.0 ;
      RECT  1254600.0 2151600.0 1255800.0 2152800.0 ;
      RECT  1254600.0 2158800.0 1255800.0 2160000.0 ;
      RECT  1257000.0 2158800.0 1258200.0 2160000.0 ;
      RECT  1257000.0 2158800.0 1258200.0 2160000.0 ;
      RECT  1254600.0 2158800.0 1255800.0 2160000.0 ;
      RECT  1257000.0 2158800.0 1258200.0 2160000.0 ;
      RECT  1259400.0 2158800.0 1260600.0 2160000.0 ;
      RECT  1259400.0 2158800.0 1260600.0 2160000.0 ;
      RECT  1257000.0 2158800.0 1258200.0 2160000.0 ;
      RECT  1256700.0 2153850.0 1255500.0 2155050.0 ;
      RECT  1257000.0 2164200.0 1258200.0 2165400.0 ;
      RECT  1254600.0 2151600.0 1255800.0 2152800.0 ;
      RECT  1257000.0 2151600.0 1258200.0 2152800.0 ;
      RECT  1254600.0 2158800.0 1255800.0 2160000.0 ;
      RECT  1259400.0 2158800.0 1260600.0 2160000.0 ;
      RECT  1251600.0 2154000.0 1261800.0 2154900.0 ;
      RECT  1251600.0 2165100.0 1261800.0 2166000.0 ;
      RECT  1267200.0 2158800.0 1268400.0 2166000.0 ;
      RECT  1264800.0 2151600.0 1266000.0 2152800.0 ;
      RECT  1267200.0 2151600.0 1268400.0 2152800.0 ;
      RECT  1267200.0 2151600.0 1268400.0 2152800.0 ;
      RECT  1264800.0 2151600.0 1266000.0 2152800.0 ;
      RECT  1264800.0 2158800.0 1266000.0 2160000.0 ;
      RECT  1267200.0 2158800.0 1268400.0 2160000.0 ;
      RECT  1267200.0 2158800.0 1268400.0 2160000.0 ;
      RECT  1264800.0 2158800.0 1266000.0 2160000.0 ;
      RECT  1267200.0 2158800.0 1268400.0 2160000.0 ;
      RECT  1269600.0 2158800.0 1270800.0 2160000.0 ;
      RECT  1269600.0 2158800.0 1270800.0 2160000.0 ;
      RECT  1267200.0 2158800.0 1268400.0 2160000.0 ;
      RECT  1266900.0 2153850.0 1265700.0 2155050.0 ;
      RECT  1267200.0 2164200.0 1268400.0 2165400.0 ;
      RECT  1264800.0 2151600.0 1266000.0 2152800.0 ;
      RECT  1267200.0 2151600.0 1268400.0 2152800.0 ;
      RECT  1264800.0 2158800.0 1266000.0 2160000.0 ;
      RECT  1269600.0 2158800.0 1270800.0 2160000.0 ;
      RECT  1261800.0 2154000.0 1272000.0 2154900.0 ;
      RECT  1261800.0 2165100.0 1272000.0 2166000.0 ;
      RECT  1277400.0 2158800.0 1278600.0 2166000.0 ;
      RECT  1275000.0 2151600.0 1276200.0 2152800.0 ;
      RECT  1277400.0 2151600.0 1278600.0 2152800.0 ;
      RECT  1277400.0 2151600.0 1278600.0 2152800.0 ;
      RECT  1275000.0 2151600.0 1276200.0 2152800.0 ;
      RECT  1275000.0 2158800.0 1276200.0 2160000.0 ;
      RECT  1277400.0 2158800.0 1278600.0 2160000.0 ;
      RECT  1277400.0 2158800.0 1278600.0 2160000.0 ;
      RECT  1275000.0 2158800.0 1276200.0 2160000.0 ;
      RECT  1277400.0 2158800.0 1278600.0 2160000.0 ;
      RECT  1279800.0 2158800.0 1281000.0 2160000.0 ;
      RECT  1279800.0 2158800.0 1281000.0 2160000.0 ;
      RECT  1277400.0 2158800.0 1278600.0 2160000.0 ;
      RECT  1277100.0 2153850.0 1275900.0 2155050.0 ;
      RECT  1277400.0 2164200.0 1278600.0 2165400.0 ;
      RECT  1275000.0 2151600.0 1276200.0 2152800.0 ;
      RECT  1277400.0 2151600.0 1278600.0 2152800.0 ;
      RECT  1275000.0 2158800.0 1276200.0 2160000.0 ;
      RECT  1279800.0 2158800.0 1281000.0 2160000.0 ;
      RECT  1272000.0 2154000.0 1282200.0 2154900.0 ;
      RECT  1272000.0 2165100.0 1282200.0 2166000.0 ;
      RECT  1287600.0 2158800.0 1288800.0 2166000.0 ;
      RECT  1285200.0 2151600.0 1286400.0 2152800.0 ;
      RECT  1287600.0 2151600.0 1288800.0 2152800.0 ;
      RECT  1287600.0 2151600.0 1288800.0 2152800.0 ;
      RECT  1285200.0 2151600.0 1286400.0 2152800.0 ;
      RECT  1285200.0 2158800.0 1286400.0 2160000.0 ;
      RECT  1287600.0 2158800.0 1288800.0 2160000.0 ;
      RECT  1287600.0 2158800.0 1288800.0 2160000.0 ;
      RECT  1285200.0 2158800.0 1286400.0 2160000.0 ;
      RECT  1287600.0 2158800.0 1288800.0 2160000.0 ;
      RECT  1290000.0 2158800.0 1291200.0 2160000.0 ;
      RECT  1290000.0 2158800.0 1291200.0 2160000.0 ;
      RECT  1287600.0 2158800.0 1288800.0 2160000.0 ;
      RECT  1287300.0 2153850.0 1286100.0 2155050.0 ;
      RECT  1287600.0 2164200.0 1288800.0 2165400.0 ;
      RECT  1285200.0 2151600.0 1286400.0 2152800.0 ;
      RECT  1287600.0 2151600.0 1288800.0 2152800.0 ;
      RECT  1285200.0 2158800.0 1286400.0 2160000.0 ;
      RECT  1290000.0 2158800.0 1291200.0 2160000.0 ;
      RECT  1282200.0 2154000.0 1292400.0 2154900.0 ;
      RECT  1282200.0 2165100.0 1292400.0 2166000.0 ;
      RECT  1297800.0 2158800.0 1299000.0 2166000.0 ;
      RECT  1295400.0 2151600.0 1296600.0 2152800.0 ;
      RECT  1297800.0 2151600.0 1299000.0 2152800.0 ;
      RECT  1297800.0 2151600.0 1299000.0 2152800.0 ;
      RECT  1295400.0 2151600.0 1296600.0 2152800.0 ;
      RECT  1295400.0 2158800.0 1296600.0 2160000.0 ;
      RECT  1297800.0 2158800.0 1299000.0 2160000.0 ;
      RECT  1297800.0 2158800.0 1299000.0 2160000.0 ;
      RECT  1295400.0 2158800.0 1296600.0 2160000.0 ;
      RECT  1297800.0 2158800.0 1299000.0 2160000.0 ;
      RECT  1300200.0 2158800.0 1301400.0 2160000.0 ;
      RECT  1300200.0 2158800.0 1301400.0 2160000.0 ;
      RECT  1297800.0 2158800.0 1299000.0 2160000.0 ;
      RECT  1297500.0 2153850.0 1296300.0 2155050.0 ;
      RECT  1297800.0 2164200.0 1299000.0 2165400.0 ;
      RECT  1295400.0 2151600.0 1296600.0 2152800.0 ;
      RECT  1297800.0 2151600.0 1299000.0 2152800.0 ;
      RECT  1295400.0 2158800.0 1296600.0 2160000.0 ;
      RECT  1300200.0 2158800.0 1301400.0 2160000.0 ;
      RECT  1292400.0 2154000.0 1302600.0 2154900.0 ;
      RECT  1292400.0 2165100.0 1302600.0 2166000.0 ;
      RECT  1308000.0 2158800.0 1309200.0 2166000.0 ;
      RECT  1305600.0 2151600.0 1306800.0 2152800.0 ;
      RECT  1308000.0 2151600.0 1309200.0 2152800.0 ;
      RECT  1308000.0 2151600.0 1309200.0 2152800.0 ;
      RECT  1305600.0 2151600.0 1306800.0 2152800.0 ;
      RECT  1305600.0 2158800.0 1306800.0 2160000.0 ;
      RECT  1308000.0 2158800.0 1309200.0 2160000.0 ;
      RECT  1308000.0 2158800.0 1309200.0 2160000.0 ;
      RECT  1305600.0 2158800.0 1306800.0 2160000.0 ;
      RECT  1308000.0 2158800.0 1309200.0 2160000.0 ;
      RECT  1310400.0 2158800.0 1311600.0 2160000.0 ;
      RECT  1310400.0 2158800.0 1311600.0 2160000.0 ;
      RECT  1308000.0 2158800.0 1309200.0 2160000.0 ;
      RECT  1307700.0 2153850.0 1306500.0 2155050.0 ;
      RECT  1308000.0 2164200.0 1309200.0 2165400.0 ;
      RECT  1305600.0 2151600.0 1306800.0 2152800.0 ;
      RECT  1308000.0 2151600.0 1309200.0 2152800.0 ;
      RECT  1305600.0 2158800.0 1306800.0 2160000.0 ;
      RECT  1310400.0 2158800.0 1311600.0 2160000.0 ;
      RECT  1302600.0 2154000.0 1312800.0 2154900.0 ;
      RECT  1302600.0 2165100.0 1312800.0 2166000.0 ;
      RECT  1318200.0 2158800.0 1319400.0 2166000.0 ;
      RECT  1315800.0 2151600.0 1317000.0 2152800.0 ;
      RECT  1318200.0 2151600.0 1319400.0 2152800.0 ;
      RECT  1318200.0 2151600.0 1319400.0 2152800.0 ;
      RECT  1315800.0 2151600.0 1317000.0 2152800.0 ;
      RECT  1315800.0 2158800.0 1317000.0 2160000.0 ;
      RECT  1318200.0 2158800.0 1319400.0 2160000.0 ;
      RECT  1318200.0 2158800.0 1319400.0 2160000.0 ;
      RECT  1315800.0 2158800.0 1317000.0 2160000.0 ;
      RECT  1318200.0 2158800.0 1319400.0 2160000.0 ;
      RECT  1320600.0 2158800.0 1321800.0 2160000.0 ;
      RECT  1320600.0 2158800.0 1321800.0 2160000.0 ;
      RECT  1318200.0 2158800.0 1319400.0 2160000.0 ;
      RECT  1317900.0 2153850.0 1316700.0 2155050.0 ;
      RECT  1318200.0 2164200.0 1319400.0 2165400.0 ;
      RECT  1315800.0 2151600.0 1317000.0 2152800.0 ;
      RECT  1318200.0 2151600.0 1319400.0 2152800.0 ;
      RECT  1315800.0 2158800.0 1317000.0 2160000.0 ;
      RECT  1320600.0 2158800.0 1321800.0 2160000.0 ;
      RECT  1312800.0 2154000.0 1323000.0 2154900.0 ;
      RECT  1312800.0 2165100.0 1323000.0 2166000.0 ;
      RECT  1328400.0 2158800.0 1329600.0 2166000.0 ;
      RECT  1326000.0 2151600.0 1327200.0 2152800.0 ;
      RECT  1328400.0 2151600.0 1329600.0 2152800.0 ;
      RECT  1328400.0 2151600.0 1329600.0 2152800.0 ;
      RECT  1326000.0 2151600.0 1327200.0 2152800.0 ;
      RECT  1326000.0 2158800.0 1327200.0 2160000.0 ;
      RECT  1328400.0 2158800.0 1329600.0 2160000.0 ;
      RECT  1328400.0 2158800.0 1329600.0 2160000.0 ;
      RECT  1326000.0 2158800.0 1327200.0 2160000.0 ;
      RECT  1328400.0 2158800.0 1329600.0 2160000.0 ;
      RECT  1330800.0 2158800.0 1332000.0 2160000.0 ;
      RECT  1330800.0 2158800.0 1332000.0 2160000.0 ;
      RECT  1328400.0 2158800.0 1329600.0 2160000.0 ;
      RECT  1328100.0 2153850.0 1326900.0 2155050.0 ;
      RECT  1328400.0 2164200.0 1329600.0 2165400.0 ;
      RECT  1326000.0 2151600.0 1327200.0 2152800.0 ;
      RECT  1328400.0 2151600.0 1329600.0 2152800.0 ;
      RECT  1326000.0 2158800.0 1327200.0 2160000.0 ;
      RECT  1330800.0 2158800.0 1332000.0 2160000.0 ;
      RECT  1323000.0 2154000.0 1333200.0 2154900.0 ;
      RECT  1323000.0 2165100.0 1333200.0 2166000.0 ;
      RECT  1338600.0 2158800.0 1339800.0 2166000.0 ;
      RECT  1336200.0 2151600.0 1337400.0 2152800.0 ;
      RECT  1338600.0 2151600.0 1339800.0 2152800.0 ;
      RECT  1338600.0 2151600.0 1339800.0 2152800.0 ;
      RECT  1336200.0 2151600.0 1337400.0 2152800.0 ;
      RECT  1336200.0 2158800.0 1337400.0 2160000.0 ;
      RECT  1338600.0 2158800.0 1339800.0 2160000.0 ;
      RECT  1338600.0 2158800.0 1339800.0 2160000.0 ;
      RECT  1336200.0 2158800.0 1337400.0 2160000.0 ;
      RECT  1338600.0 2158800.0 1339800.0 2160000.0 ;
      RECT  1341000.0 2158800.0 1342200.0 2160000.0 ;
      RECT  1341000.0 2158800.0 1342200.0 2160000.0 ;
      RECT  1338600.0 2158800.0 1339800.0 2160000.0 ;
      RECT  1338300.0 2153850.0 1337100.0 2155050.0 ;
      RECT  1338600.0 2164200.0 1339800.0 2165400.0 ;
      RECT  1336200.0 2151600.0 1337400.0 2152800.0 ;
      RECT  1338600.0 2151600.0 1339800.0 2152800.0 ;
      RECT  1336200.0 2158800.0 1337400.0 2160000.0 ;
      RECT  1341000.0 2158800.0 1342200.0 2160000.0 ;
      RECT  1333200.0 2154000.0 1343400.0 2154900.0 ;
      RECT  1333200.0 2165100.0 1343400.0 2166000.0 ;
      RECT  1348800.0 2158800.0 1350000.0 2166000.0 ;
      RECT  1346400.0 2151600.0 1347600.0 2152800.0 ;
      RECT  1348800.0 2151600.0 1350000.0 2152800.0 ;
      RECT  1348800.0 2151600.0 1350000.0 2152800.0 ;
      RECT  1346400.0 2151600.0 1347600.0 2152800.0 ;
      RECT  1346400.0 2158800.0 1347600.0 2160000.0 ;
      RECT  1348800.0 2158800.0 1350000.0 2160000.0 ;
      RECT  1348800.0 2158800.0 1350000.0 2160000.0 ;
      RECT  1346400.0 2158800.0 1347600.0 2160000.0 ;
      RECT  1348800.0 2158800.0 1350000.0 2160000.0 ;
      RECT  1351200.0 2158800.0 1352400.0 2160000.0 ;
      RECT  1351200.0 2158800.0 1352400.0 2160000.0 ;
      RECT  1348800.0 2158800.0 1350000.0 2160000.0 ;
      RECT  1348500.0 2153850.0 1347300.0 2155050.0 ;
      RECT  1348800.0 2164200.0 1350000.0 2165400.0 ;
      RECT  1346400.0 2151600.0 1347600.0 2152800.0 ;
      RECT  1348800.0 2151600.0 1350000.0 2152800.0 ;
      RECT  1346400.0 2158800.0 1347600.0 2160000.0 ;
      RECT  1351200.0 2158800.0 1352400.0 2160000.0 ;
      RECT  1343400.0 2154000.0 1353600.0 2154900.0 ;
      RECT  1343400.0 2165100.0 1353600.0 2166000.0 ;
      RECT  1359000.0 2158800.0 1360200.0 2166000.0 ;
      RECT  1356600.0 2151600.0 1357800.0 2152800.0 ;
      RECT  1359000.0 2151600.0 1360200.0 2152800.0 ;
      RECT  1359000.0 2151600.0 1360200.0 2152800.0 ;
      RECT  1356600.0 2151600.0 1357800.0 2152800.0 ;
      RECT  1356600.0 2158800.0 1357800.0 2160000.0 ;
      RECT  1359000.0 2158800.0 1360200.0 2160000.0 ;
      RECT  1359000.0 2158800.0 1360200.0 2160000.0 ;
      RECT  1356600.0 2158800.0 1357800.0 2160000.0 ;
      RECT  1359000.0 2158800.0 1360200.0 2160000.0 ;
      RECT  1361400.0 2158800.0 1362600.0 2160000.0 ;
      RECT  1361400.0 2158800.0 1362600.0 2160000.0 ;
      RECT  1359000.0 2158800.0 1360200.0 2160000.0 ;
      RECT  1358700.0 2153850.0 1357500.0 2155050.0 ;
      RECT  1359000.0 2164200.0 1360200.0 2165400.0 ;
      RECT  1356600.0 2151600.0 1357800.0 2152800.0 ;
      RECT  1359000.0 2151600.0 1360200.0 2152800.0 ;
      RECT  1356600.0 2158800.0 1357800.0 2160000.0 ;
      RECT  1361400.0 2158800.0 1362600.0 2160000.0 ;
      RECT  1353600.0 2154000.0 1363800.0 2154900.0 ;
      RECT  1353600.0 2165100.0 1363800.0 2166000.0 ;
      RECT  1369200.0 2158800.0 1370400.0 2166000.0 ;
      RECT  1366800.0 2151600.0 1368000.0 2152800.0 ;
      RECT  1369200.0 2151600.0 1370400.0 2152800.0 ;
      RECT  1369200.0 2151600.0 1370400.0 2152800.0 ;
      RECT  1366800.0 2151600.0 1368000.0 2152800.0 ;
      RECT  1366800.0 2158800.0 1368000.0 2160000.0 ;
      RECT  1369200.0 2158800.0 1370400.0 2160000.0 ;
      RECT  1369200.0 2158800.0 1370400.0 2160000.0 ;
      RECT  1366800.0 2158800.0 1368000.0 2160000.0 ;
      RECT  1369200.0 2158800.0 1370400.0 2160000.0 ;
      RECT  1371600.0 2158800.0 1372800.0 2160000.0 ;
      RECT  1371600.0 2158800.0 1372800.0 2160000.0 ;
      RECT  1369200.0 2158800.0 1370400.0 2160000.0 ;
      RECT  1368900.0 2153850.0 1367700.0 2155050.0 ;
      RECT  1369200.0 2164200.0 1370400.0 2165400.0 ;
      RECT  1366800.0 2151600.0 1368000.0 2152800.0 ;
      RECT  1369200.0 2151600.0 1370400.0 2152800.0 ;
      RECT  1366800.0 2158800.0 1368000.0 2160000.0 ;
      RECT  1371600.0 2158800.0 1372800.0 2160000.0 ;
      RECT  1363800.0 2154000.0 1374000.0 2154900.0 ;
      RECT  1363800.0 2165100.0 1374000.0 2166000.0 ;
      RECT  1379400.0 2158800.0 1380600.0 2166000.0 ;
      RECT  1377000.0 2151600.0 1378200.0 2152800.0 ;
      RECT  1379400.0 2151600.0 1380600.0 2152800.0 ;
      RECT  1379400.0 2151600.0 1380600.0 2152800.0 ;
      RECT  1377000.0 2151600.0 1378200.0 2152800.0 ;
      RECT  1377000.0 2158800.0 1378200.0 2160000.0 ;
      RECT  1379400.0 2158800.0 1380600.0 2160000.0 ;
      RECT  1379400.0 2158800.0 1380600.0 2160000.0 ;
      RECT  1377000.0 2158800.0 1378200.0 2160000.0 ;
      RECT  1379400.0 2158800.0 1380600.0 2160000.0 ;
      RECT  1381800.0 2158800.0 1383000.0 2160000.0 ;
      RECT  1381800.0 2158800.0 1383000.0 2160000.0 ;
      RECT  1379400.0 2158800.0 1380600.0 2160000.0 ;
      RECT  1379100.0 2153850.0 1377900.0 2155050.0 ;
      RECT  1379400.0 2164200.0 1380600.0 2165400.0 ;
      RECT  1377000.0 2151600.0 1378200.0 2152800.0 ;
      RECT  1379400.0 2151600.0 1380600.0 2152800.0 ;
      RECT  1377000.0 2158800.0 1378200.0 2160000.0 ;
      RECT  1381800.0 2158800.0 1383000.0 2160000.0 ;
      RECT  1374000.0 2154000.0 1384200.0 2154900.0 ;
      RECT  1374000.0 2165100.0 1384200.0 2166000.0 ;
      RECT  1389600.0 2158800.0 1390800.0 2166000.0 ;
      RECT  1387200.0 2151600.0 1388400.0 2152800.0 ;
      RECT  1389600.0 2151600.0 1390800.0 2152800.0 ;
      RECT  1389600.0 2151600.0 1390800.0 2152800.0 ;
      RECT  1387200.0 2151600.0 1388400.0 2152800.0 ;
      RECT  1387200.0 2158800.0 1388400.0 2160000.0 ;
      RECT  1389600.0 2158800.0 1390800.0 2160000.0 ;
      RECT  1389600.0 2158800.0 1390800.0 2160000.0 ;
      RECT  1387200.0 2158800.0 1388400.0 2160000.0 ;
      RECT  1389600.0 2158800.0 1390800.0 2160000.0 ;
      RECT  1392000.0 2158800.0 1393200.0 2160000.0 ;
      RECT  1392000.0 2158800.0 1393200.0 2160000.0 ;
      RECT  1389600.0 2158800.0 1390800.0 2160000.0 ;
      RECT  1389300.0 2153850.0 1388100.0 2155050.0 ;
      RECT  1389600.0 2164200.0 1390800.0 2165400.0 ;
      RECT  1387200.0 2151600.0 1388400.0 2152800.0 ;
      RECT  1389600.0 2151600.0 1390800.0 2152800.0 ;
      RECT  1387200.0 2158800.0 1388400.0 2160000.0 ;
      RECT  1392000.0 2158800.0 1393200.0 2160000.0 ;
      RECT  1384200.0 2154000.0 1394400.0 2154900.0 ;
      RECT  1384200.0 2165100.0 1394400.0 2166000.0 ;
      RECT  1399800.0 2158800.0 1401000.0 2166000.0 ;
      RECT  1397400.0 2151600.0 1398600.0 2152800.0 ;
      RECT  1399800.0 2151600.0 1401000.0 2152800.0 ;
      RECT  1399800.0 2151600.0 1401000.0 2152800.0 ;
      RECT  1397400.0 2151600.0 1398600.0 2152800.0 ;
      RECT  1397400.0 2158800.0 1398600.0 2160000.0 ;
      RECT  1399800.0 2158800.0 1401000.0 2160000.0 ;
      RECT  1399800.0 2158800.0 1401000.0 2160000.0 ;
      RECT  1397400.0 2158800.0 1398600.0 2160000.0 ;
      RECT  1399800.0 2158800.0 1401000.0 2160000.0 ;
      RECT  1402200.0 2158800.0 1403400.0 2160000.0 ;
      RECT  1402200.0 2158800.0 1403400.0 2160000.0 ;
      RECT  1399800.0 2158800.0 1401000.0 2160000.0 ;
      RECT  1399500.0 2153850.0 1398300.0 2155050.0 ;
      RECT  1399800.0 2164200.0 1401000.0 2165400.0 ;
      RECT  1397400.0 2151600.0 1398600.0 2152800.0 ;
      RECT  1399800.0 2151600.0 1401000.0 2152800.0 ;
      RECT  1397400.0 2158800.0 1398600.0 2160000.0 ;
      RECT  1402200.0 2158800.0 1403400.0 2160000.0 ;
      RECT  1394400.0 2154000.0 1404600.0 2154900.0 ;
      RECT  1394400.0 2165100.0 1404600.0 2166000.0 ;
      RECT  1410000.0 2158800.0 1411200.0 2166000.0 ;
      RECT  1407600.0 2151600.0 1408800.0 2152800.0 ;
      RECT  1410000.0 2151600.0 1411200.0 2152800.0 ;
      RECT  1410000.0 2151600.0 1411200.0 2152800.0 ;
      RECT  1407600.0 2151600.0 1408800.0 2152800.0 ;
      RECT  1407600.0 2158800.0 1408800.0 2160000.0 ;
      RECT  1410000.0 2158800.0 1411200.0 2160000.0 ;
      RECT  1410000.0 2158800.0 1411200.0 2160000.0 ;
      RECT  1407600.0 2158800.0 1408800.0 2160000.0 ;
      RECT  1410000.0 2158800.0 1411200.0 2160000.0 ;
      RECT  1412400.0 2158800.0 1413600.0 2160000.0 ;
      RECT  1412400.0 2158800.0 1413600.0 2160000.0 ;
      RECT  1410000.0 2158800.0 1411200.0 2160000.0 ;
      RECT  1409700.0 2153850.0 1408500.0 2155050.0 ;
      RECT  1410000.0 2164200.0 1411200.0 2165400.0 ;
      RECT  1407600.0 2151600.0 1408800.0 2152800.0 ;
      RECT  1410000.0 2151600.0 1411200.0 2152800.0 ;
      RECT  1407600.0 2158800.0 1408800.0 2160000.0 ;
      RECT  1412400.0 2158800.0 1413600.0 2160000.0 ;
      RECT  1404600.0 2154000.0 1414800.0 2154900.0 ;
      RECT  1404600.0 2165100.0 1414800.0 2166000.0 ;
      RECT  1420200.0 2158800.0 1421400.0 2166000.0 ;
      RECT  1417800.0 2151600.0 1419000.0 2152800.0 ;
      RECT  1420200.0 2151600.0 1421400.0 2152800.0 ;
      RECT  1420200.0 2151600.0 1421400.0 2152800.0 ;
      RECT  1417800.0 2151600.0 1419000.0 2152800.0 ;
      RECT  1417800.0 2158800.0 1419000.0 2160000.0 ;
      RECT  1420200.0 2158800.0 1421400.0 2160000.0 ;
      RECT  1420200.0 2158800.0 1421400.0 2160000.0 ;
      RECT  1417800.0 2158800.0 1419000.0 2160000.0 ;
      RECT  1420200.0 2158800.0 1421400.0 2160000.0 ;
      RECT  1422600.0 2158800.0 1423800.0 2160000.0 ;
      RECT  1422600.0 2158800.0 1423800.0 2160000.0 ;
      RECT  1420200.0 2158800.0 1421400.0 2160000.0 ;
      RECT  1419900.0 2153850.0 1418700.0 2155050.0 ;
      RECT  1420200.0 2164200.0 1421400.0 2165400.0 ;
      RECT  1417800.0 2151600.0 1419000.0 2152800.0 ;
      RECT  1420200.0 2151600.0 1421400.0 2152800.0 ;
      RECT  1417800.0 2158800.0 1419000.0 2160000.0 ;
      RECT  1422600.0 2158800.0 1423800.0 2160000.0 ;
      RECT  1414800.0 2154000.0 1425000.0 2154900.0 ;
      RECT  1414800.0 2165100.0 1425000.0 2166000.0 ;
      RECT  1430400.0 2158800.0 1431600.0 2166000.0 ;
      RECT  1428000.0 2151600.0 1429200.0 2152800.0 ;
      RECT  1430400.0 2151600.0 1431600.0 2152800.0 ;
      RECT  1430400.0 2151600.0 1431600.0 2152800.0 ;
      RECT  1428000.0 2151600.0 1429200.0 2152800.0 ;
      RECT  1428000.0 2158800.0 1429200.0 2160000.0 ;
      RECT  1430400.0 2158800.0 1431600.0 2160000.0 ;
      RECT  1430400.0 2158800.0 1431600.0 2160000.0 ;
      RECT  1428000.0 2158800.0 1429200.0 2160000.0 ;
      RECT  1430400.0 2158800.0 1431600.0 2160000.0 ;
      RECT  1432800.0 2158800.0 1434000.0 2160000.0 ;
      RECT  1432800.0 2158800.0 1434000.0 2160000.0 ;
      RECT  1430400.0 2158800.0 1431600.0 2160000.0 ;
      RECT  1430100.0 2153850.0 1428900.0 2155050.0 ;
      RECT  1430400.0 2164200.0 1431600.0 2165400.0 ;
      RECT  1428000.0 2151600.0 1429200.0 2152800.0 ;
      RECT  1430400.0 2151600.0 1431600.0 2152800.0 ;
      RECT  1428000.0 2158800.0 1429200.0 2160000.0 ;
      RECT  1432800.0 2158800.0 1434000.0 2160000.0 ;
      RECT  1425000.0 2154000.0 1435200.0 2154900.0 ;
      RECT  1425000.0 2165100.0 1435200.0 2166000.0 ;
      RECT  1440600.0 2158800.0 1441800.0 2166000.0 ;
      RECT  1438200.0 2151600.0 1439400.0 2152800.0 ;
      RECT  1440600.0 2151600.0 1441800.0 2152800.0 ;
      RECT  1440600.0 2151600.0 1441800.0 2152800.0 ;
      RECT  1438200.0 2151600.0 1439400.0 2152800.0 ;
      RECT  1438200.0 2158800.0 1439400.0 2160000.0 ;
      RECT  1440600.0 2158800.0 1441800.0 2160000.0 ;
      RECT  1440600.0 2158800.0 1441800.0 2160000.0 ;
      RECT  1438200.0 2158800.0 1439400.0 2160000.0 ;
      RECT  1440600.0 2158800.0 1441800.0 2160000.0 ;
      RECT  1443000.0 2158800.0 1444200.0 2160000.0 ;
      RECT  1443000.0 2158800.0 1444200.0 2160000.0 ;
      RECT  1440600.0 2158800.0 1441800.0 2160000.0 ;
      RECT  1440300.0 2153850.0 1439100.0 2155050.0 ;
      RECT  1440600.0 2164200.0 1441800.0 2165400.0 ;
      RECT  1438200.0 2151600.0 1439400.0 2152800.0 ;
      RECT  1440600.0 2151600.0 1441800.0 2152800.0 ;
      RECT  1438200.0 2158800.0 1439400.0 2160000.0 ;
      RECT  1443000.0 2158800.0 1444200.0 2160000.0 ;
      RECT  1435200.0 2154000.0 1445400.0 2154900.0 ;
      RECT  1435200.0 2165100.0 1445400.0 2166000.0 ;
      RECT  1450800.0 2158800.0 1452000.0 2166000.0 ;
      RECT  1448400.0 2151600.0 1449600.0 2152800.0 ;
      RECT  1450800.0 2151600.0 1452000.0 2152800.0 ;
      RECT  1450800.0 2151600.0 1452000.0 2152800.0 ;
      RECT  1448400.0 2151600.0 1449600.0 2152800.0 ;
      RECT  1448400.0 2158800.0 1449600.0 2160000.0 ;
      RECT  1450800.0 2158800.0 1452000.0 2160000.0 ;
      RECT  1450800.0 2158800.0 1452000.0 2160000.0 ;
      RECT  1448400.0 2158800.0 1449600.0 2160000.0 ;
      RECT  1450800.0 2158800.0 1452000.0 2160000.0 ;
      RECT  1453200.0 2158800.0 1454400.0 2160000.0 ;
      RECT  1453200.0 2158800.0 1454400.0 2160000.0 ;
      RECT  1450800.0 2158800.0 1452000.0 2160000.0 ;
      RECT  1450500.0 2153850.0 1449300.0 2155050.0 ;
      RECT  1450800.0 2164200.0 1452000.0 2165400.0 ;
      RECT  1448400.0 2151600.0 1449600.0 2152800.0 ;
      RECT  1450800.0 2151600.0 1452000.0 2152800.0 ;
      RECT  1448400.0 2158800.0 1449600.0 2160000.0 ;
      RECT  1453200.0 2158800.0 1454400.0 2160000.0 ;
      RECT  1445400.0 2154000.0 1455600.0 2154900.0 ;
      RECT  1445400.0 2165100.0 1455600.0 2166000.0 ;
      RECT  1461000.0 2158800.0 1462200.0 2166000.0 ;
      RECT  1458600.0 2151600.0 1459800.0 2152800.0 ;
      RECT  1461000.0 2151600.0 1462200.0 2152800.0 ;
      RECT  1461000.0 2151600.0 1462200.0 2152800.0 ;
      RECT  1458600.0 2151600.0 1459800.0 2152800.0 ;
      RECT  1458600.0 2158800.0 1459800.0 2160000.0 ;
      RECT  1461000.0 2158800.0 1462200.0 2160000.0 ;
      RECT  1461000.0 2158800.0 1462200.0 2160000.0 ;
      RECT  1458600.0 2158800.0 1459800.0 2160000.0 ;
      RECT  1461000.0 2158800.0 1462200.0 2160000.0 ;
      RECT  1463400.0 2158800.0 1464600.0 2160000.0 ;
      RECT  1463400.0 2158800.0 1464600.0 2160000.0 ;
      RECT  1461000.0 2158800.0 1462200.0 2160000.0 ;
      RECT  1460700.0 2153850.0 1459500.0 2155050.0 ;
      RECT  1461000.0 2164200.0 1462200.0 2165400.0 ;
      RECT  1458600.0 2151600.0 1459800.0 2152800.0 ;
      RECT  1461000.0 2151600.0 1462200.0 2152800.0 ;
      RECT  1458600.0 2158800.0 1459800.0 2160000.0 ;
      RECT  1463400.0 2158800.0 1464600.0 2160000.0 ;
      RECT  1455600.0 2154000.0 1465800.0 2154900.0 ;
      RECT  1455600.0 2165100.0 1465800.0 2166000.0 ;
      RECT  1471200.0 2158800.0 1472400.0 2166000.0 ;
      RECT  1468800.0 2151600.0 1470000.0 2152800.0 ;
      RECT  1471200.0 2151600.0 1472400.0 2152800.0 ;
      RECT  1471200.0 2151600.0 1472400.0 2152800.0 ;
      RECT  1468800.0 2151600.0 1470000.0 2152800.0 ;
      RECT  1468800.0 2158800.0 1470000.0 2160000.0 ;
      RECT  1471200.0 2158800.0 1472400.0 2160000.0 ;
      RECT  1471200.0 2158800.0 1472400.0 2160000.0 ;
      RECT  1468800.0 2158800.0 1470000.0 2160000.0 ;
      RECT  1471200.0 2158800.0 1472400.0 2160000.0 ;
      RECT  1473600.0 2158800.0 1474800.0 2160000.0 ;
      RECT  1473600.0 2158800.0 1474800.0 2160000.0 ;
      RECT  1471200.0 2158800.0 1472400.0 2160000.0 ;
      RECT  1470900.0 2153850.0 1469700.0 2155050.0 ;
      RECT  1471200.0 2164200.0 1472400.0 2165400.0 ;
      RECT  1468800.0 2151600.0 1470000.0 2152800.0 ;
      RECT  1471200.0 2151600.0 1472400.0 2152800.0 ;
      RECT  1468800.0 2158800.0 1470000.0 2160000.0 ;
      RECT  1473600.0 2158800.0 1474800.0 2160000.0 ;
      RECT  1465800.0 2154000.0 1476000.0 2154900.0 ;
      RECT  1465800.0 2165100.0 1476000.0 2166000.0 ;
      RECT  1481400.0 2158800.0 1482600.0 2166000.0 ;
      RECT  1479000.0 2151600.0 1480200.0 2152800.0 ;
      RECT  1481400.0 2151600.0 1482600.0 2152800.0 ;
      RECT  1481400.0 2151600.0 1482600.0 2152800.0 ;
      RECT  1479000.0 2151600.0 1480200.0 2152800.0 ;
      RECT  1479000.0 2158800.0 1480200.0 2160000.0 ;
      RECT  1481400.0 2158800.0 1482600.0 2160000.0 ;
      RECT  1481400.0 2158800.0 1482600.0 2160000.0 ;
      RECT  1479000.0 2158800.0 1480200.0 2160000.0 ;
      RECT  1481400.0 2158800.0 1482600.0 2160000.0 ;
      RECT  1483800.0 2158800.0 1485000.0 2160000.0 ;
      RECT  1483800.0 2158800.0 1485000.0 2160000.0 ;
      RECT  1481400.0 2158800.0 1482600.0 2160000.0 ;
      RECT  1481100.0 2153850.0 1479900.0 2155050.0 ;
      RECT  1481400.0 2164200.0 1482600.0 2165400.0 ;
      RECT  1479000.0 2151600.0 1480200.0 2152800.0 ;
      RECT  1481400.0 2151600.0 1482600.0 2152800.0 ;
      RECT  1479000.0 2158800.0 1480200.0 2160000.0 ;
      RECT  1483800.0 2158800.0 1485000.0 2160000.0 ;
      RECT  1476000.0 2154000.0 1486200.0 2154900.0 ;
      RECT  1476000.0 2165100.0 1486200.0 2166000.0 ;
      RECT  1491600.0 2158800.0 1492800.0 2166000.0 ;
      RECT  1489200.0 2151600.0 1490400.0 2152800.0 ;
      RECT  1491600.0 2151600.0 1492800.0 2152800.0 ;
      RECT  1491600.0 2151600.0 1492800.0 2152800.0 ;
      RECT  1489200.0 2151600.0 1490400.0 2152800.0 ;
      RECT  1489200.0 2158800.0 1490400.0 2160000.0 ;
      RECT  1491600.0 2158800.0 1492800.0 2160000.0 ;
      RECT  1491600.0 2158800.0 1492800.0 2160000.0 ;
      RECT  1489200.0 2158800.0 1490400.0 2160000.0 ;
      RECT  1491600.0 2158800.0 1492800.0 2160000.0 ;
      RECT  1494000.0 2158800.0 1495200.0 2160000.0 ;
      RECT  1494000.0 2158800.0 1495200.0 2160000.0 ;
      RECT  1491600.0 2158800.0 1492800.0 2160000.0 ;
      RECT  1491300.0 2153850.0 1490100.0 2155050.0 ;
      RECT  1491600.0 2164200.0 1492800.0 2165400.0 ;
      RECT  1489200.0 2151600.0 1490400.0 2152800.0 ;
      RECT  1491600.0 2151600.0 1492800.0 2152800.0 ;
      RECT  1489200.0 2158800.0 1490400.0 2160000.0 ;
      RECT  1494000.0 2158800.0 1495200.0 2160000.0 ;
      RECT  1486200.0 2154000.0 1496400.0 2154900.0 ;
      RECT  1486200.0 2165100.0 1496400.0 2166000.0 ;
      RECT  1501800.0 2158800.0 1503000.0 2166000.0 ;
      RECT  1499400.0 2151600.0 1500600.0 2152800.0 ;
      RECT  1501800.0 2151600.0 1503000.0 2152800.0 ;
      RECT  1501800.0 2151600.0 1503000.0 2152800.0 ;
      RECT  1499400.0 2151600.0 1500600.0 2152800.0 ;
      RECT  1499400.0 2158800.0 1500600.0 2160000.0 ;
      RECT  1501800.0 2158800.0 1503000.0 2160000.0 ;
      RECT  1501800.0 2158800.0 1503000.0 2160000.0 ;
      RECT  1499400.0 2158800.0 1500600.0 2160000.0 ;
      RECT  1501800.0 2158800.0 1503000.0 2160000.0 ;
      RECT  1504200.0 2158800.0 1505400.0 2160000.0 ;
      RECT  1504200.0 2158800.0 1505400.0 2160000.0 ;
      RECT  1501800.0 2158800.0 1503000.0 2160000.0 ;
      RECT  1501500.0 2153850.0 1500300.0 2155050.0 ;
      RECT  1501800.0 2164200.0 1503000.0 2165400.0 ;
      RECT  1499400.0 2151600.0 1500600.0 2152800.0 ;
      RECT  1501800.0 2151600.0 1503000.0 2152800.0 ;
      RECT  1499400.0 2158800.0 1500600.0 2160000.0 ;
      RECT  1504200.0 2158800.0 1505400.0 2160000.0 ;
      RECT  1496400.0 2154000.0 1506600.0 2154900.0 ;
      RECT  1496400.0 2165100.0 1506600.0 2166000.0 ;
      RECT  1512000.0 2158800.0 1513200.0 2166000.0 ;
      RECT  1509600.0 2151600.0 1510800.0 2152800.0 ;
      RECT  1512000.0 2151600.0 1513200.0 2152800.0 ;
      RECT  1512000.0 2151600.0 1513200.0 2152800.0 ;
      RECT  1509600.0 2151600.0 1510800.0 2152800.0 ;
      RECT  1509600.0 2158800.0 1510800.0 2160000.0 ;
      RECT  1512000.0 2158800.0 1513200.0 2160000.0 ;
      RECT  1512000.0 2158800.0 1513200.0 2160000.0 ;
      RECT  1509600.0 2158800.0 1510800.0 2160000.0 ;
      RECT  1512000.0 2158800.0 1513200.0 2160000.0 ;
      RECT  1514400.0 2158800.0 1515600.0 2160000.0 ;
      RECT  1514400.0 2158800.0 1515600.0 2160000.0 ;
      RECT  1512000.0 2158800.0 1513200.0 2160000.0 ;
      RECT  1511700.0 2153850.0 1510500.0 2155050.0 ;
      RECT  1512000.0 2164200.0 1513200.0 2165400.0 ;
      RECT  1509600.0 2151600.0 1510800.0 2152800.0 ;
      RECT  1512000.0 2151600.0 1513200.0 2152800.0 ;
      RECT  1509600.0 2158800.0 1510800.0 2160000.0 ;
      RECT  1514400.0 2158800.0 1515600.0 2160000.0 ;
      RECT  1506600.0 2154000.0 1516800.0 2154900.0 ;
      RECT  1506600.0 2165100.0 1516800.0 2166000.0 ;
      RECT  1522200.0 2158800.0 1523400.0 2166000.0 ;
      RECT  1519800.0 2151600.0 1521000.0 2152800.0 ;
      RECT  1522200.0 2151600.0 1523400.0 2152800.0 ;
      RECT  1522200.0 2151600.0 1523400.0 2152800.0 ;
      RECT  1519800.0 2151600.0 1521000.0 2152800.0 ;
      RECT  1519800.0 2158800.0 1521000.0 2160000.0 ;
      RECT  1522200.0 2158800.0 1523400.0 2160000.0 ;
      RECT  1522200.0 2158800.0 1523400.0 2160000.0 ;
      RECT  1519800.0 2158800.0 1521000.0 2160000.0 ;
      RECT  1522200.0 2158800.0 1523400.0 2160000.0 ;
      RECT  1524600.0 2158800.0 1525800.0 2160000.0 ;
      RECT  1524600.0 2158800.0 1525800.0 2160000.0 ;
      RECT  1522200.0 2158800.0 1523400.0 2160000.0 ;
      RECT  1521900.0 2153850.0 1520700.0 2155050.0 ;
      RECT  1522200.0 2164200.0 1523400.0 2165400.0 ;
      RECT  1519800.0 2151600.0 1521000.0 2152800.0 ;
      RECT  1522200.0 2151600.0 1523400.0 2152800.0 ;
      RECT  1519800.0 2158800.0 1521000.0 2160000.0 ;
      RECT  1524600.0 2158800.0 1525800.0 2160000.0 ;
      RECT  1516800.0 2154000.0 1527000.0 2154900.0 ;
      RECT  1516800.0 2165100.0 1527000.0 2166000.0 ;
      RECT  221400.0 2154000.0 1527000.0 2154900.0 ;
      RECT  221400.0 2165100.0 1527000.0 2166000.0 ;
      RECT  224400.0 342750.0 256200.0 343650.0 ;
      RECT  227400.0 340650.0 259200.0 341550.0 ;
      RECT  265200.0 342750.0 297000.0 343650.0 ;
      RECT  268200.0 340650.0 300000.0 341550.0 ;
      RECT  306000.0 342750.0 337800.0 343650.0 ;
      RECT  309000.0 340650.0 340800.0 341550.0 ;
      RECT  346800.0 342750.0 378600.0 343650.0 ;
      RECT  349800.0 340650.0 381600.0 341550.0 ;
      RECT  387600.0 342750.0 419400.0 343650.0 ;
      RECT  390600.0 340650.0 422400.0 341550.0 ;
      RECT  428400.0 342750.0 460200.0 343650.0 ;
      RECT  431400.0 340650.0 463200.0 341550.0 ;
      RECT  469200.0 342750.0 501000.0 343650.0 ;
      RECT  472200.0 340650.0 504000.0 341550.0 ;
      RECT  510000.0 342750.0 541800.0 343650.0 ;
      RECT  513000.0 340650.0 544800.0 341550.0 ;
      RECT  550800.0 342750.0 582600.0 343650.0 ;
      RECT  553800.0 340650.0 585600.0 341550.0 ;
      RECT  591600.0 342750.0 623400.0 343650.0 ;
      RECT  594600.0 340650.0 626400.0 341550.0 ;
      RECT  632400.0 342750.0 664200.0 343650.0 ;
      RECT  635400.0 340650.0 667200.0 341550.0 ;
      RECT  673200.0 342750.0 705000.0 343650.0 ;
      RECT  676200.0 340650.0 708000.0 341550.0 ;
      RECT  714000.0 342750.0 745800.0 343650.0 ;
      RECT  717000.0 340650.0 748800.0 341550.0 ;
      RECT  754800.0 342750.0 786600.0 343650.0 ;
      RECT  757800.0 340650.0 789600.0 341550.0 ;
      RECT  795600.0 342750.0 827400.0 343650.0 ;
      RECT  798600.0 340650.0 830400.0 341550.0 ;
      RECT  836400.0 342750.0 868200.0 343650.0 ;
      RECT  839400.0 340650.0 871200.0 341550.0 ;
      RECT  877200.0 342750.0 909000.0 343650.0 ;
      RECT  880200.0 340650.0 912000.0 341550.0 ;
      RECT  918000.0 342750.0 949800.0 343650.0 ;
      RECT  921000.0 340650.0 952800.0 341550.0 ;
      RECT  958800.0 342750.0 990600.0 343650.0 ;
      RECT  961800.0 340650.0 993600.0 341550.0 ;
      RECT  999600.0 342750.0 1031400.0 343650.0 ;
      RECT  1002600.0 340650.0 1034400.0 341550.0 ;
      RECT  1040400.0 342750.0 1072200.0 343650.0 ;
      RECT  1043400.0 340650.0 1075200.0 341550.0 ;
      RECT  1081200.0 342750.0 1113000.0 343650.0 ;
      RECT  1084200.0 340650.0 1116000.0 341550.0 ;
      RECT  1122000.0 342750.0 1153800.0 343650.0 ;
      RECT  1125000.0 340650.0 1156800.0 341550.0 ;
      RECT  1162800.0 342750.0 1194600.0 343650.0 ;
      RECT  1165800.0 340650.0 1197600.0 341550.0 ;
      RECT  1203600.0 342750.0 1235400.0 343650.0 ;
      RECT  1206600.0 340650.0 1238400.0 341550.0 ;
      RECT  1244400.0 342750.0 1276200.0 343650.0 ;
      RECT  1247400.0 340650.0 1279200.0 341550.0 ;
      RECT  1285200.0 342750.0 1317000.0 343650.0 ;
      RECT  1288200.0 340650.0 1320000.0 341550.0 ;
      RECT  1326000.0 342750.0 1357800.0 343650.0 ;
      RECT  1329000.0 340650.0 1360800.0 341550.0 ;
      RECT  1366800.0 342750.0 1398600.0 343650.0 ;
      RECT  1369800.0 340650.0 1401600.0 341550.0 ;
      RECT  1407600.0 342750.0 1439400.0 343650.0 ;
      RECT  1410600.0 340650.0 1442400.0 341550.0 ;
      RECT  1448400.0 342750.0 1480200.0 343650.0 ;
      RECT  1451400.0 340650.0 1483200.0 341550.0 ;
      RECT  1489200.0 342750.0 1521000.0 343650.0 ;
      RECT  1492200.0 340650.0 1524000.0 341550.0 ;
      RECT  227250.0 376500.0 228150.0 377400.0 ;
      RECT  224400.0 376500.0 227700.0 377400.0 ;
      RECT  227250.0 370350.0 228150.0 376950.0 ;
      RECT  224850.0 354600.0 225750.0 355500.0 ;
      RECT  225300.0 354600.0 227850.0 355500.0 ;
      RECT  224850.0 355050.0 225750.0 359850.0 ;
      RECT  224700.0 359250.0 225900.0 360450.0 ;
      RECT  227100.0 359250.0 228300.0 360450.0 ;
      RECT  227100.0 359250.0 228300.0 360450.0 ;
      RECT  224700.0 359250.0 225900.0 360450.0 ;
      RECT  224700.0 369750.0 225900.0 370950.0 ;
      RECT  227100.0 369750.0 228300.0 370950.0 ;
      RECT  227100.0 369750.0 228300.0 370950.0 ;
      RECT  224700.0 369750.0 225900.0 370950.0 ;
      RECT  224250.0 376350.0 225450.0 377550.0 ;
      RECT  227250.0 354450.0 228450.0 355650.0 ;
      RECT  224700.0 369750.0 225900.0 370950.0 ;
      RECT  227100.0 359250.0 228300.0 360450.0 ;
      RECT  231000.0 357450.0 232200.0 358650.0 ;
      RECT  231000.0 357450.0 232200.0 358650.0 ;
      RECT  237450.0 376500.0 238350.0 377400.0 ;
      RECT  234600.0 376500.0 237900.0 377400.0 ;
      RECT  237450.0 370350.0 238350.0 376950.0 ;
      RECT  235050.0 354600.0 235950.0 355500.0 ;
      RECT  235500.0 354600.0 238050.0 355500.0 ;
      RECT  235050.0 355050.0 235950.0 359850.0 ;
      RECT  234900.0 359250.0 236100.0 360450.0 ;
      RECT  237300.0 359250.0 238500.0 360450.0 ;
      RECT  237300.0 359250.0 238500.0 360450.0 ;
      RECT  234900.0 359250.0 236100.0 360450.0 ;
      RECT  234900.0 369750.0 236100.0 370950.0 ;
      RECT  237300.0 369750.0 238500.0 370950.0 ;
      RECT  237300.0 369750.0 238500.0 370950.0 ;
      RECT  234900.0 369750.0 236100.0 370950.0 ;
      RECT  234450.0 376350.0 235650.0 377550.0 ;
      RECT  237450.0 354450.0 238650.0 355650.0 ;
      RECT  234900.0 369750.0 236100.0 370950.0 ;
      RECT  237300.0 359250.0 238500.0 360450.0 ;
      RECT  241200.0 357450.0 242400.0 358650.0 ;
      RECT  241200.0 357450.0 242400.0 358650.0 ;
      RECT  247650.0 376500.0 248550.0 377400.0 ;
      RECT  244800.0 376500.0 248100.0 377400.0 ;
      RECT  247650.0 370350.0 248550.0 376950.0 ;
      RECT  245250.0 354600.0 246150.0 355500.0 ;
      RECT  245700.0 354600.0 248250.0 355500.0 ;
      RECT  245250.0 355050.0 246150.0 359850.0 ;
      RECT  245100.0 359250.0 246300.0 360450.0 ;
      RECT  247500.0 359250.0 248700.0 360450.0 ;
      RECT  247500.0 359250.0 248700.0 360450.0 ;
      RECT  245100.0 359250.0 246300.0 360450.0 ;
      RECT  245100.0 369750.0 246300.0 370950.0 ;
      RECT  247500.0 369750.0 248700.0 370950.0 ;
      RECT  247500.0 369750.0 248700.0 370950.0 ;
      RECT  245100.0 369750.0 246300.0 370950.0 ;
      RECT  244650.0 376350.0 245850.0 377550.0 ;
      RECT  247650.0 354450.0 248850.0 355650.0 ;
      RECT  245100.0 369750.0 246300.0 370950.0 ;
      RECT  247500.0 359250.0 248700.0 360450.0 ;
      RECT  251400.0 357450.0 252600.0 358650.0 ;
      RECT  251400.0 357450.0 252600.0 358650.0 ;
      RECT  257850.0 376500.0 258750.0 377400.0 ;
      RECT  255000.0 376500.0 258300.0 377400.0 ;
      RECT  257850.0 370350.0 258750.0 376950.0 ;
      RECT  255450.0 354600.0 256350.0 355500.0 ;
      RECT  255900.0 354600.0 258450.0 355500.0 ;
      RECT  255450.0 355050.0 256350.0 359850.0 ;
      RECT  255300.0 359250.0 256500.0 360450.0 ;
      RECT  257700.0 359250.0 258900.0 360450.0 ;
      RECT  257700.0 359250.0 258900.0 360450.0 ;
      RECT  255300.0 359250.0 256500.0 360450.0 ;
      RECT  255300.0 369750.0 256500.0 370950.0 ;
      RECT  257700.0 369750.0 258900.0 370950.0 ;
      RECT  257700.0 369750.0 258900.0 370950.0 ;
      RECT  255300.0 369750.0 256500.0 370950.0 ;
      RECT  254850.0 376350.0 256050.0 377550.0 ;
      RECT  257850.0 354450.0 259050.0 355650.0 ;
      RECT  255300.0 369750.0 256500.0 370950.0 ;
      RECT  257700.0 359250.0 258900.0 360450.0 ;
      RECT  261600.0 357450.0 262800.0 358650.0 ;
      RECT  261600.0 357450.0 262800.0 358650.0 ;
      RECT  268050.0 376500.0 268950.0 377400.0 ;
      RECT  265200.0 376500.0 268500.0 377400.0 ;
      RECT  268050.0 370350.0 268950.0 376950.0 ;
      RECT  265650.0 354600.0 266550.0 355500.0 ;
      RECT  266100.0 354600.0 268650.0 355500.0 ;
      RECT  265650.0 355050.0 266550.0 359850.0 ;
      RECT  265500.0 359250.0 266700.0 360450.0 ;
      RECT  267900.0 359250.0 269100.0 360450.0 ;
      RECT  267900.0 359250.0 269100.0 360450.0 ;
      RECT  265500.0 359250.0 266700.0 360450.0 ;
      RECT  265500.0 369750.0 266700.0 370950.0 ;
      RECT  267900.0 369750.0 269100.0 370950.0 ;
      RECT  267900.0 369750.0 269100.0 370950.0 ;
      RECT  265500.0 369750.0 266700.0 370950.0 ;
      RECT  265050.0 376350.0 266250.0 377550.0 ;
      RECT  268050.0 354450.0 269250.0 355650.0 ;
      RECT  265500.0 369750.0 266700.0 370950.0 ;
      RECT  267900.0 359250.0 269100.0 360450.0 ;
      RECT  271800.0 357450.0 273000.0 358650.0 ;
      RECT  271800.0 357450.0 273000.0 358650.0 ;
      RECT  278250.0 376500.0 279150.0 377400.0 ;
      RECT  275400.0 376500.0 278700.0 377400.0 ;
      RECT  278250.0 370350.0 279150.0 376950.0 ;
      RECT  275850.0 354600.0 276750.0 355500.0 ;
      RECT  276300.0 354600.0 278850.0 355500.0 ;
      RECT  275850.0 355050.0 276750.0 359850.0 ;
      RECT  275700.0 359250.0 276900.0 360450.0 ;
      RECT  278100.0 359250.0 279300.0 360450.0 ;
      RECT  278100.0 359250.0 279300.0 360450.0 ;
      RECT  275700.0 359250.0 276900.0 360450.0 ;
      RECT  275700.0 369750.0 276900.0 370950.0 ;
      RECT  278100.0 369750.0 279300.0 370950.0 ;
      RECT  278100.0 369750.0 279300.0 370950.0 ;
      RECT  275700.0 369750.0 276900.0 370950.0 ;
      RECT  275250.0 376350.0 276450.0 377550.0 ;
      RECT  278250.0 354450.0 279450.0 355650.0 ;
      RECT  275700.0 369750.0 276900.0 370950.0 ;
      RECT  278100.0 359250.0 279300.0 360450.0 ;
      RECT  282000.0 357450.0 283200.0 358650.0 ;
      RECT  282000.0 357450.0 283200.0 358650.0 ;
      RECT  288450.0 376500.0 289350.0 377400.0 ;
      RECT  285600.0 376500.0 288900.0 377400.0 ;
      RECT  288450.0 370350.0 289350.0 376950.0 ;
      RECT  286050.0 354600.0 286950.0 355500.0 ;
      RECT  286500.0 354600.0 289050.0 355500.0 ;
      RECT  286050.0 355050.0 286950.0 359850.0 ;
      RECT  285900.0 359250.0 287100.0 360450.0 ;
      RECT  288300.0 359250.0 289500.0 360450.0 ;
      RECT  288300.0 359250.0 289500.0 360450.0 ;
      RECT  285900.0 359250.0 287100.0 360450.0 ;
      RECT  285900.0 369750.0 287100.0 370950.0 ;
      RECT  288300.0 369750.0 289500.0 370950.0 ;
      RECT  288300.0 369750.0 289500.0 370950.0 ;
      RECT  285900.0 369750.0 287100.0 370950.0 ;
      RECT  285450.0 376350.0 286650.0 377550.0 ;
      RECT  288450.0 354450.0 289650.0 355650.0 ;
      RECT  285900.0 369750.0 287100.0 370950.0 ;
      RECT  288300.0 359250.0 289500.0 360450.0 ;
      RECT  292200.0 357450.0 293400.0 358650.0 ;
      RECT  292200.0 357450.0 293400.0 358650.0 ;
      RECT  298650.0 376500.0 299550.0 377400.0 ;
      RECT  295800.0 376500.0 299100.0 377400.0 ;
      RECT  298650.0 370350.0 299550.0 376950.0 ;
      RECT  296250.0 354600.0 297150.0 355500.0 ;
      RECT  296700.0 354600.0 299250.0 355500.0 ;
      RECT  296250.0 355050.0 297150.0 359850.0 ;
      RECT  296100.0 359250.0 297300.0 360450.0 ;
      RECT  298500.0 359250.0 299700.0 360450.0 ;
      RECT  298500.0 359250.0 299700.0 360450.0 ;
      RECT  296100.0 359250.0 297300.0 360450.0 ;
      RECT  296100.0 369750.0 297300.0 370950.0 ;
      RECT  298500.0 369750.0 299700.0 370950.0 ;
      RECT  298500.0 369750.0 299700.0 370950.0 ;
      RECT  296100.0 369750.0 297300.0 370950.0 ;
      RECT  295650.0 376350.0 296850.0 377550.0 ;
      RECT  298650.0 354450.0 299850.0 355650.0 ;
      RECT  296100.0 369750.0 297300.0 370950.0 ;
      RECT  298500.0 359250.0 299700.0 360450.0 ;
      RECT  302400.0 357450.0 303600.0 358650.0 ;
      RECT  302400.0 357450.0 303600.0 358650.0 ;
      RECT  308850.0 376500.0 309750.0 377400.0 ;
      RECT  306000.0 376500.0 309300.0 377400.0 ;
      RECT  308850.0 370350.0 309750.0 376950.0 ;
      RECT  306450.0 354600.0 307350.0 355500.0 ;
      RECT  306900.0 354600.0 309450.0 355500.0 ;
      RECT  306450.0 355050.0 307350.0 359850.0 ;
      RECT  306300.0 359250.0 307500.0 360450.0 ;
      RECT  308700.0 359250.0 309900.0 360450.0 ;
      RECT  308700.0 359250.0 309900.0 360450.0 ;
      RECT  306300.0 359250.0 307500.0 360450.0 ;
      RECT  306300.0 369750.0 307500.0 370950.0 ;
      RECT  308700.0 369750.0 309900.0 370950.0 ;
      RECT  308700.0 369750.0 309900.0 370950.0 ;
      RECT  306300.0 369750.0 307500.0 370950.0 ;
      RECT  305850.0 376350.0 307050.0 377550.0 ;
      RECT  308850.0 354450.0 310050.0 355650.0 ;
      RECT  306300.0 369750.0 307500.0 370950.0 ;
      RECT  308700.0 359250.0 309900.0 360450.0 ;
      RECT  312600.0 357450.0 313800.0 358650.0 ;
      RECT  312600.0 357450.0 313800.0 358650.0 ;
      RECT  319050.0 376500.0 319950.0 377400.0 ;
      RECT  316200.0 376500.0 319500.0 377400.0 ;
      RECT  319050.0 370350.0 319950.0 376950.0 ;
      RECT  316650.0 354600.0 317550.0 355500.0 ;
      RECT  317100.0 354600.0 319650.0 355500.0 ;
      RECT  316650.0 355050.0 317550.0 359850.0 ;
      RECT  316500.0 359250.0 317700.0 360450.0 ;
      RECT  318900.0 359250.0 320100.0 360450.0 ;
      RECT  318900.0 359250.0 320100.0 360450.0 ;
      RECT  316500.0 359250.0 317700.0 360450.0 ;
      RECT  316500.0 369750.0 317700.0 370950.0 ;
      RECT  318900.0 369750.0 320100.0 370950.0 ;
      RECT  318900.0 369750.0 320100.0 370950.0 ;
      RECT  316500.0 369750.0 317700.0 370950.0 ;
      RECT  316050.0 376350.0 317250.0 377550.0 ;
      RECT  319050.0 354450.0 320250.0 355650.0 ;
      RECT  316500.0 369750.0 317700.0 370950.0 ;
      RECT  318900.0 359250.0 320100.0 360450.0 ;
      RECT  322800.0 357450.0 324000.0 358650.0 ;
      RECT  322800.0 357450.0 324000.0 358650.0 ;
      RECT  329250.0 376500.0 330150.0 377400.0 ;
      RECT  326400.0 376500.0 329700.0 377400.0 ;
      RECT  329250.0 370350.0 330150.0 376950.0 ;
      RECT  326850.0 354600.0 327750.0 355500.0 ;
      RECT  327300.0 354600.0 329850.0 355500.0 ;
      RECT  326850.0 355050.0 327750.0 359850.0 ;
      RECT  326700.0 359250.0 327900.0 360450.0 ;
      RECT  329100.0 359250.0 330300.0 360450.0 ;
      RECT  329100.0 359250.0 330300.0 360450.0 ;
      RECT  326700.0 359250.0 327900.0 360450.0 ;
      RECT  326700.0 369750.0 327900.0 370950.0 ;
      RECT  329100.0 369750.0 330300.0 370950.0 ;
      RECT  329100.0 369750.0 330300.0 370950.0 ;
      RECT  326700.0 369750.0 327900.0 370950.0 ;
      RECT  326250.0 376350.0 327450.0 377550.0 ;
      RECT  329250.0 354450.0 330450.0 355650.0 ;
      RECT  326700.0 369750.0 327900.0 370950.0 ;
      RECT  329100.0 359250.0 330300.0 360450.0 ;
      RECT  333000.0 357450.0 334200.0 358650.0 ;
      RECT  333000.0 357450.0 334200.0 358650.0 ;
      RECT  339450.0 376500.0 340350.0 377400.0 ;
      RECT  336600.0 376500.0 339900.0 377400.0 ;
      RECT  339450.0 370350.0 340350.0 376950.0 ;
      RECT  337050.0 354600.0 337950.0 355500.0 ;
      RECT  337500.0 354600.0 340050.0 355500.0 ;
      RECT  337050.0 355050.0 337950.0 359850.0 ;
      RECT  336900.0 359250.0 338100.0 360450.0 ;
      RECT  339300.0 359250.0 340500.0 360450.0 ;
      RECT  339300.0 359250.0 340500.0 360450.0 ;
      RECT  336900.0 359250.0 338100.0 360450.0 ;
      RECT  336900.0 369750.0 338100.0 370950.0 ;
      RECT  339300.0 369750.0 340500.0 370950.0 ;
      RECT  339300.0 369750.0 340500.0 370950.0 ;
      RECT  336900.0 369750.0 338100.0 370950.0 ;
      RECT  336450.0 376350.0 337650.0 377550.0 ;
      RECT  339450.0 354450.0 340650.0 355650.0 ;
      RECT  336900.0 369750.0 338100.0 370950.0 ;
      RECT  339300.0 359250.0 340500.0 360450.0 ;
      RECT  343200.0 357450.0 344400.0 358650.0 ;
      RECT  343200.0 357450.0 344400.0 358650.0 ;
      RECT  349650.0 376500.0 350550.0 377400.0 ;
      RECT  346800.0 376500.0 350100.0 377400.0 ;
      RECT  349650.0 370350.0 350550.0 376950.0 ;
      RECT  347250.0 354600.0 348150.0 355500.0 ;
      RECT  347700.0 354600.0 350250.0 355500.0 ;
      RECT  347250.0 355050.0 348150.0 359850.0 ;
      RECT  347100.0 359250.0 348300.0 360450.0 ;
      RECT  349500.0 359250.0 350700.0 360450.0 ;
      RECT  349500.0 359250.0 350700.0 360450.0 ;
      RECT  347100.0 359250.0 348300.0 360450.0 ;
      RECT  347100.0 369750.0 348300.0 370950.0 ;
      RECT  349500.0 369750.0 350700.0 370950.0 ;
      RECT  349500.0 369750.0 350700.0 370950.0 ;
      RECT  347100.0 369750.0 348300.0 370950.0 ;
      RECT  346650.0 376350.0 347850.0 377550.0 ;
      RECT  349650.0 354450.0 350850.0 355650.0 ;
      RECT  347100.0 369750.0 348300.0 370950.0 ;
      RECT  349500.0 359250.0 350700.0 360450.0 ;
      RECT  353400.0 357450.0 354600.0 358650.0 ;
      RECT  353400.0 357450.0 354600.0 358650.0 ;
      RECT  359850.0 376500.0 360750.0 377400.0 ;
      RECT  357000.0 376500.0 360300.0 377400.0 ;
      RECT  359850.0 370350.0 360750.0 376950.0 ;
      RECT  357450.0 354600.0 358350.0 355500.0 ;
      RECT  357900.0 354600.0 360450.0 355500.0 ;
      RECT  357450.0 355050.0 358350.0 359850.0 ;
      RECT  357300.0 359250.0 358500.0 360450.0 ;
      RECT  359700.0 359250.0 360900.0 360450.0 ;
      RECT  359700.0 359250.0 360900.0 360450.0 ;
      RECT  357300.0 359250.0 358500.0 360450.0 ;
      RECT  357300.0 369750.0 358500.0 370950.0 ;
      RECT  359700.0 369750.0 360900.0 370950.0 ;
      RECT  359700.0 369750.0 360900.0 370950.0 ;
      RECT  357300.0 369750.0 358500.0 370950.0 ;
      RECT  356850.0 376350.0 358050.0 377550.0 ;
      RECT  359850.0 354450.0 361050.0 355650.0 ;
      RECT  357300.0 369750.0 358500.0 370950.0 ;
      RECT  359700.0 359250.0 360900.0 360450.0 ;
      RECT  363600.0 357450.0 364800.0 358650.0 ;
      RECT  363600.0 357450.0 364800.0 358650.0 ;
      RECT  370050.0 376500.0 370950.0 377400.0 ;
      RECT  367200.0 376500.0 370500.0 377400.0 ;
      RECT  370050.0 370350.0 370950.0 376950.0 ;
      RECT  367650.0 354600.0 368550.0 355500.0 ;
      RECT  368100.0 354600.0 370650.0 355500.0 ;
      RECT  367650.0 355050.0 368550.0 359850.0 ;
      RECT  367500.0 359250.0 368700.0 360450.0 ;
      RECT  369900.0 359250.0 371100.0 360450.0 ;
      RECT  369900.0 359250.0 371100.0 360450.0 ;
      RECT  367500.0 359250.0 368700.0 360450.0 ;
      RECT  367500.0 369750.0 368700.0 370950.0 ;
      RECT  369900.0 369750.0 371100.0 370950.0 ;
      RECT  369900.0 369750.0 371100.0 370950.0 ;
      RECT  367500.0 369750.0 368700.0 370950.0 ;
      RECT  367050.0 376350.0 368250.0 377550.0 ;
      RECT  370050.0 354450.0 371250.0 355650.0 ;
      RECT  367500.0 369750.0 368700.0 370950.0 ;
      RECT  369900.0 359250.0 371100.0 360450.0 ;
      RECT  373800.0 357450.0 375000.0 358650.0 ;
      RECT  373800.0 357450.0 375000.0 358650.0 ;
      RECT  380250.0 376500.0 381150.0 377400.0 ;
      RECT  377400.0 376500.0 380700.0 377400.0 ;
      RECT  380250.0 370350.0 381150.0 376950.0 ;
      RECT  377850.0 354600.0 378750.0 355500.0 ;
      RECT  378300.0 354600.0 380850.0 355500.0 ;
      RECT  377850.0 355050.0 378750.0 359850.0 ;
      RECT  377700.0 359250.0 378900.0 360450.0 ;
      RECT  380100.0 359250.0 381300.0 360450.0 ;
      RECT  380100.0 359250.0 381300.0 360450.0 ;
      RECT  377700.0 359250.0 378900.0 360450.0 ;
      RECT  377700.0 369750.0 378900.0 370950.0 ;
      RECT  380100.0 369750.0 381300.0 370950.0 ;
      RECT  380100.0 369750.0 381300.0 370950.0 ;
      RECT  377700.0 369750.0 378900.0 370950.0 ;
      RECT  377250.0 376350.0 378450.0 377550.0 ;
      RECT  380250.0 354450.0 381450.0 355650.0 ;
      RECT  377700.0 369750.0 378900.0 370950.0 ;
      RECT  380100.0 359250.0 381300.0 360450.0 ;
      RECT  384000.0 357450.0 385200.0 358650.0 ;
      RECT  384000.0 357450.0 385200.0 358650.0 ;
      RECT  390450.0 376500.0 391350.0 377400.0 ;
      RECT  387600.0 376500.0 390900.0 377400.0 ;
      RECT  390450.0 370350.0 391350.0 376950.0 ;
      RECT  388050.0 354600.0 388950.0 355500.0 ;
      RECT  388500.0 354600.0 391050.0 355500.0 ;
      RECT  388050.0 355050.0 388950.0 359850.0 ;
      RECT  387900.0 359250.0 389100.0 360450.0 ;
      RECT  390300.0 359250.0 391500.0 360450.0 ;
      RECT  390300.0 359250.0 391500.0 360450.0 ;
      RECT  387900.0 359250.0 389100.0 360450.0 ;
      RECT  387900.0 369750.0 389100.0 370950.0 ;
      RECT  390300.0 369750.0 391500.0 370950.0 ;
      RECT  390300.0 369750.0 391500.0 370950.0 ;
      RECT  387900.0 369750.0 389100.0 370950.0 ;
      RECT  387450.0 376350.0 388650.0 377550.0 ;
      RECT  390450.0 354450.0 391650.0 355650.0 ;
      RECT  387900.0 369750.0 389100.0 370950.0 ;
      RECT  390300.0 359250.0 391500.0 360450.0 ;
      RECT  394200.0 357450.0 395400.0 358650.0 ;
      RECT  394200.0 357450.0 395400.0 358650.0 ;
      RECT  400650.0 376500.0 401550.0 377400.0 ;
      RECT  397800.0 376500.0 401100.0 377400.0 ;
      RECT  400650.0 370350.0 401550.0 376950.0 ;
      RECT  398250.0 354600.0 399150.0 355500.0 ;
      RECT  398700.0 354600.0 401250.0 355500.0 ;
      RECT  398250.0 355050.0 399150.0 359850.0 ;
      RECT  398100.0 359250.0 399300.0 360450.0 ;
      RECT  400500.0 359250.0 401700.0 360450.0 ;
      RECT  400500.0 359250.0 401700.0 360450.0 ;
      RECT  398100.0 359250.0 399300.0 360450.0 ;
      RECT  398100.0 369750.0 399300.0 370950.0 ;
      RECT  400500.0 369750.0 401700.0 370950.0 ;
      RECT  400500.0 369750.0 401700.0 370950.0 ;
      RECT  398100.0 369750.0 399300.0 370950.0 ;
      RECT  397650.0 376350.0 398850.0 377550.0 ;
      RECT  400650.0 354450.0 401850.0 355650.0 ;
      RECT  398100.0 369750.0 399300.0 370950.0 ;
      RECT  400500.0 359250.0 401700.0 360450.0 ;
      RECT  404400.0 357450.0 405600.0 358650.0 ;
      RECT  404400.0 357450.0 405600.0 358650.0 ;
      RECT  410850.0 376500.0 411750.0 377400.0 ;
      RECT  408000.0 376500.0 411300.0 377400.0 ;
      RECT  410850.0 370350.0 411750.0 376950.0 ;
      RECT  408450.0 354600.0 409350.0 355500.0 ;
      RECT  408900.0 354600.0 411450.0 355500.0 ;
      RECT  408450.0 355050.0 409350.0 359850.0 ;
      RECT  408300.0 359250.0 409500.0 360450.0 ;
      RECT  410700.0 359250.0 411900.0 360450.0 ;
      RECT  410700.0 359250.0 411900.0 360450.0 ;
      RECT  408300.0 359250.0 409500.0 360450.0 ;
      RECT  408300.0 369750.0 409500.0 370950.0 ;
      RECT  410700.0 369750.0 411900.0 370950.0 ;
      RECT  410700.0 369750.0 411900.0 370950.0 ;
      RECT  408300.0 369750.0 409500.0 370950.0 ;
      RECT  407850.0 376350.0 409050.0 377550.0 ;
      RECT  410850.0 354450.0 412050.0 355650.0 ;
      RECT  408300.0 369750.0 409500.0 370950.0 ;
      RECT  410700.0 359250.0 411900.0 360450.0 ;
      RECT  414600.0 357450.0 415800.0 358650.0 ;
      RECT  414600.0 357450.0 415800.0 358650.0 ;
      RECT  421050.0 376500.0 421950.0 377400.0 ;
      RECT  418200.0 376500.0 421500.0 377400.0 ;
      RECT  421050.0 370350.0 421950.0 376950.0 ;
      RECT  418650.0 354600.0 419550.0 355500.0 ;
      RECT  419100.0 354600.0 421650.0 355500.0 ;
      RECT  418650.0 355050.0 419550.0 359850.0 ;
      RECT  418500.0 359250.0 419700.0 360450.0 ;
      RECT  420900.0 359250.0 422100.0 360450.0 ;
      RECT  420900.0 359250.0 422100.0 360450.0 ;
      RECT  418500.0 359250.0 419700.0 360450.0 ;
      RECT  418500.0 369750.0 419700.0 370950.0 ;
      RECT  420900.0 369750.0 422100.0 370950.0 ;
      RECT  420900.0 369750.0 422100.0 370950.0 ;
      RECT  418500.0 369750.0 419700.0 370950.0 ;
      RECT  418050.0 376350.0 419250.0 377550.0 ;
      RECT  421050.0 354450.0 422250.0 355650.0 ;
      RECT  418500.0 369750.0 419700.0 370950.0 ;
      RECT  420900.0 359250.0 422100.0 360450.0 ;
      RECT  424800.0 357450.0 426000.0 358650.0 ;
      RECT  424800.0 357450.0 426000.0 358650.0 ;
      RECT  431250.0 376500.0 432150.0 377400.0 ;
      RECT  428400.0 376500.0 431700.0 377400.0 ;
      RECT  431250.0 370350.0 432150.0 376950.0 ;
      RECT  428850.0 354600.0 429750.0 355500.0 ;
      RECT  429300.0 354600.0 431850.0 355500.0 ;
      RECT  428850.0 355050.0 429750.0 359850.0 ;
      RECT  428700.0 359250.0 429900.0 360450.0 ;
      RECT  431100.0 359250.0 432300.0 360450.0 ;
      RECT  431100.0 359250.0 432300.0 360450.0 ;
      RECT  428700.0 359250.0 429900.0 360450.0 ;
      RECT  428700.0 369750.0 429900.0 370950.0 ;
      RECT  431100.0 369750.0 432300.0 370950.0 ;
      RECT  431100.0 369750.0 432300.0 370950.0 ;
      RECT  428700.0 369750.0 429900.0 370950.0 ;
      RECT  428250.0 376350.0 429450.0 377550.0 ;
      RECT  431250.0 354450.0 432450.0 355650.0 ;
      RECT  428700.0 369750.0 429900.0 370950.0 ;
      RECT  431100.0 359250.0 432300.0 360450.0 ;
      RECT  435000.0 357450.0 436200.0 358650.0 ;
      RECT  435000.0 357450.0 436200.0 358650.0 ;
      RECT  441450.0 376500.0 442350.0 377400.0 ;
      RECT  438600.0 376500.0 441900.0 377400.0 ;
      RECT  441450.0 370350.0 442350.0 376950.0 ;
      RECT  439050.0 354600.0 439950.0 355500.0 ;
      RECT  439500.0 354600.0 442050.0 355500.0 ;
      RECT  439050.0 355050.0 439950.0 359850.0 ;
      RECT  438900.0 359250.0 440100.0 360450.0 ;
      RECT  441300.0 359250.0 442500.0 360450.0 ;
      RECT  441300.0 359250.0 442500.0 360450.0 ;
      RECT  438900.0 359250.0 440100.0 360450.0 ;
      RECT  438900.0 369750.0 440100.0 370950.0 ;
      RECT  441300.0 369750.0 442500.0 370950.0 ;
      RECT  441300.0 369750.0 442500.0 370950.0 ;
      RECT  438900.0 369750.0 440100.0 370950.0 ;
      RECT  438450.0 376350.0 439650.0 377550.0 ;
      RECT  441450.0 354450.0 442650.0 355650.0 ;
      RECT  438900.0 369750.0 440100.0 370950.0 ;
      RECT  441300.0 359250.0 442500.0 360450.0 ;
      RECT  445200.0 357450.0 446400.0 358650.0 ;
      RECT  445200.0 357450.0 446400.0 358650.0 ;
      RECT  451650.0 376500.0 452550.0 377400.0 ;
      RECT  448800.0 376500.0 452100.0 377400.0 ;
      RECT  451650.0 370350.0 452550.0 376950.0 ;
      RECT  449250.0 354600.0 450150.0 355500.0 ;
      RECT  449700.0 354600.0 452250.0 355500.0 ;
      RECT  449250.0 355050.0 450150.0 359850.0 ;
      RECT  449100.0 359250.0 450300.0 360450.0 ;
      RECT  451500.0 359250.0 452700.0 360450.0 ;
      RECT  451500.0 359250.0 452700.0 360450.0 ;
      RECT  449100.0 359250.0 450300.0 360450.0 ;
      RECT  449100.0 369750.0 450300.0 370950.0 ;
      RECT  451500.0 369750.0 452700.0 370950.0 ;
      RECT  451500.0 369750.0 452700.0 370950.0 ;
      RECT  449100.0 369750.0 450300.0 370950.0 ;
      RECT  448650.0 376350.0 449850.0 377550.0 ;
      RECT  451650.0 354450.0 452850.0 355650.0 ;
      RECT  449100.0 369750.0 450300.0 370950.0 ;
      RECT  451500.0 359250.0 452700.0 360450.0 ;
      RECT  455400.0 357450.0 456600.0 358650.0 ;
      RECT  455400.0 357450.0 456600.0 358650.0 ;
      RECT  461850.0 376500.0 462750.0 377400.0 ;
      RECT  459000.0 376500.0 462300.0 377400.0 ;
      RECT  461850.0 370350.0 462750.0 376950.0 ;
      RECT  459450.0 354600.0 460350.0 355500.0 ;
      RECT  459900.0 354600.0 462450.0 355500.0 ;
      RECT  459450.0 355050.0 460350.0 359850.0 ;
      RECT  459300.0 359250.0 460500.0 360450.0 ;
      RECT  461700.0 359250.0 462900.0 360450.0 ;
      RECT  461700.0 359250.0 462900.0 360450.0 ;
      RECT  459300.0 359250.0 460500.0 360450.0 ;
      RECT  459300.0 369750.0 460500.0 370950.0 ;
      RECT  461700.0 369750.0 462900.0 370950.0 ;
      RECT  461700.0 369750.0 462900.0 370950.0 ;
      RECT  459300.0 369750.0 460500.0 370950.0 ;
      RECT  458850.0 376350.0 460050.0 377550.0 ;
      RECT  461850.0 354450.0 463050.0 355650.0 ;
      RECT  459300.0 369750.0 460500.0 370950.0 ;
      RECT  461700.0 359250.0 462900.0 360450.0 ;
      RECT  465600.0 357450.0 466800.0 358650.0 ;
      RECT  465600.0 357450.0 466800.0 358650.0 ;
      RECT  472050.0 376500.0 472950.0 377400.0 ;
      RECT  469200.0 376500.0 472500.0 377400.0 ;
      RECT  472050.0 370350.0 472950.0 376950.0 ;
      RECT  469650.0 354600.0 470550.0 355500.0 ;
      RECT  470100.0 354600.0 472650.0 355500.0 ;
      RECT  469650.0 355050.0 470550.0 359850.0 ;
      RECT  469500.0 359250.0 470700.0 360450.0 ;
      RECT  471900.0 359250.0 473100.0 360450.0 ;
      RECT  471900.0 359250.0 473100.0 360450.0 ;
      RECT  469500.0 359250.0 470700.0 360450.0 ;
      RECT  469500.0 369750.0 470700.0 370950.0 ;
      RECT  471900.0 369750.0 473100.0 370950.0 ;
      RECT  471900.0 369750.0 473100.0 370950.0 ;
      RECT  469500.0 369750.0 470700.0 370950.0 ;
      RECT  469050.0 376350.0 470250.0 377550.0 ;
      RECT  472050.0 354450.0 473250.0 355650.0 ;
      RECT  469500.0 369750.0 470700.0 370950.0 ;
      RECT  471900.0 359250.0 473100.0 360450.0 ;
      RECT  475800.0 357450.0 477000.0 358650.0 ;
      RECT  475800.0 357450.0 477000.0 358650.0 ;
      RECT  482250.0 376500.0 483150.0 377400.0 ;
      RECT  479400.0 376500.0 482700.0 377400.0 ;
      RECT  482250.0 370350.0 483150.0 376950.0 ;
      RECT  479850.0 354600.0 480750.0 355500.0 ;
      RECT  480300.0 354600.0 482850.0 355500.0 ;
      RECT  479850.0 355050.0 480750.0 359850.0 ;
      RECT  479700.0 359250.0 480900.0 360450.0 ;
      RECT  482100.0 359250.0 483300.0 360450.0 ;
      RECT  482100.0 359250.0 483300.0 360450.0 ;
      RECT  479700.0 359250.0 480900.0 360450.0 ;
      RECT  479700.0 369750.0 480900.0 370950.0 ;
      RECT  482100.0 369750.0 483300.0 370950.0 ;
      RECT  482100.0 369750.0 483300.0 370950.0 ;
      RECT  479700.0 369750.0 480900.0 370950.0 ;
      RECT  479250.0 376350.0 480450.0 377550.0 ;
      RECT  482250.0 354450.0 483450.0 355650.0 ;
      RECT  479700.0 369750.0 480900.0 370950.0 ;
      RECT  482100.0 359250.0 483300.0 360450.0 ;
      RECT  486000.0 357450.0 487200.0 358650.0 ;
      RECT  486000.0 357450.0 487200.0 358650.0 ;
      RECT  492450.0 376500.0 493350.0 377400.0 ;
      RECT  489600.0 376500.0 492900.0 377400.0 ;
      RECT  492450.0 370350.0 493350.0 376950.0 ;
      RECT  490050.0 354600.0 490950.0 355500.0 ;
      RECT  490500.0 354600.0 493050.0 355500.0 ;
      RECT  490050.0 355050.0 490950.0 359850.0 ;
      RECT  489900.0 359250.0 491100.0 360450.0 ;
      RECT  492300.0 359250.0 493500.0 360450.0 ;
      RECT  492300.0 359250.0 493500.0 360450.0 ;
      RECT  489900.0 359250.0 491100.0 360450.0 ;
      RECT  489900.0 369750.0 491100.0 370950.0 ;
      RECT  492300.0 369750.0 493500.0 370950.0 ;
      RECT  492300.0 369750.0 493500.0 370950.0 ;
      RECT  489900.0 369750.0 491100.0 370950.0 ;
      RECT  489450.0 376350.0 490650.0 377550.0 ;
      RECT  492450.0 354450.0 493650.0 355650.0 ;
      RECT  489900.0 369750.0 491100.0 370950.0 ;
      RECT  492300.0 359250.0 493500.0 360450.0 ;
      RECT  496200.0 357450.0 497400.0 358650.0 ;
      RECT  496200.0 357450.0 497400.0 358650.0 ;
      RECT  502650.0 376500.0 503550.0 377400.0 ;
      RECT  499800.0 376500.0 503100.0 377400.0 ;
      RECT  502650.0 370350.0 503550.0 376950.0 ;
      RECT  500250.0 354600.0 501150.0 355500.0 ;
      RECT  500700.0 354600.0 503250.0 355500.0 ;
      RECT  500250.0 355050.0 501150.0 359850.0 ;
      RECT  500100.0 359250.0 501300.0 360450.0 ;
      RECT  502500.0 359250.0 503700.0 360450.0 ;
      RECT  502500.0 359250.0 503700.0 360450.0 ;
      RECT  500100.0 359250.0 501300.0 360450.0 ;
      RECT  500100.0 369750.0 501300.0 370950.0 ;
      RECT  502500.0 369750.0 503700.0 370950.0 ;
      RECT  502500.0 369750.0 503700.0 370950.0 ;
      RECT  500100.0 369750.0 501300.0 370950.0 ;
      RECT  499650.0 376350.0 500850.0 377550.0 ;
      RECT  502650.0 354450.0 503850.0 355650.0 ;
      RECT  500100.0 369750.0 501300.0 370950.0 ;
      RECT  502500.0 359250.0 503700.0 360450.0 ;
      RECT  506400.0 357450.0 507600.0 358650.0 ;
      RECT  506400.0 357450.0 507600.0 358650.0 ;
      RECT  512850.0 376500.0 513750.0 377400.0 ;
      RECT  510000.0 376500.0 513300.0 377400.0 ;
      RECT  512850.0 370350.0 513750.0 376950.0 ;
      RECT  510450.0 354600.0 511350.0 355500.0 ;
      RECT  510900.0 354600.0 513450.0 355500.0 ;
      RECT  510450.0 355050.0 511350.0 359850.0 ;
      RECT  510300.0 359250.0 511500.0 360450.0 ;
      RECT  512700.0 359250.0 513900.0 360450.0 ;
      RECT  512700.0 359250.0 513900.0 360450.0 ;
      RECT  510300.0 359250.0 511500.0 360450.0 ;
      RECT  510300.0 369750.0 511500.0 370950.0 ;
      RECT  512700.0 369750.0 513900.0 370950.0 ;
      RECT  512700.0 369750.0 513900.0 370950.0 ;
      RECT  510300.0 369750.0 511500.0 370950.0 ;
      RECT  509850.0 376350.0 511050.0 377550.0 ;
      RECT  512850.0 354450.0 514050.0 355650.0 ;
      RECT  510300.0 369750.0 511500.0 370950.0 ;
      RECT  512700.0 359250.0 513900.0 360450.0 ;
      RECT  516600.0 357450.0 517800.0 358650.0 ;
      RECT  516600.0 357450.0 517800.0 358650.0 ;
      RECT  523050.0 376500.0 523950.0 377400.0 ;
      RECT  520200.0 376500.0 523500.0 377400.0 ;
      RECT  523050.0 370350.0 523950.0 376950.0 ;
      RECT  520650.0 354600.0 521550.0 355500.0 ;
      RECT  521100.0 354600.0 523650.0 355500.0 ;
      RECT  520650.0 355050.0 521550.0 359850.0 ;
      RECT  520500.0 359250.0 521700.0 360450.0 ;
      RECT  522900.0 359250.0 524100.0 360450.0 ;
      RECT  522900.0 359250.0 524100.0 360450.0 ;
      RECT  520500.0 359250.0 521700.0 360450.0 ;
      RECT  520500.0 369750.0 521700.0 370950.0 ;
      RECT  522900.0 369750.0 524100.0 370950.0 ;
      RECT  522900.0 369750.0 524100.0 370950.0 ;
      RECT  520500.0 369750.0 521700.0 370950.0 ;
      RECT  520050.0 376350.0 521250.0 377550.0 ;
      RECT  523050.0 354450.0 524250.0 355650.0 ;
      RECT  520500.0 369750.0 521700.0 370950.0 ;
      RECT  522900.0 359250.0 524100.0 360450.0 ;
      RECT  526800.0 357450.0 528000.0 358650.0 ;
      RECT  526800.0 357450.0 528000.0 358650.0 ;
      RECT  533250.0 376500.0 534150.0 377400.0 ;
      RECT  530400.0 376500.0 533700.0 377400.0 ;
      RECT  533250.0 370350.0 534150.0 376950.0 ;
      RECT  530850.0 354600.0 531750.0 355500.0 ;
      RECT  531300.0 354600.0 533850.0 355500.0 ;
      RECT  530850.0 355050.0 531750.0 359850.0 ;
      RECT  530700.0 359250.0 531900.0 360450.0 ;
      RECT  533100.0 359250.0 534300.0 360450.0 ;
      RECT  533100.0 359250.0 534300.0 360450.0 ;
      RECT  530700.0 359250.0 531900.0 360450.0 ;
      RECT  530700.0 369750.0 531900.0 370950.0 ;
      RECT  533100.0 369750.0 534300.0 370950.0 ;
      RECT  533100.0 369750.0 534300.0 370950.0 ;
      RECT  530700.0 369750.0 531900.0 370950.0 ;
      RECT  530250.0 376350.0 531450.0 377550.0 ;
      RECT  533250.0 354450.0 534450.0 355650.0 ;
      RECT  530700.0 369750.0 531900.0 370950.0 ;
      RECT  533100.0 359250.0 534300.0 360450.0 ;
      RECT  537000.0 357450.0 538200.0 358650.0 ;
      RECT  537000.0 357450.0 538200.0 358650.0 ;
      RECT  543450.0 376500.0 544350.0 377400.0 ;
      RECT  540600.0 376500.0 543900.0 377400.0 ;
      RECT  543450.0 370350.0 544350.0 376950.0 ;
      RECT  541050.0 354600.0 541950.0 355500.0 ;
      RECT  541500.0 354600.0 544050.0 355500.0 ;
      RECT  541050.0 355050.0 541950.0 359850.0 ;
      RECT  540900.0 359250.0 542100.0 360450.0 ;
      RECT  543300.0 359250.0 544500.0 360450.0 ;
      RECT  543300.0 359250.0 544500.0 360450.0 ;
      RECT  540900.0 359250.0 542100.0 360450.0 ;
      RECT  540900.0 369750.0 542100.0 370950.0 ;
      RECT  543300.0 369750.0 544500.0 370950.0 ;
      RECT  543300.0 369750.0 544500.0 370950.0 ;
      RECT  540900.0 369750.0 542100.0 370950.0 ;
      RECT  540450.0 376350.0 541650.0 377550.0 ;
      RECT  543450.0 354450.0 544650.0 355650.0 ;
      RECT  540900.0 369750.0 542100.0 370950.0 ;
      RECT  543300.0 359250.0 544500.0 360450.0 ;
      RECT  547200.0 357450.0 548400.0 358650.0 ;
      RECT  547200.0 357450.0 548400.0 358650.0 ;
      RECT  553650.0 376500.0 554550.0 377400.0 ;
      RECT  550800.0 376500.0 554100.0 377400.0 ;
      RECT  553650.0 370350.0 554550.0 376950.0 ;
      RECT  551250.0 354600.0 552150.0 355500.0 ;
      RECT  551700.0 354600.0 554250.0 355500.0 ;
      RECT  551250.0 355050.0 552150.0 359850.0 ;
      RECT  551100.0 359250.0 552300.0 360450.0 ;
      RECT  553500.0 359250.0 554700.0 360450.0 ;
      RECT  553500.0 359250.0 554700.0 360450.0 ;
      RECT  551100.0 359250.0 552300.0 360450.0 ;
      RECT  551100.0 369750.0 552300.0 370950.0 ;
      RECT  553500.0 369750.0 554700.0 370950.0 ;
      RECT  553500.0 369750.0 554700.0 370950.0 ;
      RECT  551100.0 369750.0 552300.0 370950.0 ;
      RECT  550650.0 376350.0 551850.0 377550.0 ;
      RECT  553650.0 354450.0 554850.0 355650.0 ;
      RECT  551100.0 369750.0 552300.0 370950.0 ;
      RECT  553500.0 359250.0 554700.0 360450.0 ;
      RECT  557400.0 357450.0 558600.0 358650.0 ;
      RECT  557400.0 357450.0 558600.0 358650.0 ;
      RECT  563850.0 376500.0 564750.0 377400.0 ;
      RECT  561000.0 376500.0 564300.0 377400.0 ;
      RECT  563850.0 370350.0 564750.0 376950.0 ;
      RECT  561450.0 354600.0 562350.0 355500.0 ;
      RECT  561900.0 354600.0 564450.0 355500.0 ;
      RECT  561450.0 355050.0 562350.0 359850.0 ;
      RECT  561300.0 359250.0 562500.0 360450.0 ;
      RECT  563700.0 359250.0 564900.0 360450.0 ;
      RECT  563700.0 359250.0 564900.0 360450.0 ;
      RECT  561300.0 359250.0 562500.0 360450.0 ;
      RECT  561300.0 369750.0 562500.0 370950.0 ;
      RECT  563700.0 369750.0 564900.0 370950.0 ;
      RECT  563700.0 369750.0 564900.0 370950.0 ;
      RECT  561300.0 369750.0 562500.0 370950.0 ;
      RECT  560850.0 376350.0 562050.0 377550.0 ;
      RECT  563850.0 354450.0 565050.0 355650.0 ;
      RECT  561300.0 369750.0 562500.0 370950.0 ;
      RECT  563700.0 359250.0 564900.0 360450.0 ;
      RECT  567600.0 357450.0 568800.0 358650.0 ;
      RECT  567600.0 357450.0 568800.0 358650.0 ;
      RECT  574050.0 376500.0 574950.0 377400.0 ;
      RECT  571200.0 376500.0 574500.0 377400.0 ;
      RECT  574050.0 370350.0 574950.0 376950.0 ;
      RECT  571650.0 354600.0 572550.0 355500.0 ;
      RECT  572100.0 354600.0 574650.0 355500.0 ;
      RECT  571650.0 355050.0 572550.0 359850.0 ;
      RECT  571500.0 359250.0 572700.0 360450.0 ;
      RECT  573900.0 359250.0 575100.0 360450.0 ;
      RECT  573900.0 359250.0 575100.0 360450.0 ;
      RECT  571500.0 359250.0 572700.0 360450.0 ;
      RECT  571500.0 369750.0 572700.0 370950.0 ;
      RECT  573900.0 369750.0 575100.0 370950.0 ;
      RECT  573900.0 369750.0 575100.0 370950.0 ;
      RECT  571500.0 369750.0 572700.0 370950.0 ;
      RECT  571050.0 376350.0 572250.0 377550.0 ;
      RECT  574050.0 354450.0 575250.0 355650.0 ;
      RECT  571500.0 369750.0 572700.0 370950.0 ;
      RECT  573900.0 359250.0 575100.0 360450.0 ;
      RECT  577800.0 357450.0 579000.0 358650.0 ;
      RECT  577800.0 357450.0 579000.0 358650.0 ;
      RECT  584250.0 376500.0 585150.0 377400.0 ;
      RECT  581400.0 376500.0 584700.0 377400.0 ;
      RECT  584250.0 370350.0 585150.0 376950.0 ;
      RECT  581850.0 354600.0 582750.0 355500.0 ;
      RECT  582300.0 354600.0 584850.0 355500.0 ;
      RECT  581850.0 355050.0 582750.0 359850.0 ;
      RECT  581700.0 359250.0 582900.0 360450.0 ;
      RECT  584100.0 359250.0 585300.0 360450.0 ;
      RECT  584100.0 359250.0 585300.0 360450.0 ;
      RECT  581700.0 359250.0 582900.0 360450.0 ;
      RECT  581700.0 369750.0 582900.0 370950.0 ;
      RECT  584100.0 369750.0 585300.0 370950.0 ;
      RECT  584100.0 369750.0 585300.0 370950.0 ;
      RECT  581700.0 369750.0 582900.0 370950.0 ;
      RECT  581250.0 376350.0 582450.0 377550.0 ;
      RECT  584250.0 354450.0 585450.0 355650.0 ;
      RECT  581700.0 369750.0 582900.0 370950.0 ;
      RECT  584100.0 359250.0 585300.0 360450.0 ;
      RECT  588000.0 357450.0 589200.0 358650.0 ;
      RECT  588000.0 357450.0 589200.0 358650.0 ;
      RECT  594450.0 376500.0 595350.0 377400.0 ;
      RECT  591600.0 376500.0 594900.0 377400.0 ;
      RECT  594450.0 370350.0 595350.0 376950.0 ;
      RECT  592050.0 354600.0 592950.0 355500.0 ;
      RECT  592500.0 354600.0 595050.0 355500.0 ;
      RECT  592050.0 355050.0 592950.0 359850.0 ;
      RECT  591900.0 359250.0 593100.0 360450.0 ;
      RECT  594300.0 359250.0 595500.0 360450.0 ;
      RECT  594300.0 359250.0 595500.0 360450.0 ;
      RECT  591900.0 359250.0 593100.0 360450.0 ;
      RECT  591900.0 369750.0 593100.0 370950.0 ;
      RECT  594300.0 369750.0 595500.0 370950.0 ;
      RECT  594300.0 369750.0 595500.0 370950.0 ;
      RECT  591900.0 369750.0 593100.0 370950.0 ;
      RECT  591450.0 376350.0 592650.0 377550.0 ;
      RECT  594450.0 354450.0 595650.0 355650.0 ;
      RECT  591900.0 369750.0 593100.0 370950.0 ;
      RECT  594300.0 359250.0 595500.0 360450.0 ;
      RECT  598200.0 357450.0 599400.0 358650.0 ;
      RECT  598200.0 357450.0 599400.0 358650.0 ;
      RECT  604650.0 376500.0 605550.0 377400.0 ;
      RECT  601800.0 376500.0 605100.0 377400.0 ;
      RECT  604650.0 370350.0 605550.0 376950.0 ;
      RECT  602250.0 354600.0 603150.0 355500.0 ;
      RECT  602700.0 354600.0 605250.0 355500.0 ;
      RECT  602250.0 355050.0 603150.0 359850.0 ;
      RECT  602100.0 359250.0 603300.0 360450.0 ;
      RECT  604500.0 359250.0 605700.0 360450.0 ;
      RECT  604500.0 359250.0 605700.0 360450.0 ;
      RECT  602100.0 359250.0 603300.0 360450.0 ;
      RECT  602100.0 369750.0 603300.0 370950.0 ;
      RECT  604500.0 369750.0 605700.0 370950.0 ;
      RECT  604500.0 369750.0 605700.0 370950.0 ;
      RECT  602100.0 369750.0 603300.0 370950.0 ;
      RECT  601650.0 376350.0 602850.0 377550.0 ;
      RECT  604650.0 354450.0 605850.0 355650.0 ;
      RECT  602100.0 369750.0 603300.0 370950.0 ;
      RECT  604500.0 359250.0 605700.0 360450.0 ;
      RECT  608400.0 357450.0 609600.0 358650.0 ;
      RECT  608400.0 357450.0 609600.0 358650.0 ;
      RECT  614850.0 376500.0 615750.0 377400.0 ;
      RECT  612000.0 376500.0 615300.0 377400.0 ;
      RECT  614850.0 370350.0 615750.0 376950.0 ;
      RECT  612450.0 354600.0 613350.0 355500.0 ;
      RECT  612900.0 354600.0 615450.0 355500.0 ;
      RECT  612450.0 355050.0 613350.0 359850.0 ;
      RECT  612300.0 359250.0 613500.0 360450.0 ;
      RECT  614700.0 359250.0 615900.0 360450.0 ;
      RECT  614700.0 359250.0 615900.0 360450.0 ;
      RECT  612300.0 359250.0 613500.0 360450.0 ;
      RECT  612300.0 369750.0 613500.0 370950.0 ;
      RECT  614700.0 369750.0 615900.0 370950.0 ;
      RECT  614700.0 369750.0 615900.0 370950.0 ;
      RECT  612300.0 369750.0 613500.0 370950.0 ;
      RECT  611850.0 376350.0 613050.0 377550.0 ;
      RECT  614850.0 354450.0 616050.0 355650.0 ;
      RECT  612300.0 369750.0 613500.0 370950.0 ;
      RECT  614700.0 359250.0 615900.0 360450.0 ;
      RECT  618600.0 357450.0 619800.0 358650.0 ;
      RECT  618600.0 357450.0 619800.0 358650.0 ;
      RECT  625050.0 376500.0 625950.0 377400.0 ;
      RECT  622200.0 376500.0 625500.0 377400.0 ;
      RECT  625050.0 370350.0 625950.0 376950.0 ;
      RECT  622650.0 354600.0 623550.0 355500.0 ;
      RECT  623100.0 354600.0 625650.0 355500.0 ;
      RECT  622650.0 355050.0 623550.0 359850.0 ;
      RECT  622500.0 359250.0 623700.0 360450.0 ;
      RECT  624900.0 359250.0 626100.0 360450.0 ;
      RECT  624900.0 359250.0 626100.0 360450.0 ;
      RECT  622500.0 359250.0 623700.0 360450.0 ;
      RECT  622500.0 369750.0 623700.0 370950.0 ;
      RECT  624900.0 369750.0 626100.0 370950.0 ;
      RECT  624900.0 369750.0 626100.0 370950.0 ;
      RECT  622500.0 369750.0 623700.0 370950.0 ;
      RECT  622050.0 376350.0 623250.0 377550.0 ;
      RECT  625050.0 354450.0 626250.0 355650.0 ;
      RECT  622500.0 369750.0 623700.0 370950.0 ;
      RECT  624900.0 359250.0 626100.0 360450.0 ;
      RECT  628800.0 357450.0 630000.0 358650.0 ;
      RECT  628800.0 357450.0 630000.0 358650.0 ;
      RECT  635250.0 376500.0 636150.0 377400.0 ;
      RECT  632400.0 376500.0 635700.0 377400.0 ;
      RECT  635250.0 370350.0 636150.0 376950.0 ;
      RECT  632850.0 354600.0 633750.0 355500.0 ;
      RECT  633300.0 354600.0 635850.0 355500.0 ;
      RECT  632850.0 355050.0 633750.0 359850.0 ;
      RECT  632700.0 359250.0 633900.0 360450.0 ;
      RECT  635100.0 359250.0 636300.0 360450.0 ;
      RECT  635100.0 359250.0 636300.0 360450.0 ;
      RECT  632700.0 359250.0 633900.0 360450.0 ;
      RECT  632700.0 369750.0 633900.0 370950.0 ;
      RECT  635100.0 369750.0 636300.0 370950.0 ;
      RECT  635100.0 369750.0 636300.0 370950.0 ;
      RECT  632700.0 369750.0 633900.0 370950.0 ;
      RECT  632250.0 376350.0 633450.0 377550.0 ;
      RECT  635250.0 354450.0 636450.0 355650.0 ;
      RECT  632700.0 369750.0 633900.0 370950.0 ;
      RECT  635100.0 359250.0 636300.0 360450.0 ;
      RECT  639000.0 357450.0 640200.0 358650.0 ;
      RECT  639000.0 357450.0 640200.0 358650.0 ;
      RECT  645450.0 376500.0 646350.0 377400.0 ;
      RECT  642600.0 376500.0 645900.0 377400.0 ;
      RECT  645450.0 370350.0 646350.0 376950.0 ;
      RECT  643050.0 354600.0 643950.0 355500.0 ;
      RECT  643500.0 354600.0 646050.0 355500.0 ;
      RECT  643050.0 355050.0 643950.0 359850.0 ;
      RECT  642900.0 359250.0 644100.0 360450.0 ;
      RECT  645300.0 359250.0 646500.0 360450.0 ;
      RECT  645300.0 359250.0 646500.0 360450.0 ;
      RECT  642900.0 359250.0 644100.0 360450.0 ;
      RECT  642900.0 369750.0 644100.0 370950.0 ;
      RECT  645300.0 369750.0 646500.0 370950.0 ;
      RECT  645300.0 369750.0 646500.0 370950.0 ;
      RECT  642900.0 369750.0 644100.0 370950.0 ;
      RECT  642450.0 376350.0 643650.0 377550.0 ;
      RECT  645450.0 354450.0 646650.0 355650.0 ;
      RECT  642900.0 369750.0 644100.0 370950.0 ;
      RECT  645300.0 359250.0 646500.0 360450.0 ;
      RECT  649200.0 357450.0 650400.0 358650.0 ;
      RECT  649200.0 357450.0 650400.0 358650.0 ;
      RECT  655650.0 376500.0 656550.0 377400.0 ;
      RECT  652800.0 376500.0 656100.0 377400.0 ;
      RECT  655650.0 370350.0 656550.0 376950.0 ;
      RECT  653250.0 354600.0 654150.0 355500.0 ;
      RECT  653700.0 354600.0 656250.0 355500.0 ;
      RECT  653250.0 355050.0 654150.0 359850.0 ;
      RECT  653100.0 359250.0 654300.0 360450.0 ;
      RECT  655500.0 359250.0 656700.0 360450.0 ;
      RECT  655500.0 359250.0 656700.0 360450.0 ;
      RECT  653100.0 359250.0 654300.0 360450.0 ;
      RECT  653100.0 369750.0 654300.0 370950.0 ;
      RECT  655500.0 369750.0 656700.0 370950.0 ;
      RECT  655500.0 369750.0 656700.0 370950.0 ;
      RECT  653100.0 369750.0 654300.0 370950.0 ;
      RECT  652650.0 376350.0 653850.0 377550.0 ;
      RECT  655650.0 354450.0 656850.0 355650.0 ;
      RECT  653100.0 369750.0 654300.0 370950.0 ;
      RECT  655500.0 359250.0 656700.0 360450.0 ;
      RECT  659400.0 357450.0 660600.0 358650.0 ;
      RECT  659400.0 357450.0 660600.0 358650.0 ;
      RECT  665850.0 376500.0 666750.0 377400.0 ;
      RECT  663000.0 376500.0 666300.0 377400.0 ;
      RECT  665850.0 370350.0 666750.0 376950.0 ;
      RECT  663450.0 354600.0 664350.0 355500.0 ;
      RECT  663900.0 354600.0 666450.0 355500.0 ;
      RECT  663450.0 355050.0 664350.0 359850.0 ;
      RECT  663300.0 359250.0 664500.0 360450.0 ;
      RECT  665700.0 359250.0 666900.0 360450.0 ;
      RECT  665700.0 359250.0 666900.0 360450.0 ;
      RECT  663300.0 359250.0 664500.0 360450.0 ;
      RECT  663300.0 369750.0 664500.0 370950.0 ;
      RECT  665700.0 369750.0 666900.0 370950.0 ;
      RECT  665700.0 369750.0 666900.0 370950.0 ;
      RECT  663300.0 369750.0 664500.0 370950.0 ;
      RECT  662850.0 376350.0 664050.0 377550.0 ;
      RECT  665850.0 354450.0 667050.0 355650.0 ;
      RECT  663300.0 369750.0 664500.0 370950.0 ;
      RECT  665700.0 359250.0 666900.0 360450.0 ;
      RECT  669600.0 357450.0 670800.0 358650.0 ;
      RECT  669600.0 357450.0 670800.0 358650.0 ;
      RECT  676050.0 376500.0 676950.0 377400.0 ;
      RECT  673200.0 376500.0 676500.0 377400.0 ;
      RECT  676050.0 370350.0 676950.0 376950.0 ;
      RECT  673650.0 354600.0 674550.0 355500.0 ;
      RECT  674100.0 354600.0 676650.0 355500.0 ;
      RECT  673650.0 355050.0 674550.0 359850.0 ;
      RECT  673500.0 359250.0 674700.0 360450.0 ;
      RECT  675900.0 359250.0 677100.0 360450.0 ;
      RECT  675900.0 359250.0 677100.0 360450.0 ;
      RECT  673500.0 359250.0 674700.0 360450.0 ;
      RECT  673500.0 369750.0 674700.0 370950.0 ;
      RECT  675900.0 369750.0 677100.0 370950.0 ;
      RECT  675900.0 369750.0 677100.0 370950.0 ;
      RECT  673500.0 369750.0 674700.0 370950.0 ;
      RECT  673050.0 376350.0 674250.0 377550.0 ;
      RECT  676050.0 354450.0 677250.0 355650.0 ;
      RECT  673500.0 369750.0 674700.0 370950.0 ;
      RECT  675900.0 359250.0 677100.0 360450.0 ;
      RECT  679800.0 357450.0 681000.0 358650.0 ;
      RECT  679800.0 357450.0 681000.0 358650.0 ;
      RECT  686250.0 376500.0 687150.0 377400.0 ;
      RECT  683400.0 376500.0 686700.0 377400.0 ;
      RECT  686250.0 370350.0 687150.0 376950.0 ;
      RECT  683850.0 354600.0 684750.0 355500.0 ;
      RECT  684300.0 354600.0 686850.0 355500.0 ;
      RECT  683850.0 355050.0 684750.0 359850.0 ;
      RECT  683700.0 359250.0 684900.0 360450.0 ;
      RECT  686100.0 359250.0 687300.0 360450.0 ;
      RECT  686100.0 359250.0 687300.0 360450.0 ;
      RECT  683700.0 359250.0 684900.0 360450.0 ;
      RECT  683700.0 369750.0 684900.0 370950.0 ;
      RECT  686100.0 369750.0 687300.0 370950.0 ;
      RECT  686100.0 369750.0 687300.0 370950.0 ;
      RECT  683700.0 369750.0 684900.0 370950.0 ;
      RECT  683250.0 376350.0 684450.0 377550.0 ;
      RECT  686250.0 354450.0 687450.0 355650.0 ;
      RECT  683700.0 369750.0 684900.0 370950.0 ;
      RECT  686100.0 359250.0 687300.0 360450.0 ;
      RECT  690000.0 357450.0 691200.0 358650.0 ;
      RECT  690000.0 357450.0 691200.0 358650.0 ;
      RECT  696450.0 376500.0 697350.0 377400.0 ;
      RECT  693600.0 376500.0 696900.0 377400.0 ;
      RECT  696450.0 370350.0 697350.0 376950.0 ;
      RECT  694050.0 354600.0 694950.0 355500.0 ;
      RECT  694500.0 354600.0 697050.0 355500.0 ;
      RECT  694050.0 355050.0 694950.0 359850.0 ;
      RECT  693900.0 359250.0 695100.0 360450.0 ;
      RECT  696300.0 359250.0 697500.0 360450.0 ;
      RECT  696300.0 359250.0 697500.0 360450.0 ;
      RECT  693900.0 359250.0 695100.0 360450.0 ;
      RECT  693900.0 369750.0 695100.0 370950.0 ;
      RECT  696300.0 369750.0 697500.0 370950.0 ;
      RECT  696300.0 369750.0 697500.0 370950.0 ;
      RECT  693900.0 369750.0 695100.0 370950.0 ;
      RECT  693450.0 376350.0 694650.0 377550.0 ;
      RECT  696450.0 354450.0 697650.0 355650.0 ;
      RECT  693900.0 369750.0 695100.0 370950.0 ;
      RECT  696300.0 359250.0 697500.0 360450.0 ;
      RECT  700200.0 357450.0 701400.0 358650.0 ;
      RECT  700200.0 357450.0 701400.0 358650.0 ;
      RECT  706650.0 376500.0 707550.0 377400.0 ;
      RECT  703800.0 376500.0 707100.0 377400.0 ;
      RECT  706650.0 370350.0 707550.0 376950.0 ;
      RECT  704250.0 354600.0 705150.0 355500.0 ;
      RECT  704700.0 354600.0 707250.0 355500.0 ;
      RECT  704250.0 355050.0 705150.0 359850.0 ;
      RECT  704100.0 359250.0 705300.0 360450.0 ;
      RECT  706500.0 359250.0 707700.0 360450.0 ;
      RECT  706500.0 359250.0 707700.0 360450.0 ;
      RECT  704100.0 359250.0 705300.0 360450.0 ;
      RECT  704100.0 369750.0 705300.0 370950.0 ;
      RECT  706500.0 369750.0 707700.0 370950.0 ;
      RECT  706500.0 369750.0 707700.0 370950.0 ;
      RECT  704100.0 369750.0 705300.0 370950.0 ;
      RECT  703650.0 376350.0 704850.0 377550.0 ;
      RECT  706650.0 354450.0 707850.0 355650.0 ;
      RECT  704100.0 369750.0 705300.0 370950.0 ;
      RECT  706500.0 359250.0 707700.0 360450.0 ;
      RECT  710400.0 357450.0 711600.0 358650.0 ;
      RECT  710400.0 357450.0 711600.0 358650.0 ;
      RECT  716850.0 376500.0 717750.0 377400.0 ;
      RECT  714000.0 376500.0 717300.0 377400.0 ;
      RECT  716850.0 370350.0 717750.0 376950.0 ;
      RECT  714450.0 354600.0 715350.0 355500.0 ;
      RECT  714900.0 354600.0 717450.0 355500.0 ;
      RECT  714450.0 355050.0 715350.0 359850.0 ;
      RECT  714300.0 359250.0 715500.0 360450.0 ;
      RECT  716700.0 359250.0 717900.0 360450.0 ;
      RECT  716700.0 359250.0 717900.0 360450.0 ;
      RECT  714300.0 359250.0 715500.0 360450.0 ;
      RECT  714300.0 369750.0 715500.0 370950.0 ;
      RECT  716700.0 369750.0 717900.0 370950.0 ;
      RECT  716700.0 369750.0 717900.0 370950.0 ;
      RECT  714300.0 369750.0 715500.0 370950.0 ;
      RECT  713850.0 376350.0 715050.0 377550.0 ;
      RECT  716850.0 354450.0 718050.0 355650.0 ;
      RECT  714300.0 369750.0 715500.0 370950.0 ;
      RECT  716700.0 359250.0 717900.0 360450.0 ;
      RECT  720600.0 357450.0 721800.0 358650.0 ;
      RECT  720600.0 357450.0 721800.0 358650.0 ;
      RECT  727050.0 376500.0 727950.0 377400.0 ;
      RECT  724200.0 376500.0 727500.0 377400.0 ;
      RECT  727050.0 370350.0 727950.0 376950.0 ;
      RECT  724650.0 354600.0 725550.0 355500.0 ;
      RECT  725100.0 354600.0 727650.0 355500.0 ;
      RECT  724650.0 355050.0 725550.0 359850.0 ;
      RECT  724500.0 359250.0 725700.0 360450.0 ;
      RECT  726900.0 359250.0 728100.0 360450.0 ;
      RECT  726900.0 359250.0 728100.0 360450.0 ;
      RECT  724500.0 359250.0 725700.0 360450.0 ;
      RECT  724500.0 369750.0 725700.0 370950.0 ;
      RECT  726900.0 369750.0 728100.0 370950.0 ;
      RECT  726900.0 369750.0 728100.0 370950.0 ;
      RECT  724500.0 369750.0 725700.0 370950.0 ;
      RECT  724050.0 376350.0 725250.0 377550.0 ;
      RECT  727050.0 354450.0 728250.0 355650.0 ;
      RECT  724500.0 369750.0 725700.0 370950.0 ;
      RECT  726900.0 359250.0 728100.0 360450.0 ;
      RECT  730800.0 357450.0 732000.0 358650.0 ;
      RECT  730800.0 357450.0 732000.0 358650.0 ;
      RECT  737250.0 376500.0 738150.0 377400.0 ;
      RECT  734400.0 376500.0 737700.0 377400.0 ;
      RECT  737250.0 370350.0 738150.0 376950.0 ;
      RECT  734850.0 354600.0 735750.0 355500.0 ;
      RECT  735300.0 354600.0 737850.0 355500.0 ;
      RECT  734850.0 355050.0 735750.0 359850.0 ;
      RECT  734700.0 359250.0 735900.0 360450.0 ;
      RECT  737100.0 359250.0 738300.0 360450.0 ;
      RECT  737100.0 359250.0 738300.0 360450.0 ;
      RECT  734700.0 359250.0 735900.0 360450.0 ;
      RECT  734700.0 369750.0 735900.0 370950.0 ;
      RECT  737100.0 369750.0 738300.0 370950.0 ;
      RECT  737100.0 369750.0 738300.0 370950.0 ;
      RECT  734700.0 369750.0 735900.0 370950.0 ;
      RECT  734250.0 376350.0 735450.0 377550.0 ;
      RECT  737250.0 354450.0 738450.0 355650.0 ;
      RECT  734700.0 369750.0 735900.0 370950.0 ;
      RECT  737100.0 359250.0 738300.0 360450.0 ;
      RECT  741000.0 357450.0 742200.0 358650.0 ;
      RECT  741000.0 357450.0 742200.0 358650.0 ;
      RECT  747450.0 376500.0 748350.0 377400.0 ;
      RECT  744600.0 376500.0 747900.0 377400.0 ;
      RECT  747450.0 370350.0 748350.0 376950.0 ;
      RECT  745050.0 354600.0 745950.0 355500.0 ;
      RECT  745500.0 354600.0 748050.0 355500.0 ;
      RECT  745050.0 355050.0 745950.0 359850.0 ;
      RECT  744900.0 359250.0 746100.0 360450.0 ;
      RECT  747300.0 359250.0 748500.0 360450.0 ;
      RECT  747300.0 359250.0 748500.0 360450.0 ;
      RECT  744900.0 359250.0 746100.0 360450.0 ;
      RECT  744900.0 369750.0 746100.0 370950.0 ;
      RECT  747300.0 369750.0 748500.0 370950.0 ;
      RECT  747300.0 369750.0 748500.0 370950.0 ;
      RECT  744900.0 369750.0 746100.0 370950.0 ;
      RECT  744450.0 376350.0 745650.0 377550.0 ;
      RECT  747450.0 354450.0 748650.0 355650.0 ;
      RECT  744900.0 369750.0 746100.0 370950.0 ;
      RECT  747300.0 359250.0 748500.0 360450.0 ;
      RECT  751200.0 357450.0 752400.0 358650.0 ;
      RECT  751200.0 357450.0 752400.0 358650.0 ;
      RECT  757650.0 376500.0 758550.0 377400.0 ;
      RECT  754800.0 376500.0 758100.0 377400.0 ;
      RECT  757650.0 370350.0 758550.0 376950.0 ;
      RECT  755250.0 354600.0 756150.0 355500.0 ;
      RECT  755700.0 354600.0 758250.0 355500.0 ;
      RECT  755250.0 355050.0 756150.0 359850.0 ;
      RECT  755100.0 359250.0 756300.0 360450.0 ;
      RECT  757500.0 359250.0 758700.0 360450.0 ;
      RECT  757500.0 359250.0 758700.0 360450.0 ;
      RECT  755100.0 359250.0 756300.0 360450.0 ;
      RECT  755100.0 369750.0 756300.0 370950.0 ;
      RECT  757500.0 369750.0 758700.0 370950.0 ;
      RECT  757500.0 369750.0 758700.0 370950.0 ;
      RECT  755100.0 369750.0 756300.0 370950.0 ;
      RECT  754650.0 376350.0 755850.0 377550.0 ;
      RECT  757650.0 354450.0 758850.0 355650.0 ;
      RECT  755100.0 369750.0 756300.0 370950.0 ;
      RECT  757500.0 359250.0 758700.0 360450.0 ;
      RECT  761400.0 357450.0 762600.0 358650.0 ;
      RECT  761400.0 357450.0 762600.0 358650.0 ;
      RECT  767850.0 376500.0 768750.0 377400.0 ;
      RECT  765000.0 376500.0 768300.0 377400.0 ;
      RECT  767850.0 370350.0 768750.0 376950.0 ;
      RECT  765450.0 354600.0 766350.0 355500.0 ;
      RECT  765900.0 354600.0 768450.0 355500.0 ;
      RECT  765450.0 355050.0 766350.0 359850.0 ;
      RECT  765300.0 359250.0 766500.0 360450.0 ;
      RECT  767700.0 359250.0 768900.0 360450.0 ;
      RECT  767700.0 359250.0 768900.0 360450.0 ;
      RECT  765300.0 359250.0 766500.0 360450.0 ;
      RECT  765300.0 369750.0 766500.0 370950.0 ;
      RECT  767700.0 369750.0 768900.0 370950.0 ;
      RECT  767700.0 369750.0 768900.0 370950.0 ;
      RECT  765300.0 369750.0 766500.0 370950.0 ;
      RECT  764850.0 376350.0 766050.0 377550.0 ;
      RECT  767850.0 354450.0 769050.0 355650.0 ;
      RECT  765300.0 369750.0 766500.0 370950.0 ;
      RECT  767700.0 359250.0 768900.0 360450.0 ;
      RECT  771600.0 357450.0 772800.0 358650.0 ;
      RECT  771600.0 357450.0 772800.0 358650.0 ;
      RECT  778050.0 376500.0 778950.0 377400.0 ;
      RECT  775200.0 376500.0 778500.0 377400.0 ;
      RECT  778050.0 370350.0 778950.0 376950.0 ;
      RECT  775650.0 354600.0 776550.0 355500.0 ;
      RECT  776100.0 354600.0 778650.0 355500.0 ;
      RECT  775650.0 355050.0 776550.0 359850.0 ;
      RECT  775500.0 359250.0 776700.0 360450.0 ;
      RECT  777900.0 359250.0 779100.0 360450.0 ;
      RECT  777900.0 359250.0 779100.0 360450.0 ;
      RECT  775500.0 359250.0 776700.0 360450.0 ;
      RECT  775500.0 369750.0 776700.0 370950.0 ;
      RECT  777900.0 369750.0 779100.0 370950.0 ;
      RECT  777900.0 369750.0 779100.0 370950.0 ;
      RECT  775500.0 369750.0 776700.0 370950.0 ;
      RECT  775050.0 376350.0 776250.0 377550.0 ;
      RECT  778050.0 354450.0 779250.0 355650.0 ;
      RECT  775500.0 369750.0 776700.0 370950.0 ;
      RECT  777900.0 359250.0 779100.0 360450.0 ;
      RECT  781800.0 357450.0 783000.0 358650.0 ;
      RECT  781800.0 357450.0 783000.0 358650.0 ;
      RECT  788250.0 376500.0 789150.0 377400.0 ;
      RECT  785400.0 376500.0 788700.0 377400.0 ;
      RECT  788250.0 370350.0 789150.0 376950.0 ;
      RECT  785850.0 354600.0 786750.0 355500.0 ;
      RECT  786300.0 354600.0 788850.0 355500.0 ;
      RECT  785850.0 355050.0 786750.0 359850.0 ;
      RECT  785700.0 359250.0 786900.0 360450.0 ;
      RECT  788100.0 359250.0 789300.0 360450.0 ;
      RECT  788100.0 359250.0 789300.0 360450.0 ;
      RECT  785700.0 359250.0 786900.0 360450.0 ;
      RECT  785700.0 369750.0 786900.0 370950.0 ;
      RECT  788100.0 369750.0 789300.0 370950.0 ;
      RECT  788100.0 369750.0 789300.0 370950.0 ;
      RECT  785700.0 369750.0 786900.0 370950.0 ;
      RECT  785250.0 376350.0 786450.0 377550.0 ;
      RECT  788250.0 354450.0 789450.0 355650.0 ;
      RECT  785700.0 369750.0 786900.0 370950.0 ;
      RECT  788100.0 359250.0 789300.0 360450.0 ;
      RECT  792000.0 357450.0 793200.0 358650.0 ;
      RECT  792000.0 357450.0 793200.0 358650.0 ;
      RECT  798450.0 376500.0 799350.0 377400.0 ;
      RECT  795600.0 376500.0 798900.0 377400.0 ;
      RECT  798450.0 370350.0 799350.0 376950.0 ;
      RECT  796050.0 354600.0 796950.0 355500.0 ;
      RECT  796500.0 354600.0 799050.0 355500.0 ;
      RECT  796050.0 355050.0 796950.0 359850.0 ;
      RECT  795900.0 359250.0 797100.0 360450.0 ;
      RECT  798300.0 359250.0 799500.0 360450.0 ;
      RECT  798300.0 359250.0 799500.0 360450.0 ;
      RECT  795900.0 359250.0 797100.0 360450.0 ;
      RECT  795900.0 369750.0 797100.0 370950.0 ;
      RECT  798300.0 369750.0 799500.0 370950.0 ;
      RECT  798300.0 369750.0 799500.0 370950.0 ;
      RECT  795900.0 369750.0 797100.0 370950.0 ;
      RECT  795450.0 376350.0 796650.0 377550.0 ;
      RECT  798450.0 354450.0 799650.0 355650.0 ;
      RECT  795900.0 369750.0 797100.0 370950.0 ;
      RECT  798300.0 359250.0 799500.0 360450.0 ;
      RECT  802200.0 357450.0 803400.0 358650.0 ;
      RECT  802200.0 357450.0 803400.0 358650.0 ;
      RECT  808650.0 376500.0 809550.0 377400.0 ;
      RECT  805800.0 376500.0 809100.0 377400.0 ;
      RECT  808650.0 370350.0 809550.0 376950.0 ;
      RECT  806250.0 354600.0 807150.0 355500.0 ;
      RECT  806700.0 354600.0 809250.0 355500.0 ;
      RECT  806250.0 355050.0 807150.0 359850.0 ;
      RECT  806100.0 359250.0 807300.0 360450.0 ;
      RECT  808500.0 359250.0 809700.0 360450.0 ;
      RECT  808500.0 359250.0 809700.0 360450.0 ;
      RECT  806100.0 359250.0 807300.0 360450.0 ;
      RECT  806100.0 369750.0 807300.0 370950.0 ;
      RECT  808500.0 369750.0 809700.0 370950.0 ;
      RECT  808500.0 369750.0 809700.0 370950.0 ;
      RECT  806100.0 369750.0 807300.0 370950.0 ;
      RECT  805650.0 376350.0 806850.0 377550.0 ;
      RECT  808650.0 354450.0 809850.0 355650.0 ;
      RECT  806100.0 369750.0 807300.0 370950.0 ;
      RECT  808500.0 359250.0 809700.0 360450.0 ;
      RECT  812400.0 357450.0 813600.0 358650.0 ;
      RECT  812400.0 357450.0 813600.0 358650.0 ;
      RECT  818850.0 376500.0 819750.0 377400.0 ;
      RECT  816000.0 376500.0 819300.0 377400.0 ;
      RECT  818850.0 370350.0 819750.0 376950.0 ;
      RECT  816450.0 354600.0 817350.0 355500.0 ;
      RECT  816900.0 354600.0 819450.0 355500.0 ;
      RECT  816450.0 355050.0 817350.0 359850.0 ;
      RECT  816300.0 359250.0 817500.0 360450.0 ;
      RECT  818700.0 359250.0 819900.0 360450.0 ;
      RECT  818700.0 359250.0 819900.0 360450.0 ;
      RECT  816300.0 359250.0 817500.0 360450.0 ;
      RECT  816300.0 369750.0 817500.0 370950.0 ;
      RECT  818700.0 369750.0 819900.0 370950.0 ;
      RECT  818700.0 369750.0 819900.0 370950.0 ;
      RECT  816300.0 369750.0 817500.0 370950.0 ;
      RECT  815850.0 376350.0 817050.0 377550.0 ;
      RECT  818850.0 354450.0 820050.0 355650.0 ;
      RECT  816300.0 369750.0 817500.0 370950.0 ;
      RECT  818700.0 359250.0 819900.0 360450.0 ;
      RECT  822600.0 357450.0 823800.0 358650.0 ;
      RECT  822600.0 357450.0 823800.0 358650.0 ;
      RECT  829050.0 376500.0 829950.0 377400.0 ;
      RECT  826200.0 376500.0 829500.0 377400.0 ;
      RECT  829050.0 370350.0 829950.0 376950.0 ;
      RECT  826650.0 354600.0 827550.0 355500.0 ;
      RECT  827100.0 354600.0 829650.0 355500.0 ;
      RECT  826650.0 355050.0 827550.0 359850.0 ;
      RECT  826500.0 359250.0 827700.0 360450.0 ;
      RECT  828900.0 359250.0 830100.0 360450.0 ;
      RECT  828900.0 359250.0 830100.0 360450.0 ;
      RECT  826500.0 359250.0 827700.0 360450.0 ;
      RECT  826500.0 369750.0 827700.0 370950.0 ;
      RECT  828900.0 369750.0 830100.0 370950.0 ;
      RECT  828900.0 369750.0 830100.0 370950.0 ;
      RECT  826500.0 369750.0 827700.0 370950.0 ;
      RECT  826050.0 376350.0 827250.0 377550.0 ;
      RECT  829050.0 354450.0 830250.0 355650.0 ;
      RECT  826500.0 369750.0 827700.0 370950.0 ;
      RECT  828900.0 359250.0 830100.0 360450.0 ;
      RECT  832800.0 357450.0 834000.0 358650.0 ;
      RECT  832800.0 357450.0 834000.0 358650.0 ;
      RECT  839250.0 376500.0 840150.0 377400.0 ;
      RECT  836400.0 376500.0 839700.0 377400.0 ;
      RECT  839250.0 370350.0 840150.0 376950.0 ;
      RECT  836850.0 354600.0 837750.0 355500.0 ;
      RECT  837300.0 354600.0 839850.0 355500.0 ;
      RECT  836850.0 355050.0 837750.0 359850.0 ;
      RECT  836700.0 359250.0 837900.0 360450.0 ;
      RECT  839100.0 359250.0 840300.0 360450.0 ;
      RECT  839100.0 359250.0 840300.0 360450.0 ;
      RECT  836700.0 359250.0 837900.0 360450.0 ;
      RECT  836700.0 369750.0 837900.0 370950.0 ;
      RECT  839100.0 369750.0 840300.0 370950.0 ;
      RECT  839100.0 369750.0 840300.0 370950.0 ;
      RECT  836700.0 369750.0 837900.0 370950.0 ;
      RECT  836250.0 376350.0 837450.0 377550.0 ;
      RECT  839250.0 354450.0 840450.0 355650.0 ;
      RECT  836700.0 369750.0 837900.0 370950.0 ;
      RECT  839100.0 359250.0 840300.0 360450.0 ;
      RECT  843000.0 357450.0 844200.0 358650.0 ;
      RECT  843000.0 357450.0 844200.0 358650.0 ;
      RECT  849450.0 376500.0 850350.0 377400.0 ;
      RECT  846600.0 376500.0 849900.0 377400.0 ;
      RECT  849450.0 370350.0 850350.0 376950.0 ;
      RECT  847050.0 354600.0 847950.0 355500.0 ;
      RECT  847500.0 354600.0 850050.0 355500.0 ;
      RECT  847050.0 355050.0 847950.0 359850.0 ;
      RECT  846900.0 359250.0 848100.0 360450.0 ;
      RECT  849300.0 359250.0 850500.0 360450.0 ;
      RECT  849300.0 359250.0 850500.0 360450.0 ;
      RECT  846900.0 359250.0 848100.0 360450.0 ;
      RECT  846900.0 369750.0 848100.0 370950.0 ;
      RECT  849300.0 369750.0 850500.0 370950.0 ;
      RECT  849300.0 369750.0 850500.0 370950.0 ;
      RECT  846900.0 369750.0 848100.0 370950.0 ;
      RECT  846450.0 376350.0 847650.0 377550.0 ;
      RECT  849450.0 354450.0 850650.0 355650.0 ;
      RECT  846900.0 369750.0 848100.0 370950.0 ;
      RECT  849300.0 359250.0 850500.0 360450.0 ;
      RECT  853200.0 357450.0 854400.0 358650.0 ;
      RECT  853200.0 357450.0 854400.0 358650.0 ;
      RECT  859650.0 376500.0 860550.0 377400.0 ;
      RECT  856800.0 376500.0 860100.0 377400.0 ;
      RECT  859650.0 370350.0 860550.0 376950.0 ;
      RECT  857250.0 354600.0 858150.0 355500.0 ;
      RECT  857700.0 354600.0 860250.0 355500.0 ;
      RECT  857250.0 355050.0 858150.0 359850.0 ;
      RECT  857100.0 359250.0 858300.0 360450.0 ;
      RECT  859500.0 359250.0 860700.0 360450.0 ;
      RECT  859500.0 359250.0 860700.0 360450.0 ;
      RECT  857100.0 359250.0 858300.0 360450.0 ;
      RECT  857100.0 369750.0 858300.0 370950.0 ;
      RECT  859500.0 369750.0 860700.0 370950.0 ;
      RECT  859500.0 369750.0 860700.0 370950.0 ;
      RECT  857100.0 369750.0 858300.0 370950.0 ;
      RECT  856650.0 376350.0 857850.0 377550.0 ;
      RECT  859650.0 354450.0 860850.0 355650.0 ;
      RECT  857100.0 369750.0 858300.0 370950.0 ;
      RECT  859500.0 359250.0 860700.0 360450.0 ;
      RECT  863400.0 357450.0 864600.0 358650.0 ;
      RECT  863400.0 357450.0 864600.0 358650.0 ;
      RECT  869850.0 376500.0 870750.0 377400.0 ;
      RECT  867000.0 376500.0 870300.0 377400.0 ;
      RECT  869850.0 370350.0 870750.0 376950.0 ;
      RECT  867450.0 354600.0 868350.0 355500.0 ;
      RECT  867900.0 354600.0 870450.0 355500.0 ;
      RECT  867450.0 355050.0 868350.0 359850.0 ;
      RECT  867300.0 359250.0 868500.0 360450.0 ;
      RECT  869700.0 359250.0 870900.0 360450.0 ;
      RECT  869700.0 359250.0 870900.0 360450.0 ;
      RECT  867300.0 359250.0 868500.0 360450.0 ;
      RECT  867300.0 369750.0 868500.0 370950.0 ;
      RECT  869700.0 369750.0 870900.0 370950.0 ;
      RECT  869700.0 369750.0 870900.0 370950.0 ;
      RECT  867300.0 369750.0 868500.0 370950.0 ;
      RECT  866850.0 376350.0 868050.0 377550.0 ;
      RECT  869850.0 354450.0 871050.0 355650.0 ;
      RECT  867300.0 369750.0 868500.0 370950.0 ;
      RECT  869700.0 359250.0 870900.0 360450.0 ;
      RECT  873600.0 357450.0 874800.0 358650.0 ;
      RECT  873600.0 357450.0 874800.0 358650.0 ;
      RECT  880050.0 376500.0 880950.0 377400.0 ;
      RECT  877200.0 376500.0 880500.0 377400.0 ;
      RECT  880050.0 370350.0 880950.0 376950.0 ;
      RECT  877650.0 354600.0 878550.0 355500.0 ;
      RECT  878100.0 354600.0 880650.0 355500.0 ;
      RECT  877650.0 355050.0 878550.0 359850.0 ;
      RECT  877500.0 359250.0 878700.0 360450.0 ;
      RECT  879900.0 359250.0 881100.0 360450.0 ;
      RECT  879900.0 359250.0 881100.0 360450.0 ;
      RECT  877500.0 359250.0 878700.0 360450.0 ;
      RECT  877500.0 369750.0 878700.0 370950.0 ;
      RECT  879900.0 369750.0 881100.0 370950.0 ;
      RECT  879900.0 369750.0 881100.0 370950.0 ;
      RECT  877500.0 369750.0 878700.0 370950.0 ;
      RECT  877050.0 376350.0 878250.0 377550.0 ;
      RECT  880050.0 354450.0 881250.0 355650.0 ;
      RECT  877500.0 369750.0 878700.0 370950.0 ;
      RECT  879900.0 359250.0 881100.0 360450.0 ;
      RECT  883800.0 357450.0 885000.0 358650.0 ;
      RECT  883800.0 357450.0 885000.0 358650.0 ;
      RECT  890250.0 376500.0 891150.0 377400.0 ;
      RECT  887400.0 376500.0 890700.0 377400.0 ;
      RECT  890250.0 370350.0 891150.0 376950.0 ;
      RECT  887850.0 354600.0 888750.0 355500.0 ;
      RECT  888300.0 354600.0 890850.0 355500.0 ;
      RECT  887850.0 355050.0 888750.0 359850.0 ;
      RECT  887700.0 359250.0 888900.0 360450.0 ;
      RECT  890100.0 359250.0 891300.0 360450.0 ;
      RECT  890100.0 359250.0 891300.0 360450.0 ;
      RECT  887700.0 359250.0 888900.0 360450.0 ;
      RECT  887700.0 369750.0 888900.0 370950.0 ;
      RECT  890100.0 369750.0 891300.0 370950.0 ;
      RECT  890100.0 369750.0 891300.0 370950.0 ;
      RECT  887700.0 369750.0 888900.0 370950.0 ;
      RECT  887250.0 376350.0 888450.0 377550.0 ;
      RECT  890250.0 354450.0 891450.0 355650.0 ;
      RECT  887700.0 369750.0 888900.0 370950.0 ;
      RECT  890100.0 359250.0 891300.0 360450.0 ;
      RECT  894000.0 357450.0 895200.0 358650.0 ;
      RECT  894000.0 357450.0 895200.0 358650.0 ;
      RECT  900450.0 376500.0 901350.0 377400.0 ;
      RECT  897600.0 376500.0 900900.0 377400.0 ;
      RECT  900450.0 370350.0 901350.0 376950.0 ;
      RECT  898050.0 354600.0 898950.0 355500.0 ;
      RECT  898500.0 354600.0 901050.0 355500.0 ;
      RECT  898050.0 355050.0 898950.0 359850.0 ;
      RECT  897900.0 359250.0 899100.0 360450.0 ;
      RECT  900300.0 359250.0 901500.0 360450.0 ;
      RECT  900300.0 359250.0 901500.0 360450.0 ;
      RECT  897900.0 359250.0 899100.0 360450.0 ;
      RECT  897900.0 369750.0 899100.0 370950.0 ;
      RECT  900300.0 369750.0 901500.0 370950.0 ;
      RECT  900300.0 369750.0 901500.0 370950.0 ;
      RECT  897900.0 369750.0 899100.0 370950.0 ;
      RECT  897450.0 376350.0 898650.0 377550.0 ;
      RECT  900450.0 354450.0 901650.0 355650.0 ;
      RECT  897900.0 369750.0 899100.0 370950.0 ;
      RECT  900300.0 359250.0 901500.0 360450.0 ;
      RECT  904200.0 357450.0 905400.0 358650.0 ;
      RECT  904200.0 357450.0 905400.0 358650.0 ;
      RECT  910650.0 376500.0 911550.0 377400.0 ;
      RECT  907800.0 376500.0 911100.0 377400.0 ;
      RECT  910650.0 370350.0 911550.0 376950.0 ;
      RECT  908250.0 354600.0 909150.0 355500.0 ;
      RECT  908700.0 354600.0 911250.0 355500.0 ;
      RECT  908250.0 355050.0 909150.0 359850.0 ;
      RECT  908100.0 359250.0 909300.0 360450.0 ;
      RECT  910500.0 359250.0 911700.0 360450.0 ;
      RECT  910500.0 359250.0 911700.0 360450.0 ;
      RECT  908100.0 359250.0 909300.0 360450.0 ;
      RECT  908100.0 369750.0 909300.0 370950.0 ;
      RECT  910500.0 369750.0 911700.0 370950.0 ;
      RECT  910500.0 369750.0 911700.0 370950.0 ;
      RECT  908100.0 369750.0 909300.0 370950.0 ;
      RECT  907650.0 376350.0 908850.0 377550.0 ;
      RECT  910650.0 354450.0 911850.0 355650.0 ;
      RECT  908100.0 369750.0 909300.0 370950.0 ;
      RECT  910500.0 359250.0 911700.0 360450.0 ;
      RECT  914400.0 357450.0 915600.0 358650.0 ;
      RECT  914400.0 357450.0 915600.0 358650.0 ;
      RECT  920850.0 376500.0 921750.0 377400.0 ;
      RECT  918000.0 376500.0 921300.0 377400.0 ;
      RECT  920850.0 370350.0 921750.0 376950.0 ;
      RECT  918450.0 354600.0 919350.0 355500.0 ;
      RECT  918900.0 354600.0 921450.0 355500.0 ;
      RECT  918450.0 355050.0 919350.0 359850.0 ;
      RECT  918300.0 359250.0 919500.0 360450.0 ;
      RECT  920700.0 359250.0 921900.0 360450.0 ;
      RECT  920700.0 359250.0 921900.0 360450.0 ;
      RECT  918300.0 359250.0 919500.0 360450.0 ;
      RECT  918300.0 369750.0 919500.0 370950.0 ;
      RECT  920700.0 369750.0 921900.0 370950.0 ;
      RECT  920700.0 369750.0 921900.0 370950.0 ;
      RECT  918300.0 369750.0 919500.0 370950.0 ;
      RECT  917850.0 376350.0 919050.0 377550.0 ;
      RECT  920850.0 354450.0 922050.0 355650.0 ;
      RECT  918300.0 369750.0 919500.0 370950.0 ;
      RECT  920700.0 359250.0 921900.0 360450.0 ;
      RECT  924600.0 357450.0 925800.0 358650.0 ;
      RECT  924600.0 357450.0 925800.0 358650.0 ;
      RECT  931050.0 376500.0 931950.0 377400.0 ;
      RECT  928200.0 376500.0 931500.0 377400.0 ;
      RECT  931050.0 370350.0 931950.0 376950.0 ;
      RECT  928650.0 354600.0 929550.0 355500.0 ;
      RECT  929100.0 354600.0 931650.0 355500.0 ;
      RECT  928650.0 355050.0 929550.0 359850.0 ;
      RECT  928500.0 359250.0 929700.0 360450.0 ;
      RECT  930900.0 359250.0 932100.0 360450.0 ;
      RECT  930900.0 359250.0 932100.0 360450.0 ;
      RECT  928500.0 359250.0 929700.0 360450.0 ;
      RECT  928500.0 369750.0 929700.0 370950.0 ;
      RECT  930900.0 369750.0 932100.0 370950.0 ;
      RECT  930900.0 369750.0 932100.0 370950.0 ;
      RECT  928500.0 369750.0 929700.0 370950.0 ;
      RECT  928050.0 376350.0 929250.0 377550.0 ;
      RECT  931050.0 354450.0 932250.0 355650.0 ;
      RECT  928500.0 369750.0 929700.0 370950.0 ;
      RECT  930900.0 359250.0 932100.0 360450.0 ;
      RECT  934800.0 357450.0 936000.0 358650.0 ;
      RECT  934800.0 357450.0 936000.0 358650.0 ;
      RECT  941250.0 376500.0 942150.0 377400.0 ;
      RECT  938400.0 376500.0 941700.0 377400.0 ;
      RECT  941250.0 370350.0 942150.0 376950.0 ;
      RECT  938850.0 354600.0 939750.0 355500.0 ;
      RECT  939300.0 354600.0 941850.0 355500.0 ;
      RECT  938850.0 355050.0 939750.0 359850.0 ;
      RECT  938700.0 359250.0 939900.0 360450.0 ;
      RECT  941100.0 359250.0 942300.0 360450.0 ;
      RECT  941100.0 359250.0 942300.0 360450.0 ;
      RECT  938700.0 359250.0 939900.0 360450.0 ;
      RECT  938700.0 369750.0 939900.0 370950.0 ;
      RECT  941100.0 369750.0 942300.0 370950.0 ;
      RECT  941100.0 369750.0 942300.0 370950.0 ;
      RECT  938700.0 369750.0 939900.0 370950.0 ;
      RECT  938250.0 376350.0 939450.0 377550.0 ;
      RECT  941250.0 354450.0 942450.0 355650.0 ;
      RECT  938700.0 369750.0 939900.0 370950.0 ;
      RECT  941100.0 359250.0 942300.0 360450.0 ;
      RECT  945000.0 357450.0 946200.0 358650.0 ;
      RECT  945000.0 357450.0 946200.0 358650.0 ;
      RECT  951450.0 376500.0 952350.0 377400.0 ;
      RECT  948600.0 376500.0 951900.0 377400.0 ;
      RECT  951450.0 370350.0 952350.0 376950.0 ;
      RECT  949050.0 354600.0 949950.0 355500.0 ;
      RECT  949500.0 354600.0 952050.0 355500.0 ;
      RECT  949050.0 355050.0 949950.0 359850.0 ;
      RECT  948900.0 359250.0 950100.0 360450.0 ;
      RECT  951300.0 359250.0 952500.0 360450.0 ;
      RECT  951300.0 359250.0 952500.0 360450.0 ;
      RECT  948900.0 359250.0 950100.0 360450.0 ;
      RECT  948900.0 369750.0 950100.0 370950.0 ;
      RECT  951300.0 369750.0 952500.0 370950.0 ;
      RECT  951300.0 369750.0 952500.0 370950.0 ;
      RECT  948900.0 369750.0 950100.0 370950.0 ;
      RECT  948450.0 376350.0 949650.0 377550.0 ;
      RECT  951450.0 354450.0 952650.0 355650.0 ;
      RECT  948900.0 369750.0 950100.0 370950.0 ;
      RECT  951300.0 359250.0 952500.0 360450.0 ;
      RECT  955200.0 357450.0 956400.0 358650.0 ;
      RECT  955200.0 357450.0 956400.0 358650.0 ;
      RECT  961650.0 376500.0 962550.0 377400.0 ;
      RECT  958800.0 376500.0 962100.0 377400.0 ;
      RECT  961650.0 370350.0 962550.0 376950.0 ;
      RECT  959250.0 354600.0 960150.0 355500.0 ;
      RECT  959700.0 354600.0 962250.0 355500.0 ;
      RECT  959250.0 355050.0 960150.0 359850.0 ;
      RECT  959100.0 359250.0 960300.0 360450.0 ;
      RECT  961500.0 359250.0 962700.0 360450.0 ;
      RECT  961500.0 359250.0 962700.0 360450.0 ;
      RECT  959100.0 359250.0 960300.0 360450.0 ;
      RECT  959100.0 369750.0 960300.0 370950.0 ;
      RECT  961500.0 369750.0 962700.0 370950.0 ;
      RECT  961500.0 369750.0 962700.0 370950.0 ;
      RECT  959100.0 369750.0 960300.0 370950.0 ;
      RECT  958650.0 376350.0 959850.0 377550.0 ;
      RECT  961650.0 354450.0 962850.0 355650.0 ;
      RECT  959100.0 369750.0 960300.0 370950.0 ;
      RECT  961500.0 359250.0 962700.0 360450.0 ;
      RECT  965400.0 357450.0 966600.0 358650.0 ;
      RECT  965400.0 357450.0 966600.0 358650.0 ;
      RECT  971850.0 376500.0 972750.0 377400.0 ;
      RECT  969000.0 376500.0 972300.0 377400.0 ;
      RECT  971850.0 370350.0 972750.0 376950.0 ;
      RECT  969450.0 354600.0 970350.0 355500.0 ;
      RECT  969900.0 354600.0 972450.0 355500.0 ;
      RECT  969450.0 355050.0 970350.0 359850.0 ;
      RECT  969300.0 359250.0 970500.0 360450.0 ;
      RECT  971700.0 359250.0 972900.0 360450.0 ;
      RECT  971700.0 359250.0 972900.0 360450.0 ;
      RECT  969300.0 359250.0 970500.0 360450.0 ;
      RECT  969300.0 369750.0 970500.0 370950.0 ;
      RECT  971700.0 369750.0 972900.0 370950.0 ;
      RECT  971700.0 369750.0 972900.0 370950.0 ;
      RECT  969300.0 369750.0 970500.0 370950.0 ;
      RECT  968850.0 376350.0 970050.0 377550.0 ;
      RECT  971850.0 354450.0 973050.0 355650.0 ;
      RECT  969300.0 369750.0 970500.0 370950.0 ;
      RECT  971700.0 359250.0 972900.0 360450.0 ;
      RECT  975600.0 357450.0 976800.0 358650.0 ;
      RECT  975600.0 357450.0 976800.0 358650.0 ;
      RECT  982050.0 376500.0 982950.0 377400.0 ;
      RECT  979200.0 376500.0 982500.0 377400.0 ;
      RECT  982050.0 370350.0 982950.0 376950.0 ;
      RECT  979650.0 354600.0 980550.0 355500.0 ;
      RECT  980100.0 354600.0 982650.0 355500.0 ;
      RECT  979650.0 355050.0 980550.0 359850.0 ;
      RECT  979500.0 359250.0 980700.0 360450.0 ;
      RECT  981900.0 359250.0 983100.0 360450.0 ;
      RECT  981900.0 359250.0 983100.0 360450.0 ;
      RECT  979500.0 359250.0 980700.0 360450.0 ;
      RECT  979500.0 369750.0 980700.0 370950.0 ;
      RECT  981900.0 369750.0 983100.0 370950.0 ;
      RECT  981900.0 369750.0 983100.0 370950.0 ;
      RECT  979500.0 369750.0 980700.0 370950.0 ;
      RECT  979050.0 376350.0 980250.0 377550.0 ;
      RECT  982050.0 354450.0 983250.0 355650.0 ;
      RECT  979500.0 369750.0 980700.0 370950.0 ;
      RECT  981900.0 359250.0 983100.0 360450.0 ;
      RECT  985800.0 357450.0 987000.0 358650.0 ;
      RECT  985800.0 357450.0 987000.0 358650.0 ;
      RECT  992250.0 376500.0 993150.0 377400.0 ;
      RECT  989400.0 376500.0 992700.0 377400.0 ;
      RECT  992250.0 370350.0 993150.0 376950.0 ;
      RECT  989850.0 354600.0 990750.0 355500.0 ;
      RECT  990300.0 354600.0 992850.0 355500.0 ;
      RECT  989850.0 355050.0 990750.0 359850.0 ;
      RECT  989700.0 359250.0 990900.0 360450.0 ;
      RECT  992100.0 359250.0 993300.0 360450.0 ;
      RECT  992100.0 359250.0 993300.0 360450.0 ;
      RECT  989700.0 359250.0 990900.0 360450.0 ;
      RECT  989700.0 369750.0 990900.0 370950.0 ;
      RECT  992100.0 369750.0 993300.0 370950.0 ;
      RECT  992100.0 369750.0 993300.0 370950.0 ;
      RECT  989700.0 369750.0 990900.0 370950.0 ;
      RECT  989250.0 376350.0 990450.0 377550.0 ;
      RECT  992250.0 354450.0 993450.0 355650.0 ;
      RECT  989700.0 369750.0 990900.0 370950.0 ;
      RECT  992100.0 359250.0 993300.0 360450.0 ;
      RECT  996000.0 357450.0 997200.0 358650.0 ;
      RECT  996000.0 357450.0 997200.0 358650.0 ;
      RECT  1002450.0 376500.0 1003350.0 377400.0 ;
      RECT  999600.0 376500.0 1002900.0 377400.0 ;
      RECT  1002450.0 370350.0 1003350.0 376950.0 ;
      RECT  1000050.0 354600.0 1000950.0 355500.0 ;
      RECT  1000500.0 354600.0 1003050.0 355500.0 ;
      RECT  1000050.0 355050.0 1000950.0 359850.0 ;
      RECT  999900.0 359250.0 1001100.0 360450.0 ;
      RECT  1002300.0 359250.0 1003500.0 360450.0 ;
      RECT  1002300.0 359250.0 1003500.0 360450.0 ;
      RECT  999900.0 359250.0 1001100.0 360450.0 ;
      RECT  999900.0 369750.0 1001100.0 370950.0 ;
      RECT  1002300.0 369750.0 1003500.0 370950.0 ;
      RECT  1002300.0 369750.0 1003500.0 370950.0 ;
      RECT  999900.0 369750.0 1001100.0 370950.0 ;
      RECT  999450.0 376350.0 1000650.0 377550.0 ;
      RECT  1002450.0 354450.0 1003650.0 355650.0 ;
      RECT  999900.0 369750.0 1001100.0 370950.0 ;
      RECT  1002300.0 359250.0 1003500.0 360450.0 ;
      RECT  1006200.0 357450.0 1007400.0 358650.0 ;
      RECT  1006200.0 357450.0 1007400.0 358650.0 ;
      RECT  1012650.0 376500.0 1013550.0 377400.0 ;
      RECT  1009800.0 376500.0 1013100.0 377400.0 ;
      RECT  1012650.0 370350.0 1013550.0 376950.0 ;
      RECT  1010250.0 354600.0 1011150.0 355500.0 ;
      RECT  1010700.0 354600.0 1013250.0 355500.0 ;
      RECT  1010250.0 355050.0 1011150.0 359850.0 ;
      RECT  1010100.0 359250.0 1011300.0 360450.0 ;
      RECT  1012500.0 359250.0 1013700.0 360450.0 ;
      RECT  1012500.0 359250.0 1013700.0 360450.0 ;
      RECT  1010100.0 359250.0 1011300.0 360450.0 ;
      RECT  1010100.0 369750.0 1011300.0 370950.0 ;
      RECT  1012500.0 369750.0 1013700.0 370950.0 ;
      RECT  1012500.0 369750.0 1013700.0 370950.0 ;
      RECT  1010100.0 369750.0 1011300.0 370950.0 ;
      RECT  1009650.0 376350.0 1010850.0 377550.0 ;
      RECT  1012650.0 354450.0 1013850.0 355650.0 ;
      RECT  1010100.0 369750.0 1011300.0 370950.0 ;
      RECT  1012500.0 359250.0 1013700.0 360450.0 ;
      RECT  1016400.0 357450.0 1017600.0 358650.0 ;
      RECT  1016400.0 357450.0 1017600.0 358650.0 ;
      RECT  1022850.0 376500.0 1023750.0 377400.0 ;
      RECT  1020000.0 376500.0 1023300.0 377400.0 ;
      RECT  1022850.0 370350.0 1023750.0 376950.0 ;
      RECT  1020450.0 354600.0 1021350.0 355500.0 ;
      RECT  1020900.0 354600.0 1023450.0 355500.0 ;
      RECT  1020450.0 355050.0 1021350.0 359850.0 ;
      RECT  1020300.0 359250.0 1021500.0 360450.0 ;
      RECT  1022700.0 359250.0 1023900.0 360450.0 ;
      RECT  1022700.0 359250.0 1023900.0 360450.0 ;
      RECT  1020300.0 359250.0 1021500.0 360450.0 ;
      RECT  1020300.0 369750.0 1021500.0 370950.0 ;
      RECT  1022700.0 369750.0 1023900.0 370950.0 ;
      RECT  1022700.0 369750.0 1023900.0 370950.0 ;
      RECT  1020300.0 369750.0 1021500.0 370950.0 ;
      RECT  1019850.0 376350.0 1021050.0 377550.0 ;
      RECT  1022850.0 354450.0 1024050.0 355650.0 ;
      RECT  1020300.0 369750.0 1021500.0 370950.0 ;
      RECT  1022700.0 359250.0 1023900.0 360450.0 ;
      RECT  1026600.0 357450.0 1027800.0 358650.0 ;
      RECT  1026600.0 357450.0 1027800.0 358650.0 ;
      RECT  1033050.0 376500.0 1033950.0 377400.0 ;
      RECT  1030200.0 376500.0 1033500.0 377400.0 ;
      RECT  1033050.0 370350.0 1033950.0 376950.0 ;
      RECT  1030650.0 354600.0 1031550.0 355500.0 ;
      RECT  1031100.0 354600.0 1033650.0 355500.0 ;
      RECT  1030650.0 355050.0 1031550.0 359850.0 ;
      RECT  1030500.0 359250.0 1031700.0 360450.0 ;
      RECT  1032900.0 359250.0 1034100.0 360450.0 ;
      RECT  1032900.0 359250.0 1034100.0 360450.0 ;
      RECT  1030500.0 359250.0 1031700.0 360450.0 ;
      RECT  1030500.0 369750.0 1031700.0 370950.0 ;
      RECT  1032900.0 369750.0 1034100.0 370950.0 ;
      RECT  1032900.0 369750.0 1034100.0 370950.0 ;
      RECT  1030500.0 369750.0 1031700.0 370950.0 ;
      RECT  1030050.0 376350.0 1031250.0 377550.0 ;
      RECT  1033050.0 354450.0 1034250.0 355650.0 ;
      RECT  1030500.0 369750.0 1031700.0 370950.0 ;
      RECT  1032900.0 359250.0 1034100.0 360450.0 ;
      RECT  1036800.0 357450.0 1038000.0 358650.0 ;
      RECT  1036800.0 357450.0 1038000.0 358650.0 ;
      RECT  1043250.0 376500.0 1044150.0 377400.0 ;
      RECT  1040400.0 376500.0 1043700.0 377400.0 ;
      RECT  1043250.0 370350.0 1044150.0 376950.0 ;
      RECT  1040850.0 354600.0 1041750.0 355500.0 ;
      RECT  1041300.0 354600.0 1043850.0 355500.0 ;
      RECT  1040850.0 355050.0 1041750.0 359850.0 ;
      RECT  1040700.0 359250.0 1041900.0 360450.0 ;
      RECT  1043100.0 359250.0 1044300.0 360450.0 ;
      RECT  1043100.0 359250.0 1044300.0 360450.0 ;
      RECT  1040700.0 359250.0 1041900.0 360450.0 ;
      RECT  1040700.0 369750.0 1041900.0 370950.0 ;
      RECT  1043100.0 369750.0 1044300.0 370950.0 ;
      RECT  1043100.0 369750.0 1044300.0 370950.0 ;
      RECT  1040700.0 369750.0 1041900.0 370950.0 ;
      RECT  1040250.0 376350.0 1041450.0 377550.0 ;
      RECT  1043250.0 354450.0 1044450.0 355650.0 ;
      RECT  1040700.0 369750.0 1041900.0 370950.0 ;
      RECT  1043100.0 359250.0 1044300.0 360450.0 ;
      RECT  1047000.0 357450.0 1048200.0 358650.0 ;
      RECT  1047000.0 357450.0 1048200.0 358650.0 ;
      RECT  1053450.0 376500.0 1054350.0 377400.0 ;
      RECT  1050600.0 376500.0 1053900.0 377400.0 ;
      RECT  1053450.0 370350.0 1054350.0 376950.0 ;
      RECT  1051050.0 354600.0 1051950.0 355500.0 ;
      RECT  1051500.0 354600.0 1054050.0 355500.0 ;
      RECT  1051050.0 355050.0 1051950.0 359850.0 ;
      RECT  1050900.0 359250.0 1052100.0 360450.0 ;
      RECT  1053300.0 359250.0 1054500.0 360450.0 ;
      RECT  1053300.0 359250.0 1054500.0 360450.0 ;
      RECT  1050900.0 359250.0 1052100.0 360450.0 ;
      RECT  1050900.0 369750.0 1052100.0 370950.0 ;
      RECT  1053300.0 369750.0 1054500.0 370950.0 ;
      RECT  1053300.0 369750.0 1054500.0 370950.0 ;
      RECT  1050900.0 369750.0 1052100.0 370950.0 ;
      RECT  1050450.0 376350.0 1051650.0 377550.0 ;
      RECT  1053450.0 354450.0 1054650.0 355650.0 ;
      RECT  1050900.0 369750.0 1052100.0 370950.0 ;
      RECT  1053300.0 359250.0 1054500.0 360450.0 ;
      RECT  1057200.0 357450.0 1058400.0 358650.0 ;
      RECT  1057200.0 357450.0 1058400.0 358650.0 ;
      RECT  1063650.0 376500.0 1064550.0 377400.0 ;
      RECT  1060800.0 376500.0 1064100.0 377400.0 ;
      RECT  1063650.0 370350.0 1064550.0 376950.0 ;
      RECT  1061250.0 354600.0 1062150.0 355500.0 ;
      RECT  1061700.0 354600.0 1064250.0 355500.0 ;
      RECT  1061250.0 355050.0 1062150.0 359850.0 ;
      RECT  1061100.0 359250.0 1062300.0 360450.0 ;
      RECT  1063500.0 359250.0 1064700.0 360450.0 ;
      RECT  1063500.0 359250.0 1064700.0 360450.0 ;
      RECT  1061100.0 359250.0 1062300.0 360450.0 ;
      RECT  1061100.0 369750.0 1062300.0 370950.0 ;
      RECT  1063500.0 369750.0 1064700.0 370950.0 ;
      RECT  1063500.0 369750.0 1064700.0 370950.0 ;
      RECT  1061100.0 369750.0 1062300.0 370950.0 ;
      RECT  1060650.0 376350.0 1061850.0 377550.0 ;
      RECT  1063650.0 354450.0 1064850.0 355650.0 ;
      RECT  1061100.0 369750.0 1062300.0 370950.0 ;
      RECT  1063500.0 359250.0 1064700.0 360450.0 ;
      RECT  1067400.0 357450.0 1068600.0 358650.0 ;
      RECT  1067400.0 357450.0 1068600.0 358650.0 ;
      RECT  1073850.0 376500.0 1074750.0 377400.0 ;
      RECT  1071000.0 376500.0 1074300.0 377400.0 ;
      RECT  1073850.0 370350.0 1074750.0 376950.0 ;
      RECT  1071450.0 354600.0 1072350.0 355500.0 ;
      RECT  1071900.0 354600.0 1074450.0 355500.0 ;
      RECT  1071450.0 355050.0 1072350.0 359850.0 ;
      RECT  1071300.0 359250.0 1072500.0 360450.0 ;
      RECT  1073700.0 359250.0 1074900.0 360450.0 ;
      RECT  1073700.0 359250.0 1074900.0 360450.0 ;
      RECT  1071300.0 359250.0 1072500.0 360450.0 ;
      RECT  1071300.0 369750.0 1072500.0 370950.0 ;
      RECT  1073700.0 369750.0 1074900.0 370950.0 ;
      RECT  1073700.0 369750.0 1074900.0 370950.0 ;
      RECT  1071300.0 369750.0 1072500.0 370950.0 ;
      RECT  1070850.0 376350.0 1072050.0 377550.0 ;
      RECT  1073850.0 354450.0 1075050.0 355650.0 ;
      RECT  1071300.0 369750.0 1072500.0 370950.0 ;
      RECT  1073700.0 359250.0 1074900.0 360450.0 ;
      RECT  1077600.0 357450.0 1078800.0 358650.0 ;
      RECT  1077600.0 357450.0 1078800.0 358650.0 ;
      RECT  1084050.0 376500.0 1084950.0 377400.0 ;
      RECT  1081200.0 376500.0 1084500.0 377400.0 ;
      RECT  1084050.0 370350.0 1084950.0 376950.0 ;
      RECT  1081650.0 354600.0 1082550.0 355500.0 ;
      RECT  1082100.0 354600.0 1084650.0 355500.0 ;
      RECT  1081650.0 355050.0 1082550.0 359850.0 ;
      RECT  1081500.0 359250.0 1082700.0 360450.0 ;
      RECT  1083900.0 359250.0 1085100.0 360450.0 ;
      RECT  1083900.0 359250.0 1085100.0 360450.0 ;
      RECT  1081500.0 359250.0 1082700.0 360450.0 ;
      RECT  1081500.0 369750.0 1082700.0 370950.0 ;
      RECT  1083900.0 369750.0 1085100.0 370950.0 ;
      RECT  1083900.0 369750.0 1085100.0 370950.0 ;
      RECT  1081500.0 369750.0 1082700.0 370950.0 ;
      RECT  1081050.0 376350.0 1082250.0 377550.0 ;
      RECT  1084050.0 354450.0 1085250.0 355650.0 ;
      RECT  1081500.0 369750.0 1082700.0 370950.0 ;
      RECT  1083900.0 359250.0 1085100.0 360450.0 ;
      RECT  1087800.0 357450.0 1089000.0 358650.0 ;
      RECT  1087800.0 357450.0 1089000.0 358650.0 ;
      RECT  1094250.0 376500.0 1095150.0 377400.0 ;
      RECT  1091400.0 376500.0 1094700.0 377400.0 ;
      RECT  1094250.0 370350.0 1095150.0 376950.0 ;
      RECT  1091850.0 354600.0 1092750.0 355500.0 ;
      RECT  1092300.0 354600.0 1094850.0 355500.0 ;
      RECT  1091850.0 355050.0 1092750.0 359850.0 ;
      RECT  1091700.0 359250.0 1092900.0 360450.0 ;
      RECT  1094100.0 359250.0 1095300.0 360450.0 ;
      RECT  1094100.0 359250.0 1095300.0 360450.0 ;
      RECT  1091700.0 359250.0 1092900.0 360450.0 ;
      RECT  1091700.0 369750.0 1092900.0 370950.0 ;
      RECT  1094100.0 369750.0 1095300.0 370950.0 ;
      RECT  1094100.0 369750.0 1095300.0 370950.0 ;
      RECT  1091700.0 369750.0 1092900.0 370950.0 ;
      RECT  1091250.0 376350.0 1092450.0 377550.0 ;
      RECT  1094250.0 354450.0 1095450.0 355650.0 ;
      RECT  1091700.0 369750.0 1092900.0 370950.0 ;
      RECT  1094100.0 359250.0 1095300.0 360450.0 ;
      RECT  1098000.0 357450.0 1099200.0 358650.0 ;
      RECT  1098000.0 357450.0 1099200.0 358650.0 ;
      RECT  1104450.0 376500.0 1105350.0 377400.0 ;
      RECT  1101600.0 376500.0 1104900.0 377400.0 ;
      RECT  1104450.0 370350.0 1105350.0 376950.0 ;
      RECT  1102050.0 354600.0 1102950.0 355500.0 ;
      RECT  1102500.0 354600.0 1105050.0 355500.0 ;
      RECT  1102050.0 355050.0 1102950.0 359850.0 ;
      RECT  1101900.0 359250.0 1103100.0 360450.0 ;
      RECT  1104300.0 359250.0 1105500.0 360450.0 ;
      RECT  1104300.0 359250.0 1105500.0 360450.0 ;
      RECT  1101900.0 359250.0 1103100.0 360450.0 ;
      RECT  1101900.0 369750.0 1103100.0 370950.0 ;
      RECT  1104300.0 369750.0 1105500.0 370950.0 ;
      RECT  1104300.0 369750.0 1105500.0 370950.0 ;
      RECT  1101900.0 369750.0 1103100.0 370950.0 ;
      RECT  1101450.0 376350.0 1102650.0 377550.0 ;
      RECT  1104450.0 354450.0 1105650.0 355650.0 ;
      RECT  1101900.0 369750.0 1103100.0 370950.0 ;
      RECT  1104300.0 359250.0 1105500.0 360450.0 ;
      RECT  1108200.0 357450.0 1109400.0 358650.0 ;
      RECT  1108200.0 357450.0 1109400.0 358650.0 ;
      RECT  1114650.0 376500.0 1115550.0 377400.0 ;
      RECT  1111800.0 376500.0 1115100.0 377400.0 ;
      RECT  1114650.0 370350.0 1115550.0 376950.0 ;
      RECT  1112250.0 354600.0 1113150.0 355500.0 ;
      RECT  1112700.0 354600.0 1115250.0 355500.0 ;
      RECT  1112250.0 355050.0 1113150.0 359850.0 ;
      RECT  1112100.0 359250.0 1113300.0 360450.0 ;
      RECT  1114500.0 359250.0 1115700.0 360450.0 ;
      RECT  1114500.0 359250.0 1115700.0 360450.0 ;
      RECT  1112100.0 359250.0 1113300.0 360450.0 ;
      RECT  1112100.0 369750.0 1113300.0 370950.0 ;
      RECT  1114500.0 369750.0 1115700.0 370950.0 ;
      RECT  1114500.0 369750.0 1115700.0 370950.0 ;
      RECT  1112100.0 369750.0 1113300.0 370950.0 ;
      RECT  1111650.0 376350.0 1112850.0 377550.0 ;
      RECT  1114650.0 354450.0 1115850.0 355650.0 ;
      RECT  1112100.0 369750.0 1113300.0 370950.0 ;
      RECT  1114500.0 359250.0 1115700.0 360450.0 ;
      RECT  1118400.0 357450.0 1119600.0 358650.0 ;
      RECT  1118400.0 357450.0 1119600.0 358650.0 ;
      RECT  1124850.0 376500.0 1125750.0 377400.0 ;
      RECT  1122000.0 376500.0 1125300.0 377400.0 ;
      RECT  1124850.0 370350.0 1125750.0 376950.0 ;
      RECT  1122450.0 354600.0 1123350.0 355500.0 ;
      RECT  1122900.0 354600.0 1125450.0 355500.0 ;
      RECT  1122450.0 355050.0 1123350.0 359850.0 ;
      RECT  1122300.0 359250.0 1123500.0 360450.0 ;
      RECT  1124700.0 359250.0 1125900.0 360450.0 ;
      RECT  1124700.0 359250.0 1125900.0 360450.0 ;
      RECT  1122300.0 359250.0 1123500.0 360450.0 ;
      RECT  1122300.0 369750.0 1123500.0 370950.0 ;
      RECT  1124700.0 369750.0 1125900.0 370950.0 ;
      RECT  1124700.0 369750.0 1125900.0 370950.0 ;
      RECT  1122300.0 369750.0 1123500.0 370950.0 ;
      RECT  1121850.0 376350.0 1123050.0 377550.0 ;
      RECT  1124850.0 354450.0 1126050.0 355650.0 ;
      RECT  1122300.0 369750.0 1123500.0 370950.0 ;
      RECT  1124700.0 359250.0 1125900.0 360450.0 ;
      RECT  1128600.0 357450.0 1129800.0 358650.0 ;
      RECT  1128600.0 357450.0 1129800.0 358650.0 ;
      RECT  1135050.0 376500.0 1135950.0 377400.0 ;
      RECT  1132200.0 376500.0 1135500.0 377400.0 ;
      RECT  1135050.0 370350.0 1135950.0 376950.0 ;
      RECT  1132650.0 354600.0 1133550.0 355500.0 ;
      RECT  1133100.0 354600.0 1135650.0 355500.0 ;
      RECT  1132650.0 355050.0 1133550.0 359850.0 ;
      RECT  1132500.0 359250.0 1133700.0 360450.0 ;
      RECT  1134900.0 359250.0 1136100.0 360450.0 ;
      RECT  1134900.0 359250.0 1136100.0 360450.0 ;
      RECT  1132500.0 359250.0 1133700.0 360450.0 ;
      RECT  1132500.0 369750.0 1133700.0 370950.0 ;
      RECT  1134900.0 369750.0 1136100.0 370950.0 ;
      RECT  1134900.0 369750.0 1136100.0 370950.0 ;
      RECT  1132500.0 369750.0 1133700.0 370950.0 ;
      RECT  1132050.0 376350.0 1133250.0 377550.0 ;
      RECT  1135050.0 354450.0 1136250.0 355650.0 ;
      RECT  1132500.0 369750.0 1133700.0 370950.0 ;
      RECT  1134900.0 359250.0 1136100.0 360450.0 ;
      RECT  1138800.0 357450.0 1140000.0 358650.0 ;
      RECT  1138800.0 357450.0 1140000.0 358650.0 ;
      RECT  1145250.0 376500.0 1146150.0 377400.0 ;
      RECT  1142400.0 376500.0 1145700.0 377400.0 ;
      RECT  1145250.0 370350.0 1146150.0 376950.0 ;
      RECT  1142850.0 354600.0 1143750.0 355500.0 ;
      RECT  1143300.0 354600.0 1145850.0 355500.0 ;
      RECT  1142850.0 355050.0 1143750.0 359850.0 ;
      RECT  1142700.0 359250.0 1143900.0 360450.0 ;
      RECT  1145100.0 359250.0 1146300.0 360450.0 ;
      RECT  1145100.0 359250.0 1146300.0 360450.0 ;
      RECT  1142700.0 359250.0 1143900.0 360450.0 ;
      RECT  1142700.0 369750.0 1143900.0 370950.0 ;
      RECT  1145100.0 369750.0 1146300.0 370950.0 ;
      RECT  1145100.0 369750.0 1146300.0 370950.0 ;
      RECT  1142700.0 369750.0 1143900.0 370950.0 ;
      RECT  1142250.0 376350.0 1143450.0 377550.0 ;
      RECT  1145250.0 354450.0 1146450.0 355650.0 ;
      RECT  1142700.0 369750.0 1143900.0 370950.0 ;
      RECT  1145100.0 359250.0 1146300.0 360450.0 ;
      RECT  1149000.0 357450.0 1150200.0 358650.0 ;
      RECT  1149000.0 357450.0 1150200.0 358650.0 ;
      RECT  1155450.0 376500.0 1156350.0 377400.0 ;
      RECT  1152600.0 376500.0 1155900.0 377400.0 ;
      RECT  1155450.0 370350.0 1156350.0 376950.0 ;
      RECT  1153050.0 354600.0 1153950.0 355500.0 ;
      RECT  1153500.0 354600.0 1156050.0 355500.0 ;
      RECT  1153050.0 355050.0 1153950.0 359850.0 ;
      RECT  1152900.0 359250.0 1154100.0 360450.0 ;
      RECT  1155300.0 359250.0 1156500.0 360450.0 ;
      RECT  1155300.0 359250.0 1156500.0 360450.0 ;
      RECT  1152900.0 359250.0 1154100.0 360450.0 ;
      RECT  1152900.0 369750.0 1154100.0 370950.0 ;
      RECT  1155300.0 369750.0 1156500.0 370950.0 ;
      RECT  1155300.0 369750.0 1156500.0 370950.0 ;
      RECT  1152900.0 369750.0 1154100.0 370950.0 ;
      RECT  1152450.0 376350.0 1153650.0 377550.0 ;
      RECT  1155450.0 354450.0 1156650.0 355650.0 ;
      RECT  1152900.0 369750.0 1154100.0 370950.0 ;
      RECT  1155300.0 359250.0 1156500.0 360450.0 ;
      RECT  1159200.0 357450.0 1160400.0 358650.0 ;
      RECT  1159200.0 357450.0 1160400.0 358650.0 ;
      RECT  1165650.0 376500.0 1166550.0 377400.0 ;
      RECT  1162800.0 376500.0 1166100.0 377400.0 ;
      RECT  1165650.0 370350.0 1166550.0 376950.0 ;
      RECT  1163250.0 354600.0 1164150.0 355500.0 ;
      RECT  1163700.0 354600.0 1166250.0 355500.0 ;
      RECT  1163250.0 355050.0 1164150.0 359850.0 ;
      RECT  1163100.0 359250.0 1164300.0 360450.0 ;
      RECT  1165500.0 359250.0 1166700.0 360450.0 ;
      RECT  1165500.0 359250.0 1166700.0 360450.0 ;
      RECT  1163100.0 359250.0 1164300.0 360450.0 ;
      RECT  1163100.0 369750.0 1164300.0 370950.0 ;
      RECT  1165500.0 369750.0 1166700.0 370950.0 ;
      RECT  1165500.0 369750.0 1166700.0 370950.0 ;
      RECT  1163100.0 369750.0 1164300.0 370950.0 ;
      RECT  1162650.0 376350.0 1163850.0 377550.0 ;
      RECT  1165650.0 354450.0 1166850.0 355650.0 ;
      RECT  1163100.0 369750.0 1164300.0 370950.0 ;
      RECT  1165500.0 359250.0 1166700.0 360450.0 ;
      RECT  1169400.0 357450.0 1170600.0 358650.0 ;
      RECT  1169400.0 357450.0 1170600.0 358650.0 ;
      RECT  1175850.0 376500.0 1176750.0 377400.0 ;
      RECT  1173000.0 376500.0 1176300.0 377400.0 ;
      RECT  1175850.0 370350.0 1176750.0 376950.0 ;
      RECT  1173450.0 354600.0 1174350.0 355500.0 ;
      RECT  1173900.0 354600.0 1176450.0 355500.0 ;
      RECT  1173450.0 355050.0 1174350.0 359850.0 ;
      RECT  1173300.0 359250.0 1174500.0 360450.0 ;
      RECT  1175700.0 359250.0 1176900.0 360450.0 ;
      RECT  1175700.0 359250.0 1176900.0 360450.0 ;
      RECT  1173300.0 359250.0 1174500.0 360450.0 ;
      RECT  1173300.0 369750.0 1174500.0 370950.0 ;
      RECT  1175700.0 369750.0 1176900.0 370950.0 ;
      RECT  1175700.0 369750.0 1176900.0 370950.0 ;
      RECT  1173300.0 369750.0 1174500.0 370950.0 ;
      RECT  1172850.0 376350.0 1174050.0 377550.0 ;
      RECT  1175850.0 354450.0 1177050.0 355650.0 ;
      RECT  1173300.0 369750.0 1174500.0 370950.0 ;
      RECT  1175700.0 359250.0 1176900.0 360450.0 ;
      RECT  1179600.0 357450.0 1180800.0 358650.0 ;
      RECT  1179600.0 357450.0 1180800.0 358650.0 ;
      RECT  1186050.0 376500.0 1186950.0 377400.0 ;
      RECT  1183200.0 376500.0 1186500.0 377400.0 ;
      RECT  1186050.0 370350.0 1186950.0 376950.0 ;
      RECT  1183650.0 354600.0 1184550.0 355500.0 ;
      RECT  1184100.0 354600.0 1186650.0 355500.0 ;
      RECT  1183650.0 355050.0 1184550.0 359850.0 ;
      RECT  1183500.0 359250.0 1184700.0 360450.0 ;
      RECT  1185900.0 359250.0 1187100.0 360450.0 ;
      RECT  1185900.0 359250.0 1187100.0 360450.0 ;
      RECT  1183500.0 359250.0 1184700.0 360450.0 ;
      RECT  1183500.0 369750.0 1184700.0 370950.0 ;
      RECT  1185900.0 369750.0 1187100.0 370950.0 ;
      RECT  1185900.0 369750.0 1187100.0 370950.0 ;
      RECT  1183500.0 369750.0 1184700.0 370950.0 ;
      RECT  1183050.0 376350.0 1184250.0 377550.0 ;
      RECT  1186050.0 354450.0 1187250.0 355650.0 ;
      RECT  1183500.0 369750.0 1184700.0 370950.0 ;
      RECT  1185900.0 359250.0 1187100.0 360450.0 ;
      RECT  1189800.0 357450.0 1191000.0 358650.0 ;
      RECT  1189800.0 357450.0 1191000.0 358650.0 ;
      RECT  1196250.0 376500.0 1197150.0 377400.0 ;
      RECT  1193400.0 376500.0 1196700.0 377400.0 ;
      RECT  1196250.0 370350.0 1197150.0 376950.0 ;
      RECT  1193850.0 354600.0 1194750.0 355500.0 ;
      RECT  1194300.0 354600.0 1196850.0 355500.0 ;
      RECT  1193850.0 355050.0 1194750.0 359850.0 ;
      RECT  1193700.0 359250.0 1194900.0 360450.0 ;
      RECT  1196100.0 359250.0 1197300.0 360450.0 ;
      RECT  1196100.0 359250.0 1197300.0 360450.0 ;
      RECT  1193700.0 359250.0 1194900.0 360450.0 ;
      RECT  1193700.0 369750.0 1194900.0 370950.0 ;
      RECT  1196100.0 369750.0 1197300.0 370950.0 ;
      RECT  1196100.0 369750.0 1197300.0 370950.0 ;
      RECT  1193700.0 369750.0 1194900.0 370950.0 ;
      RECT  1193250.0 376350.0 1194450.0 377550.0 ;
      RECT  1196250.0 354450.0 1197450.0 355650.0 ;
      RECT  1193700.0 369750.0 1194900.0 370950.0 ;
      RECT  1196100.0 359250.0 1197300.0 360450.0 ;
      RECT  1200000.0 357450.0 1201200.0 358650.0 ;
      RECT  1200000.0 357450.0 1201200.0 358650.0 ;
      RECT  1206450.0 376500.0 1207350.0 377400.0 ;
      RECT  1203600.0 376500.0 1206900.0 377400.0 ;
      RECT  1206450.0 370350.0 1207350.0 376950.0 ;
      RECT  1204050.0 354600.0 1204950.0 355500.0 ;
      RECT  1204500.0 354600.0 1207050.0 355500.0 ;
      RECT  1204050.0 355050.0 1204950.0 359850.0 ;
      RECT  1203900.0 359250.0 1205100.0 360450.0 ;
      RECT  1206300.0 359250.0 1207500.0 360450.0 ;
      RECT  1206300.0 359250.0 1207500.0 360450.0 ;
      RECT  1203900.0 359250.0 1205100.0 360450.0 ;
      RECT  1203900.0 369750.0 1205100.0 370950.0 ;
      RECT  1206300.0 369750.0 1207500.0 370950.0 ;
      RECT  1206300.0 369750.0 1207500.0 370950.0 ;
      RECT  1203900.0 369750.0 1205100.0 370950.0 ;
      RECT  1203450.0 376350.0 1204650.0 377550.0 ;
      RECT  1206450.0 354450.0 1207650.0 355650.0 ;
      RECT  1203900.0 369750.0 1205100.0 370950.0 ;
      RECT  1206300.0 359250.0 1207500.0 360450.0 ;
      RECT  1210200.0 357450.0 1211400.0 358650.0 ;
      RECT  1210200.0 357450.0 1211400.0 358650.0 ;
      RECT  1216650.0 376500.0 1217550.0 377400.0 ;
      RECT  1213800.0 376500.0 1217100.0 377400.0 ;
      RECT  1216650.0 370350.0 1217550.0 376950.0 ;
      RECT  1214250.0 354600.0 1215150.0 355500.0 ;
      RECT  1214700.0 354600.0 1217250.0 355500.0 ;
      RECT  1214250.0 355050.0 1215150.0 359850.0 ;
      RECT  1214100.0 359250.0 1215300.0 360450.0 ;
      RECT  1216500.0 359250.0 1217700.0 360450.0 ;
      RECT  1216500.0 359250.0 1217700.0 360450.0 ;
      RECT  1214100.0 359250.0 1215300.0 360450.0 ;
      RECT  1214100.0 369750.0 1215300.0 370950.0 ;
      RECT  1216500.0 369750.0 1217700.0 370950.0 ;
      RECT  1216500.0 369750.0 1217700.0 370950.0 ;
      RECT  1214100.0 369750.0 1215300.0 370950.0 ;
      RECT  1213650.0 376350.0 1214850.0 377550.0 ;
      RECT  1216650.0 354450.0 1217850.0 355650.0 ;
      RECT  1214100.0 369750.0 1215300.0 370950.0 ;
      RECT  1216500.0 359250.0 1217700.0 360450.0 ;
      RECT  1220400.0 357450.0 1221600.0 358650.0 ;
      RECT  1220400.0 357450.0 1221600.0 358650.0 ;
      RECT  1226850.0 376500.0 1227750.0 377400.0 ;
      RECT  1224000.0 376500.0 1227300.0 377400.0 ;
      RECT  1226850.0 370350.0 1227750.0 376950.0 ;
      RECT  1224450.0 354600.0 1225350.0 355500.0 ;
      RECT  1224900.0 354600.0 1227450.0 355500.0 ;
      RECT  1224450.0 355050.0 1225350.0 359850.0 ;
      RECT  1224300.0 359250.0 1225500.0 360450.0 ;
      RECT  1226700.0 359250.0 1227900.0 360450.0 ;
      RECT  1226700.0 359250.0 1227900.0 360450.0 ;
      RECT  1224300.0 359250.0 1225500.0 360450.0 ;
      RECT  1224300.0 369750.0 1225500.0 370950.0 ;
      RECT  1226700.0 369750.0 1227900.0 370950.0 ;
      RECT  1226700.0 369750.0 1227900.0 370950.0 ;
      RECT  1224300.0 369750.0 1225500.0 370950.0 ;
      RECT  1223850.0 376350.0 1225050.0 377550.0 ;
      RECT  1226850.0 354450.0 1228050.0 355650.0 ;
      RECT  1224300.0 369750.0 1225500.0 370950.0 ;
      RECT  1226700.0 359250.0 1227900.0 360450.0 ;
      RECT  1230600.0 357450.0 1231800.0 358650.0 ;
      RECT  1230600.0 357450.0 1231800.0 358650.0 ;
      RECT  1237050.0 376500.0 1237950.0 377400.0 ;
      RECT  1234200.0 376500.0 1237500.0 377400.0 ;
      RECT  1237050.0 370350.0 1237950.0 376950.0 ;
      RECT  1234650.0 354600.0 1235550.0 355500.0 ;
      RECT  1235100.0 354600.0 1237650.0 355500.0 ;
      RECT  1234650.0 355050.0 1235550.0 359850.0 ;
      RECT  1234500.0 359250.0 1235700.0 360450.0 ;
      RECT  1236900.0 359250.0 1238100.0 360450.0 ;
      RECT  1236900.0 359250.0 1238100.0 360450.0 ;
      RECT  1234500.0 359250.0 1235700.0 360450.0 ;
      RECT  1234500.0 369750.0 1235700.0 370950.0 ;
      RECT  1236900.0 369750.0 1238100.0 370950.0 ;
      RECT  1236900.0 369750.0 1238100.0 370950.0 ;
      RECT  1234500.0 369750.0 1235700.0 370950.0 ;
      RECT  1234050.0 376350.0 1235250.0 377550.0 ;
      RECT  1237050.0 354450.0 1238250.0 355650.0 ;
      RECT  1234500.0 369750.0 1235700.0 370950.0 ;
      RECT  1236900.0 359250.0 1238100.0 360450.0 ;
      RECT  1240800.0 357450.0 1242000.0 358650.0 ;
      RECT  1240800.0 357450.0 1242000.0 358650.0 ;
      RECT  1247250.0 376500.0 1248150.0 377400.0 ;
      RECT  1244400.0 376500.0 1247700.0 377400.0 ;
      RECT  1247250.0 370350.0 1248150.0 376950.0 ;
      RECT  1244850.0 354600.0 1245750.0 355500.0 ;
      RECT  1245300.0 354600.0 1247850.0 355500.0 ;
      RECT  1244850.0 355050.0 1245750.0 359850.0 ;
      RECT  1244700.0 359250.0 1245900.0 360450.0 ;
      RECT  1247100.0 359250.0 1248300.0 360450.0 ;
      RECT  1247100.0 359250.0 1248300.0 360450.0 ;
      RECT  1244700.0 359250.0 1245900.0 360450.0 ;
      RECT  1244700.0 369750.0 1245900.0 370950.0 ;
      RECT  1247100.0 369750.0 1248300.0 370950.0 ;
      RECT  1247100.0 369750.0 1248300.0 370950.0 ;
      RECT  1244700.0 369750.0 1245900.0 370950.0 ;
      RECT  1244250.0 376350.0 1245450.0 377550.0 ;
      RECT  1247250.0 354450.0 1248450.0 355650.0 ;
      RECT  1244700.0 369750.0 1245900.0 370950.0 ;
      RECT  1247100.0 359250.0 1248300.0 360450.0 ;
      RECT  1251000.0 357450.0 1252200.0 358650.0 ;
      RECT  1251000.0 357450.0 1252200.0 358650.0 ;
      RECT  1257450.0 376500.0 1258350.0 377400.0 ;
      RECT  1254600.0 376500.0 1257900.0 377400.0 ;
      RECT  1257450.0 370350.0 1258350.0 376950.0 ;
      RECT  1255050.0 354600.0 1255950.0 355500.0 ;
      RECT  1255500.0 354600.0 1258050.0 355500.0 ;
      RECT  1255050.0 355050.0 1255950.0 359850.0 ;
      RECT  1254900.0 359250.0 1256100.0 360450.0 ;
      RECT  1257300.0 359250.0 1258500.0 360450.0 ;
      RECT  1257300.0 359250.0 1258500.0 360450.0 ;
      RECT  1254900.0 359250.0 1256100.0 360450.0 ;
      RECT  1254900.0 369750.0 1256100.0 370950.0 ;
      RECT  1257300.0 369750.0 1258500.0 370950.0 ;
      RECT  1257300.0 369750.0 1258500.0 370950.0 ;
      RECT  1254900.0 369750.0 1256100.0 370950.0 ;
      RECT  1254450.0 376350.0 1255650.0 377550.0 ;
      RECT  1257450.0 354450.0 1258650.0 355650.0 ;
      RECT  1254900.0 369750.0 1256100.0 370950.0 ;
      RECT  1257300.0 359250.0 1258500.0 360450.0 ;
      RECT  1261200.0 357450.0 1262400.0 358650.0 ;
      RECT  1261200.0 357450.0 1262400.0 358650.0 ;
      RECT  1267650.0 376500.0 1268550.0 377400.0 ;
      RECT  1264800.0 376500.0 1268100.0 377400.0 ;
      RECT  1267650.0 370350.0 1268550.0 376950.0 ;
      RECT  1265250.0 354600.0 1266150.0 355500.0 ;
      RECT  1265700.0 354600.0 1268250.0 355500.0 ;
      RECT  1265250.0 355050.0 1266150.0 359850.0 ;
      RECT  1265100.0 359250.0 1266300.0 360450.0 ;
      RECT  1267500.0 359250.0 1268700.0 360450.0 ;
      RECT  1267500.0 359250.0 1268700.0 360450.0 ;
      RECT  1265100.0 359250.0 1266300.0 360450.0 ;
      RECT  1265100.0 369750.0 1266300.0 370950.0 ;
      RECT  1267500.0 369750.0 1268700.0 370950.0 ;
      RECT  1267500.0 369750.0 1268700.0 370950.0 ;
      RECT  1265100.0 369750.0 1266300.0 370950.0 ;
      RECT  1264650.0 376350.0 1265850.0 377550.0 ;
      RECT  1267650.0 354450.0 1268850.0 355650.0 ;
      RECT  1265100.0 369750.0 1266300.0 370950.0 ;
      RECT  1267500.0 359250.0 1268700.0 360450.0 ;
      RECT  1271400.0 357450.0 1272600.0 358650.0 ;
      RECT  1271400.0 357450.0 1272600.0 358650.0 ;
      RECT  1277850.0 376500.0 1278750.0 377400.0 ;
      RECT  1275000.0 376500.0 1278300.0 377400.0 ;
      RECT  1277850.0 370350.0 1278750.0 376950.0 ;
      RECT  1275450.0 354600.0 1276350.0 355500.0 ;
      RECT  1275900.0 354600.0 1278450.0 355500.0 ;
      RECT  1275450.0 355050.0 1276350.0 359850.0 ;
      RECT  1275300.0 359250.0 1276500.0 360450.0 ;
      RECT  1277700.0 359250.0 1278900.0 360450.0 ;
      RECT  1277700.0 359250.0 1278900.0 360450.0 ;
      RECT  1275300.0 359250.0 1276500.0 360450.0 ;
      RECT  1275300.0 369750.0 1276500.0 370950.0 ;
      RECT  1277700.0 369750.0 1278900.0 370950.0 ;
      RECT  1277700.0 369750.0 1278900.0 370950.0 ;
      RECT  1275300.0 369750.0 1276500.0 370950.0 ;
      RECT  1274850.0 376350.0 1276050.0 377550.0 ;
      RECT  1277850.0 354450.0 1279050.0 355650.0 ;
      RECT  1275300.0 369750.0 1276500.0 370950.0 ;
      RECT  1277700.0 359250.0 1278900.0 360450.0 ;
      RECT  1281600.0 357450.0 1282800.0 358650.0 ;
      RECT  1281600.0 357450.0 1282800.0 358650.0 ;
      RECT  1288050.0 376500.0 1288950.0 377400.0 ;
      RECT  1285200.0 376500.0 1288500.0 377400.0 ;
      RECT  1288050.0 370350.0 1288950.0 376950.0 ;
      RECT  1285650.0 354600.0 1286550.0 355500.0 ;
      RECT  1286100.0 354600.0 1288650.0 355500.0 ;
      RECT  1285650.0 355050.0 1286550.0 359850.0 ;
      RECT  1285500.0 359250.0 1286700.0 360450.0 ;
      RECT  1287900.0 359250.0 1289100.0 360450.0 ;
      RECT  1287900.0 359250.0 1289100.0 360450.0 ;
      RECT  1285500.0 359250.0 1286700.0 360450.0 ;
      RECT  1285500.0 369750.0 1286700.0 370950.0 ;
      RECT  1287900.0 369750.0 1289100.0 370950.0 ;
      RECT  1287900.0 369750.0 1289100.0 370950.0 ;
      RECT  1285500.0 369750.0 1286700.0 370950.0 ;
      RECT  1285050.0 376350.0 1286250.0 377550.0 ;
      RECT  1288050.0 354450.0 1289250.0 355650.0 ;
      RECT  1285500.0 369750.0 1286700.0 370950.0 ;
      RECT  1287900.0 359250.0 1289100.0 360450.0 ;
      RECT  1291800.0 357450.0 1293000.0 358650.0 ;
      RECT  1291800.0 357450.0 1293000.0 358650.0 ;
      RECT  1298250.0 376500.0 1299150.0 377400.0 ;
      RECT  1295400.0 376500.0 1298700.0 377400.0 ;
      RECT  1298250.0 370350.0 1299150.0 376950.0 ;
      RECT  1295850.0 354600.0 1296750.0 355500.0 ;
      RECT  1296300.0 354600.0 1298850.0 355500.0 ;
      RECT  1295850.0 355050.0 1296750.0 359850.0 ;
      RECT  1295700.0 359250.0 1296900.0 360450.0 ;
      RECT  1298100.0 359250.0 1299300.0 360450.0 ;
      RECT  1298100.0 359250.0 1299300.0 360450.0 ;
      RECT  1295700.0 359250.0 1296900.0 360450.0 ;
      RECT  1295700.0 369750.0 1296900.0 370950.0 ;
      RECT  1298100.0 369750.0 1299300.0 370950.0 ;
      RECT  1298100.0 369750.0 1299300.0 370950.0 ;
      RECT  1295700.0 369750.0 1296900.0 370950.0 ;
      RECT  1295250.0 376350.0 1296450.0 377550.0 ;
      RECT  1298250.0 354450.0 1299450.0 355650.0 ;
      RECT  1295700.0 369750.0 1296900.0 370950.0 ;
      RECT  1298100.0 359250.0 1299300.0 360450.0 ;
      RECT  1302000.0 357450.0 1303200.0 358650.0 ;
      RECT  1302000.0 357450.0 1303200.0 358650.0 ;
      RECT  1308450.0 376500.0 1309350.0 377400.0 ;
      RECT  1305600.0 376500.0 1308900.0 377400.0 ;
      RECT  1308450.0 370350.0 1309350.0 376950.0 ;
      RECT  1306050.0 354600.0 1306950.0 355500.0 ;
      RECT  1306500.0 354600.0 1309050.0 355500.0 ;
      RECT  1306050.0 355050.0 1306950.0 359850.0 ;
      RECT  1305900.0 359250.0 1307100.0 360450.0 ;
      RECT  1308300.0 359250.0 1309500.0 360450.0 ;
      RECT  1308300.0 359250.0 1309500.0 360450.0 ;
      RECT  1305900.0 359250.0 1307100.0 360450.0 ;
      RECT  1305900.0 369750.0 1307100.0 370950.0 ;
      RECT  1308300.0 369750.0 1309500.0 370950.0 ;
      RECT  1308300.0 369750.0 1309500.0 370950.0 ;
      RECT  1305900.0 369750.0 1307100.0 370950.0 ;
      RECT  1305450.0 376350.0 1306650.0 377550.0 ;
      RECT  1308450.0 354450.0 1309650.0 355650.0 ;
      RECT  1305900.0 369750.0 1307100.0 370950.0 ;
      RECT  1308300.0 359250.0 1309500.0 360450.0 ;
      RECT  1312200.0 357450.0 1313400.0 358650.0 ;
      RECT  1312200.0 357450.0 1313400.0 358650.0 ;
      RECT  1318650.0 376500.0 1319550.0 377400.0 ;
      RECT  1315800.0 376500.0 1319100.0 377400.0 ;
      RECT  1318650.0 370350.0 1319550.0 376950.0 ;
      RECT  1316250.0 354600.0 1317150.0 355500.0 ;
      RECT  1316700.0 354600.0 1319250.0 355500.0 ;
      RECT  1316250.0 355050.0 1317150.0 359850.0 ;
      RECT  1316100.0 359250.0 1317300.0 360450.0 ;
      RECT  1318500.0 359250.0 1319700.0 360450.0 ;
      RECT  1318500.0 359250.0 1319700.0 360450.0 ;
      RECT  1316100.0 359250.0 1317300.0 360450.0 ;
      RECT  1316100.0 369750.0 1317300.0 370950.0 ;
      RECT  1318500.0 369750.0 1319700.0 370950.0 ;
      RECT  1318500.0 369750.0 1319700.0 370950.0 ;
      RECT  1316100.0 369750.0 1317300.0 370950.0 ;
      RECT  1315650.0 376350.0 1316850.0 377550.0 ;
      RECT  1318650.0 354450.0 1319850.0 355650.0 ;
      RECT  1316100.0 369750.0 1317300.0 370950.0 ;
      RECT  1318500.0 359250.0 1319700.0 360450.0 ;
      RECT  1322400.0 357450.0 1323600.0 358650.0 ;
      RECT  1322400.0 357450.0 1323600.0 358650.0 ;
      RECT  1328850.0 376500.0 1329750.0 377400.0 ;
      RECT  1326000.0 376500.0 1329300.0 377400.0 ;
      RECT  1328850.0 370350.0 1329750.0 376950.0 ;
      RECT  1326450.0 354600.0 1327350.0 355500.0 ;
      RECT  1326900.0 354600.0 1329450.0 355500.0 ;
      RECT  1326450.0 355050.0 1327350.0 359850.0 ;
      RECT  1326300.0 359250.0 1327500.0 360450.0 ;
      RECT  1328700.0 359250.0 1329900.0 360450.0 ;
      RECT  1328700.0 359250.0 1329900.0 360450.0 ;
      RECT  1326300.0 359250.0 1327500.0 360450.0 ;
      RECT  1326300.0 369750.0 1327500.0 370950.0 ;
      RECT  1328700.0 369750.0 1329900.0 370950.0 ;
      RECT  1328700.0 369750.0 1329900.0 370950.0 ;
      RECT  1326300.0 369750.0 1327500.0 370950.0 ;
      RECT  1325850.0 376350.0 1327050.0 377550.0 ;
      RECT  1328850.0 354450.0 1330050.0 355650.0 ;
      RECT  1326300.0 369750.0 1327500.0 370950.0 ;
      RECT  1328700.0 359250.0 1329900.0 360450.0 ;
      RECT  1332600.0 357450.0 1333800.0 358650.0 ;
      RECT  1332600.0 357450.0 1333800.0 358650.0 ;
      RECT  1339050.0 376500.0 1339950.0 377400.0 ;
      RECT  1336200.0 376500.0 1339500.0 377400.0 ;
      RECT  1339050.0 370350.0 1339950.0 376950.0 ;
      RECT  1336650.0 354600.0 1337550.0 355500.0 ;
      RECT  1337100.0 354600.0 1339650.0 355500.0 ;
      RECT  1336650.0 355050.0 1337550.0 359850.0 ;
      RECT  1336500.0 359250.0 1337700.0 360450.0 ;
      RECT  1338900.0 359250.0 1340100.0 360450.0 ;
      RECT  1338900.0 359250.0 1340100.0 360450.0 ;
      RECT  1336500.0 359250.0 1337700.0 360450.0 ;
      RECT  1336500.0 369750.0 1337700.0 370950.0 ;
      RECT  1338900.0 369750.0 1340100.0 370950.0 ;
      RECT  1338900.0 369750.0 1340100.0 370950.0 ;
      RECT  1336500.0 369750.0 1337700.0 370950.0 ;
      RECT  1336050.0 376350.0 1337250.0 377550.0 ;
      RECT  1339050.0 354450.0 1340250.0 355650.0 ;
      RECT  1336500.0 369750.0 1337700.0 370950.0 ;
      RECT  1338900.0 359250.0 1340100.0 360450.0 ;
      RECT  1342800.0 357450.0 1344000.0 358650.0 ;
      RECT  1342800.0 357450.0 1344000.0 358650.0 ;
      RECT  1349250.0 376500.0 1350150.0 377400.0 ;
      RECT  1346400.0 376500.0 1349700.0 377400.0 ;
      RECT  1349250.0 370350.0 1350150.0 376950.0 ;
      RECT  1346850.0 354600.0 1347750.0 355500.0 ;
      RECT  1347300.0 354600.0 1349850.0 355500.0 ;
      RECT  1346850.0 355050.0 1347750.0 359850.0 ;
      RECT  1346700.0 359250.0 1347900.0 360450.0 ;
      RECT  1349100.0 359250.0 1350300.0 360450.0 ;
      RECT  1349100.0 359250.0 1350300.0 360450.0 ;
      RECT  1346700.0 359250.0 1347900.0 360450.0 ;
      RECT  1346700.0 369750.0 1347900.0 370950.0 ;
      RECT  1349100.0 369750.0 1350300.0 370950.0 ;
      RECT  1349100.0 369750.0 1350300.0 370950.0 ;
      RECT  1346700.0 369750.0 1347900.0 370950.0 ;
      RECT  1346250.0 376350.0 1347450.0 377550.0 ;
      RECT  1349250.0 354450.0 1350450.0 355650.0 ;
      RECT  1346700.0 369750.0 1347900.0 370950.0 ;
      RECT  1349100.0 359250.0 1350300.0 360450.0 ;
      RECT  1353000.0 357450.0 1354200.0 358650.0 ;
      RECT  1353000.0 357450.0 1354200.0 358650.0 ;
      RECT  1359450.0 376500.0 1360350.0 377400.0 ;
      RECT  1356600.0 376500.0 1359900.0 377400.0 ;
      RECT  1359450.0 370350.0 1360350.0 376950.0 ;
      RECT  1357050.0 354600.0 1357950.0 355500.0 ;
      RECT  1357500.0 354600.0 1360050.0 355500.0 ;
      RECT  1357050.0 355050.0 1357950.0 359850.0 ;
      RECT  1356900.0 359250.0 1358100.0 360450.0 ;
      RECT  1359300.0 359250.0 1360500.0 360450.0 ;
      RECT  1359300.0 359250.0 1360500.0 360450.0 ;
      RECT  1356900.0 359250.0 1358100.0 360450.0 ;
      RECT  1356900.0 369750.0 1358100.0 370950.0 ;
      RECT  1359300.0 369750.0 1360500.0 370950.0 ;
      RECT  1359300.0 369750.0 1360500.0 370950.0 ;
      RECT  1356900.0 369750.0 1358100.0 370950.0 ;
      RECT  1356450.0 376350.0 1357650.0 377550.0 ;
      RECT  1359450.0 354450.0 1360650.0 355650.0 ;
      RECT  1356900.0 369750.0 1358100.0 370950.0 ;
      RECT  1359300.0 359250.0 1360500.0 360450.0 ;
      RECT  1363200.0 357450.0 1364400.0 358650.0 ;
      RECT  1363200.0 357450.0 1364400.0 358650.0 ;
      RECT  1369650.0 376500.0 1370550.0 377400.0 ;
      RECT  1366800.0 376500.0 1370100.0 377400.0 ;
      RECT  1369650.0 370350.0 1370550.0 376950.0 ;
      RECT  1367250.0 354600.0 1368150.0 355500.0 ;
      RECT  1367700.0 354600.0 1370250.0 355500.0 ;
      RECT  1367250.0 355050.0 1368150.0 359850.0 ;
      RECT  1367100.0 359250.0 1368300.0 360450.0 ;
      RECT  1369500.0 359250.0 1370700.0 360450.0 ;
      RECT  1369500.0 359250.0 1370700.0 360450.0 ;
      RECT  1367100.0 359250.0 1368300.0 360450.0 ;
      RECT  1367100.0 369750.0 1368300.0 370950.0 ;
      RECT  1369500.0 369750.0 1370700.0 370950.0 ;
      RECT  1369500.0 369750.0 1370700.0 370950.0 ;
      RECT  1367100.0 369750.0 1368300.0 370950.0 ;
      RECT  1366650.0 376350.0 1367850.0 377550.0 ;
      RECT  1369650.0 354450.0 1370850.0 355650.0 ;
      RECT  1367100.0 369750.0 1368300.0 370950.0 ;
      RECT  1369500.0 359250.0 1370700.0 360450.0 ;
      RECT  1373400.0 357450.0 1374600.0 358650.0 ;
      RECT  1373400.0 357450.0 1374600.0 358650.0 ;
      RECT  1379850.0 376500.0 1380750.0 377400.0 ;
      RECT  1377000.0 376500.0 1380300.0 377400.0 ;
      RECT  1379850.0 370350.0 1380750.0 376950.0 ;
      RECT  1377450.0 354600.0 1378350.0 355500.0 ;
      RECT  1377900.0 354600.0 1380450.0 355500.0 ;
      RECT  1377450.0 355050.0 1378350.0 359850.0 ;
      RECT  1377300.0 359250.0 1378500.0 360450.0 ;
      RECT  1379700.0 359250.0 1380900.0 360450.0 ;
      RECT  1379700.0 359250.0 1380900.0 360450.0 ;
      RECT  1377300.0 359250.0 1378500.0 360450.0 ;
      RECT  1377300.0 369750.0 1378500.0 370950.0 ;
      RECT  1379700.0 369750.0 1380900.0 370950.0 ;
      RECT  1379700.0 369750.0 1380900.0 370950.0 ;
      RECT  1377300.0 369750.0 1378500.0 370950.0 ;
      RECT  1376850.0 376350.0 1378050.0 377550.0 ;
      RECT  1379850.0 354450.0 1381050.0 355650.0 ;
      RECT  1377300.0 369750.0 1378500.0 370950.0 ;
      RECT  1379700.0 359250.0 1380900.0 360450.0 ;
      RECT  1383600.0 357450.0 1384800.0 358650.0 ;
      RECT  1383600.0 357450.0 1384800.0 358650.0 ;
      RECT  1390050.0 376500.0 1390950.0 377400.0 ;
      RECT  1387200.0 376500.0 1390500.0 377400.0 ;
      RECT  1390050.0 370350.0 1390950.0 376950.0 ;
      RECT  1387650.0 354600.0 1388550.0 355500.0 ;
      RECT  1388100.0 354600.0 1390650.0 355500.0 ;
      RECT  1387650.0 355050.0 1388550.0 359850.0 ;
      RECT  1387500.0 359250.0 1388700.0 360450.0 ;
      RECT  1389900.0 359250.0 1391100.0 360450.0 ;
      RECT  1389900.0 359250.0 1391100.0 360450.0 ;
      RECT  1387500.0 359250.0 1388700.0 360450.0 ;
      RECT  1387500.0 369750.0 1388700.0 370950.0 ;
      RECT  1389900.0 369750.0 1391100.0 370950.0 ;
      RECT  1389900.0 369750.0 1391100.0 370950.0 ;
      RECT  1387500.0 369750.0 1388700.0 370950.0 ;
      RECT  1387050.0 376350.0 1388250.0 377550.0 ;
      RECT  1390050.0 354450.0 1391250.0 355650.0 ;
      RECT  1387500.0 369750.0 1388700.0 370950.0 ;
      RECT  1389900.0 359250.0 1391100.0 360450.0 ;
      RECT  1393800.0 357450.0 1395000.0 358650.0 ;
      RECT  1393800.0 357450.0 1395000.0 358650.0 ;
      RECT  1400250.0 376500.0 1401150.0 377400.0 ;
      RECT  1397400.0 376500.0 1400700.0 377400.0 ;
      RECT  1400250.0 370350.0 1401150.0 376950.0 ;
      RECT  1397850.0 354600.0 1398750.0 355500.0 ;
      RECT  1398300.0 354600.0 1400850.0 355500.0 ;
      RECT  1397850.0 355050.0 1398750.0 359850.0 ;
      RECT  1397700.0 359250.0 1398900.0 360450.0 ;
      RECT  1400100.0 359250.0 1401300.0 360450.0 ;
      RECT  1400100.0 359250.0 1401300.0 360450.0 ;
      RECT  1397700.0 359250.0 1398900.0 360450.0 ;
      RECT  1397700.0 369750.0 1398900.0 370950.0 ;
      RECT  1400100.0 369750.0 1401300.0 370950.0 ;
      RECT  1400100.0 369750.0 1401300.0 370950.0 ;
      RECT  1397700.0 369750.0 1398900.0 370950.0 ;
      RECT  1397250.0 376350.0 1398450.0 377550.0 ;
      RECT  1400250.0 354450.0 1401450.0 355650.0 ;
      RECT  1397700.0 369750.0 1398900.0 370950.0 ;
      RECT  1400100.0 359250.0 1401300.0 360450.0 ;
      RECT  1404000.0 357450.0 1405200.0 358650.0 ;
      RECT  1404000.0 357450.0 1405200.0 358650.0 ;
      RECT  1410450.0 376500.0 1411350.0 377400.0 ;
      RECT  1407600.0 376500.0 1410900.0 377400.0 ;
      RECT  1410450.0 370350.0 1411350.0 376950.0 ;
      RECT  1408050.0 354600.0 1408950.0 355500.0 ;
      RECT  1408500.0 354600.0 1411050.0 355500.0 ;
      RECT  1408050.0 355050.0 1408950.0 359850.0 ;
      RECT  1407900.0 359250.0 1409100.0 360450.0 ;
      RECT  1410300.0 359250.0 1411500.0 360450.0 ;
      RECT  1410300.0 359250.0 1411500.0 360450.0 ;
      RECT  1407900.0 359250.0 1409100.0 360450.0 ;
      RECT  1407900.0 369750.0 1409100.0 370950.0 ;
      RECT  1410300.0 369750.0 1411500.0 370950.0 ;
      RECT  1410300.0 369750.0 1411500.0 370950.0 ;
      RECT  1407900.0 369750.0 1409100.0 370950.0 ;
      RECT  1407450.0 376350.0 1408650.0 377550.0 ;
      RECT  1410450.0 354450.0 1411650.0 355650.0 ;
      RECT  1407900.0 369750.0 1409100.0 370950.0 ;
      RECT  1410300.0 359250.0 1411500.0 360450.0 ;
      RECT  1414200.0 357450.0 1415400.0 358650.0 ;
      RECT  1414200.0 357450.0 1415400.0 358650.0 ;
      RECT  1420650.0 376500.0 1421550.0 377400.0 ;
      RECT  1417800.0 376500.0 1421100.0 377400.0 ;
      RECT  1420650.0 370350.0 1421550.0 376950.0 ;
      RECT  1418250.0 354600.0 1419150.0 355500.0 ;
      RECT  1418700.0 354600.0 1421250.0 355500.0 ;
      RECT  1418250.0 355050.0 1419150.0 359850.0 ;
      RECT  1418100.0 359250.0 1419300.0 360450.0 ;
      RECT  1420500.0 359250.0 1421700.0 360450.0 ;
      RECT  1420500.0 359250.0 1421700.0 360450.0 ;
      RECT  1418100.0 359250.0 1419300.0 360450.0 ;
      RECT  1418100.0 369750.0 1419300.0 370950.0 ;
      RECT  1420500.0 369750.0 1421700.0 370950.0 ;
      RECT  1420500.0 369750.0 1421700.0 370950.0 ;
      RECT  1418100.0 369750.0 1419300.0 370950.0 ;
      RECT  1417650.0 376350.0 1418850.0 377550.0 ;
      RECT  1420650.0 354450.0 1421850.0 355650.0 ;
      RECT  1418100.0 369750.0 1419300.0 370950.0 ;
      RECT  1420500.0 359250.0 1421700.0 360450.0 ;
      RECT  1424400.0 357450.0 1425600.0 358650.0 ;
      RECT  1424400.0 357450.0 1425600.0 358650.0 ;
      RECT  1430850.0 376500.0 1431750.0 377400.0 ;
      RECT  1428000.0 376500.0 1431300.0 377400.0 ;
      RECT  1430850.0 370350.0 1431750.0 376950.0 ;
      RECT  1428450.0 354600.0 1429350.0 355500.0 ;
      RECT  1428900.0 354600.0 1431450.0 355500.0 ;
      RECT  1428450.0 355050.0 1429350.0 359850.0 ;
      RECT  1428300.0 359250.0 1429500.0 360450.0 ;
      RECT  1430700.0 359250.0 1431900.0 360450.0 ;
      RECT  1430700.0 359250.0 1431900.0 360450.0 ;
      RECT  1428300.0 359250.0 1429500.0 360450.0 ;
      RECT  1428300.0 369750.0 1429500.0 370950.0 ;
      RECT  1430700.0 369750.0 1431900.0 370950.0 ;
      RECT  1430700.0 369750.0 1431900.0 370950.0 ;
      RECT  1428300.0 369750.0 1429500.0 370950.0 ;
      RECT  1427850.0 376350.0 1429050.0 377550.0 ;
      RECT  1430850.0 354450.0 1432050.0 355650.0 ;
      RECT  1428300.0 369750.0 1429500.0 370950.0 ;
      RECT  1430700.0 359250.0 1431900.0 360450.0 ;
      RECT  1434600.0 357450.0 1435800.0 358650.0 ;
      RECT  1434600.0 357450.0 1435800.0 358650.0 ;
      RECT  1441050.0 376500.0 1441950.0 377400.0 ;
      RECT  1438200.0 376500.0 1441500.0 377400.0 ;
      RECT  1441050.0 370350.0 1441950.0 376950.0 ;
      RECT  1438650.0 354600.0 1439550.0 355500.0 ;
      RECT  1439100.0 354600.0 1441650.0 355500.0 ;
      RECT  1438650.0 355050.0 1439550.0 359850.0 ;
      RECT  1438500.0 359250.0 1439700.0 360450.0 ;
      RECT  1440900.0 359250.0 1442100.0 360450.0 ;
      RECT  1440900.0 359250.0 1442100.0 360450.0 ;
      RECT  1438500.0 359250.0 1439700.0 360450.0 ;
      RECT  1438500.0 369750.0 1439700.0 370950.0 ;
      RECT  1440900.0 369750.0 1442100.0 370950.0 ;
      RECT  1440900.0 369750.0 1442100.0 370950.0 ;
      RECT  1438500.0 369750.0 1439700.0 370950.0 ;
      RECT  1438050.0 376350.0 1439250.0 377550.0 ;
      RECT  1441050.0 354450.0 1442250.0 355650.0 ;
      RECT  1438500.0 369750.0 1439700.0 370950.0 ;
      RECT  1440900.0 359250.0 1442100.0 360450.0 ;
      RECT  1444800.0 357450.0 1446000.0 358650.0 ;
      RECT  1444800.0 357450.0 1446000.0 358650.0 ;
      RECT  1451250.0 376500.0 1452150.0 377400.0 ;
      RECT  1448400.0 376500.0 1451700.0 377400.0 ;
      RECT  1451250.0 370350.0 1452150.0 376950.0 ;
      RECT  1448850.0 354600.0 1449750.0 355500.0 ;
      RECT  1449300.0 354600.0 1451850.0 355500.0 ;
      RECT  1448850.0 355050.0 1449750.0 359850.0 ;
      RECT  1448700.0 359250.0 1449900.0 360450.0 ;
      RECT  1451100.0 359250.0 1452300.0 360450.0 ;
      RECT  1451100.0 359250.0 1452300.0 360450.0 ;
      RECT  1448700.0 359250.0 1449900.0 360450.0 ;
      RECT  1448700.0 369750.0 1449900.0 370950.0 ;
      RECT  1451100.0 369750.0 1452300.0 370950.0 ;
      RECT  1451100.0 369750.0 1452300.0 370950.0 ;
      RECT  1448700.0 369750.0 1449900.0 370950.0 ;
      RECT  1448250.0 376350.0 1449450.0 377550.0 ;
      RECT  1451250.0 354450.0 1452450.0 355650.0 ;
      RECT  1448700.0 369750.0 1449900.0 370950.0 ;
      RECT  1451100.0 359250.0 1452300.0 360450.0 ;
      RECT  1455000.0 357450.0 1456200.0 358650.0 ;
      RECT  1455000.0 357450.0 1456200.0 358650.0 ;
      RECT  1461450.0 376500.0 1462350.0 377400.0 ;
      RECT  1458600.0 376500.0 1461900.0 377400.0 ;
      RECT  1461450.0 370350.0 1462350.0 376950.0 ;
      RECT  1459050.0 354600.0 1459950.0 355500.0 ;
      RECT  1459500.0 354600.0 1462050.0 355500.0 ;
      RECT  1459050.0 355050.0 1459950.0 359850.0 ;
      RECT  1458900.0 359250.0 1460100.0 360450.0 ;
      RECT  1461300.0 359250.0 1462500.0 360450.0 ;
      RECT  1461300.0 359250.0 1462500.0 360450.0 ;
      RECT  1458900.0 359250.0 1460100.0 360450.0 ;
      RECT  1458900.0 369750.0 1460100.0 370950.0 ;
      RECT  1461300.0 369750.0 1462500.0 370950.0 ;
      RECT  1461300.0 369750.0 1462500.0 370950.0 ;
      RECT  1458900.0 369750.0 1460100.0 370950.0 ;
      RECT  1458450.0 376350.0 1459650.0 377550.0 ;
      RECT  1461450.0 354450.0 1462650.0 355650.0 ;
      RECT  1458900.0 369750.0 1460100.0 370950.0 ;
      RECT  1461300.0 359250.0 1462500.0 360450.0 ;
      RECT  1465200.0 357450.0 1466400.0 358650.0 ;
      RECT  1465200.0 357450.0 1466400.0 358650.0 ;
      RECT  1471650.0 376500.0 1472550.0 377400.0 ;
      RECT  1468800.0 376500.0 1472100.0 377400.0 ;
      RECT  1471650.0 370350.0 1472550.0 376950.0 ;
      RECT  1469250.0 354600.0 1470150.0 355500.0 ;
      RECT  1469700.0 354600.0 1472250.0 355500.0 ;
      RECT  1469250.0 355050.0 1470150.0 359850.0 ;
      RECT  1469100.0 359250.0 1470300.0 360450.0 ;
      RECT  1471500.0 359250.0 1472700.0 360450.0 ;
      RECT  1471500.0 359250.0 1472700.0 360450.0 ;
      RECT  1469100.0 359250.0 1470300.0 360450.0 ;
      RECT  1469100.0 369750.0 1470300.0 370950.0 ;
      RECT  1471500.0 369750.0 1472700.0 370950.0 ;
      RECT  1471500.0 369750.0 1472700.0 370950.0 ;
      RECT  1469100.0 369750.0 1470300.0 370950.0 ;
      RECT  1468650.0 376350.0 1469850.0 377550.0 ;
      RECT  1471650.0 354450.0 1472850.0 355650.0 ;
      RECT  1469100.0 369750.0 1470300.0 370950.0 ;
      RECT  1471500.0 359250.0 1472700.0 360450.0 ;
      RECT  1475400.0 357450.0 1476600.0 358650.0 ;
      RECT  1475400.0 357450.0 1476600.0 358650.0 ;
      RECT  1481850.0 376500.0 1482750.0 377400.0 ;
      RECT  1479000.0 376500.0 1482300.0 377400.0 ;
      RECT  1481850.0 370350.0 1482750.0 376950.0 ;
      RECT  1479450.0 354600.0 1480350.0 355500.0 ;
      RECT  1479900.0 354600.0 1482450.0 355500.0 ;
      RECT  1479450.0 355050.0 1480350.0 359850.0 ;
      RECT  1479300.0 359250.0 1480500.0 360450.0 ;
      RECT  1481700.0 359250.0 1482900.0 360450.0 ;
      RECT  1481700.0 359250.0 1482900.0 360450.0 ;
      RECT  1479300.0 359250.0 1480500.0 360450.0 ;
      RECT  1479300.0 369750.0 1480500.0 370950.0 ;
      RECT  1481700.0 369750.0 1482900.0 370950.0 ;
      RECT  1481700.0 369750.0 1482900.0 370950.0 ;
      RECT  1479300.0 369750.0 1480500.0 370950.0 ;
      RECT  1478850.0 376350.0 1480050.0 377550.0 ;
      RECT  1481850.0 354450.0 1483050.0 355650.0 ;
      RECT  1479300.0 369750.0 1480500.0 370950.0 ;
      RECT  1481700.0 359250.0 1482900.0 360450.0 ;
      RECT  1485600.0 357450.0 1486800.0 358650.0 ;
      RECT  1485600.0 357450.0 1486800.0 358650.0 ;
      RECT  1492050.0 376500.0 1492950.0 377400.0 ;
      RECT  1489200.0 376500.0 1492500.0 377400.0 ;
      RECT  1492050.0 370350.0 1492950.0 376950.0 ;
      RECT  1489650.0 354600.0 1490550.0 355500.0 ;
      RECT  1490100.0 354600.0 1492650.0 355500.0 ;
      RECT  1489650.0 355050.0 1490550.0 359850.0 ;
      RECT  1489500.0 359250.0 1490700.0 360450.0 ;
      RECT  1491900.0 359250.0 1493100.0 360450.0 ;
      RECT  1491900.0 359250.0 1493100.0 360450.0 ;
      RECT  1489500.0 359250.0 1490700.0 360450.0 ;
      RECT  1489500.0 369750.0 1490700.0 370950.0 ;
      RECT  1491900.0 369750.0 1493100.0 370950.0 ;
      RECT  1491900.0 369750.0 1493100.0 370950.0 ;
      RECT  1489500.0 369750.0 1490700.0 370950.0 ;
      RECT  1489050.0 376350.0 1490250.0 377550.0 ;
      RECT  1492050.0 354450.0 1493250.0 355650.0 ;
      RECT  1489500.0 369750.0 1490700.0 370950.0 ;
      RECT  1491900.0 359250.0 1493100.0 360450.0 ;
      RECT  1495800.0 357450.0 1497000.0 358650.0 ;
      RECT  1495800.0 357450.0 1497000.0 358650.0 ;
      RECT  1502250.0 376500.0 1503150.0 377400.0 ;
      RECT  1499400.0 376500.0 1502700.0 377400.0 ;
      RECT  1502250.0 370350.0 1503150.0 376950.0 ;
      RECT  1499850.0 354600.0 1500750.0 355500.0 ;
      RECT  1500300.0 354600.0 1502850.0 355500.0 ;
      RECT  1499850.0 355050.0 1500750.0 359850.0 ;
      RECT  1499700.0 359250.0 1500900.0 360450.0 ;
      RECT  1502100.0 359250.0 1503300.0 360450.0 ;
      RECT  1502100.0 359250.0 1503300.0 360450.0 ;
      RECT  1499700.0 359250.0 1500900.0 360450.0 ;
      RECT  1499700.0 369750.0 1500900.0 370950.0 ;
      RECT  1502100.0 369750.0 1503300.0 370950.0 ;
      RECT  1502100.0 369750.0 1503300.0 370950.0 ;
      RECT  1499700.0 369750.0 1500900.0 370950.0 ;
      RECT  1499250.0 376350.0 1500450.0 377550.0 ;
      RECT  1502250.0 354450.0 1503450.0 355650.0 ;
      RECT  1499700.0 369750.0 1500900.0 370950.0 ;
      RECT  1502100.0 359250.0 1503300.0 360450.0 ;
      RECT  1506000.0 357450.0 1507200.0 358650.0 ;
      RECT  1506000.0 357450.0 1507200.0 358650.0 ;
      RECT  1512450.0 376500.0 1513350.0 377400.0 ;
      RECT  1509600.0 376500.0 1512900.0 377400.0 ;
      RECT  1512450.0 370350.0 1513350.0 376950.0 ;
      RECT  1510050.0 354600.0 1510950.0 355500.0 ;
      RECT  1510500.0 354600.0 1513050.0 355500.0 ;
      RECT  1510050.0 355050.0 1510950.0 359850.0 ;
      RECT  1509900.0 359250.0 1511100.0 360450.0 ;
      RECT  1512300.0 359250.0 1513500.0 360450.0 ;
      RECT  1512300.0 359250.0 1513500.0 360450.0 ;
      RECT  1509900.0 359250.0 1511100.0 360450.0 ;
      RECT  1509900.0 369750.0 1511100.0 370950.0 ;
      RECT  1512300.0 369750.0 1513500.0 370950.0 ;
      RECT  1512300.0 369750.0 1513500.0 370950.0 ;
      RECT  1509900.0 369750.0 1511100.0 370950.0 ;
      RECT  1509450.0 376350.0 1510650.0 377550.0 ;
      RECT  1512450.0 354450.0 1513650.0 355650.0 ;
      RECT  1509900.0 369750.0 1511100.0 370950.0 ;
      RECT  1512300.0 359250.0 1513500.0 360450.0 ;
      RECT  1516200.0 357450.0 1517400.0 358650.0 ;
      RECT  1516200.0 357450.0 1517400.0 358650.0 ;
      RECT  1522650.0 376500.0 1523550.0 377400.0 ;
      RECT  1519800.0 376500.0 1523100.0 377400.0 ;
      RECT  1522650.0 370350.0 1523550.0 376950.0 ;
      RECT  1520250.0 354600.0 1521150.0 355500.0 ;
      RECT  1520700.0 354600.0 1523250.0 355500.0 ;
      RECT  1520250.0 355050.0 1521150.0 359850.0 ;
      RECT  1520100.0 359250.0 1521300.0 360450.0 ;
      RECT  1522500.0 359250.0 1523700.0 360450.0 ;
      RECT  1522500.0 359250.0 1523700.0 360450.0 ;
      RECT  1520100.0 359250.0 1521300.0 360450.0 ;
      RECT  1520100.0 369750.0 1521300.0 370950.0 ;
      RECT  1522500.0 369750.0 1523700.0 370950.0 ;
      RECT  1522500.0 369750.0 1523700.0 370950.0 ;
      RECT  1520100.0 369750.0 1521300.0 370950.0 ;
      RECT  1519650.0 376350.0 1520850.0 377550.0 ;
      RECT  1522650.0 354450.0 1523850.0 355650.0 ;
      RECT  1520100.0 369750.0 1521300.0 370950.0 ;
      RECT  1522500.0 359250.0 1523700.0 360450.0 ;
      RECT  1526400.0 357450.0 1527600.0 358650.0 ;
      RECT  1526400.0 357450.0 1527600.0 358650.0 ;
      RECT  227100.0 351150.0 225900.0 352350.0 ;
      RECT  237300.0 349050.0 236100.0 350250.0 ;
      RECT  247500.0 346950.0 246300.0 348150.0 ;
      RECT  257700.0 344850.0 256500.0 346050.0 ;
      RECT  267900.0 351150.0 266700.0 352350.0 ;
      RECT  278100.0 349050.0 276900.0 350250.0 ;
      RECT  288300.0 346950.0 287100.0 348150.0 ;
      RECT  298500.0 344850.0 297300.0 346050.0 ;
      RECT  308700.0 351150.0 307500.0 352350.0 ;
      RECT  318900.0 349050.0 317700.0 350250.0 ;
      RECT  329100.0 346950.0 327900.0 348150.0 ;
      RECT  339300.0 344850.0 338100.0 346050.0 ;
      RECT  349500.0 351150.0 348300.0 352350.0 ;
      RECT  359700.0 349050.0 358500.0 350250.0 ;
      RECT  369900.0 346950.0 368700.0 348150.0 ;
      RECT  380100.0 344850.0 378900.0 346050.0 ;
      RECT  390300.0 351150.0 389100.0 352350.0 ;
      RECT  400500.0 349050.0 399300.0 350250.0 ;
      RECT  410700.0 346950.0 409500.0 348150.0 ;
      RECT  420900.0 344850.0 419700.0 346050.0 ;
      RECT  431100.0 351150.0 429900.0 352350.0 ;
      RECT  441300.0 349050.0 440100.0 350250.0 ;
      RECT  451500.0 346950.0 450300.0 348150.0 ;
      RECT  461700.0 344850.0 460500.0 346050.0 ;
      RECT  471900.0 351150.0 470700.0 352350.0 ;
      RECT  482100.0 349050.0 480900.0 350250.0 ;
      RECT  492300.0 346950.0 491100.0 348150.0 ;
      RECT  502500.0 344850.0 501300.0 346050.0 ;
      RECT  512700.0 351150.0 511500.0 352350.0 ;
      RECT  522900.0 349050.0 521700.0 350250.0 ;
      RECT  533100.0 346950.0 531900.0 348150.0 ;
      RECT  543300.0 344850.0 542100.0 346050.0 ;
      RECT  553500.0 351150.0 552300.0 352350.0 ;
      RECT  563700.0 349050.0 562500.0 350250.0 ;
      RECT  573900.0 346950.0 572700.0 348150.0 ;
      RECT  584100.0 344850.0 582900.0 346050.0 ;
      RECT  594300.0 351150.0 593100.0 352350.0 ;
      RECT  604500.0 349050.0 603300.0 350250.0 ;
      RECT  614700.0 346950.0 613500.0 348150.0 ;
      RECT  624900.0 344850.0 623700.0 346050.0 ;
      RECT  635100.0 351150.0 633900.0 352350.0 ;
      RECT  645300.0 349050.0 644100.0 350250.0 ;
      RECT  655500.0 346950.0 654300.0 348150.0 ;
      RECT  665700.0 344850.0 664500.0 346050.0 ;
      RECT  675900.0 351150.0 674700.0 352350.0 ;
      RECT  686100.0 349050.0 684900.0 350250.0 ;
      RECT  696300.0 346950.0 695100.0 348150.0 ;
      RECT  706500.0 344850.0 705300.0 346050.0 ;
      RECT  716700.0 351150.0 715500.0 352350.0 ;
      RECT  726900.0 349050.0 725700.0 350250.0 ;
      RECT  737100.0 346950.0 735900.0 348150.0 ;
      RECT  747300.0 344850.0 746100.0 346050.0 ;
      RECT  757500.0 351150.0 756300.0 352350.0 ;
      RECT  767700.0 349050.0 766500.0 350250.0 ;
      RECT  777900.0 346950.0 776700.0 348150.0 ;
      RECT  788100.0 344850.0 786900.0 346050.0 ;
      RECT  798300.0 351150.0 797100.0 352350.0 ;
      RECT  808500.0 349050.0 807300.0 350250.0 ;
      RECT  818700.0 346950.0 817500.0 348150.0 ;
      RECT  828900.0 344850.0 827700.0 346050.0 ;
      RECT  839100.0 351150.0 837900.0 352350.0 ;
      RECT  849300.0 349050.0 848100.0 350250.0 ;
      RECT  859500.0 346950.0 858300.0 348150.0 ;
      RECT  869700.0 344850.0 868500.0 346050.0 ;
      RECT  879900.0 351150.0 878700.0 352350.0 ;
      RECT  890100.0 349050.0 888900.0 350250.0 ;
      RECT  900300.0 346950.0 899100.0 348150.0 ;
      RECT  910500.0 344850.0 909300.0 346050.0 ;
      RECT  920700.0 351150.0 919500.0 352350.0 ;
      RECT  930900.0 349050.0 929700.0 350250.0 ;
      RECT  941100.0 346950.0 939900.0 348150.0 ;
      RECT  951300.0 344850.0 950100.0 346050.0 ;
      RECT  961500.0 351150.0 960300.0 352350.0 ;
      RECT  971700.0 349050.0 970500.0 350250.0 ;
      RECT  981900.0 346950.0 980700.0 348150.0 ;
      RECT  992100.0 344850.0 990900.0 346050.0 ;
      RECT  1002300.0 351150.0 1001100.0 352350.0 ;
      RECT  1012500.0 349050.0 1011300.0 350250.0 ;
      RECT  1022700.0 346950.0 1021500.0 348150.0 ;
      RECT  1032900.0 344850.0 1031700.0 346050.0 ;
      RECT  1043100.0 351150.0 1041900.0 352350.0 ;
      RECT  1053300.0 349050.0 1052100.0 350250.0 ;
      RECT  1063500.0 346950.0 1062300.0 348150.0 ;
      RECT  1073700.0 344850.0 1072500.0 346050.0 ;
      RECT  1083900.0 351150.0 1082700.0 352350.0 ;
      RECT  1094100.0 349050.0 1092900.0 350250.0 ;
      RECT  1104300.0 346950.0 1103100.0 348150.0 ;
      RECT  1114500.0 344850.0 1113300.0 346050.0 ;
      RECT  1124700.0 351150.0 1123500.0 352350.0 ;
      RECT  1134900.0 349050.0 1133700.0 350250.0 ;
      RECT  1145100.0 346950.0 1143900.0 348150.0 ;
      RECT  1155300.0 344850.0 1154100.0 346050.0 ;
      RECT  1165500.0 351150.0 1164300.0 352350.0 ;
      RECT  1175700.0 349050.0 1174500.0 350250.0 ;
      RECT  1185900.0 346950.0 1184700.0 348150.0 ;
      RECT  1196100.0 344850.0 1194900.0 346050.0 ;
      RECT  1206300.0 351150.0 1205100.0 352350.0 ;
      RECT  1216500.0 349050.0 1215300.0 350250.0 ;
      RECT  1226700.0 346950.0 1225500.0 348150.0 ;
      RECT  1236900.0 344850.0 1235700.0 346050.0 ;
      RECT  1247100.0 351150.0 1245900.0 352350.0 ;
      RECT  1257300.0 349050.0 1256100.0 350250.0 ;
      RECT  1267500.0 346950.0 1266300.0 348150.0 ;
      RECT  1277700.0 344850.0 1276500.0 346050.0 ;
      RECT  1287900.0 351150.0 1286700.0 352350.0 ;
      RECT  1298100.0 349050.0 1296900.0 350250.0 ;
      RECT  1308300.0 346950.0 1307100.0 348150.0 ;
      RECT  1318500.0 344850.0 1317300.0 346050.0 ;
      RECT  1328700.0 351150.0 1327500.0 352350.0 ;
      RECT  1338900.0 349050.0 1337700.0 350250.0 ;
      RECT  1349100.0 346950.0 1347900.0 348150.0 ;
      RECT  1359300.0 344850.0 1358100.0 346050.0 ;
      RECT  1369500.0 351150.0 1368300.0 352350.0 ;
      RECT  1379700.0 349050.0 1378500.0 350250.0 ;
      RECT  1389900.0 346950.0 1388700.0 348150.0 ;
      RECT  1400100.0 344850.0 1398900.0 346050.0 ;
      RECT  1410300.0 351150.0 1409100.0 352350.0 ;
      RECT  1420500.0 349050.0 1419300.0 350250.0 ;
      RECT  1430700.0 346950.0 1429500.0 348150.0 ;
      RECT  1440900.0 344850.0 1439700.0 346050.0 ;
      RECT  1451100.0 351150.0 1449900.0 352350.0 ;
      RECT  1461300.0 349050.0 1460100.0 350250.0 ;
      RECT  1471500.0 346950.0 1470300.0 348150.0 ;
      RECT  1481700.0 344850.0 1480500.0 346050.0 ;
      RECT  1491900.0 351150.0 1490700.0 352350.0 ;
      RECT  1502100.0 349050.0 1500900.0 350250.0 ;
      RECT  1512300.0 346950.0 1511100.0 348150.0 ;
      RECT  1522500.0 344850.0 1521300.0 346050.0 ;
      RECT  225600.0 342750.0 224400.0 343950.0 ;
      RECT  227400.0 340650.0 226200.0 341850.0 ;
      RECT  235800.0 342750.0 234600.0 343950.0 ;
      RECT  237600.0 340650.0 236400.0 341850.0 ;
      RECT  246000.0 342750.0 244800.0 343950.0 ;
      RECT  247800.0 340650.0 246600.0 341850.0 ;
      RECT  256200.0 342750.0 255000.0 343950.0 ;
      RECT  258000.0 340650.0 256800.0 341850.0 ;
      RECT  266400.0 342750.0 265200.0 343950.0 ;
      RECT  268200.0 340650.0 267000.0 341850.0 ;
      RECT  276600.0 342750.0 275400.0 343950.0 ;
      RECT  278400.0 340650.0 277200.0 341850.0 ;
      RECT  286800.0 342750.0 285600.0 343950.0 ;
      RECT  288600.0 340650.0 287400.0 341850.0 ;
      RECT  297000.0 342750.0 295800.0 343950.0 ;
      RECT  298800.0 340650.0 297600.0 341850.0 ;
      RECT  307200.0 342750.0 306000.0 343950.0 ;
      RECT  309000.0 340650.0 307800.0 341850.0 ;
      RECT  317400.0 342750.0 316200.0 343950.0 ;
      RECT  319200.0 340650.0 318000.0 341850.0 ;
      RECT  327600.0 342750.0 326400.0 343950.0 ;
      RECT  329400.0 340650.0 328200.0 341850.0 ;
      RECT  337800.0 342750.0 336600.0 343950.0 ;
      RECT  339600.0 340650.0 338400.0 341850.0 ;
      RECT  348000.0 342750.0 346800.0 343950.0 ;
      RECT  349800.0 340650.0 348600.0 341850.0 ;
      RECT  358200.0 342750.0 357000.0 343950.0 ;
      RECT  360000.0 340650.0 358800.0 341850.0 ;
      RECT  368400.0 342750.0 367200.0 343950.0 ;
      RECT  370200.0 340650.0 369000.0 341850.0 ;
      RECT  378600.0 342750.0 377400.0 343950.0 ;
      RECT  380400.0 340650.0 379200.0 341850.0 ;
      RECT  388800.0 342750.0 387600.0 343950.0 ;
      RECT  390600.0 340650.0 389400.0 341850.0 ;
      RECT  399000.0 342750.0 397800.0 343950.0 ;
      RECT  400800.0 340650.0 399600.0 341850.0 ;
      RECT  409200.0 342750.0 408000.0 343950.0 ;
      RECT  411000.0 340650.0 409800.0 341850.0 ;
      RECT  419400.0 342750.0 418200.0 343950.0 ;
      RECT  421200.0 340650.0 420000.0 341850.0 ;
      RECT  429600.0 342750.0 428400.0 343950.0 ;
      RECT  431400.0 340650.0 430200.0 341850.0 ;
      RECT  439800.0 342750.0 438600.0 343950.0 ;
      RECT  441600.0 340650.0 440400.0 341850.0 ;
      RECT  450000.0 342750.0 448800.0 343950.0 ;
      RECT  451800.0 340650.0 450600.0 341850.0 ;
      RECT  460200.0 342750.0 459000.0 343950.0 ;
      RECT  462000.0 340650.0 460800.0 341850.0 ;
      RECT  470400.0 342750.0 469200.0 343950.0 ;
      RECT  472200.0 340650.0 471000.0 341850.0 ;
      RECT  480600.0 342750.0 479400.0 343950.0 ;
      RECT  482400.0 340650.0 481200.0 341850.0 ;
      RECT  490800.0 342750.0 489600.0 343950.0 ;
      RECT  492600.0 340650.0 491400.0 341850.0 ;
      RECT  501000.0 342750.0 499800.0 343950.0 ;
      RECT  502800.0 340650.0 501600.0 341850.0 ;
      RECT  511200.0 342750.0 510000.0 343950.0 ;
      RECT  513000.0 340650.0 511800.0 341850.0 ;
      RECT  521400.0 342750.0 520200.0 343950.0 ;
      RECT  523200.0 340650.0 522000.0 341850.0 ;
      RECT  531600.0 342750.0 530400.0 343950.0 ;
      RECT  533400.0 340650.0 532200.0 341850.0 ;
      RECT  541800.0 342750.0 540600.0 343950.0 ;
      RECT  543600.0 340650.0 542400.0 341850.0 ;
      RECT  552000.0 342750.0 550800.0 343950.0 ;
      RECT  553800.0 340650.0 552600.0 341850.0 ;
      RECT  562200.0 342750.0 561000.0 343950.0 ;
      RECT  564000.0 340650.0 562800.0 341850.0 ;
      RECT  572400.0 342750.0 571200.0 343950.0 ;
      RECT  574200.0 340650.0 573000.0 341850.0 ;
      RECT  582600.0 342750.0 581400.0 343950.0 ;
      RECT  584400.0 340650.0 583200.0 341850.0 ;
      RECT  592800.0 342750.0 591600.0 343950.0 ;
      RECT  594600.0 340650.0 593400.0 341850.0 ;
      RECT  603000.0 342750.0 601800.0 343950.0 ;
      RECT  604800.0 340650.0 603600.0 341850.0 ;
      RECT  613200.0 342750.0 612000.0 343950.0 ;
      RECT  615000.0 340650.0 613800.0 341850.0 ;
      RECT  623400.0 342750.0 622200.0 343950.0 ;
      RECT  625200.0 340650.0 624000.0 341850.0 ;
      RECT  633600.0 342750.0 632400.0 343950.0 ;
      RECT  635400.0 340650.0 634200.0 341850.0 ;
      RECT  643800.0 342750.0 642600.0 343950.0 ;
      RECT  645600.0 340650.0 644400.0 341850.0 ;
      RECT  654000.0 342750.0 652800.0 343950.0 ;
      RECT  655800.0 340650.0 654600.0 341850.0 ;
      RECT  664200.0 342750.0 663000.0 343950.0 ;
      RECT  666000.0 340650.0 664800.0 341850.0 ;
      RECT  674400.0 342750.0 673200.0 343950.0 ;
      RECT  676200.0 340650.0 675000.0 341850.0 ;
      RECT  684600.0 342750.0 683400.0 343950.0 ;
      RECT  686400.0 340650.0 685200.0 341850.0 ;
      RECT  694800.0 342750.0 693600.0 343950.0 ;
      RECT  696600.0 340650.0 695400.0 341850.0 ;
      RECT  705000.0 342750.0 703800.0 343950.0 ;
      RECT  706800.0 340650.0 705600.0 341850.0 ;
      RECT  715200.0 342750.0 714000.0 343950.0 ;
      RECT  717000.0 340650.0 715800.0 341850.0 ;
      RECT  725400.0 342750.0 724200.0 343950.0 ;
      RECT  727200.0 340650.0 726000.0 341850.0 ;
      RECT  735600.0 342750.0 734400.0 343950.0 ;
      RECT  737400.0 340650.0 736200.0 341850.0 ;
      RECT  745800.0 342750.0 744600.0 343950.0 ;
      RECT  747600.0 340650.0 746400.0 341850.0 ;
      RECT  756000.0 342750.0 754800.0 343950.0 ;
      RECT  757800.0 340650.0 756600.0 341850.0 ;
      RECT  766200.0 342750.0 765000.0 343950.0 ;
      RECT  768000.0 340650.0 766800.0 341850.0 ;
      RECT  776400.0 342750.0 775200.0 343950.0 ;
      RECT  778200.0 340650.0 777000.0 341850.0 ;
      RECT  786600.0 342750.0 785400.0 343950.0 ;
      RECT  788400.0 340650.0 787200.0 341850.0 ;
      RECT  796800.0 342750.0 795600.0 343950.0 ;
      RECT  798600.0 340650.0 797400.0 341850.0 ;
      RECT  807000.0 342750.0 805800.0 343950.0 ;
      RECT  808800.0 340650.0 807600.0 341850.0 ;
      RECT  817200.0 342750.0 816000.0 343950.0 ;
      RECT  819000.0 340650.0 817800.0 341850.0 ;
      RECT  827400.0 342750.0 826200.0 343950.0 ;
      RECT  829200.0 340650.0 828000.0 341850.0 ;
      RECT  837600.0 342750.0 836400.0 343950.0 ;
      RECT  839400.0 340650.0 838200.0 341850.0 ;
      RECT  847800.0 342750.0 846600.0 343950.0 ;
      RECT  849600.0 340650.0 848400.0 341850.0 ;
      RECT  858000.0 342750.0 856800.0 343950.0 ;
      RECT  859800.0 340650.0 858600.0 341850.0 ;
      RECT  868200.0 342750.0 867000.0 343950.0 ;
      RECT  870000.0 340650.0 868800.0 341850.0 ;
      RECT  878400.0 342750.0 877200.0 343950.0 ;
      RECT  880200.0 340650.0 879000.0 341850.0 ;
      RECT  888600.0 342750.0 887400.0 343950.0 ;
      RECT  890400.0 340650.0 889200.0 341850.0 ;
      RECT  898800.0 342750.0 897600.0 343950.0 ;
      RECT  900600.0 340650.0 899400.0 341850.0 ;
      RECT  909000.0 342750.0 907800.0 343950.0 ;
      RECT  910800.0 340650.0 909600.0 341850.0 ;
      RECT  919200.0 342750.0 918000.0 343950.0 ;
      RECT  921000.0 340650.0 919800.0 341850.0 ;
      RECT  929400.0 342750.0 928200.0 343950.0 ;
      RECT  931200.0 340650.0 930000.0 341850.0 ;
      RECT  939600.0 342750.0 938400.0 343950.0 ;
      RECT  941400.0 340650.0 940200.0 341850.0 ;
      RECT  949800.0 342750.0 948600.0 343950.0 ;
      RECT  951600.0 340650.0 950400.0 341850.0 ;
      RECT  960000.0 342750.0 958800.0 343950.0 ;
      RECT  961800.0 340650.0 960600.0 341850.0 ;
      RECT  970200.0 342750.0 969000.0 343950.0 ;
      RECT  972000.0 340650.0 970800.0 341850.0 ;
      RECT  980400.0 342750.0 979200.0 343950.0 ;
      RECT  982200.0 340650.0 981000.0 341850.0 ;
      RECT  990600.0 342750.0 989400.0 343950.0 ;
      RECT  992400.0 340650.0 991200.0 341850.0 ;
      RECT  1000800.0 342750.0 999600.0 343950.0 ;
      RECT  1002600.0 340650.0 1001400.0 341850.0 ;
      RECT  1011000.0 342750.0 1009800.0 343950.0 ;
      RECT  1012800.0 340650.0 1011600.0 341850.0 ;
      RECT  1021200.0 342750.0 1020000.0 343950.0 ;
      RECT  1023000.0 340650.0 1021800.0 341850.0 ;
      RECT  1031400.0 342750.0 1030200.0 343950.0 ;
      RECT  1033200.0 340650.0 1032000.0 341850.0 ;
      RECT  1041600.0 342750.0 1040400.0 343950.0 ;
      RECT  1043400.0 340650.0 1042200.0 341850.0 ;
      RECT  1051800.0 342750.0 1050600.0 343950.0 ;
      RECT  1053600.0 340650.0 1052400.0 341850.0 ;
      RECT  1062000.0 342750.0 1060800.0 343950.0 ;
      RECT  1063800.0 340650.0 1062600.0 341850.0 ;
      RECT  1072200.0 342750.0 1071000.0 343950.0 ;
      RECT  1074000.0 340650.0 1072800.0 341850.0 ;
      RECT  1082400.0 342750.0 1081200.0 343950.0 ;
      RECT  1084200.0 340650.0 1083000.0 341850.0 ;
      RECT  1092600.0 342750.0 1091400.0 343950.0 ;
      RECT  1094400.0 340650.0 1093200.0 341850.0 ;
      RECT  1102800.0 342750.0 1101600.0 343950.0 ;
      RECT  1104600.0 340650.0 1103400.0 341850.0 ;
      RECT  1113000.0 342750.0 1111800.0 343950.0 ;
      RECT  1114800.0 340650.0 1113600.0 341850.0 ;
      RECT  1123200.0 342750.0 1122000.0 343950.0 ;
      RECT  1125000.0 340650.0 1123800.0 341850.0 ;
      RECT  1133400.0 342750.0 1132200.0 343950.0 ;
      RECT  1135200.0 340650.0 1134000.0 341850.0 ;
      RECT  1143600.0 342750.0 1142400.0 343950.0 ;
      RECT  1145400.0 340650.0 1144200.0 341850.0 ;
      RECT  1153800.0 342750.0 1152600.0 343950.0 ;
      RECT  1155600.0 340650.0 1154400.0 341850.0 ;
      RECT  1164000.0 342750.0 1162800.0 343950.0 ;
      RECT  1165800.0 340650.0 1164600.0 341850.0 ;
      RECT  1174200.0 342750.0 1173000.0 343950.0 ;
      RECT  1176000.0 340650.0 1174800.0 341850.0 ;
      RECT  1184400.0 342750.0 1183200.0 343950.0 ;
      RECT  1186200.0 340650.0 1185000.0 341850.0 ;
      RECT  1194600.0 342750.0 1193400.0 343950.0 ;
      RECT  1196400.0 340650.0 1195200.0 341850.0 ;
      RECT  1204800.0 342750.0 1203600.0 343950.0 ;
      RECT  1206600.0 340650.0 1205400.0 341850.0 ;
      RECT  1215000.0 342750.0 1213800.0 343950.0 ;
      RECT  1216800.0 340650.0 1215600.0 341850.0 ;
      RECT  1225200.0 342750.0 1224000.0 343950.0 ;
      RECT  1227000.0 340650.0 1225800.0 341850.0 ;
      RECT  1235400.0 342750.0 1234200.0 343950.0 ;
      RECT  1237200.0 340650.0 1236000.0 341850.0 ;
      RECT  1245600.0 342750.0 1244400.0 343950.0 ;
      RECT  1247400.0 340650.0 1246200.0 341850.0 ;
      RECT  1255800.0 342750.0 1254600.0 343950.0 ;
      RECT  1257600.0 340650.0 1256400.0 341850.0 ;
      RECT  1266000.0 342750.0 1264800.0 343950.0 ;
      RECT  1267800.0 340650.0 1266600.0 341850.0 ;
      RECT  1276200.0 342750.0 1275000.0 343950.0 ;
      RECT  1278000.0 340650.0 1276800.0 341850.0 ;
      RECT  1286400.0 342750.0 1285200.0 343950.0 ;
      RECT  1288200.0 340650.0 1287000.0 341850.0 ;
      RECT  1296600.0 342750.0 1295400.0 343950.0 ;
      RECT  1298400.0 340650.0 1297200.0 341850.0 ;
      RECT  1306800.0 342750.0 1305600.0 343950.0 ;
      RECT  1308600.0 340650.0 1307400.0 341850.0 ;
      RECT  1317000.0 342750.0 1315800.0 343950.0 ;
      RECT  1318800.0 340650.0 1317600.0 341850.0 ;
      RECT  1327200.0 342750.0 1326000.0 343950.0 ;
      RECT  1329000.0 340650.0 1327800.0 341850.0 ;
      RECT  1337400.0 342750.0 1336200.0 343950.0 ;
      RECT  1339200.0 340650.0 1338000.0 341850.0 ;
      RECT  1347600.0 342750.0 1346400.0 343950.0 ;
      RECT  1349400.0 340650.0 1348200.0 341850.0 ;
      RECT  1357800.0 342750.0 1356600.0 343950.0 ;
      RECT  1359600.0 340650.0 1358400.0 341850.0 ;
      RECT  1368000.0 342750.0 1366800.0 343950.0 ;
      RECT  1369800.0 340650.0 1368600.0 341850.0 ;
      RECT  1378200.0 342750.0 1377000.0 343950.0 ;
      RECT  1380000.0 340650.0 1378800.0 341850.0 ;
      RECT  1388400.0 342750.0 1387200.0 343950.0 ;
      RECT  1390200.0 340650.0 1389000.0 341850.0 ;
      RECT  1398600.0 342750.0 1397400.0 343950.0 ;
      RECT  1400400.0 340650.0 1399200.0 341850.0 ;
      RECT  1408800.0 342750.0 1407600.0 343950.0 ;
      RECT  1410600.0 340650.0 1409400.0 341850.0 ;
      RECT  1419000.0 342750.0 1417800.0 343950.0 ;
      RECT  1420800.0 340650.0 1419600.0 341850.0 ;
      RECT  1429200.0 342750.0 1428000.0 343950.0 ;
      RECT  1431000.0 340650.0 1429800.0 341850.0 ;
      RECT  1439400.0 342750.0 1438200.0 343950.0 ;
      RECT  1441200.0 340650.0 1440000.0 341850.0 ;
      RECT  1449600.0 342750.0 1448400.0 343950.0 ;
      RECT  1451400.0 340650.0 1450200.0 341850.0 ;
      RECT  1459800.0 342750.0 1458600.0 343950.0 ;
      RECT  1461600.0 340650.0 1460400.0 341850.0 ;
      RECT  1470000.0 342750.0 1468800.0 343950.0 ;
      RECT  1471800.0 340650.0 1470600.0 341850.0 ;
      RECT  1480200.0 342750.0 1479000.0 343950.0 ;
      RECT  1482000.0 340650.0 1480800.0 341850.0 ;
      RECT  1490400.0 342750.0 1489200.0 343950.0 ;
      RECT  1492200.0 340650.0 1491000.0 341850.0 ;
      RECT  1500600.0 342750.0 1499400.0 343950.0 ;
      RECT  1502400.0 340650.0 1501200.0 341850.0 ;
      RECT  1510800.0 342750.0 1509600.0 343950.0 ;
      RECT  1512600.0 340650.0 1511400.0 341850.0 ;
      RECT  1521000.0 342750.0 1519800.0 343950.0 ;
      RECT  1522800.0 340650.0 1521600.0 341850.0 ;
      RECT  221400.0 351150.0 1527000.0 352350.0 ;
      RECT  221400.0 349050.0 1527000.0 350250.0 ;
      RECT  221400.0 346950.0 1527000.0 348150.0 ;
      RECT  221400.0 344850.0 1527000.0 346050.0 ;
      RECT  113550.0 6750.0 114450.0 7650.0 ;
      RECT  113550.0 11250.0 114450.0 12150.0 ;
      RECT  109350.0 6750.0 114000.0 7650.0 ;
      RECT  113550.0 7200.0 114450.0 11700.0 ;
      RECT  114000.0 11250.0 116550.0 12150.0 ;
      RECT  97950.0 6750.0 105900.0 7650.0 ;
      RECT  113550.0 21150.0 114450.0 22050.0 ;
      RECT  113550.0 25050.0 114450.0 25950.0 ;
      RECT  109350.0 21150.0 114000.0 22050.0 ;
      RECT  113550.0 21600.0 114450.0 25500.0 ;
      RECT  114000.0 25050.0 119550.0 25950.0 ;
      RECT  100950.0 21150.0 105900.0 22050.0 ;
      RECT  97950.0 29850.0 122550.0 30750.0 ;
      RECT  100950.0 43650.0 125550.0 44550.0 ;
      RECT  116550.0 7950.0 130500.0 8850.0 ;
      RECT  119550.0 5250.0 133500.0 6150.0 ;
      RECT  122550.0 19950.0 130500.0 20850.0 ;
      RECT  119550.0 22650.0 133500.0 23550.0 ;
      RECT  116550.0 35550.0 130500.0 36450.0 ;
      RECT  125550.0 32850.0 133500.0 33750.0 ;
      RECT  122550.0 47550.0 130500.0 48450.0 ;
      RECT  125550.0 50250.0 133500.0 51150.0 ;
      RECT  139950.0 7950.0 140850.0 8850.0 ;
      RECT  139950.0 6750.0 140850.0 7650.0 ;
      RECT  135900.0 7950.0 140400.0 8850.0 ;
      RECT  139950.0 7200.0 140850.0 8400.0 ;
      RECT  140400.0 6750.0 144900.0 7650.0 ;
      RECT  139950.0 19950.0 140850.0 20850.0 ;
      RECT  139950.0 21150.0 140850.0 22050.0 ;
      RECT  135900.0 19950.0 140400.0 20850.0 ;
      RECT  139950.0 20400.0 140850.0 21600.0 ;
      RECT  140400.0 21150.0 144900.0 22050.0 ;
      RECT  139950.0 35550.0 140850.0 36450.0 ;
      RECT  139950.0 34350.0 140850.0 35250.0 ;
      RECT  135900.0 35550.0 140400.0 36450.0 ;
      RECT  139950.0 34800.0 140850.0 36000.0 ;
      RECT  140400.0 34350.0 144900.0 35250.0 ;
      RECT  139950.0 47550.0 140850.0 48450.0 ;
      RECT  139950.0 48750.0 140850.0 49650.0 ;
      RECT  135900.0 47550.0 140400.0 48450.0 ;
      RECT  139950.0 48000.0 140850.0 49200.0 ;
      RECT  140400.0 48750.0 144900.0 49650.0 ;
      RECT  110100.0 12450.0 111300.0 14400.0 ;
      RECT  110100.0 600.0 111300.0 2550.0 ;
      RECT  105300.0 1950.0 106500.0 150.0 ;
      RECT  105300.0 11250.0 106500.0 14850.0 ;
      RECT  108000.0 1950.0 108900.0 11250.0 ;
      RECT  105300.0 11250.0 106500.0 12450.0 ;
      RECT  107700.0 11250.0 108900.0 12450.0 ;
      RECT  107700.0 11250.0 108900.0 12450.0 ;
      RECT  105300.0 11250.0 106500.0 12450.0 ;
      RECT  105300.0 1950.0 106500.0 3150.0 ;
      RECT  107700.0 1950.0 108900.0 3150.0 ;
      RECT  107700.0 1950.0 108900.0 3150.0 ;
      RECT  105300.0 1950.0 106500.0 3150.0 ;
      RECT  110100.0 11850.0 111300.0 13050.0 ;
      RECT  110100.0 1950.0 111300.0 3150.0 ;
      RECT  105900.0 6600.0 107100.0 7800.0 ;
      RECT  105900.0 6600.0 107100.0 7800.0 ;
      RECT  108450.0 6750.0 109350.0 7650.0 ;
      RECT  103500.0 13950.0 113100.0 14850.0 ;
      RECT  103500.0 150.0 113100.0 1050.0 ;
      RECT  110100.0 16350.0 111300.0 14400.0 ;
      RECT  110100.0 28200.0 111300.0 26250.0 ;
      RECT  105300.0 26850.0 106500.0 28650.0 ;
      RECT  105300.0 17550.0 106500.0 13950.0 ;
      RECT  108000.0 26850.0 108900.0 17550.0 ;
      RECT  105300.0 17550.0 106500.0 16350.0 ;
      RECT  107700.0 17550.0 108900.0 16350.0 ;
      RECT  107700.0 17550.0 108900.0 16350.0 ;
      RECT  105300.0 17550.0 106500.0 16350.0 ;
      RECT  105300.0 26850.0 106500.0 25650.0 ;
      RECT  107700.0 26850.0 108900.0 25650.0 ;
      RECT  107700.0 26850.0 108900.0 25650.0 ;
      RECT  105300.0 26850.0 106500.0 25650.0 ;
      RECT  110100.0 16950.0 111300.0 15750.0 ;
      RECT  110100.0 26850.0 111300.0 25650.0 ;
      RECT  105900.0 22200.0 107100.0 21000.0 ;
      RECT  105900.0 22200.0 107100.0 21000.0 ;
      RECT  108450.0 22050.0 109350.0 21150.0 ;
      RECT  103500.0 14850.0 113100.0 13950.0 ;
      RECT  103500.0 28650.0 113100.0 27750.0 ;
      RECT  149100.0 12450.0 150300.0 14400.0 ;
      RECT  149100.0 600.0 150300.0 2550.0 ;
      RECT  144300.0 1950.0 145500.0 150.0 ;
      RECT  144300.0 11250.0 145500.0 14850.0 ;
      RECT  147000.0 1950.0 147900.0 11250.0 ;
      RECT  144300.0 11250.0 145500.0 12450.0 ;
      RECT  146700.0 11250.0 147900.0 12450.0 ;
      RECT  146700.0 11250.0 147900.0 12450.0 ;
      RECT  144300.0 11250.0 145500.0 12450.0 ;
      RECT  144300.0 1950.0 145500.0 3150.0 ;
      RECT  146700.0 1950.0 147900.0 3150.0 ;
      RECT  146700.0 1950.0 147900.0 3150.0 ;
      RECT  144300.0 1950.0 145500.0 3150.0 ;
      RECT  149100.0 11850.0 150300.0 13050.0 ;
      RECT  149100.0 1950.0 150300.0 3150.0 ;
      RECT  144900.0 6600.0 146100.0 7800.0 ;
      RECT  144900.0 6600.0 146100.0 7800.0 ;
      RECT  147450.0 6750.0 148350.0 7650.0 ;
      RECT  142500.0 13950.0 152100.0 14850.0 ;
      RECT  142500.0 150.0 152100.0 1050.0 ;
      RECT  149100.0 16350.0 150300.0 14400.0 ;
      RECT  149100.0 28200.0 150300.0 26250.0 ;
      RECT  144300.0 26850.0 145500.0 28650.0 ;
      RECT  144300.0 17550.0 145500.0 13950.0 ;
      RECT  147000.0 26850.0 147900.0 17550.0 ;
      RECT  144300.0 17550.0 145500.0 16350.0 ;
      RECT  146700.0 17550.0 147900.0 16350.0 ;
      RECT  146700.0 17550.0 147900.0 16350.0 ;
      RECT  144300.0 17550.0 145500.0 16350.0 ;
      RECT  144300.0 26850.0 145500.0 25650.0 ;
      RECT  146700.0 26850.0 147900.0 25650.0 ;
      RECT  146700.0 26850.0 147900.0 25650.0 ;
      RECT  144300.0 26850.0 145500.0 25650.0 ;
      RECT  149100.0 16950.0 150300.0 15750.0 ;
      RECT  149100.0 26850.0 150300.0 25650.0 ;
      RECT  144900.0 22200.0 146100.0 21000.0 ;
      RECT  144900.0 22200.0 146100.0 21000.0 ;
      RECT  147450.0 22050.0 148350.0 21150.0 ;
      RECT  142500.0 14850.0 152100.0 13950.0 ;
      RECT  142500.0 28650.0 152100.0 27750.0 ;
      RECT  149100.0 40050.0 150300.0 42000.0 ;
      RECT  149100.0 28200.0 150300.0 30150.0 ;
      RECT  144300.0 29550.0 145500.0 27750.0 ;
      RECT  144300.0 38850.0 145500.0 42450.0 ;
      RECT  147000.0 29550.0 147900.0 38850.0 ;
      RECT  144300.0 38850.0 145500.0 40050.0 ;
      RECT  146700.0 38850.0 147900.0 40050.0 ;
      RECT  146700.0 38850.0 147900.0 40050.0 ;
      RECT  144300.0 38850.0 145500.0 40050.0 ;
      RECT  144300.0 29550.0 145500.0 30750.0 ;
      RECT  146700.0 29550.0 147900.0 30750.0 ;
      RECT  146700.0 29550.0 147900.0 30750.0 ;
      RECT  144300.0 29550.0 145500.0 30750.0 ;
      RECT  149100.0 39450.0 150300.0 40650.0 ;
      RECT  149100.0 29550.0 150300.0 30750.0 ;
      RECT  144900.0 34200.0 146100.0 35400.0 ;
      RECT  144900.0 34200.0 146100.0 35400.0 ;
      RECT  147450.0 34350.0 148350.0 35250.0 ;
      RECT  142500.0 41550.0 152100.0 42450.0 ;
      RECT  142500.0 27750.0 152100.0 28650.0 ;
      RECT  149100.0 43950.0 150300.0 42000.0 ;
      RECT  149100.0 55800.0 150300.0 53850.0 ;
      RECT  144300.0 54450.0 145500.0 56250.0 ;
      RECT  144300.0 45150.0 145500.0 41550.0 ;
      RECT  147000.0 54450.0 147900.0 45150.0 ;
      RECT  144300.0 45150.0 145500.0 43950.0 ;
      RECT  146700.0 45150.0 147900.0 43950.0 ;
      RECT  146700.0 45150.0 147900.0 43950.0 ;
      RECT  144300.0 45150.0 145500.0 43950.0 ;
      RECT  144300.0 54450.0 145500.0 53250.0 ;
      RECT  146700.0 54450.0 147900.0 53250.0 ;
      RECT  146700.0 54450.0 147900.0 53250.0 ;
      RECT  144300.0 54450.0 145500.0 53250.0 ;
      RECT  149100.0 44550.0 150300.0 43350.0 ;
      RECT  149100.0 54450.0 150300.0 53250.0 ;
      RECT  144900.0 49800.0 146100.0 48600.0 ;
      RECT  144900.0 49800.0 146100.0 48600.0 ;
      RECT  147450.0 49650.0 148350.0 48750.0 ;
      RECT  142500.0 42450.0 152100.0 41550.0 ;
      RECT  142500.0 56250.0 152100.0 55350.0 ;
      RECT  129900.0 2550.0 131100.0 150.0 ;
      RECT  129900.0 11250.0 131100.0 14850.0 ;
      RECT  134700.0 11250.0 135900.0 14850.0 ;
      RECT  137100.0 12450.0 138300.0 14400.0 ;
      RECT  137100.0 600.0 138300.0 2550.0 ;
      RECT  129900.0 11250.0 131100.0 12450.0 ;
      RECT  132300.0 11250.0 133500.0 12450.0 ;
      RECT  132300.0 11250.0 133500.0 12450.0 ;
      RECT  129900.0 11250.0 131100.0 12450.0 ;
      RECT  132300.0 11250.0 133500.0 12450.0 ;
      RECT  134700.0 11250.0 135900.0 12450.0 ;
      RECT  134700.0 11250.0 135900.0 12450.0 ;
      RECT  132300.0 11250.0 133500.0 12450.0 ;
      RECT  129900.0 2550.0 131100.0 3750.0 ;
      RECT  132300.0 2550.0 133500.0 3750.0 ;
      RECT  132300.0 2550.0 133500.0 3750.0 ;
      RECT  129900.0 2550.0 131100.0 3750.0 ;
      RECT  132300.0 2550.0 133500.0 3750.0 ;
      RECT  134700.0 2550.0 135900.0 3750.0 ;
      RECT  134700.0 2550.0 135900.0 3750.0 ;
      RECT  132300.0 2550.0 133500.0 3750.0 ;
      RECT  137100.0 11850.0 138300.0 13050.0 ;
      RECT  137100.0 1950.0 138300.0 3150.0 ;
      RECT  134700.0 5100.0 133500.0 6300.0 ;
      RECT  131700.0 7800.0 130500.0 9000.0 ;
      RECT  132300.0 11250.0 133500.0 12450.0 ;
      RECT  134700.0 2550.0 135900.0 3750.0 ;
      RECT  135900.0 7800.0 134700.0 9000.0 ;
      RECT  130500.0 7800.0 131700.0 9000.0 ;
      RECT  133500.0 5100.0 134700.0 6300.0 ;
      RECT  134700.0 7800.0 135900.0 9000.0 ;
      RECT  128100.0 13950.0 142500.0 14850.0 ;
      RECT  128100.0 150.0 142500.0 1050.0 ;
      RECT  129900.0 26250.0 131100.0 28650.0 ;
      RECT  129900.0 17550.0 131100.0 13950.0 ;
      RECT  134700.0 17550.0 135900.0 13950.0 ;
      RECT  137100.0 16350.0 138300.0 14400.0 ;
      RECT  137100.0 28200.0 138300.0 26250.0 ;
      RECT  129900.0 17550.0 131100.0 16350.0 ;
      RECT  132300.0 17550.0 133500.0 16350.0 ;
      RECT  132300.0 17550.0 133500.0 16350.0 ;
      RECT  129900.0 17550.0 131100.0 16350.0 ;
      RECT  132300.0 17550.0 133500.0 16350.0 ;
      RECT  134700.0 17550.0 135900.0 16350.0 ;
      RECT  134700.0 17550.0 135900.0 16350.0 ;
      RECT  132300.0 17550.0 133500.0 16350.0 ;
      RECT  129900.0 26250.0 131100.0 25050.0 ;
      RECT  132300.0 26250.0 133500.0 25050.0 ;
      RECT  132300.0 26250.0 133500.0 25050.0 ;
      RECT  129900.0 26250.0 131100.0 25050.0 ;
      RECT  132300.0 26250.0 133500.0 25050.0 ;
      RECT  134700.0 26250.0 135900.0 25050.0 ;
      RECT  134700.0 26250.0 135900.0 25050.0 ;
      RECT  132300.0 26250.0 133500.0 25050.0 ;
      RECT  137100.0 16950.0 138300.0 15750.0 ;
      RECT  137100.0 26850.0 138300.0 25650.0 ;
      RECT  134700.0 23700.0 133500.0 22500.0 ;
      RECT  131700.0 21000.0 130500.0 19800.0 ;
      RECT  132300.0 17550.0 133500.0 16350.0 ;
      RECT  134700.0 26250.0 135900.0 25050.0 ;
      RECT  135900.0 21000.0 134700.0 19800.0 ;
      RECT  130500.0 21000.0 131700.0 19800.0 ;
      RECT  133500.0 23700.0 134700.0 22500.0 ;
      RECT  134700.0 21000.0 135900.0 19800.0 ;
      RECT  128100.0 14850.0 142500.0 13950.0 ;
      RECT  128100.0 28650.0 142500.0 27750.0 ;
      RECT  129900.0 30150.0 131100.0 27750.0 ;
      RECT  129900.0 38850.0 131100.0 42450.0 ;
      RECT  134700.0 38850.0 135900.0 42450.0 ;
      RECT  137100.0 40050.0 138300.0 42000.0 ;
      RECT  137100.0 28200.0 138300.0 30150.0 ;
      RECT  129900.0 38850.0 131100.0 40050.0 ;
      RECT  132300.0 38850.0 133500.0 40050.0 ;
      RECT  132300.0 38850.0 133500.0 40050.0 ;
      RECT  129900.0 38850.0 131100.0 40050.0 ;
      RECT  132300.0 38850.0 133500.0 40050.0 ;
      RECT  134700.0 38850.0 135900.0 40050.0 ;
      RECT  134700.0 38850.0 135900.0 40050.0 ;
      RECT  132300.0 38850.0 133500.0 40050.0 ;
      RECT  129900.0 30150.0 131100.0 31350.0 ;
      RECT  132300.0 30150.0 133500.0 31350.0 ;
      RECT  132300.0 30150.0 133500.0 31350.0 ;
      RECT  129900.0 30150.0 131100.0 31350.0 ;
      RECT  132300.0 30150.0 133500.0 31350.0 ;
      RECT  134700.0 30150.0 135900.0 31350.0 ;
      RECT  134700.0 30150.0 135900.0 31350.0 ;
      RECT  132300.0 30150.0 133500.0 31350.0 ;
      RECT  137100.0 39450.0 138300.0 40650.0 ;
      RECT  137100.0 29550.0 138300.0 30750.0 ;
      RECT  134700.0 32700.0 133500.0 33900.0 ;
      RECT  131700.0 35400.0 130500.0 36600.0 ;
      RECT  132300.0 38850.0 133500.0 40050.0 ;
      RECT  134700.0 30150.0 135900.0 31350.0 ;
      RECT  135900.0 35400.0 134700.0 36600.0 ;
      RECT  130500.0 35400.0 131700.0 36600.0 ;
      RECT  133500.0 32700.0 134700.0 33900.0 ;
      RECT  134700.0 35400.0 135900.0 36600.0 ;
      RECT  128100.0 41550.0 142500.0 42450.0 ;
      RECT  128100.0 27750.0 142500.0 28650.0 ;
      RECT  129900.0 53850.0 131100.0 56250.0 ;
      RECT  129900.0 45150.0 131100.0 41550.0 ;
      RECT  134700.0 45150.0 135900.0 41550.0 ;
      RECT  137100.0 43950.0 138300.0 42000.0 ;
      RECT  137100.0 55800.0 138300.0 53850.0 ;
      RECT  129900.0 45150.0 131100.0 43950.0 ;
      RECT  132300.0 45150.0 133500.0 43950.0 ;
      RECT  132300.0 45150.0 133500.0 43950.0 ;
      RECT  129900.0 45150.0 131100.0 43950.0 ;
      RECT  132300.0 45150.0 133500.0 43950.0 ;
      RECT  134700.0 45150.0 135900.0 43950.0 ;
      RECT  134700.0 45150.0 135900.0 43950.0 ;
      RECT  132300.0 45150.0 133500.0 43950.0 ;
      RECT  129900.0 53850.0 131100.0 52650.0 ;
      RECT  132300.0 53850.0 133500.0 52650.0 ;
      RECT  132300.0 53850.0 133500.0 52650.0 ;
      RECT  129900.0 53850.0 131100.0 52650.0 ;
      RECT  132300.0 53850.0 133500.0 52650.0 ;
      RECT  134700.0 53850.0 135900.0 52650.0 ;
      RECT  134700.0 53850.0 135900.0 52650.0 ;
      RECT  132300.0 53850.0 133500.0 52650.0 ;
      RECT  137100.0 44550.0 138300.0 43350.0 ;
      RECT  137100.0 54450.0 138300.0 53250.0 ;
      RECT  134700.0 51300.0 133500.0 50100.0 ;
      RECT  131700.0 48600.0 130500.0 47400.0 ;
      RECT  132300.0 45150.0 133500.0 43950.0 ;
      RECT  134700.0 53850.0 135900.0 52650.0 ;
      RECT  135900.0 48600.0 134700.0 47400.0 ;
      RECT  130500.0 48600.0 131700.0 47400.0 ;
      RECT  133500.0 51300.0 134700.0 50100.0 ;
      RECT  134700.0 48600.0 135900.0 47400.0 ;
      RECT  128100.0 42450.0 142500.0 41550.0 ;
      RECT  128100.0 56250.0 142500.0 55350.0 ;
      RECT  117150.0 11100.0 115950.0 12300.0 ;
      RECT  98550.0 6600.0 97350.0 7800.0 ;
      RECT  120150.0 24900.0 118950.0 26100.0 ;
      RECT  101550.0 21000.0 100350.0 22200.0 ;
      RECT  98550.0 29700.0 97350.0 30900.0 ;
      RECT  123150.0 29700.0 121950.0 30900.0 ;
      RECT  101550.0 43500.0 100350.0 44700.0 ;
      RECT  126150.0 43500.0 124950.0 44700.0 ;
      RECT  117150.0 7800.0 115950.0 9000.0 ;
      RECT  120150.0 5100.0 118950.0 6300.0 ;
      RECT  123150.0 19800.0 121950.0 21000.0 ;
      RECT  120150.0 22500.0 118950.0 23700.0 ;
      RECT  117150.0 35400.0 115950.0 36600.0 ;
      RECT  126150.0 32700.0 124950.0 33900.0 ;
      RECT  123150.0 47400.0 121950.0 48600.0 ;
      RECT  126150.0 50100.0 124950.0 51300.0 ;
      RECT  148350.0 6750.0 152100.0 7650.0 ;
      RECT  148350.0 21150.0 152100.0 22050.0 ;
      RECT  148350.0 34350.0 152100.0 35250.0 ;
      RECT  148350.0 48750.0 152100.0 49650.0 ;
      RECT  97500.0 13950.0 152100.0 14850.0 ;
      RECT  97500.0 41550.0 152100.0 42450.0 ;
      RECT  97500.0 150.0 152100.0 1050.0 ;
      RECT  97500.0 27750.0 152100.0 28650.0 ;
      RECT  97500.0 55350.0 152100.0 56250.0 ;
      RECT  221400.0 289650.0 231600.0 338550.0 ;
      RECT  262200.0 289650.0 272400.0 338550.0 ;
      RECT  303000.0 289650.0 313200.0 338550.0 ;
      RECT  343800.0 289650.0 354000.0 338550.0 ;
      RECT  384600.0 289650.0 394800.0 338550.0 ;
      RECT  425400.0 289650.0 435600.0 338550.0 ;
      RECT  466200.0 289650.0 476400.0 338550.0 ;
      RECT  507000.0 289650.0 517200.0 338550.0 ;
      RECT  547800.0 289650.0 558000.0 338550.0 ;
      RECT  588600.0 289650.0 598800.0 338550.0 ;
      RECT  629400.0 289650.0 639600.0 338550.0 ;
      RECT  670200.0 289650.0 680400.0 338550.0 ;
      RECT  711000.0 289650.0 721200.0 338550.0 ;
      RECT  751800.0 289650.0 762000.0 338550.0 ;
      RECT  792600.0 289650.0 802800.0 338550.0 ;
      RECT  833400.0 289650.0 843600.0 338550.0 ;
      RECT  874200.0 289650.0 884400.0 338550.0 ;
      RECT  915000.0 289650.0 925200.0 338550.0 ;
      RECT  955800.0 289650.0 966000.0 338550.0 ;
      RECT  996600.0 289650.0 1006800.0 338550.0 ;
      RECT  1037400.0 289650.0 1047600.0 338550.0 ;
      RECT  1078200.0 289650.0 1088400.0 338550.0 ;
      RECT  1119000.0 289650.0 1129200.0 338550.0 ;
      RECT  1159800.0 289650.0 1170000.0 338550.0 ;
      RECT  1200600.0 289650.0 1210800.0 338550.0 ;
      RECT  1241400.0 289650.0 1251600.0 338550.0 ;
      RECT  1282200.0 289650.0 1292400.0 338550.0 ;
      RECT  1323000.0 289650.0 1333200.0 338550.0 ;
      RECT  1363800.0 289650.0 1374000.0 338550.0 ;
      RECT  1404600.0 289650.0 1414800.0 338550.0 ;
      RECT  1445400.0 289650.0 1455600.0 338550.0 ;
      RECT  1486200.0 289650.0 1496400.0 338550.0 ;
      RECT  221400.0 334350.0 1527000.0 335250.0 ;
      RECT  221400.0 307050.0 1527000.0 307950.0 ;
      RECT  221400.0 332250.0 1527000.0 333150.0 ;
      RECT  221400.0 229050.0 231600.0 289650.0 ;
      RECT  262200.0 229050.0 272400.0 289650.0 ;
      RECT  303000.0 229050.0 313200.0 289650.0 ;
      RECT  343800.0 229050.0 354000.0 289650.0 ;
      RECT  384600.0 229050.0 394800.0 289650.0 ;
      RECT  425400.0 229050.0 435600.0 289650.0 ;
      RECT  466200.0 229050.0 476400.0 289650.0 ;
      RECT  507000.0 229050.0 517200.0 289650.0 ;
      RECT  547800.0 229050.0 558000.0 289650.0 ;
      RECT  588600.0 229050.0 598800.0 289650.0 ;
      RECT  629400.0 229050.0 639600.0 289650.0 ;
      RECT  670200.0 229050.0 680400.0 289650.0 ;
      RECT  711000.0 229050.0 721200.0 289650.0 ;
      RECT  751800.0 229050.0 762000.0 289650.0 ;
      RECT  792600.0 229050.0 802800.0 289650.0 ;
      RECT  833400.0 229050.0 843600.0 289650.0 ;
      RECT  874200.0 229050.0 884400.0 289650.0 ;
      RECT  915000.0 229050.0 925200.0 289650.0 ;
      RECT  955800.0 229050.0 966000.0 289650.0 ;
      RECT  996600.0 229050.0 1006800.0 289650.0 ;
      RECT  1037400.0 229050.0 1047600.0 289650.0 ;
      RECT  1078200.0 229050.0 1088400.0 289650.0 ;
      RECT  1119000.0 229050.0 1129200.0 289650.0 ;
      RECT  1159800.0 229050.0 1170000.0 289650.0 ;
      RECT  1200600.0 229050.0 1210800.0 289650.0 ;
      RECT  1241400.0 229050.0 1251600.0 289650.0 ;
      RECT  1282200.0 229050.0 1292400.0 289650.0 ;
      RECT  1323000.0 229050.0 1333200.0 289650.0 ;
      RECT  1363800.0 229050.0 1374000.0 289650.0 ;
      RECT  1404600.0 229050.0 1414800.0 289650.0 ;
      RECT  1445400.0 229050.0 1455600.0 289650.0 ;
      RECT  1486200.0 229050.0 1496400.0 289650.0 ;
      RECT  221400.0 236250.0 1527000.0 237150.0 ;
      RECT  221400.0 238350.0 1527000.0 239250.0 ;
      RECT  221400.0 234150.0 1527000.0 235050.0 ;
      RECT  221400.0 169050.0 231600.0 229050.0 ;
      RECT  262200.0 169050.0 272400.0 229050.0 ;
      RECT  303000.0 169050.0 313200.0 229050.0 ;
      RECT  343800.0 169050.0 354000.0 229050.0 ;
      RECT  384600.0 169050.0 394800.0 229050.0 ;
      RECT  425400.0 169050.0 435600.0 229050.0 ;
      RECT  466200.0 169050.0 476400.0 229050.0 ;
      RECT  507000.0 169050.0 517200.0 229050.0 ;
      RECT  547800.0 169050.0 558000.0 229050.0 ;
      RECT  588600.0 169050.0 598800.0 229050.0 ;
      RECT  629400.0 169050.0 639600.0 229050.0 ;
      RECT  670200.0 169050.0 680400.0 229050.0 ;
      RECT  711000.0 169050.0 721200.0 229050.0 ;
      RECT  751800.0 169050.0 762000.0 229050.0 ;
      RECT  792600.0 169050.0 802800.0 229050.0 ;
      RECT  833400.0 169050.0 843600.0 229050.0 ;
      RECT  874200.0 169050.0 884400.0 229050.0 ;
      RECT  915000.0 169050.0 925200.0 229050.0 ;
      RECT  955800.0 169050.0 966000.0 229050.0 ;
      RECT  996600.0 169050.0 1006800.0 229050.0 ;
      RECT  1037400.0 169050.0 1047600.0 229050.0 ;
      RECT  1078200.0 169050.0 1088400.0 229050.0 ;
      RECT  1119000.0 169050.0 1129200.0 229050.0 ;
      RECT  1159800.0 169050.0 1170000.0 229050.0 ;
      RECT  1200600.0 169050.0 1210800.0 229050.0 ;
      RECT  1241400.0 169050.0 1251600.0 229050.0 ;
      RECT  1282200.0 169050.0 1292400.0 229050.0 ;
      RECT  1323000.0 169050.0 1333200.0 229050.0 ;
      RECT  1363800.0 169050.0 1374000.0 229050.0 ;
      RECT  1404600.0 169050.0 1414800.0 229050.0 ;
      RECT  1445400.0 169050.0 1455600.0 229050.0 ;
      RECT  1486200.0 169050.0 1496400.0 229050.0 ;
      RECT  221400.0 171450.0 1527000.0 172350.0 ;
      RECT  221400.0 225450.0 1527000.0 226350.0 ;
      RECT  221400.0 169050.0 231600.0 147150.0 ;
      RECT  262200.0 169050.0 272400.0 147150.0 ;
      RECT  303000.0 169050.0 313200.0 147150.0 ;
      RECT  343800.0 169050.0 354000.0 147150.0 ;
      RECT  384600.0 169050.0 394800.0 147150.0 ;
      RECT  425400.0 169050.0 435600.0 147150.0 ;
      RECT  466200.0 169050.0 476400.0 147150.0 ;
      RECT  507000.0 169050.0 517200.0 147150.0 ;
      RECT  547800.0 169050.0 558000.0 147150.0 ;
      RECT  588600.0 169050.0 598800.0 147150.0 ;
      RECT  629400.0 169050.0 639600.0 147150.0 ;
      RECT  670200.0 169050.0 680400.0 147150.0 ;
      RECT  711000.0 169050.0 721200.0 147150.0 ;
      RECT  751800.0 169050.0 762000.0 147150.0 ;
      RECT  792600.0 169050.0 802800.0 147150.0 ;
      RECT  833400.0 169050.0 843600.0 147150.0 ;
      RECT  874200.0 169050.0 884400.0 147150.0 ;
      RECT  915000.0 169050.0 925200.0 147150.0 ;
      RECT  955800.0 169050.0 966000.0 147150.0 ;
      RECT  996600.0 169050.0 1006800.0 147150.0 ;
      RECT  1037400.0 169050.0 1047600.0 147150.0 ;
      RECT  1078200.0 169050.0 1088400.0 147150.0 ;
      RECT  1119000.0 169050.0 1129200.0 147150.0 ;
      RECT  1159800.0 169050.0 1170000.0 147150.0 ;
      RECT  1200600.0 169050.0 1210800.0 147150.0 ;
      RECT  1241400.0 169050.0 1251600.0 147150.0 ;
      RECT  1282200.0 169050.0 1292400.0 147150.0 ;
      RECT  1323000.0 169050.0 1333200.0 147150.0 ;
      RECT  1363800.0 169050.0 1374000.0 147150.0 ;
      RECT  1404600.0 169050.0 1414800.0 147150.0 ;
      RECT  1445400.0 169050.0 1455600.0 147150.0 ;
      RECT  1486200.0 169050.0 1496400.0 147150.0 ;
      RECT  221400.0 165450.0 1496400.0 164550.0 ;
      RECT  221400.0 167850.0 1496400.0 166950.0 ;
      RECT  221400.0 149550.0 1496400.0 148650.0 ;
      RECT  221400.0 163350.0 1496400.0 162450.0 ;
      RECT  106350.0 387300.0 107250.0 388200.0 ;
      RECT  106350.0 385350.0 107250.0 386250.0 ;
      RECT  102900.0 387300.0 106800.0 388200.0 ;
      RECT  106350.0 385800.0 107250.0 387750.0 ;
      RECT  106800.0 385350.0 110700.0 386250.0 ;
      RECT  106350.0 397800.0 107250.0 398700.0 ;
      RECT  106350.0 399750.0 107250.0 400650.0 ;
      RECT  102900.0 397800.0 106800.0 398700.0 ;
      RECT  106350.0 398250.0 107250.0 400200.0 ;
      RECT  106800.0 399750.0 110700.0 400650.0 ;
      RECT  106350.0 414900.0 107250.0 415800.0 ;
      RECT  106350.0 412950.0 107250.0 413850.0 ;
      RECT  102900.0 414900.0 106800.0 415800.0 ;
      RECT  106350.0 413400.0 107250.0 415350.0 ;
      RECT  106800.0 412950.0 110700.0 413850.0 ;
      RECT  106350.0 425400.0 107250.0 426300.0 ;
      RECT  106350.0 427350.0 107250.0 428250.0 ;
      RECT  102900.0 425400.0 106800.0 426300.0 ;
      RECT  106350.0 425850.0 107250.0 427800.0 ;
      RECT  106800.0 427350.0 110700.0 428250.0 ;
      RECT  106350.0 442500.0 107250.0 443400.0 ;
      RECT  106350.0 440550.0 107250.0 441450.0 ;
      RECT  102900.0 442500.0 106800.0 443400.0 ;
      RECT  106350.0 441000.0 107250.0 442950.0 ;
      RECT  106800.0 440550.0 110700.0 441450.0 ;
      RECT  106350.0 453000.0 107250.0 453900.0 ;
      RECT  106350.0 454950.0 107250.0 455850.0 ;
      RECT  102900.0 453000.0 106800.0 453900.0 ;
      RECT  106350.0 453450.0 107250.0 455400.0 ;
      RECT  106800.0 454950.0 110700.0 455850.0 ;
      RECT  106350.0 470100.0 107250.0 471000.0 ;
      RECT  106350.0 468150.0 107250.0 469050.0 ;
      RECT  102900.0 470100.0 106800.0 471000.0 ;
      RECT  106350.0 468600.0 107250.0 470550.0 ;
      RECT  106800.0 468150.0 110700.0 469050.0 ;
      RECT  106350.0 480600.0 107250.0 481500.0 ;
      RECT  106350.0 482550.0 107250.0 483450.0 ;
      RECT  102900.0 480600.0 106800.0 481500.0 ;
      RECT  106350.0 481050.0 107250.0 483000.0 ;
      RECT  106800.0 482550.0 110700.0 483450.0 ;
      RECT  106350.0 497700.0 107250.0 498600.0 ;
      RECT  106350.0 495750.0 107250.0 496650.0 ;
      RECT  102900.0 497700.0 106800.0 498600.0 ;
      RECT  106350.0 496200.0 107250.0 498150.0 ;
      RECT  106800.0 495750.0 110700.0 496650.0 ;
      RECT  106350.0 508200.0 107250.0 509100.0 ;
      RECT  106350.0 510150.0 107250.0 511050.0 ;
      RECT  102900.0 508200.0 106800.0 509100.0 ;
      RECT  106350.0 508650.0 107250.0 510600.0 ;
      RECT  106800.0 510150.0 110700.0 511050.0 ;
      RECT  106350.0 525300.0 107250.0 526200.0 ;
      RECT  106350.0 523350.0 107250.0 524250.0 ;
      RECT  102900.0 525300.0 106800.0 526200.0 ;
      RECT  106350.0 523800.0 107250.0 525750.0 ;
      RECT  106800.0 523350.0 110700.0 524250.0 ;
      RECT  106350.0 535800.0 107250.0 536700.0 ;
      RECT  106350.0 537750.0 107250.0 538650.0 ;
      RECT  102900.0 535800.0 106800.0 536700.0 ;
      RECT  106350.0 536250.0 107250.0 538200.0 ;
      RECT  106800.0 537750.0 110700.0 538650.0 ;
      RECT  106350.0 552900.0 107250.0 553800.0 ;
      RECT  106350.0 550950.0 107250.0 551850.0 ;
      RECT  102900.0 552900.0 106800.0 553800.0 ;
      RECT  106350.0 551400.0 107250.0 553350.0 ;
      RECT  106800.0 550950.0 110700.0 551850.0 ;
      RECT  106350.0 563400.0 107250.0 564300.0 ;
      RECT  106350.0 565350.0 107250.0 566250.0 ;
      RECT  102900.0 563400.0 106800.0 564300.0 ;
      RECT  106350.0 563850.0 107250.0 565800.0 ;
      RECT  106800.0 565350.0 110700.0 566250.0 ;
      RECT  106350.0 580500.0 107250.0 581400.0 ;
      RECT  106350.0 578550.0 107250.0 579450.0 ;
      RECT  102900.0 580500.0 106800.0 581400.0 ;
      RECT  106350.0 579000.0 107250.0 580950.0 ;
      RECT  106800.0 578550.0 110700.0 579450.0 ;
      RECT  106350.0 591000.0 107250.0 591900.0 ;
      RECT  106350.0 592950.0 107250.0 593850.0 ;
      RECT  102900.0 591000.0 106800.0 591900.0 ;
      RECT  106350.0 591450.0 107250.0 593400.0 ;
      RECT  106800.0 592950.0 110700.0 593850.0 ;
      RECT  106350.0 608100.0 107250.0 609000.0 ;
      RECT  106350.0 606150.0 107250.0 607050.0 ;
      RECT  102900.0 608100.0 106800.0 609000.0 ;
      RECT  106350.0 606600.0 107250.0 608550.0 ;
      RECT  106800.0 606150.0 110700.0 607050.0 ;
      RECT  106350.0 618600.0 107250.0 619500.0 ;
      RECT  106350.0 620550.0 107250.0 621450.0 ;
      RECT  102900.0 618600.0 106800.0 619500.0 ;
      RECT  106350.0 619050.0 107250.0 621000.0 ;
      RECT  106800.0 620550.0 110700.0 621450.0 ;
      RECT  106350.0 635700.0 107250.0 636600.0 ;
      RECT  106350.0 633750.0 107250.0 634650.0 ;
      RECT  102900.0 635700.0 106800.0 636600.0 ;
      RECT  106350.0 634200.0 107250.0 636150.0 ;
      RECT  106800.0 633750.0 110700.0 634650.0 ;
      RECT  106350.0 646200.0 107250.0 647100.0 ;
      RECT  106350.0 648150.0 107250.0 649050.0 ;
      RECT  102900.0 646200.0 106800.0 647100.0 ;
      RECT  106350.0 646650.0 107250.0 648600.0 ;
      RECT  106800.0 648150.0 110700.0 649050.0 ;
      RECT  106350.0 663300.0 107250.0 664200.0 ;
      RECT  106350.0 661350.0 107250.0 662250.0 ;
      RECT  102900.0 663300.0 106800.0 664200.0 ;
      RECT  106350.0 661800.0 107250.0 663750.0 ;
      RECT  106800.0 661350.0 110700.0 662250.0 ;
      RECT  106350.0 673800.0 107250.0 674700.0 ;
      RECT  106350.0 675750.0 107250.0 676650.0 ;
      RECT  102900.0 673800.0 106800.0 674700.0 ;
      RECT  106350.0 674250.0 107250.0 676200.0 ;
      RECT  106800.0 675750.0 110700.0 676650.0 ;
      RECT  106350.0 690900.0 107250.0 691800.0 ;
      RECT  106350.0 688950.0 107250.0 689850.0 ;
      RECT  102900.0 690900.0 106800.0 691800.0 ;
      RECT  106350.0 689400.0 107250.0 691350.0 ;
      RECT  106800.0 688950.0 110700.0 689850.0 ;
      RECT  106350.0 701400.0 107250.0 702300.0 ;
      RECT  106350.0 703350.0 107250.0 704250.0 ;
      RECT  102900.0 701400.0 106800.0 702300.0 ;
      RECT  106350.0 701850.0 107250.0 703800.0 ;
      RECT  106800.0 703350.0 110700.0 704250.0 ;
      RECT  106350.0 718500.0 107250.0 719400.0 ;
      RECT  106350.0 716550.0 107250.0 717450.0 ;
      RECT  102900.0 718500.0 106800.0 719400.0 ;
      RECT  106350.0 717000.0 107250.0 718950.0 ;
      RECT  106800.0 716550.0 110700.0 717450.0 ;
      RECT  106350.0 729000.0 107250.0 729900.0 ;
      RECT  106350.0 730950.0 107250.0 731850.0 ;
      RECT  102900.0 729000.0 106800.0 729900.0 ;
      RECT  106350.0 729450.0 107250.0 731400.0 ;
      RECT  106800.0 730950.0 110700.0 731850.0 ;
      RECT  106350.0 746100.0 107250.0 747000.0 ;
      RECT  106350.0 744150.0 107250.0 745050.0 ;
      RECT  102900.0 746100.0 106800.0 747000.0 ;
      RECT  106350.0 744600.0 107250.0 746550.0 ;
      RECT  106800.0 744150.0 110700.0 745050.0 ;
      RECT  106350.0 756600.0 107250.0 757500.0 ;
      RECT  106350.0 758550.0 107250.0 759450.0 ;
      RECT  102900.0 756600.0 106800.0 757500.0 ;
      RECT  106350.0 757050.0 107250.0 759000.0 ;
      RECT  106800.0 758550.0 110700.0 759450.0 ;
      RECT  106350.0 773700.0 107250.0 774600.0 ;
      RECT  106350.0 771750.0 107250.0 772650.0 ;
      RECT  102900.0 773700.0 106800.0 774600.0 ;
      RECT  106350.0 772200.0 107250.0 774150.0 ;
      RECT  106800.0 771750.0 110700.0 772650.0 ;
      RECT  106350.0 784200.0 107250.0 785100.0 ;
      RECT  106350.0 786150.0 107250.0 787050.0 ;
      RECT  102900.0 784200.0 106800.0 785100.0 ;
      RECT  106350.0 784650.0 107250.0 786600.0 ;
      RECT  106800.0 786150.0 110700.0 787050.0 ;
      RECT  106350.0 801300.0 107250.0 802200.0 ;
      RECT  106350.0 799350.0 107250.0 800250.0 ;
      RECT  102900.0 801300.0 106800.0 802200.0 ;
      RECT  106350.0 799800.0 107250.0 801750.0 ;
      RECT  106800.0 799350.0 110700.0 800250.0 ;
      RECT  106350.0 811800.0 107250.0 812700.0 ;
      RECT  106350.0 813750.0 107250.0 814650.0 ;
      RECT  102900.0 811800.0 106800.0 812700.0 ;
      RECT  106350.0 812250.0 107250.0 814200.0 ;
      RECT  106800.0 813750.0 110700.0 814650.0 ;
      RECT  106350.0 828900.0 107250.0 829800.0 ;
      RECT  106350.0 826950.0 107250.0 827850.0 ;
      RECT  102900.0 828900.0 106800.0 829800.0 ;
      RECT  106350.0 827400.0 107250.0 829350.0 ;
      RECT  106800.0 826950.0 110700.0 827850.0 ;
      RECT  106350.0 839400.0 107250.0 840300.0 ;
      RECT  106350.0 841350.0 107250.0 842250.0 ;
      RECT  102900.0 839400.0 106800.0 840300.0 ;
      RECT  106350.0 839850.0 107250.0 841800.0 ;
      RECT  106800.0 841350.0 110700.0 842250.0 ;
      RECT  106350.0 856500.0 107250.0 857400.0 ;
      RECT  106350.0 854550.0 107250.0 855450.0 ;
      RECT  102900.0 856500.0 106800.0 857400.0 ;
      RECT  106350.0 855000.0 107250.0 856950.0 ;
      RECT  106800.0 854550.0 110700.0 855450.0 ;
      RECT  106350.0 867000.0 107250.0 867900.0 ;
      RECT  106350.0 868950.0 107250.0 869850.0 ;
      RECT  102900.0 867000.0 106800.0 867900.0 ;
      RECT  106350.0 867450.0 107250.0 869400.0 ;
      RECT  106800.0 868950.0 110700.0 869850.0 ;
      RECT  106350.0 884100.0 107250.0 885000.0 ;
      RECT  106350.0 882150.0 107250.0 883050.0 ;
      RECT  102900.0 884100.0 106800.0 885000.0 ;
      RECT  106350.0 882600.0 107250.0 884550.0 ;
      RECT  106800.0 882150.0 110700.0 883050.0 ;
      RECT  106350.0 894600.0 107250.0 895500.0 ;
      RECT  106350.0 896550.0 107250.0 897450.0 ;
      RECT  102900.0 894600.0 106800.0 895500.0 ;
      RECT  106350.0 895050.0 107250.0 897000.0 ;
      RECT  106800.0 896550.0 110700.0 897450.0 ;
      RECT  106350.0 911700.0 107250.0 912600.0 ;
      RECT  106350.0 909750.0 107250.0 910650.0 ;
      RECT  102900.0 911700.0 106800.0 912600.0 ;
      RECT  106350.0 910200.0 107250.0 912150.0 ;
      RECT  106800.0 909750.0 110700.0 910650.0 ;
      RECT  106350.0 922200.0 107250.0 923100.0 ;
      RECT  106350.0 924150.0 107250.0 925050.0 ;
      RECT  102900.0 922200.0 106800.0 923100.0 ;
      RECT  106350.0 922650.0 107250.0 924600.0 ;
      RECT  106800.0 924150.0 110700.0 925050.0 ;
      RECT  106350.0 939300.0 107250.0 940200.0 ;
      RECT  106350.0 937350.0 107250.0 938250.0 ;
      RECT  102900.0 939300.0 106800.0 940200.0 ;
      RECT  106350.0 937800.0 107250.0 939750.0 ;
      RECT  106800.0 937350.0 110700.0 938250.0 ;
      RECT  106350.0 949800.0 107250.0 950700.0 ;
      RECT  106350.0 951750.0 107250.0 952650.0 ;
      RECT  102900.0 949800.0 106800.0 950700.0 ;
      RECT  106350.0 950250.0 107250.0 952200.0 ;
      RECT  106800.0 951750.0 110700.0 952650.0 ;
      RECT  106350.0 966900.0 107250.0 967800.0 ;
      RECT  106350.0 964950.0 107250.0 965850.0 ;
      RECT  102900.0 966900.0 106800.0 967800.0 ;
      RECT  106350.0 965400.0 107250.0 967350.0 ;
      RECT  106800.0 964950.0 110700.0 965850.0 ;
      RECT  106350.0 977400.0 107250.0 978300.0 ;
      RECT  106350.0 979350.0 107250.0 980250.0 ;
      RECT  102900.0 977400.0 106800.0 978300.0 ;
      RECT  106350.0 977850.0 107250.0 979800.0 ;
      RECT  106800.0 979350.0 110700.0 980250.0 ;
      RECT  106350.0 994500.0 107250.0 995400.0 ;
      RECT  106350.0 992550.0 107250.0 993450.0 ;
      RECT  102900.0 994500.0 106800.0 995400.0 ;
      RECT  106350.0 993000.0 107250.0 994950.0 ;
      RECT  106800.0 992550.0 110700.0 993450.0 ;
      RECT  106350.0 1005000.0 107250.0 1005900.0 ;
      RECT  106350.0 1006950.0 107250.0 1007850.0 ;
      RECT  102900.0 1005000.0 106800.0 1005900.0 ;
      RECT  106350.0 1005450.0 107250.0 1007400.0 ;
      RECT  106800.0 1006950.0 110700.0 1007850.0 ;
      RECT  106350.0 1022100.0 107250.0 1023000.0 ;
      RECT  106350.0 1020150.0 107250.0 1021050.0 ;
      RECT  102900.0 1022100.0 106800.0 1023000.0 ;
      RECT  106350.0 1020600.0 107250.0 1022550.0 ;
      RECT  106800.0 1020150.0 110700.0 1021050.0 ;
      RECT  106350.0 1032600.0 107250.0 1033500.0 ;
      RECT  106350.0 1034550.0 107250.0 1035450.0 ;
      RECT  102900.0 1032600.0 106800.0 1033500.0 ;
      RECT  106350.0 1033050.0 107250.0 1035000.0 ;
      RECT  106800.0 1034550.0 110700.0 1035450.0 ;
      RECT  106350.0 1049700.0 107250.0 1050600.0 ;
      RECT  106350.0 1047750.0 107250.0 1048650.0 ;
      RECT  102900.0 1049700.0 106800.0 1050600.0 ;
      RECT  106350.0 1048200.0 107250.0 1050150.0 ;
      RECT  106800.0 1047750.0 110700.0 1048650.0 ;
      RECT  106350.0 1060200.0 107250.0 1061100.0 ;
      RECT  106350.0 1062150.0 107250.0 1063050.0 ;
      RECT  102900.0 1060200.0 106800.0 1061100.0 ;
      RECT  106350.0 1060650.0 107250.0 1062600.0 ;
      RECT  106800.0 1062150.0 110700.0 1063050.0 ;
      RECT  106350.0 1077300.0 107250.0 1078200.0 ;
      RECT  106350.0 1075350.0 107250.0 1076250.0 ;
      RECT  102900.0 1077300.0 106800.0 1078200.0 ;
      RECT  106350.0 1075800.0 107250.0 1077750.0 ;
      RECT  106800.0 1075350.0 110700.0 1076250.0 ;
      RECT  106350.0 1087800.0 107250.0 1088700.0 ;
      RECT  106350.0 1089750.0 107250.0 1090650.0 ;
      RECT  102900.0 1087800.0 106800.0 1088700.0 ;
      RECT  106350.0 1088250.0 107250.0 1090200.0 ;
      RECT  106800.0 1089750.0 110700.0 1090650.0 ;
      RECT  106350.0 1104900.0 107250.0 1105800.0 ;
      RECT  106350.0 1102950.0 107250.0 1103850.0 ;
      RECT  102900.0 1104900.0 106800.0 1105800.0 ;
      RECT  106350.0 1103400.0 107250.0 1105350.0 ;
      RECT  106800.0 1102950.0 110700.0 1103850.0 ;
      RECT  106350.0 1115400.0 107250.0 1116300.0 ;
      RECT  106350.0 1117350.0 107250.0 1118250.0 ;
      RECT  102900.0 1115400.0 106800.0 1116300.0 ;
      RECT  106350.0 1115850.0 107250.0 1117800.0 ;
      RECT  106800.0 1117350.0 110700.0 1118250.0 ;
      RECT  106350.0 1132500.0 107250.0 1133400.0 ;
      RECT  106350.0 1130550.0 107250.0 1131450.0 ;
      RECT  102900.0 1132500.0 106800.0 1133400.0 ;
      RECT  106350.0 1131000.0 107250.0 1132950.0 ;
      RECT  106800.0 1130550.0 110700.0 1131450.0 ;
      RECT  106350.0 1143000.0 107250.0 1143900.0 ;
      RECT  106350.0 1144950.0 107250.0 1145850.0 ;
      RECT  102900.0 1143000.0 106800.0 1143900.0 ;
      RECT  106350.0 1143450.0 107250.0 1145400.0 ;
      RECT  106800.0 1144950.0 110700.0 1145850.0 ;
      RECT  106350.0 1160100.0 107250.0 1161000.0 ;
      RECT  106350.0 1158150.0 107250.0 1159050.0 ;
      RECT  102900.0 1160100.0 106800.0 1161000.0 ;
      RECT  106350.0 1158600.0 107250.0 1160550.0 ;
      RECT  106800.0 1158150.0 110700.0 1159050.0 ;
      RECT  106350.0 1170600.0 107250.0 1171500.0 ;
      RECT  106350.0 1172550.0 107250.0 1173450.0 ;
      RECT  102900.0 1170600.0 106800.0 1171500.0 ;
      RECT  106350.0 1171050.0 107250.0 1173000.0 ;
      RECT  106800.0 1172550.0 110700.0 1173450.0 ;
      RECT  106350.0 1187700.0 107250.0 1188600.0 ;
      RECT  106350.0 1185750.0 107250.0 1186650.0 ;
      RECT  102900.0 1187700.0 106800.0 1188600.0 ;
      RECT  106350.0 1186200.0 107250.0 1188150.0 ;
      RECT  106800.0 1185750.0 110700.0 1186650.0 ;
      RECT  106350.0 1198200.0 107250.0 1199100.0 ;
      RECT  106350.0 1200150.0 107250.0 1201050.0 ;
      RECT  102900.0 1198200.0 106800.0 1199100.0 ;
      RECT  106350.0 1198650.0 107250.0 1200600.0 ;
      RECT  106800.0 1200150.0 110700.0 1201050.0 ;
      RECT  106350.0 1215300.0 107250.0 1216200.0 ;
      RECT  106350.0 1213350.0 107250.0 1214250.0 ;
      RECT  102900.0 1215300.0 106800.0 1216200.0 ;
      RECT  106350.0 1213800.0 107250.0 1215750.0 ;
      RECT  106800.0 1213350.0 110700.0 1214250.0 ;
      RECT  106350.0 1225800.0 107250.0 1226700.0 ;
      RECT  106350.0 1227750.0 107250.0 1228650.0 ;
      RECT  102900.0 1225800.0 106800.0 1226700.0 ;
      RECT  106350.0 1226250.0 107250.0 1228200.0 ;
      RECT  106800.0 1227750.0 110700.0 1228650.0 ;
      RECT  106350.0 1242900.0 107250.0 1243800.0 ;
      RECT  106350.0 1240950.0 107250.0 1241850.0 ;
      RECT  102900.0 1242900.0 106800.0 1243800.0 ;
      RECT  106350.0 1241400.0 107250.0 1243350.0 ;
      RECT  106800.0 1240950.0 110700.0 1241850.0 ;
      RECT  106350.0 1253400.0 107250.0 1254300.0 ;
      RECT  106350.0 1255350.0 107250.0 1256250.0 ;
      RECT  102900.0 1253400.0 106800.0 1254300.0 ;
      RECT  106350.0 1253850.0 107250.0 1255800.0 ;
      RECT  106800.0 1255350.0 110700.0 1256250.0 ;
      RECT  106350.0 1270500.0 107250.0 1271400.0 ;
      RECT  106350.0 1268550.0 107250.0 1269450.0 ;
      RECT  102900.0 1270500.0 106800.0 1271400.0 ;
      RECT  106350.0 1269000.0 107250.0 1270950.0 ;
      RECT  106800.0 1268550.0 110700.0 1269450.0 ;
      RECT  106350.0 1281000.0 107250.0 1281900.0 ;
      RECT  106350.0 1282950.0 107250.0 1283850.0 ;
      RECT  102900.0 1281000.0 106800.0 1281900.0 ;
      RECT  106350.0 1281450.0 107250.0 1283400.0 ;
      RECT  106800.0 1282950.0 110700.0 1283850.0 ;
      RECT  106350.0 1298100.0 107250.0 1299000.0 ;
      RECT  106350.0 1296150.0 107250.0 1297050.0 ;
      RECT  102900.0 1298100.0 106800.0 1299000.0 ;
      RECT  106350.0 1296600.0 107250.0 1298550.0 ;
      RECT  106800.0 1296150.0 110700.0 1297050.0 ;
      RECT  106350.0 1308600.0 107250.0 1309500.0 ;
      RECT  106350.0 1310550.0 107250.0 1311450.0 ;
      RECT  102900.0 1308600.0 106800.0 1309500.0 ;
      RECT  106350.0 1309050.0 107250.0 1311000.0 ;
      RECT  106800.0 1310550.0 110700.0 1311450.0 ;
      RECT  106350.0 1325700.0 107250.0 1326600.0 ;
      RECT  106350.0 1323750.0 107250.0 1324650.0 ;
      RECT  102900.0 1325700.0 106800.0 1326600.0 ;
      RECT  106350.0 1324200.0 107250.0 1326150.0 ;
      RECT  106800.0 1323750.0 110700.0 1324650.0 ;
      RECT  106350.0 1336200.0 107250.0 1337100.0 ;
      RECT  106350.0 1338150.0 107250.0 1339050.0 ;
      RECT  102900.0 1336200.0 106800.0 1337100.0 ;
      RECT  106350.0 1336650.0 107250.0 1338600.0 ;
      RECT  106800.0 1338150.0 110700.0 1339050.0 ;
      RECT  106350.0 1353300.0 107250.0 1354200.0 ;
      RECT  106350.0 1351350.0 107250.0 1352250.0 ;
      RECT  102900.0 1353300.0 106800.0 1354200.0 ;
      RECT  106350.0 1351800.0 107250.0 1353750.0 ;
      RECT  106800.0 1351350.0 110700.0 1352250.0 ;
      RECT  106350.0 1363800.0 107250.0 1364700.0 ;
      RECT  106350.0 1365750.0 107250.0 1366650.0 ;
      RECT  102900.0 1363800.0 106800.0 1364700.0 ;
      RECT  106350.0 1364250.0 107250.0 1366200.0 ;
      RECT  106800.0 1365750.0 110700.0 1366650.0 ;
      RECT  106350.0 1380900.0 107250.0 1381800.0 ;
      RECT  106350.0 1378950.0 107250.0 1379850.0 ;
      RECT  102900.0 1380900.0 106800.0 1381800.0 ;
      RECT  106350.0 1379400.0 107250.0 1381350.0 ;
      RECT  106800.0 1378950.0 110700.0 1379850.0 ;
      RECT  106350.0 1391400.0 107250.0 1392300.0 ;
      RECT  106350.0 1393350.0 107250.0 1394250.0 ;
      RECT  102900.0 1391400.0 106800.0 1392300.0 ;
      RECT  106350.0 1391850.0 107250.0 1393800.0 ;
      RECT  106800.0 1393350.0 110700.0 1394250.0 ;
      RECT  106350.0 1408500.0 107250.0 1409400.0 ;
      RECT  106350.0 1406550.0 107250.0 1407450.0 ;
      RECT  102900.0 1408500.0 106800.0 1409400.0 ;
      RECT  106350.0 1407000.0 107250.0 1408950.0 ;
      RECT  106800.0 1406550.0 110700.0 1407450.0 ;
      RECT  106350.0 1419000.0 107250.0 1419900.0 ;
      RECT  106350.0 1420950.0 107250.0 1421850.0 ;
      RECT  102900.0 1419000.0 106800.0 1419900.0 ;
      RECT  106350.0 1419450.0 107250.0 1421400.0 ;
      RECT  106800.0 1420950.0 110700.0 1421850.0 ;
      RECT  106350.0 1436100.0 107250.0 1437000.0 ;
      RECT  106350.0 1434150.0 107250.0 1435050.0 ;
      RECT  102900.0 1436100.0 106800.0 1437000.0 ;
      RECT  106350.0 1434600.0 107250.0 1436550.0 ;
      RECT  106800.0 1434150.0 110700.0 1435050.0 ;
      RECT  106350.0 1446600.0 107250.0 1447500.0 ;
      RECT  106350.0 1448550.0 107250.0 1449450.0 ;
      RECT  102900.0 1446600.0 106800.0 1447500.0 ;
      RECT  106350.0 1447050.0 107250.0 1449000.0 ;
      RECT  106800.0 1448550.0 110700.0 1449450.0 ;
      RECT  106350.0 1463700.0 107250.0 1464600.0 ;
      RECT  106350.0 1461750.0 107250.0 1462650.0 ;
      RECT  102900.0 1463700.0 106800.0 1464600.0 ;
      RECT  106350.0 1462200.0 107250.0 1464150.0 ;
      RECT  106800.0 1461750.0 110700.0 1462650.0 ;
      RECT  106350.0 1474200.0 107250.0 1475100.0 ;
      RECT  106350.0 1476150.0 107250.0 1477050.0 ;
      RECT  102900.0 1474200.0 106800.0 1475100.0 ;
      RECT  106350.0 1474650.0 107250.0 1476600.0 ;
      RECT  106800.0 1476150.0 110700.0 1477050.0 ;
      RECT  106350.0 1491300.0 107250.0 1492200.0 ;
      RECT  106350.0 1489350.0 107250.0 1490250.0 ;
      RECT  102900.0 1491300.0 106800.0 1492200.0 ;
      RECT  106350.0 1489800.0 107250.0 1491750.0 ;
      RECT  106800.0 1489350.0 110700.0 1490250.0 ;
      RECT  106350.0 1501800.0 107250.0 1502700.0 ;
      RECT  106350.0 1503750.0 107250.0 1504650.0 ;
      RECT  102900.0 1501800.0 106800.0 1502700.0 ;
      RECT  106350.0 1502250.0 107250.0 1504200.0 ;
      RECT  106800.0 1503750.0 110700.0 1504650.0 ;
      RECT  106350.0 1518900.0 107250.0 1519800.0 ;
      RECT  106350.0 1516950.0 107250.0 1517850.0 ;
      RECT  102900.0 1518900.0 106800.0 1519800.0 ;
      RECT  106350.0 1517400.0 107250.0 1519350.0 ;
      RECT  106800.0 1516950.0 110700.0 1517850.0 ;
      RECT  106350.0 1529400.0 107250.0 1530300.0 ;
      RECT  106350.0 1531350.0 107250.0 1532250.0 ;
      RECT  102900.0 1529400.0 106800.0 1530300.0 ;
      RECT  106350.0 1529850.0 107250.0 1531800.0 ;
      RECT  106800.0 1531350.0 110700.0 1532250.0 ;
      RECT  106350.0 1546500.0 107250.0 1547400.0 ;
      RECT  106350.0 1544550.0 107250.0 1545450.0 ;
      RECT  102900.0 1546500.0 106800.0 1547400.0 ;
      RECT  106350.0 1545000.0 107250.0 1546950.0 ;
      RECT  106800.0 1544550.0 110700.0 1545450.0 ;
      RECT  106350.0 1557000.0 107250.0 1557900.0 ;
      RECT  106350.0 1558950.0 107250.0 1559850.0 ;
      RECT  102900.0 1557000.0 106800.0 1557900.0 ;
      RECT  106350.0 1557450.0 107250.0 1559400.0 ;
      RECT  106800.0 1558950.0 110700.0 1559850.0 ;
      RECT  106350.0 1574100.0 107250.0 1575000.0 ;
      RECT  106350.0 1572150.0 107250.0 1573050.0 ;
      RECT  102900.0 1574100.0 106800.0 1575000.0 ;
      RECT  106350.0 1572600.0 107250.0 1574550.0 ;
      RECT  106800.0 1572150.0 110700.0 1573050.0 ;
      RECT  106350.0 1584600.0 107250.0 1585500.0 ;
      RECT  106350.0 1586550.0 107250.0 1587450.0 ;
      RECT  102900.0 1584600.0 106800.0 1585500.0 ;
      RECT  106350.0 1585050.0 107250.0 1587000.0 ;
      RECT  106800.0 1586550.0 110700.0 1587450.0 ;
      RECT  106350.0 1601700.0 107250.0 1602600.0 ;
      RECT  106350.0 1599750.0 107250.0 1600650.0 ;
      RECT  102900.0 1601700.0 106800.0 1602600.0 ;
      RECT  106350.0 1600200.0 107250.0 1602150.0 ;
      RECT  106800.0 1599750.0 110700.0 1600650.0 ;
      RECT  106350.0 1612200.0 107250.0 1613100.0 ;
      RECT  106350.0 1614150.0 107250.0 1615050.0 ;
      RECT  102900.0 1612200.0 106800.0 1613100.0 ;
      RECT  106350.0 1612650.0 107250.0 1614600.0 ;
      RECT  106800.0 1614150.0 110700.0 1615050.0 ;
      RECT  106350.0 1629300.0 107250.0 1630200.0 ;
      RECT  106350.0 1627350.0 107250.0 1628250.0 ;
      RECT  102900.0 1629300.0 106800.0 1630200.0 ;
      RECT  106350.0 1627800.0 107250.0 1629750.0 ;
      RECT  106800.0 1627350.0 110700.0 1628250.0 ;
      RECT  106350.0 1639800.0 107250.0 1640700.0 ;
      RECT  106350.0 1641750.0 107250.0 1642650.0 ;
      RECT  102900.0 1639800.0 106800.0 1640700.0 ;
      RECT  106350.0 1640250.0 107250.0 1642200.0 ;
      RECT  106800.0 1641750.0 110700.0 1642650.0 ;
      RECT  106350.0 1656900.0 107250.0 1657800.0 ;
      RECT  106350.0 1654950.0 107250.0 1655850.0 ;
      RECT  102900.0 1656900.0 106800.0 1657800.0 ;
      RECT  106350.0 1655400.0 107250.0 1657350.0 ;
      RECT  106800.0 1654950.0 110700.0 1655850.0 ;
      RECT  106350.0 1667400.0 107250.0 1668300.0 ;
      RECT  106350.0 1669350.0 107250.0 1670250.0 ;
      RECT  102900.0 1667400.0 106800.0 1668300.0 ;
      RECT  106350.0 1667850.0 107250.0 1669800.0 ;
      RECT  106800.0 1669350.0 110700.0 1670250.0 ;
      RECT  106350.0 1684500.0 107250.0 1685400.0 ;
      RECT  106350.0 1682550.0 107250.0 1683450.0 ;
      RECT  102900.0 1684500.0 106800.0 1685400.0 ;
      RECT  106350.0 1683000.0 107250.0 1684950.0 ;
      RECT  106800.0 1682550.0 110700.0 1683450.0 ;
      RECT  106350.0 1695000.0 107250.0 1695900.0 ;
      RECT  106350.0 1696950.0 107250.0 1697850.0 ;
      RECT  102900.0 1695000.0 106800.0 1695900.0 ;
      RECT  106350.0 1695450.0 107250.0 1697400.0 ;
      RECT  106800.0 1696950.0 110700.0 1697850.0 ;
      RECT  106350.0 1712100.0 107250.0 1713000.0 ;
      RECT  106350.0 1710150.0 107250.0 1711050.0 ;
      RECT  102900.0 1712100.0 106800.0 1713000.0 ;
      RECT  106350.0 1710600.0 107250.0 1712550.0 ;
      RECT  106800.0 1710150.0 110700.0 1711050.0 ;
      RECT  106350.0 1722600.0 107250.0 1723500.0 ;
      RECT  106350.0 1724550.0 107250.0 1725450.0 ;
      RECT  102900.0 1722600.0 106800.0 1723500.0 ;
      RECT  106350.0 1723050.0 107250.0 1725000.0 ;
      RECT  106800.0 1724550.0 110700.0 1725450.0 ;
      RECT  106350.0 1739700.0 107250.0 1740600.0 ;
      RECT  106350.0 1737750.0 107250.0 1738650.0 ;
      RECT  102900.0 1739700.0 106800.0 1740600.0 ;
      RECT  106350.0 1738200.0 107250.0 1740150.0 ;
      RECT  106800.0 1737750.0 110700.0 1738650.0 ;
      RECT  106350.0 1750200.0 107250.0 1751100.0 ;
      RECT  106350.0 1752150.0 107250.0 1753050.0 ;
      RECT  102900.0 1750200.0 106800.0 1751100.0 ;
      RECT  106350.0 1750650.0 107250.0 1752600.0 ;
      RECT  106800.0 1752150.0 110700.0 1753050.0 ;
      RECT  106350.0 1767300.0 107250.0 1768200.0 ;
      RECT  106350.0 1765350.0 107250.0 1766250.0 ;
      RECT  102900.0 1767300.0 106800.0 1768200.0 ;
      RECT  106350.0 1765800.0 107250.0 1767750.0 ;
      RECT  106800.0 1765350.0 110700.0 1766250.0 ;
      RECT  106350.0 1777800.0 107250.0 1778700.0 ;
      RECT  106350.0 1779750.0 107250.0 1780650.0 ;
      RECT  102900.0 1777800.0 106800.0 1778700.0 ;
      RECT  106350.0 1778250.0 107250.0 1780200.0 ;
      RECT  106800.0 1779750.0 110700.0 1780650.0 ;
      RECT  106350.0 1794900.0 107250.0 1795800.0 ;
      RECT  106350.0 1792950.0 107250.0 1793850.0 ;
      RECT  102900.0 1794900.0 106800.0 1795800.0 ;
      RECT  106350.0 1793400.0 107250.0 1795350.0 ;
      RECT  106800.0 1792950.0 110700.0 1793850.0 ;
      RECT  106350.0 1805400.0 107250.0 1806300.0 ;
      RECT  106350.0 1807350.0 107250.0 1808250.0 ;
      RECT  102900.0 1805400.0 106800.0 1806300.0 ;
      RECT  106350.0 1805850.0 107250.0 1807800.0 ;
      RECT  106800.0 1807350.0 110700.0 1808250.0 ;
      RECT  106350.0 1822500.0 107250.0 1823400.0 ;
      RECT  106350.0 1820550.0 107250.0 1821450.0 ;
      RECT  102900.0 1822500.0 106800.0 1823400.0 ;
      RECT  106350.0 1821000.0 107250.0 1822950.0 ;
      RECT  106800.0 1820550.0 110700.0 1821450.0 ;
      RECT  106350.0 1833000.0 107250.0 1833900.0 ;
      RECT  106350.0 1834950.0 107250.0 1835850.0 ;
      RECT  102900.0 1833000.0 106800.0 1833900.0 ;
      RECT  106350.0 1833450.0 107250.0 1835400.0 ;
      RECT  106800.0 1834950.0 110700.0 1835850.0 ;
      RECT  106350.0 1850100.0 107250.0 1851000.0 ;
      RECT  106350.0 1848150.0 107250.0 1849050.0 ;
      RECT  102900.0 1850100.0 106800.0 1851000.0 ;
      RECT  106350.0 1848600.0 107250.0 1850550.0 ;
      RECT  106800.0 1848150.0 110700.0 1849050.0 ;
      RECT  106350.0 1860600.0 107250.0 1861500.0 ;
      RECT  106350.0 1862550.0 107250.0 1863450.0 ;
      RECT  102900.0 1860600.0 106800.0 1861500.0 ;
      RECT  106350.0 1861050.0 107250.0 1863000.0 ;
      RECT  106800.0 1862550.0 110700.0 1863450.0 ;
      RECT  106350.0 1877700.0 107250.0 1878600.0 ;
      RECT  106350.0 1875750.0 107250.0 1876650.0 ;
      RECT  102900.0 1877700.0 106800.0 1878600.0 ;
      RECT  106350.0 1876200.0 107250.0 1878150.0 ;
      RECT  106800.0 1875750.0 110700.0 1876650.0 ;
      RECT  106350.0 1888200.0 107250.0 1889100.0 ;
      RECT  106350.0 1890150.0 107250.0 1891050.0 ;
      RECT  102900.0 1888200.0 106800.0 1889100.0 ;
      RECT  106350.0 1888650.0 107250.0 1890600.0 ;
      RECT  106800.0 1890150.0 110700.0 1891050.0 ;
      RECT  106350.0 1905300.0 107250.0 1906200.0 ;
      RECT  106350.0 1903350.0 107250.0 1904250.0 ;
      RECT  102900.0 1905300.0 106800.0 1906200.0 ;
      RECT  106350.0 1903800.0 107250.0 1905750.0 ;
      RECT  106800.0 1903350.0 110700.0 1904250.0 ;
      RECT  106350.0 1915800.0 107250.0 1916700.0 ;
      RECT  106350.0 1917750.0 107250.0 1918650.0 ;
      RECT  102900.0 1915800.0 106800.0 1916700.0 ;
      RECT  106350.0 1916250.0 107250.0 1918200.0 ;
      RECT  106800.0 1917750.0 110700.0 1918650.0 ;
      RECT  106350.0 1932900.0 107250.0 1933800.0 ;
      RECT  106350.0 1930950.0 107250.0 1931850.0 ;
      RECT  102900.0 1932900.0 106800.0 1933800.0 ;
      RECT  106350.0 1931400.0 107250.0 1933350.0 ;
      RECT  106800.0 1930950.0 110700.0 1931850.0 ;
      RECT  106350.0 1943400.0 107250.0 1944300.0 ;
      RECT  106350.0 1945350.0 107250.0 1946250.0 ;
      RECT  102900.0 1943400.0 106800.0 1944300.0 ;
      RECT  106350.0 1943850.0 107250.0 1945800.0 ;
      RECT  106800.0 1945350.0 110700.0 1946250.0 ;
      RECT  106350.0 1960500.0 107250.0 1961400.0 ;
      RECT  106350.0 1958550.0 107250.0 1959450.0 ;
      RECT  102900.0 1960500.0 106800.0 1961400.0 ;
      RECT  106350.0 1959000.0 107250.0 1960950.0 ;
      RECT  106800.0 1958550.0 110700.0 1959450.0 ;
      RECT  106350.0 1971000.0 107250.0 1971900.0 ;
      RECT  106350.0 1972950.0 107250.0 1973850.0 ;
      RECT  102900.0 1971000.0 106800.0 1971900.0 ;
      RECT  106350.0 1971450.0 107250.0 1973400.0 ;
      RECT  106800.0 1972950.0 110700.0 1973850.0 ;
      RECT  106350.0 1988100.0 107250.0 1989000.0 ;
      RECT  106350.0 1986150.0 107250.0 1987050.0 ;
      RECT  102900.0 1988100.0 106800.0 1989000.0 ;
      RECT  106350.0 1986600.0 107250.0 1988550.0 ;
      RECT  106800.0 1986150.0 110700.0 1987050.0 ;
      RECT  106350.0 1998600.0 107250.0 1999500.0 ;
      RECT  106350.0 2000550.0 107250.0 2001450.0 ;
      RECT  102900.0 1998600.0 106800.0 1999500.0 ;
      RECT  106350.0 1999050.0 107250.0 2001000.0 ;
      RECT  106800.0 2000550.0 110700.0 2001450.0 ;
      RECT  106350.0 2015700.0 107250.0 2016600.0 ;
      RECT  106350.0 2013750.0 107250.0 2014650.0 ;
      RECT  102900.0 2015700.0 106800.0 2016600.0 ;
      RECT  106350.0 2014200.0 107250.0 2016150.0 ;
      RECT  106800.0 2013750.0 110700.0 2014650.0 ;
      RECT  106350.0 2026200.0 107250.0 2027100.0 ;
      RECT  106350.0 2028150.0 107250.0 2029050.0 ;
      RECT  102900.0 2026200.0 106800.0 2027100.0 ;
      RECT  106350.0 2026650.0 107250.0 2028600.0 ;
      RECT  106800.0 2028150.0 110700.0 2029050.0 ;
      RECT  106350.0 2043300.0 107250.0 2044200.0 ;
      RECT  106350.0 2041350.0 107250.0 2042250.0 ;
      RECT  102900.0 2043300.0 106800.0 2044200.0 ;
      RECT  106350.0 2041800.0 107250.0 2043750.0 ;
      RECT  106800.0 2041350.0 110700.0 2042250.0 ;
      RECT  106350.0 2053800.0 107250.0 2054700.0 ;
      RECT  106350.0 2055750.0 107250.0 2056650.0 ;
      RECT  102900.0 2053800.0 106800.0 2054700.0 ;
      RECT  106350.0 2054250.0 107250.0 2056200.0 ;
      RECT  106800.0 2055750.0 110700.0 2056650.0 ;
      RECT  106350.0 2070900.0 107250.0 2071800.0 ;
      RECT  106350.0 2068950.0 107250.0 2069850.0 ;
      RECT  102900.0 2070900.0 106800.0 2071800.0 ;
      RECT  106350.0 2069400.0 107250.0 2071350.0 ;
      RECT  106800.0 2068950.0 110700.0 2069850.0 ;
      RECT  106350.0 2081400.0 107250.0 2082300.0 ;
      RECT  106350.0 2083350.0 107250.0 2084250.0 ;
      RECT  102900.0 2081400.0 106800.0 2082300.0 ;
      RECT  106350.0 2081850.0 107250.0 2083800.0 ;
      RECT  106800.0 2083350.0 110700.0 2084250.0 ;
      RECT  106350.0 2098500.0 107250.0 2099400.0 ;
      RECT  106350.0 2096550.0 107250.0 2097450.0 ;
      RECT  102900.0 2098500.0 106800.0 2099400.0 ;
      RECT  106350.0 2097000.0 107250.0 2098950.0 ;
      RECT  106800.0 2096550.0 110700.0 2097450.0 ;
      RECT  106350.0 2109000.0 107250.0 2109900.0 ;
      RECT  106350.0 2110950.0 107250.0 2111850.0 ;
      RECT  102900.0 2109000.0 106800.0 2109900.0 ;
      RECT  106350.0 2109450.0 107250.0 2111400.0 ;
      RECT  106800.0 2110950.0 110700.0 2111850.0 ;
      RECT  106350.0 2126100.0 107250.0 2127000.0 ;
      RECT  106350.0 2124150.0 107250.0 2125050.0 ;
      RECT  102900.0 2126100.0 106800.0 2127000.0 ;
      RECT  106350.0 2124600.0 107250.0 2126550.0 ;
      RECT  106800.0 2124150.0 110700.0 2125050.0 ;
      RECT  106350.0 2136600.0 107250.0 2137500.0 ;
      RECT  106350.0 2138550.0 107250.0 2139450.0 ;
      RECT  102900.0 2136600.0 106800.0 2137500.0 ;
      RECT  106350.0 2137050.0 107250.0 2139000.0 ;
      RECT  106800.0 2138550.0 110700.0 2139450.0 ;
      RECT  59550.0 164550.0 92700.0 165450.0 ;
      RECT  61650.0 178950.0 92700.0 179850.0 ;
      RECT  63750.0 192150.0 92700.0 193050.0 ;
      RECT  65850.0 206550.0 92700.0 207450.0 ;
      RECT  67950.0 219750.0 92700.0 220650.0 ;
      RECT  70050.0 234150.0 92700.0 235050.0 ;
      RECT  72150.0 247350.0 92700.0 248250.0 ;
      RECT  74250.0 261750.0 92700.0 262650.0 ;
      RECT  76350.0 274950.0 92700.0 275850.0 ;
      RECT  78450.0 289350.0 92700.0 290250.0 ;
      RECT  80550.0 302550.0 92700.0 303450.0 ;
      RECT  82650.0 316950.0 92700.0 317850.0 ;
      RECT  84750.0 330150.0 92700.0 331050.0 ;
      RECT  86850.0 344550.0 92700.0 345450.0 ;
      RECT  88950.0 357750.0 92700.0 358650.0 ;
      RECT  91050.0 372150.0 92700.0 373050.0 ;
      RECT  59550.0 387300.0 95700.0 388200.0 ;
      RECT  67950.0 385350.0 98100.0 386250.0 ;
      RECT  76350.0 383400.0 100500.0 384300.0 ;
      RECT  59550.0 397800.0 95700.0 398700.0 ;
      RECT  67950.0 399750.0 98100.0 400650.0 ;
      RECT  78450.0 401700.0 100500.0 402600.0 ;
      RECT  59550.0 414900.0 95700.0 415800.0 ;
      RECT  67950.0 412950.0 98100.0 413850.0 ;
      RECT  80550.0 411000.0 100500.0 411900.0 ;
      RECT  59550.0 425400.0 95700.0 426300.0 ;
      RECT  67950.0 427350.0 98100.0 428250.0 ;
      RECT  82650.0 429300.0 100500.0 430200.0 ;
      RECT  59550.0 442500.0 95700.0 443400.0 ;
      RECT  67950.0 440550.0 98100.0 441450.0 ;
      RECT  84750.0 438600.0 100500.0 439500.0 ;
      RECT  59550.0 453000.0 95700.0 453900.0 ;
      RECT  67950.0 454950.0 98100.0 455850.0 ;
      RECT  86850.0 456900.0 100500.0 457800.0 ;
      RECT  59550.0 470100.0 95700.0 471000.0 ;
      RECT  67950.0 468150.0 98100.0 469050.0 ;
      RECT  88950.0 466200.0 100500.0 467100.0 ;
      RECT  59550.0 480600.0 95700.0 481500.0 ;
      RECT  67950.0 482550.0 98100.0 483450.0 ;
      RECT  91050.0 484500.0 100500.0 485400.0 ;
      RECT  59550.0 497700.0 95700.0 498600.0 ;
      RECT  70050.0 495750.0 98100.0 496650.0 ;
      RECT  76350.0 493800.0 100500.0 494700.0 ;
      RECT  59550.0 508200.0 95700.0 509100.0 ;
      RECT  70050.0 510150.0 98100.0 511050.0 ;
      RECT  78450.0 512100.0 100500.0 513000.0 ;
      RECT  59550.0 525300.0 95700.0 526200.0 ;
      RECT  70050.0 523350.0 98100.0 524250.0 ;
      RECT  80550.0 521400.0 100500.0 522300.0 ;
      RECT  59550.0 535800.0 95700.0 536700.0 ;
      RECT  70050.0 537750.0 98100.0 538650.0 ;
      RECT  82650.0 539700.0 100500.0 540600.0 ;
      RECT  59550.0 552900.0 95700.0 553800.0 ;
      RECT  70050.0 550950.0 98100.0 551850.0 ;
      RECT  84750.0 549000.0 100500.0 549900.0 ;
      RECT  59550.0 563400.0 95700.0 564300.0 ;
      RECT  70050.0 565350.0 98100.0 566250.0 ;
      RECT  86850.0 567300.0 100500.0 568200.0 ;
      RECT  59550.0 580500.0 95700.0 581400.0 ;
      RECT  70050.0 578550.0 98100.0 579450.0 ;
      RECT  88950.0 576600.0 100500.0 577500.0 ;
      RECT  59550.0 591000.0 95700.0 591900.0 ;
      RECT  70050.0 592950.0 98100.0 593850.0 ;
      RECT  91050.0 594900.0 100500.0 595800.0 ;
      RECT  59550.0 608100.0 95700.0 609000.0 ;
      RECT  72150.0 606150.0 98100.0 607050.0 ;
      RECT  76350.0 604200.0 100500.0 605100.0 ;
      RECT  59550.0 618600.0 95700.0 619500.0 ;
      RECT  72150.0 620550.0 98100.0 621450.0 ;
      RECT  78450.0 622500.0 100500.0 623400.0 ;
      RECT  59550.0 635700.0 95700.0 636600.0 ;
      RECT  72150.0 633750.0 98100.0 634650.0 ;
      RECT  80550.0 631800.0 100500.0 632700.0 ;
      RECT  59550.0 646200.0 95700.0 647100.0 ;
      RECT  72150.0 648150.0 98100.0 649050.0 ;
      RECT  82650.0 650100.0 100500.0 651000.0 ;
      RECT  59550.0 663300.0 95700.0 664200.0 ;
      RECT  72150.0 661350.0 98100.0 662250.0 ;
      RECT  84750.0 659400.0 100500.0 660300.0 ;
      RECT  59550.0 673800.0 95700.0 674700.0 ;
      RECT  72150.0 675750.0 98100.0 676650.0 ;
      RECT  86850.0 677700.0 100500.0 678600.0 ;
      RECT  59550.0 690900.0 95700.0 691800.0 ;
      RECT  72150.0 688950.0 98100.0 689850.0 ;
      RECT  88950.0 687000.0 100500.0 687900.0 ;
      RECT  59550.0 701400.0 95700.0 702300.0 ;
      RECT  72150.0 703350.0 98100.0 704250.0 ;
      RECT  91050.0 705300.0 100500.0 706200.0 ;
      RECT  59550.0 718500.0 95700.0 719400.0 ;
      RECT  74250.0 716550.0 98100.0 717450.0 ;
      RECT  76350.0 714600.0 100500.0 715500.0 ;
      RECT  59550.0 729000.0 95700.0 729900.0 ;
      RECT  74250.0 730950.0 98100.0 731850.0 ;
      RECT  78450.0 732900.0 100500.0 733800.0 ;
      RECT  59550.0 746100.0 95700.0 747000.0 ;
      RECT  74250.0 744150.0 98100.0 745050.0 ;
      RECT  80550.0 742200.0 100500.0 743100.0 ;
      RECT  59550.0 756600.0 95700.0 757500.0 ;
      RECT  74250.0 758550.0 98100.0 759450.0 ;
      RECT  82650.0 760500.0 100500.0 761400.0 ;
      RECT  59550.0 773700.0 95700.0 774600.0 ;
      RECT  74250.0 771750.0 98100.0 772650.0 ;
      RECT  84750.0 769800.0 100500.0 770700.0 ;
      RECT  59550.0 784200.0 95700.0 785100.0 ;
      RECT  74250.0 786150.0 98100.0 787050.0 ;
      RECT  86850.0 788100.0 100500.0 789000.0 ;
      RECT  59550.0 801300.0 95700.0 802200.0 ;
      RECT  74250.0 799350.0 98100.0 800250.0 ;
      RECT  88950.0 797400.0 100500.0 798300.0 ;
      RECT  59550.0 811800.0 95700.0 812700.0 ;
      RECT  74250.0 813750.0 98100.0 814650.0 ;
      RECT  91050.0 815700.0 100500.0 816600.0 ;
      RECT  61650.0 828900.0 95700.0 829800.0 ;
      RECT  67950.0 826950.0 98100.0 827850.0 ;
      RECT  76350.0 825000.0 100500.0 825900.0 ;
      RECT  61650.0 839400.0 95700.0 840300.0 ;
      RECT  67950.0 841350.0 98100.0 842250.0 ;
      RECT  78450.0 843300.0 100500.0 844200.0 ;
      RECT  61650.0 856500.0 95700.0 857400.0 ;
      RECT  67950.0 854550.0 98100.0 855450.0 ;
      RECT  80550.0 852600.0 100500.0 853500.0 ;
      RECT  61650.0 867000.0 95700.0 867900.0 ;
      RECT  67950.0 868950.0 98100.0 869850.0 ;
      RECT  82650.0 870900.0 100500.0 871800.0 ;
      RECT  61650.0 884100.0 95700.0 885000.0 ;
      RECT  67950.0 882150.0 98100.0 883050.0 ;
      RECT  84750.0 880200.0 100500.0 881100.0 ;
      RECT  61650.0 894600.0 95700.0 895500.0 ;
      RECT  67950.0 896550.0 98100.0 897450.0 ;
      RECT  86850.0 898500.0 100500.0 899400.0 ;
      RECT  61650.0 911700.0 95700.0 912600.0 ;
      RECT  67950.0 909750.0 98100.0 910650.0 ;
      RECT  88950.0 907800.0 100500.0 908700.0 ;
      RECT  61650.0 922200.0 95700.0 923100.0 ;
      RECT  67950.0 924150.0 98100.0 925050.0 ;
      RECT  91050.0 926100.0 100500.0 927000.0 ;
      RECT  61650.0 939300.0 95700.0 940200.0 ;
      RECT  70050.0 937350.0 98100.0 938250.0 ;
      RECT  76350.0 935400.0 100500.0 936300.0 ;
      RECT  61650.0 949800.0 95700.0 950700.0 ;
      RECT  70050.0 951750.0 98100.0 952650.0 ;
      RECT  78450.0 953700.0 100500.0 954600.0 ;
      RECT  61650.0 966900.0 95700.0 967800.0 ;
      RECT  70050.0 964950.0 98100.0 965850.0 ;
      RECT  80550.0 963000.0 100500.0 963900.0 ;
      RECT  61650.0 977400.0 95700.0 978300.0 ;
      RECT  70050.0 979350.0 98100.0 980250.0 ;
      RECT  82650.0 981300.0 100500.0 982200.0 ;
      RECT  61650.0 994500.0 95700.0 995400.0 ;
      RECT  70050.0 992550.0 98100.0 993450.0 ;
      RECT  84750.0 990600.0 100500.0 991500.0 ;
      RECT  61650.0 1005000.0 95700.0 1005900.0 ;
      RECT  70050.0 1006950.0 98100.0 1007850.0 ;
      RECT  86850.0 1008900.0 100500.0 1009800.0 ;
      RECT  61650.0 1022100.0 95700.0 1023000.0 ;
      RECT  70050.0 1020150.0 98100.0 1021050.0 ;
      RECT  88950.0 1018200.0 100500.0 1019100.0 ;
      RECT  61650.0 1032600.0 95700.0 1033500.0 ;
      RECT  70050.0 1034550.0 98100.0 1035450.0 ;
      RECT  91050.0 1036500.0 100500.0 1037400.0 ;
      RECT  61650.0 1049700.0 95700.0 1050600.0 ;
      RECT  72150.0 1047750.0 98100.0 1048650.0 ;
      RECT  76350.0 1045800.0 100500.0 1046700.0 ;
      RECT  61650.0 1060200.0 95700.0 1061100.0 ;
      RECT  72150.0 1062150.0 98100.0 1063050.0 ;
      RECT  78450.0 1064100.0 100500.0 1065000.0 ;
      RECT  61650.0 1077300.0 95700.0 1078200.0 ;
      RECT  72150.0 1075350.0 98100.0 1076250.0 ;
      RECT  80550.0 1073400.0 100500.0 1074300.0 ;
      RECT  61650.0 1087800.0 95700.0 1088700.0 ;
      RECT  72150.0 1089750.0 98100.0 1090650.0 ;
      RECT  82650.0 1091700.0 100500.0 1092600.0 ;
      RECT  61650.0 1104900.0 95700.0 1105800.0 ;
      RECT  72150.0 1102950.0 98100.0 1103850.0 ;
      RECT  84750.0 1101000.0 100500.0 1101900.0 ;
      RECT  61650.0 1115400.0 95700.0 1116300.0 ;
      RECT  72150.0 1117350.0 98100.0 1118250.0 ;
      RECT  86850.0 1119300.0 100500.0 1120200.0 ;
      RECT  61650.0 1132500.0 95700.0 1133400.0 ;
      RECT  72150.0 1130550.0 98100.0 1131450.0 ;
      RECT  88950.0 1128600.0 100500.0 1129500.0 ;
      RECT  61650.0 1143000.0 95700.0 1143900.0 ;
      RECT  72150.0 1144950.0 98100.0 1145850.0 ;
      RECT  91050.0 1146900.0 100500.0 1147800.0 ;
      RECT  61650.0 1160100.0 95700.0 1161000.0 ;
      RECT  74250.0 1158150.0 98100.0 1159050.0 ;
      RECT  76350.0 1156200.0 100500.0 1157100.0 ;
      RECT  61650.0 1170600.0 95700.0 1171500.0 ;
      RECT  74250.0 1172550.0 98100.0 1173450.0 ;
      RECT  78450.0 1174500.0 100500.0 1175400.0 ;
      RECT  61650.0 1187700.0 95700.0 1188600.0 ;
      RECT  74250.0 1185750.0 98100.0 1186650.0 ;
      RECT  80550.0 1183800.0 100500.0 1184700.0 ;
      RECT  61650.0 1198200.0 95700.0 1199100.0 ;
      RECT  74250.0 1200150.0 98100.0 1201050.0 ;
      RECT  82650.0 1202100.0 100500.0 1203000.0 ;
      RECT  61650.0 1215300.0 95700.0 1216200.0 ;
      RECT  74250.0 1213350.0 98100.0 1214250.0 ;
      RECT  84750.0 1211400.0 100500.0 1212300.0 ;
      RECT  61650.0 1225800.0 95700.0 1226700.0 ;
      RECT  74250.0 1227750.0 98100.0 1228650.0 ;
      RECT  86850.0 1229700.0 100500.0 1230600.0 ;
      RECT  61650.0 1242900.0 95700.0 1243800.0 ;
      RECT  74250.0 1240950.0 98100.0 1241850.0 ;
      RECT  88950.0 1239000.0 100500.0 1239900.0 ;
      RECT  61650.0 1253400.0 95700.0 1254300.0 ;
      RECT  74250.0 1255350.0 98100.0 1256250.0 ;
      RECT  91050.0 1257300.0 100500.0 1258200.0 ;
      RECT  63750.0 1270500.0 95700.0 1271400.0 ;
      RECT  67950.0 1268550.0 98100.0 1269450.0 ;
      RECT  76350.0 1266600.0 100500.0 1267500.0 ;
      RECT  63750.0 1281000.0 95700.0 1281900.0 ;
      RECT  67950.0 1282950.0 98100.0 1283850.0 ;
      RECT  78450.0 1284900.0 100500.0 1285800.0 ;
      RECT  63750.0 1298100.0 95700.0 1299000.0 ;
      RECT  67950.0 1296150.0 98100.0 1297050.0 ;
      RECT  80550.0 1294200.0 100500.0 1295100.0 ;
      RECT  63750.0 1308600.0 95700.0 1309500.0 ;
      RECT  67950.0 1310550.0 98100.0 1311450.0 ;
      RECT  82650.0 1312500.0 100500.0 1313400.0 ;
      RECT  63750.0 1325700.0 95700.0 1326600.0 ;
      RECT  67950.0 1323750.0 98100.0 1324650.0 ;
      RECT  84750.0 1321800.0 100500.0 1322700.0 ;
      RECT  63750.0 1336200.0 95700.0 1337100.0 ;
      RECT  67950.0 1338150.0 98100.0 1339050.0 ;
      RECT  86850.0 1340100.0 100500.0 1341000.0 ;
      RECT  63750.0 1353300.0 95700.0 1354200.0 ;
      RECT  67950.0 1351350.0 98100.0 1352250.0 ;
      RECT  88950.0 1349400.0 100500.0 1350300.0 ;
      RECT  63750.0 1363800.0 95700.0 1364700.0 ;
      RECT  67950.0 1365750.0 98100.0 1366650.0 ;
      RECT  91050.0 1367700.0 100500.0 1368600.0 ;
      RECT  63750.0 1380900.0 95700.0 1381800.0 ;
      RECT  70050.0 1378950.0 98100.0 1379850.0 ;
      RECT  76350.0 1377000.0 100500.0 1377900.0 ;
      RECT  63750.0 1391400.0 95700.0 1392300.0 ;
      RECT  70050.0 1393350.0 98100.0 1394250.0 ;
      RECT  78450.0 1395300.0 100500.0 1396200.0 ;
      RECT  63750.0 1408500.0 95700.0 1409400.0 ;
      RECT  70050.0 1406550.0 98100.0 1407450.0 ;
      RECT  80550.0 1404600.0 100500.0 1405500.0 ;
      RECT  63750.0 1419000.0 95700.0 1419900.0 ;
      RECT  70050.0 1420950.0 98100.0 1421850.0 ;
      RECT  82650.0 1422900.0 100500.0 1423800.0 ;
      RECT  63750.0 1436100.0 95700.0 1437000.0 ;
      RECT  70050.0 1434150.0 98100.0 1435050.0 ;
      RECT  84750.0 1432200.0 100500.0 1433100.0 ;
      RECT  63750.0 1446600.0 95700.0 1447500.0 ;
      RECT  70050.0 1448550.0 98100.0 1449450.0 ;
      RECT  86850.0 1450500.0 100500.0 1451400.0 ;
      RECT  63750.0 1463700.0 95700.0 1464600.0 ;
      RECT  70050.0 1461750.0 98100.0 1462650.0 ;
      RECT  88950.0 1459800.0 100500.0 1460700.0 ;
      RECT  63750.0 1474200.0 95700.0 1475100.0 ;
      RECT  70050.0 1476150.0 98100.0 1477050.0 ;
      RECT  91050.0 1478100.0 100500.0 1479000.0 ;
      RECT  63750.0 1491300.0 95700.0 1492200.0 ;
      RECT  72150.0 1489350.0 98100.0 1490250.0 ;
      RECT  76350.0 1487400.0 100500.0 1488300.0 ;
      RECT  63750.0 1501800.0 95700.0 1502700.0 ;
      RECT  72150.0 1503750.0 98100.0 1504650.0 ;
      RECT  78450.0 1505700.0 100500.0 1506600.0 ;
      RECT  63750.0 1518900.0 95700.0 1519800.0 ;
      RECT  72150.0 1516950.0 98100.0 1517850.0 ;
      RECT  80550.0 1515000.0 100500.0 1515900.0 ;
      RECT  63750.0 1529400.0 95700.0 1530300.0 ;
      RECT  72150.0 1531350.0 98100.0 1532250.0 ;
      RECT  82650.0 1533300.0 100500.0 1534200.0 ;
      RECT  63750.0 1546500.0 95700.0 1547400.0 ;
      RECT  72150.0 1544550.0 98100.0 1545450.0 ;
      RECT  84750.0 1542600.0 100500.0 1543500.0 ;
      RECT  63750.0 1557000.0 95700.0 1557900.0 ;
      RECT  72150.0 1558950.0 98100.0 1559850.0 ;
      RECT  86850.0 1560900.0 100500.0 1561800.0 ;
      RECT  63750.0 1574100.0 95700.0 1575000.0 ;
      RECT  72150.0 1572150.0 98100.0 1573050.0 ;
      RECT  88950.0 1570200.0 100500.0 1571100.0 ;
      RECT  63750.0 1584600.0 95700.0 1585500.0 ;
      RECT  72150.0 1586550.0 98100.0 1587450.0 ;
      RECT  91050.0 1588500.0 100500.0 1589400.0 ;
      RECT  63750.0 1601700.0 95700.0 1602600.0 ;
      RECT  74250.0 1599750.0 98100.0 1600650.0 ;
      RECT  76350.0 1597800.0 100500.0 1598700.0 ;
      RECT  63750.0 1612200.0 95700.0 1613100.0 ;
      RECT  74250.0 1614150.0 98100.0 1615050.0 ;
      RECT  78450.0 1616100.0 100500.0 1617000.0 ;
      RECT  63750.0 1629300.0 95700.0 1630200.0 ;
      RECT  74250.0 1627350.0 98100.0 1628250.0 ;
      RECT  80550.0 1625400.0 100500.0 1626300.0 ;
      RECT  63750.0 1639800.0 95700.0 1640700.0 ;
      RECT  74250.0 1641750.0 98100.0 1642650.0 ;
      RECT  82650.0 1643700.0 100500.0 1644600.0 ;
      RECT  63750.0 1656900.0 95700.0 1657800.0 ;
      RECT  74250.0 1654950.0 98100.0 1655850.0 ;
      RECT  84750.0 1653000.0 100500.0 1653900.0 ;
      RECT  63750.0 1667400.0 95700.0 1668300.0 ;
      RECT  74250.0 1669350.0 98100.0 1670250.0 ;
      RECT  86850.0 1671300.0 100500.0 1672200.0 ;
      RECT  63750.0 1684500.0 95700.0 1685400.0 ;
      RECT  74250.0 1682550.0 98100.0 1683450.0 ;
      RECT  88950.0 1680600.0 100500.0 1681500.0 ;
      RECT  63750.0 1695000.0 95700.0 1695900.0 ;
      RECT  74250.0 1696950.0 98100.0 1697850.0 ;
      RECT  91050.0 1698900.0 100500.0 1699800.0 ;
      RECT  65850.0 1712100.0 95700.0 1713000.0 ;
      RECT  67950.0 1710150.0 98100.0 1711050.0 ;
      RECT  76350.0 1708200.0 100500.0 1709100.0 ;
      RECT  65850.0 1722600.0 95700.0 1723500.0 ;
      RECT  67950.0 1724550.0 98100.0 1725450.0 ;
      RECT  78450.0 1726500.0 100500.0 1727400.0 ;
      RECT  65850.0 1739700.0 95700.0 1740600.0 ;
      RECT  67950.0 1737750.0 98100.0 1738650.0 ;
      RECT  80550.0 1735800.0 100500.0 1736700.0 ;
      RECT  65850.0 1750200.0 95700.0 1751100.0 ;
      RECT  67950.0 1752150.0 98100.0 1753050.0 ;
      RECT  82650.0 1754100.0 100500.0 1755000.0 ;
      RECT  65850.0 1767300.0 95700.0 1768200.0 ;
      RECT  67950.0 1765350.0 98100.0 1766250.0 ;
      RECT  84750.0 1763400.0 100500.0 1764300.0 ;
      RECT  65850.0 1777800.0 95700.0 1778700.0 ;
      RECT  67950.0 1779750.0 98100.0 1780650.0 ;
      RECT  86850.0 1781700.0 100500.0 1782600.0 ;
      RECT  65850.0 1794900.0 95700.0 1795800.0 ;
      RECT  67950.0 1792950.0 98100.0 1793850.0 ;
      RECT  88950.0 1791000.0 100500.0 1791900.0 ;
      RECT  65850.0 1805400.0 95700.0 1806300.0 ;
      RECT  67950.0 1807350.0 98100.0 1808250.0 ;
      RECT  91050.0 1809300.0 100500.0 1810200.0 ;
      RECT  65850.0 1822500.0 95700.0 1823400.0 ;
      RECT  70050.0 1820550.0 98100.0 1821450.0 ;
      RECT  76350.0 1818600.0 100500.0 1819500.0 ;
      RECT  65850.0 1833000.0 95700.0 1833900.0 ;
      RECT  70050.0 1834950.0 98100.0 1835850.0 ;
      RECT  78450.0 1836900.0 100500.0 1837800.0 ;
      RECT  65850.0 1850100.0 95700.0 1851000.0 ;
      RECT  70050.0 1848150.0 98100.0 1849050.0 ;
      RECT  80550.0 1846200.0 100500.0 1847100.0 ;
      RECT  65850.0 1860600.0 95700.0 1861500.0 ;
      RECT  70050.0 1862550.0 98100.0 1863450.0 ;
      RECT  82650.0 1864500.0 100500.0 1865400.0 ;
      RECT  65850.0 1877700.0 95700.0 1878600.0 ;
      RECT  70050.0 1875750.0 98100.0 1876650.0 ;
      RECT  84750.0 1873800.0 100500.0 1874700.0 ;
      RECT  65850.0 1888200.0 95700.0 1889100.0 ;
      RECT  70050.0 1890150.0 98100.0 1891050.0 ;
      RECT  86850.0 1892100.0 100500.0 1893000.0 ;
      RECT  65850.0 1905300.0 95700.0 1906200.0 ;
      RECT  70050.0 1903350.0 98100.0 1904250.0 ;
      RECT  88950.0 1901400.0 100500.0 1902300.0 ;
      RECT  65850.0 1915800.0 95700.0 1916700.0 ;
      RECT  70050.0 1917750.0 98100.0 1918650.0 ;
      RECT  91050.0 1919700.0 100500.0 1920600.0 ;
      RECT  65850.0 1932900.0 95700.0 1933800.0 ;
      RECT  72150.0 1930950.0 98100.0 1931850.0 ;
      RECT  76350.0 1929000.0 100500.0 1929900.0 ;
      RECT  65850.0 1943400.0 95700.0 1944300.0 ;
      RECT  72150.0 1945350.0 98100.0 1946250.0 ;
      RECT  78450.0 1947300.0 100500.0 1948200.0 ;
      RECT  65850.0 1960500.0 95700.0 1961400.0 ;
      RECT  72150.0 1958550.0 98100.0 1959450.0 ;
      RECT  80550.0 1956600.0 100500.0 1957500.0 ;
      RECT  65850.0 1971000.0 95700.0 1971900.0 ;
      RECT  72150.0 1972950.0 98100.0 1973850.0 ;
      RECT  82650.0 1974900.0 100500.0 1975800.0 ;
      RECT  65850.0 1988100.0 95700.0 1989000.0 ;
      RECT  72150.0 1986150.0 98100.0 1987050.0 ;
      RECT  84750.0 1984200.0 100500.0 1985100.0 ;
      RECT  65850.0 1998600.0 95700.0 1999500.0 ;
      RECT  72150.0 2000550.0 98100.0 2001450.0 ;
      RECT  86850.0 2002500.0 100500.0 2003400.0 ;
      RECT  65850.0 2015700.0 95700.0 2016600.0 ;
      RECT  72150.0 2013750.0 98100.0 2014650.0 ;
      RECT  88950.0 2011800.0 100500.0 2012700.0 ;
      RECT  65850.0 2026200.0 95700.0 2027100.0 ;
      RECT  72150.0 2028150.0 98100.0 2029050.0 ;
      RECT  91050.0 2030100.0 100500.0 2031000.0 ;
      RECT  65850.0 2043300.0 95700.0 2044200.0 ;
      RECT  74250.0 2041350.0 98100.0 2042250.0 ;
      RECT  76350.0 2039400.0 100500.0 2040300.0 ;
      RECT  65850.0 2053800.0 95700.0 2054700.0 ;
      RECT  74250.0 2055750.0 98100.0 2056650.0 ;
      RECT  78450.0 2057700.0 100500.0 2058600.0 ;
      RECT  65850.0 2070900.0 95700.0 2071800.0 ;
      RECT  74250.0 2068950.0 98100.0 2069850.0 ;
      RECT  80550.0 2067000.0 100500.0 2067900.0 ;
      RECT  65850.0 2081400.0 95700.0 2082300.0 ;
      RECT  74250.0 2083350.0 98100.0 2084250.0 ;
      RECT  82650.0 2085300.0 100500.0 2086200.0 ;
      RECT  65850.0 2098500.0 95700.0 2099400.0 ;
      RECT  74250.0 2096550.0 98100.0 2097450.0 ;
      RECT  84750.0 2094600.0 100500.0 2095500.0 ;
      RECT  65850.0 2109000.0 95700.0 2109900.0 ;
      RECT  74250.0 2110950.0 98100.0 2111850.0 ;
      RECT  86850.0 2112900.0 100500.0 2113800.0 ;
      RECT  65850.0 2126100.0 95700.0 2127000.0 ;
      RECT  74250.0 2124150.0 98100.0 2125050.0 ;
      RECT  88950.0 2122200.0 100500.0 2123100.0 ;
      RECT  65850.0 2136600.0 95700.0 2137500.0 ;
      RECT  74250.0 2138550.0 98100.0 2139450.0 ;
      RECT  91050.0 2140500.0 100500.0 2141400.0 ;
      RECT  131250.0 164550.0 130350.0 165450.0 ;
      RECT  131250.0 169050.0 130350.0 169950.0 ;
      RECT  135450.0 164550.0 130800.0 165450.0 ;
      RECT  131250.0 165000.0 130350.0 169500.0 ;
      RECT  130800.0 169050.0 128250.0 169950.0 ;
      RECT  146850.0 164550.0 138900.0 165450.0 ;
      RECT  131250.0 178950.0 130350.0 179850.0 ;
      RECT  131250.0 182850.0 130350.0 183750.0 ;
      RECT  135450.0 178950.0 130800.0 179850.0 ;
      RECT  131250.0 179400.0 130350.0 183300.0 ;
      RECT  130800.0 182850.0 125250.0 183750.0 ;
      RECT  143850.0 178950.0 138900.0 179850.0 ;
      RECT  146850.0 187650.0 122250.0 188550.0 ;
      RECT  143850.0 201450.0 119250.0 202350.0 ;
      RECT  128250.0 165750.0 114300.0 166650.0 ;
      RECT  125250.0 163050.0 111300.0 163950.0 ;
      RECT  122250.0 177750.0 114300.0 178650.0 ;
      RECT  125250.0 180450.0 111300.0 181350.0 ;
      RECT  128250.0 193350.0 114300.0 194250.0 ;
      RECT  119250.0 190650.0 111300.0 191550.0 ;
      RECT  122250.0 205350.0 114300.0 206250.0 ;
      RECT  119250.0 208050.0 111300.0 208950.0 ;
      RECT  104850.0 165750.0 103950.0 166650.0 ;
      RECT  104850.0 164550.0 103950.0 165450.0 ;
      RECT  108900.0 165750.0 104400.0 166650.0 ;
      RECT  104850.0 165000.0 103950.0 166200.0 ;
      RECT  104400.0 164550.0 99900.0 165450.0 ;
      RECT  104850.0 177750.0 103950.0 178650.0 ;
      RECT  104850.0 178950.0 103950.0 179850.0 ;
      RECT  108900.0 177750.0 104400.0 178650.0 ;
      RECT  104850.0 178200.0 103950.0 179400.0 ;
      RECT  104400.0 178950.0 99900.0 179850.0 ;
      RECT  104850.0 193350.0 103950.0 194250.0 ;
      RECT  104850.0 192150.0 103950.0 193050.0 ;
      RECT  108900.0 193350.0 104400.0 194250.0 ;
      RECT  104850.0 192600.0 103950.0 193800.0 ;
      RECT  104400.0 192150.0 99900.0 193050.0 ;
      RECT  104850.0 205350.0 103950.0 206250.0 ;
      RECT  104850.0 206550.0 103950.0 207450.0 ;
      RECT  108900.0 205350.0 104400.0 206250.0 ;
      RECT  104850.0 205800.0 103950.0 207000.0 ;
      RECT  104400.0 206550.0 99900.0 207450.0 ;
      RECT  134700.0 170250.0 133500.0 172200.0 ;
      RECT  134700.0 158400.0 133500.0 160350.0 ;
      RECT  139500.0 159750.0 138300.0 157950.0 ;
      RECT  139500.0 169050.0 138300.0 172650.0 ;
      RECT  136800.0 159750.0 135900.0 169050.0 ;
      RECT  139500.0 169050.0 138300.0 170250.0 ;
      RECT  137100.0 169050.0 135900.0 170250.0 ;
      RECT  137100.0 169050.0 135900.0 170250.0 ;
      RECT  139500.0 169050.0 138300.0 170250.0 ;
      RECT  139500.0 159750.0 138300.0 160950.0 ;
      RECT  137100.0 159750.0 135900.0 160950.0 ;
      RECT  137100.0 159750.0 135900.0 160950.0 ;
      RECT  139500.0 159750.0 138300.0 160950.0 ;
      RECT  134700.0 169650.0 133500.0 170850.0 ;
      RECT  134700.0 159750.0 133500.0 160950.0 ;
      RECT  138900.0 164400.0 137700.0 165600.0 ;
      RECT  138900.0 164400.0 137700.0 165600.0 ;
      RECT  136350.0 164550.0 135450.0 165450.0 ;
      RECT  141300.0 171750.0 131700.0 172650.0 ;
      RECT  141300.0 157950.0 131700.0 158850.0 ;
      RECT  134700.0 174150.0 133500.0 172200.0 ;
      RECT  134700.0 186000.0 133500.0 184050.0 ;
      RECT  139500.0 184650.0 138300.0 186450.0 ;
      RECT  139500.0 175350.0 138300.0 171750.0 ;
      RECT  136800.0 184650.0 135900.0 175350.0 ;
      RECT  139500.0 175350.0 138300.0 174150.0 ;
      RECT  137100.0 175350.0 135900.0 174150.0 ;
      RECT  137100.0 175350.0 135900.0 174150.0 ;
      RECT  139500.0 175350.0 138300.0 174150.0 ;
      RECT  139500.0 184650.0 138300.0 183450.0 ;
      RECT  137100.0 184650.0 135900.0 183450.0 ;
      RECT  137100.0 184650.0 135900.0 183450.0 ;
      RECT  139500.0 184650.0 138300.0 183450.0 ;
      RECT  134700.0 174750.0 133500.0 173550.0 ;
      RECT  134700.0 184650.0 133500.0 183450.0 ;
      RECT  138900.0 180000.0 137700.0 178800.0 ;
      RECT  138900.0 180000.0 137700.0 178800.0 ;
      RECT  136350.0 179850.0 135450.0 178950.0 ;
      RECT  141300.0 172650.0 131700.0 171750.0 ;
      RECT  141300.0 186450.0 131700.0 185550.0 ;
      RECT  95700.0 170250.0 94500.0 172200.0 ;
      RECT  95700.0 158400.0 94500.0 160350.0 ;
      RECT  100500.0 159750.0 99300.0 157950.0 ;
      RECT  100500.0 169050.0 99300.0 172650.0 ;
      RECT  97800.0 159750.0 96900.0 169050.0 ;
      RECT  100500.0 169050.0 99300.0 170250.0 ;
      RECT  98100.0 169050.0 96900.0 170250.0 ;
      RECT  98100.0 169050.0 96900.0 170250.0 ;
      RECT  100500.0 169050.0 99300.0 170250.0 ;
      RECT  100500.0 159750.0 99300.0 160950.0 ;
      RECT  98100.0 159750.0 96900.0 160950.0 ;
      RECT  98100.0 159750.0 96900.0 160950.0 ;
      RECT  100500.0 159750.0 99300.0 160950.0 ;
      RECT  95700.0 169650.0 94500.0 170850.0 ;
      RECT  95700.0 159750.0 94500.0 160950.0 ;
      RECT  99900.0 164400.0 98700.0 165600.0 ;
      RECT  99900.0 164400.0 98700.0 165600.0 ;
      RECT  97350.0 164550.0 96450.0 165450.0 ;
      RECT  102300.0 171750.0 92700.0 172650.0 ;
      RECT  102300.0 157950.0 92700.0 158850.0 ;
      RECT  95700.0 174150.0 94500.0 172200.0 ;
      RECT  95700.0 186000.0 94500.0 184050.0 ;
      RECT  100500.0 184650.0 99300.0 186450.0 ;
      RECT  100500.0 175350.0 99300.0 171750.0 ;
      RECT  97800.0 184650.0 96900.0 175350.0 ;
      RECT  100500.0 175350.0 99300.0 174150.0 ;
      RECT  98100.0 175350.0 96900.0 174150.0 ;
      RECT  98100.0 175350.0 96900.0 174150.0 ;
      RECT  100500.0 175350.0 99300.0 174150.0 ;
      RECT  100500.0 184650.0 99300.0 183450.0 ;
      RECT  98100.0 184650.0 96900.0 183450.0 ;
      RECT  98100.0 184650.0 96900.0 183450.0 ;
      RECT  100500.0 184650.0 99300.0 183450.0 ;
      RECT  95700.0 174750.0 94500.0 173550.0 ;
      RECT  95700.0 184650.0 94500.0 183450.0 ;
      RECT  99900.0 180000.0 98700.0 178800.0 ;
      RECT  99900.0 180000.0 98700.0 178800.0 ;
      RECT  97350.0 179850.0 96450.0 178950.0 ;
      RECT  102300.0 172650.0 92700.0 171750.0 ;
      RECT  102300.0 186450.0 92700.0 185550.0 ;
      RECT  95700.0 197850.0 94500.0 199800.0 ;
      RECT  95700.0 186000.0 94500.0 187950.0 ;
      RECT  100500.0 187350.0 99300.0 185550.0 ;
      RECT  100500.0 196650.0 99300.0 200250.0 ;
      RECT  97800.0 187350.0 96900.0 196650.0 ;
      RECT  100500.0 196650.0 99300.0 197850.0 ;
      RECT  98100.0 196650.0 96900.0 197850.0 ;
      RECT  98100.0 196650.0 96900.0 197850.0 ;
      RECT  100500.0 196650.0 99300.0 197850.0 ;
      RECT  100500.0 187350.0 99300.0 188550.0 ;
      RECT  98100.0 187350.0 96900.0 188550.0 ;
      RECT  98100.0 187350.0 96900.0 188550.0 ;
      RECT  100500.0 187350.0 99300.0 188550.0 ;
      RECT  95700.0 197250.0 94500.0 198450.0 ;
      RECT  95700.0 187350.0 94500.0 188550.0 ;
      RECT  99900.0 192000.0 98700.0 193200.0 ;
      RECT  99900.0 192000.0 98700.0 193200.0 ;
      RECT  97350.0 192150.0 96450.0 193050.0 ;
      RECT  102300.0 199350.0 92700.0 200250.0 ;
      RECT  102300.0 185550.0 92700.0 186450.0 ;
      RECT  95700.0 201750.0 94500.0 199800.0 ;
      RECT  95700.0 213600.0 94500.0 211650.0 ;
      RECT  100500.0 212250.0 99300.0 214050.0 ;
      RECT  100500.0 202950.0 99300.0 199350.0 ;
      RECT  97800.0 212250.0 96900.0 202950.0 ;
      RECT  100500.0 202950.0 99300.0 201750.0 ;
      RECT  98100.0 202950.0 96900.0 201750.0 ;
      RECT  98100.0 202950.0 96900.0 201750.0 ;
      RECT  100500.0 202950.0 99300.0 201750.0 ;
      RECT  100500.0 212250.0 99300.0 211050.0 ;
      RECT  98100.0 212250.0 96900.0 211050.0 ;
      RECT  98100.0 212250.0 96900.0 211050.0 ;
      RECT  100500.0 212250.0 99300.0 211050.0 ;
      RECT  95700.0 202350.0 94500.0 201150.0 ;
      RECT  95700.0 212250.0 94500.0 211050.0 ;
      RECT  99900.0 207600.0 98700.0 206400.0 ;
      RECT  99900.0 207600.0 98700.0 206400.0 ;
      RECT  97350.0 207450.0 96450.0 206550.0 ;
      RECT  102300.0 200250.0 92700.0 199350.0 ;
      RECT  102300.0 214050.0 92700.0 213150.0 ;
      RECT  114900.0 160350.0 113700.0 157950.0 ;
      RECT  114900.0 169050.0 113700.0 172650.0 ;
      RECT  110100.0 169050.0 108900.0 172650.0 ;
      RECT  107700.0 170250.0 106500.0 172200.0 ;
      RECT  107700.0 158400.0 106500.0 160350.0 ;
      RECT  114900.0 169050.0 113700.0 170250.0 ;
      RECT  112500.0 169050.0 111300.0 170250.0 ;
      RECT  112500.0 169050.0 111300.0 170250.0 ;
      RECT  114900.0 169050.0 113700.0 170250.0 ;
      RECT  112500.0 169050.0 111300.0 170250.0 ;
      RECT  110100.0 169050.0 108900.0 170250.0 ;
      RECT  110100.0 169050.0 108900.0 170250.0 ;
      RECT  112500.0 169050.0 111300.0 170250.0 ;
      RECT  114900.0 160350.0 113700.0 161550.0 ;
      RECT  112500.0 160350.0 111300.0 161550.0 ;
      RECT  112500.0 160350.0 111300.0 161550.0 ;
      RECT  114900.0 160350.0 113700.0 161550.0 ;
      RECT  112500.0 160350.0 111300.0 161550.0 ;
      RECT  110100.0 160350.0 108900.0 161550.0 ;
      RECT  110100.0 160350.0 108900.0 161550.0 ;
      RECT  112500.0 160350.0 111300.0 161550.0 ;
      RECT  107700.0 169650.0 106500.0 170850.0 ;
      RECT  107700.0 159750.0 106500.0 160950.0 ;
      RECT  110100.0 162900.0 111300.0 164100.0 ;
      RECT  113100.0 165600.0 114300.0 166800.0 ;
      RECT  112500.0 169050.0 111300.0 170250.0 ;
      RECT  110100.0 160350.0 108900.0 161550.0 ;
      RECT  108900.0 165600.0 110100.0 166800.0 ;
      RECT  114300.0 165600.0 113100.0 166800.0 ;
      RECT  111300.0 162900.0 110100.0 164100.0 ;
      RECT  110100.0 165600.0 108900.0 166800.0 ;
      RECT  116700.0 171750.0 102300.0 172650.0 ;
      RECT  116700.0 157950.0 102300.0 158850.0 ;
      RECT  114900.0 184050.0 113700.0 186450.0 ;
      RECT  114900.0 175350.0 113700.0 171750.0 ;
      RECT  110100.0 175350.0 108900.0 171750.0 ;
      RECT  107700.0 174150.0 106500.0 172200.0 ;
      RECT  107700.0 186000.0 106500.0 184050.0 ;
      RECT  114900.0 175350.0 113700.0 174150.0 ;
      RECT  112500.0 175350.0 111300.0 174150.0 ;
      RECT  112500.0 175350.0 111300.0 174150.0 ;
      RECT  114900.0 175350.0 113700.0 174150.0 ;
      RECT  112500.0 175350.0 111300.0 174150.0 ;
      RECT  110100.0 175350.0 108900.0 174150.0 ;
      RECT  110100.0 175350.0 108900.0 174150.0 ;
      RECT  112500.0 175350.0 111300.0 174150.0 ;
      RECT  114900.0 184050.0 113700.0 182850.0 ;
      RECT  112500.0 184050.0 111300.0 182850.0 ;
      RECT  112500.0 184050.0 111300.0 182850.0 ;
      RECT  114900.0 184050.0 113700.0 182850.0 ;
      RECT  112500.0 184050.0 111300.0 182850.0 ;
      RECT  110100.0 184050.0 108900.0 182850.0 ;
      RECT  110100.0 184050.0 108900.0 182850.0 ;
      RECT  112500.0 184050.0 111300.0 182850.0 ;
      RECT  107700.0 174750.0 106500.0 173550.0 ;
      RECT  107700.0 184650.0 106500.0 183450.0 ;
      RECT  110100.0 181500.0 111300.0 180300.0 ;
      RECT  113100.0 178800.0 114300.0 177600.0 ;
      RECT  112500.0 175350.0 111300.0 174150.0 ;
      RECT  110100.0 184050.0 108900.0 182850.0 ;
      RECT  108900.0 178800.0 110100.0 177600.0 ;
      RECT  114300.0 178800.0 113100.0 177600.0 ;
      RECT  111300.0 181500.0 110100.0 180300.0 ;
      RECT  110100.0 178800.0 108900.0 177600.0 ;
      RECT  116700.0 172650.0 102300.0 171750.0 ;
      RECT  116700.0 186450.0 102300.0 185550.0 ;
      RECT  114900.0 187950.0 113700.0 185550.0 ;
      RECT  114900.0 196650.0 113700.0 200250.0 ;
      RECT  110100.0 196650.0 108900.0 200250.0 ;
      RECT  107700.0 197850.0 106500.0 199800.0 ;
      RECT  107700.0 186000.0 106500.0 187950.0 ;
      RECT  114900.0 196650.0 113700.0 197850.0 ;
      RECT  112500.0 196650.0 111300.0 197850.0 ;
      RECT  112500.0 196650.0 111300.0 197850.0 ;
      RECT  114900.0 196650.0 113700.0 197850.0 ;
      RECT  112500.0 196650.0 111300.0 197850.0 ;
      RECT  110100.0 196650.0 108900.0 197850.0 ;
      RECT  110100.0 196650.0 108900.0 197850.0 ;
      RECT  112500.0 196650.0 111300.0 197850.0 ;
      RECT  114900.0 187950.0 113700.0 189150.0 ;
      RECT  112500.0 187950.0 111300.0 189150.0 ;
      RECT  112500.0 187950.0 111300.0 189150.0 ;
      RECT  114900.0 187950.0 113700.0 189150.0 ;
      RECT  112500.0 187950.0 111300.0 189150.0 ;
      RECT  110100.0 187950.0 108900.0 189150.0 ;
      RECT  110100.0 187950.0 108900.0 189150.0 ;
      RECT  112500.0 187950.0 111300.0 189150.0 ;
      RECT  107700.0 197250.0 106500.0 198450.0 ;
      RECT  107700.0 187350.0 106500.0 188550.0 ;
      RECT  110100.0 190500.0 111300.0 191700.0 ;
      RECT  113100.0 193200.0 114300.0 194400.0 ;
      RECT  112500.0 196650.0 111300.0 197850.0 ;
      RECT  110100.0 187950.0 108900.0 189150.0 ;
      RECT  108900.0 193200.0 110100.0 194400.0 ;
      RECT  114300.0 193200.0 113100.0 194400.0 ;
      RECT  111300.0 190500.0 110100.0 191700.0 ;
      RECT  110100.0 193200.0 108900.0 194400.0 ;
      RECT  116700.0 199350.0 102300.0 200250.0 ;
      RECT  116700.0 185550.0 102300.0 186450.0 ;
      RECT  114900.0 211650.0 113700.0 214050.0 ;
      RECT  114900.0 202950.0 113700.0 199350.0 ;
      RECT  110100.0 202950.0 108900.0 199350.0 ;
      RECT  107700.0 201750.0 106500.0 199800.0 ;
      RECT  107700.0 213600.0 106500.0 211650.0 ;
      RECT  114900.0 202950.0 113700.0 201750.0 ;
      RECT  112500.0 202950.0 111300.0 201750.0 ;
      RECT  112500.0 202950.0 111300.0 201750.0 ;
      RECT  114900.0 202950.0 113700.0 201750.0 ;
      RECT  112500.0 202950.0 111300.0 201750.0 ;
      RECT  110100.0 202950.0 108900.0 201750.0 ;
      RECT  110100.0 202950.0 108900.0 201750.0 ;
      RECT  112500.0 202950.0 111300.0 201750.0 ;
      RECT  114900.0 211650.0 113700.0 210450.0 ;
      RECT  112500.0 211650.0 111300.0 210450.0 ;
      RECT  112500.0 211650.0 111300.0 210450.0 ;
      RECT  114900.0 211650.0 113700.0 210450.0 ;
      RECT  112500.0 211650.0 111300.0 210450.0 ;
      RECT  110100.0 211650.0 108900.0 210450.0 ;
      RECT  110100.0 211650.0 108900.0 210450.0 ;
      RECT  112500.0 211650.0 111300.0 210450.0 ;
      RECT  107700.0 202350.0 106500.0 201150.0 ;
      RECT  107700.0 212250.0 106500.0 211050.0 ;
      RECT  110100.0 209100.0 111300.0 207900.0 ;
      RECT  113100.0 206400.0 114300.0 205200.0 ;
      RECT  112500.0 202950.0 111300.0 201750.0 ;
      RECT  110100.0 211650.0 108900.0 210450.0 ;
      RECT  108900.0 206400.0 110100.0 205200.0 ;
      RECT  114300.0 206400.0 113100.0 205200.0 ;
      RECT  111300.0 209100.0 110100.0 207900.0 ;
      RECT  110100.0 206400.0 108900.0 205200.0 ;
      RECT  116700.0 200250.0 102300.0 199350.0 ;
      RECT  116700.0 214050.0 102300.0 213150.0 ;
      RECT  127650.0 168900.0 128850.0 170100.0 ;
      RECT  146250.0 164400.0 147450.0 165600.0 ;
      RECT  124650.0 182700.0 125850.0 183900.0 ;
      RECT  143250.0 178800.0 144450.0 180000.0 ;
      RECT  146250.0 187500.0 147450.0 188700.0 ;
      RECT  121650.0 187500.0 122850.0 188700.0 ;
      RECT  143250.0 201300.0 144450.0 202500.0 ;
      RECT  118650.0 201300.0 119850.0 202500.0 ;
      RECT  127650.0 165600.0 128850.0 166800.0 ;
      RECT  124650.0 162900.0 125850.0 164100.0 ;
      RECT  121650.0 177600.0 122850.0 178800.0 ;
      RECT  124650.0 180300.0 125850.0 181500.0 ;
      RECT  127650.0 193200.0 128850.0 194400.0 ;
      RECT  118650.0 190500.0 119850.0 191700.0 ;
      RECT  121650.0 205200.0 122850.0 206400.0 ;
      RECT  118650.0 207900.0 119850.0 209100.0 ;
      RECT  96450.0 164550.0 92700.0 165450.0 ;
      RECT  96450.0 178950.0 92700.0 179850.0 ;
      RECT  96450.0 192150.0 92700.0 193050.0 ;
      RECT  96450.0 206550.0 92700.0 207450.0 ;
      RECT  147300.0 171750.0 92700.0 172650.0 ;
      RECT  147300.0 199350.0 92700.0 200250.0 ;
      RECT  147300.0 157950.0 92700.0 158850.0 ;
      RECT  147300.0 185550.0 92700.0 186450.0 ;
      RECT  147300.0 213150.0 92700.0 214050.0 ;
      RECT  131250.0 219750.0 130350.0 220650.0 ;
      RECT  131250.0 224250.0 130350.0 225150.0 ;
      RECT  135450.0 219750.0 130800.0 220650.0 ;
      RECT  131250.0 220200.0 130350.0 224700.0 ;
      RECT  130800.0 224250.0 128250.0 225150.0 ;
      RECT  146850.0 219750.0 138900.0 220650.0 ;
      RECT  131250.0 234150.0 130350.0 235050.0 ;
      RECT  131250.0 238050.0 130350.0 238950.0 ;
      RECT  135450.0 234150.0 130800.0 235050.0 ;
      RECT  131250.0 234600.0 130350.0 238500.0 ;
      RECT  130800.0 238050.0 125250.0 238950.0 ;
      RECT  143850.0 234150.0 138900.0 235050.0 ;
      RECT  146850.0 242850.0 122250.0 243750.0 ;
      RECT  143850.0 256650.0 119250.0 257550.0 ;
      RECT  128250.0 220950.0 114300.0 221850.0 ;
      RECT  125250.0 218250.0 111300.0 219150.0 ;
      RECT  122250.0 232950.0 114300.0 233850.0 ;
      RECT  125250.0 235650.0 111300.0 236550.0 ;
      RECT  128250.0 248550.0 114300.0 249450.0 ;
      RECT  119250.0 245850.0 111300.0 246750.0 ;
      RECT  122250.0 260550.0 114300.0 261450.0 ;
      RECT  119250.0 263250.0 111300.0 264150.0 ;
      RECT  104850.0 220950.0 103950.0 221850.0 ;
      RECT  104850.0 219750.0 103950.0 220650.0 ;
      RECT  108900.0 220950.0 104400.0 221850.0 ;
      RECT  104850.0 220200.0 103950.0 221400.0 ;
      RECT  104400.0 219750.0 99900.0 220650.0 ;
      RECT  104850.0 232950.0 103950.0 233850.0 ;
      RECT  104850.0 234150.0 103950.0 235050.0 ;
      RECT  108900.0 232950.0 104400.0 233850.0 ;
      RECT  104850.0 233400.0 103950.0 234600.0 ;
      RECT  104400.0 234150.0 99900.0 235050.0 ;
      RECT  104850.0 248550.0 103950.0 249450.0 ;
      RECT  104850.0 247350.0 103950.0 248250.0 ;
      RECT  108900.0 248550.0 104400.0 249450.0 ;
      RECT  104850.0 247800.0 103950.0 249000.0 ;
      RECT  104400.0 247350.0 99900.0 248250.0 ;
      RECT  104850.0 260550.0 103950.0 261450.0 ;
      RECT  104850.0 261750.0 103950.0 262650.0 ;
      RECT  108900.0 260550.0 104400.0 261450.0 ;
      RECT  104850.0 261000.0 103950.0 262200.0 ;
      RECT  104400.0 261750.0 99900.0 262650.0 ;
      RECT  134700.0 225450.0 133500.0 227400.0 ;
      RECT  134700.0 213600.0 133500.0 215550.0 ;
      RECT  139500.0 214950.0 138300.0 213150.0 ;
      RECT  139500.0 224250.0 138300.0 227850.0 ;
      RECT  136800.0 214950.0 135900.0 224250.0 ;
      RECT  139500.0 224250.0 138300.0 225450.0 ;
      RECT  137100.0 224250.0 135900.0 225450.0 ;
      RECT  137100.0 224250.0 135900.0 225450.0 ;
      RECT  139500.0 224250.0 138300.0 225450.0 ;
      RECT  139500.0 214950.0 138300.0 216150.0 ;
      RECT  137100.0 214950.0 135900.0 216150.0 ;
      RECT  137100.0 214950.0 135900.0 216150.0 ;
      RECT  139500.0 214950.0 138300.0 216150.0 ;
      RECT  134700.0 224850.0 133500.0 226050.0 ;
      RECT  134700.0 214950.0 133500.0 216150.0 ;
      RECT  138900.0 219600.0 137700.0 220800.0 ;
      RECT  138900.0 219600.0 137700.0 220800.0 ;
      RECT  136350.0 219750.0 135450.0 220650.0 ;
      RECT  141300.0 226950.0 131700.0 227850.0 ;
      RECT  141300.0 213150.0 131700.0 214050.0 ;
      RECT  134700.0 229350.0 133500.0 227400.0 ;
      RECT  134700.0 241200.0 133500.0 239250.0 ;
      RECT  139500.0 239850.0 138300.0 241650.0 ;
      RECT  139500.0 230550.0 138300.0 226950.0 ;
      RECT  136800.0 239850.0 135900.0 230550.0 ;
      RECT  139500.0 230550.0 138300.0 229350.0 ;
      RECT  137100.0 230550.0 135900.0 229350.0 ;
      RECT  137100.0 230550.0 135900.0 229350.0 ;
      RECT  139500.0 230550.0 138300.0 229350.0 ;
      RECT  139500.0 239850.0 138300.0 238650.0 ;
      RECT  137100.0 239850.0 135900.0 238650.0 ;
      RECT  137100.0 239850.0 135900.0 238650.0 ;
      RECT  139500.0 239850.0 138300.0 238650.0 ;
      RECT  134700.0 229950.0 133500.0 228750.0 ;
      RECT  134700.0 239850.0 133500.0 238650.0 ;
      RECT  138900.0 235200.0 137700.0 234000.0 ;
      RECT  138900.0 235200.0 137700.0 234000.0 ;
      RECT  136350.0 235050.0 135450.0 234150.0 ;
      RECT  141300.0 227850.0 131700.0 226950.0 ;
      RECT  141300.0 241650.0 131700.0 240750.0 ;
      RECT  95700.0 225450.0 94500.0 227400.0 ;
      RECT  95700.0 213600.0 94500.0 215550.0 ;
      RECT  100500.0 214950.0 99300.0 213150.0 ;
      RECT  100500.0 224250.0 99300.0 227850.0 ;
      RECT  97800.0 214950.0 96900.0 224250.0 ;
      RECT  100500.0 224250.0 99300.0 225450.0 ;
      RECT  98100.0 224250.0 96900.0 225450.0 ;
      RECT  98100.0 224250.0 96900.0 225450.0 ;
      RECT  100500.0 224250.0 99300.0 225450.0 ;
      RECT  100500.0 214950.0 99300.0 216150.0 ;
      RECT  98100.0 214950.0 96900.0 216150.0 ;
      RECT  98100.0 214950.0 96900.0 216150.0 ;
      RECT  100500.0 214950.0 99300.0 216150.0 ;
      RECT  95700.0 224850.0 94500.0 226050.0 ;
      RECT  95700.0 214950.0 94500.0 216150.0 ;
      RECT  99900.0 219600.0 98700.0 220800.0 ;
      RECT  99900.0 219600.0 98700.0 220800.0 ;
      RECT  97350.0 219750.0 96450.0 220650.0 ;
      RECT  102300.0 226950.0 92700.0 227850.0 ;
      RECT  102300.0 213150.0 92700.0 214050.0 ;
      RECT  95700.0 229350.0 94500.0 227400.0 ;
      RECT  95700.0 241200.0 94500.0 239250.0 ;
      RECT  100500.0 239850.0 99300.0 241650.0 ;
      RECT  100500.0 230550.0 99300.0 226950.0 ;
      RECT  97800.0 239850.0 96900.0 230550.0 ;
      RECT  100500.0 230550.0 99300.0 229350.0 ;
      RECT  98100.0 230550.0 96900.0 229350.0 ;
      RECT  98100.0 230550.0 96900.0 229350.0 ;
      RECT  100500.0 230550.0 99300.0 229350.0 ;
      RECT  100500.0 239850.0 99300.0 238650.0 ;
      RECT  98100.0 239850.0 96900.0 238650.0 ;
      RECT  98100.0 239850.0 96900.0 238650.0 ;
      RECT  100500.0 239850.0 99300.0 238650.0 ;
      RECT  95700.0 229950.0 94500.0 228750.0 ;
      RECT  95700.0 239850.0 94500.0 238650.0 ;
      RECT  99900.0 235200.0 98700.0 234000.0 ;
      RECT  99900.0 235200.0 98700.0 234000.0 ;
      RECT  97350.0 235050.0 96450.0 234150.0 ;
      RECT  102300.0 227850.0 92700.0 226950.0 ;
      RECT  102300.0 241650.0 92700.0 240750.0 ;
      RECT  95700.0 253050.0 94500.0 255000.0 ;
      RECT  95700.0 241200.0 94500.0 243150.0 ;
      RECT  100500.0 242550.0 99300.0 240750.0 ;
      RECT  100500.0 251850.0 99300.0 255450.0 ;
      RECT  97800.0 242550.0 96900.0 251850.0 ;
      RECT  100500.0 251850.0 99300.0 253050.0 ;
      RECT  98100.0 251850.0 96900.0 253050.0 ;
      RECT  98100.0 251850.0 96900.0 253050.0 ;
      RECT  100500.0 251850.0 99300.0 253050.0 ;
      RECT  100500.0 242550.0 99300.0 243750.0 ;
      RECT  98100.0 242550.0 96900.0 243750.0 ;
      RECT  98100.0 242550.0 96900.0 243750.0 ;
      RECT  100500.0 242550.0 99300.0 243750.0 ;
      RECT  95700.0 252450.0 94500.0 253650.0 ;
      RECT  95700.0 242550.0 94500.0 243750.0 ;
      RECT  99900.0 247200.0 98700.0 248400.0 ;
      RECT  99900.0 247200.0 98700.0 248400.0 ;
      RECT  97350.0 247350.0 96450.0 248250.0 ;
      RECT  102300.0 254550.0 92700.0 255450.0 ;
      RECT  102300.0 240750.0 92700.0 241650.0 ;
      RECT  95700.0 256950.0 94500.0 255000.0 ;
      RECT  95700.0 268800.0 94500.0 266850.0 ;
      RECT  100500.0 267450.0 99300.0 269250.0 ;
      RECT  100500.0 258150.0 99300.0 254550.0 ;
      RECT  97800.0 267450.0 96900.0 258150.0 ;
      RECT  100500.0 258150.0 99300.0 256950.0 ;
      RECT  98100.0 258150.0 96900.0 256950.0 ;
      RECT  98100.0 258150.0 96900.0 256950.0 ;
      RECT  100500.0 258150.0 99300.0 256950.0 ;
      RECT  100500.0 267450.0 99300.0 266250.0 ;
      RECT  98100.0 267450.0 96900.0 266250.0 ;
      RECT  98100.0 267450.0 96900.0 266250.0 ;
      RECT  100500.0 267450.0 99300.0 266250.0 ;
      RECT  95700.0 257550.0 94500.0 256350.0 ;
      RECT  95700.0 267450.0 94500.0 266250.0 ;
      RECT  99900.0 262800.0 98700.0 261600.0 ;
      RECT  99900.0 262800.0 98700.0 261600.0 ;
      RECT  97350.0 262650.0 96450.0 261750.0 ;
      RECT  102300.0 255450.0 92700.0 254550.0 ;
      RECT  102300.0 269250.0 92700.0 268350.0 ;
      RECT  114900.0 215550.0 113700.0 213150.0 ;
      RECT  114900.0 224250.0 113700.0 227850.0 ;
      RECT  110100.0 224250.0 108900.0 227850.0 ;
      RECT  107700.0 225450.0 106500.0 227400.0 ;
      RECT  107700.0 213600.0 106500.0 215550.0 ;
      RECT  114900.0 224250.0 113700.0 225450.0 ;
      RECT  112500.0 224250.0 111300.0 225450.0 ;
      RECT  112500.0 224250.0 111300.0 225450.0 ;
      RECT  114900.0 224250.0 113700.0 225450.0 ;
      RECT  112500.0 224250.0 111300.0 225450.0 ;
      RECT  110100.0 224250.0 108900.0 225450.0 ;
      RECT  110100.0 224250.0 108900.0 225450.0 ;
      RECT  112500.0 224250.0 111300.0 225450.0 ;
      RECT  114900.0 215550.0 113700.0 216750.0 ;
      RECT  112500.0 215550.0 111300.0 216750.0 ;
      RECT  112500.0 215550.0 111300.0 216750.0 ;
      RECT  114900.0 215550.0 113700.0 216750.0 ;
      RECT  112500.0 215550.0 111300.0 216750.0 ;
      RECT  110100.0 215550.0 108900.0 216750.0 ;
      RECT  110100.0 215550.0 108900.0 216750.0 ;
      RECT  112500.0 215550.0 111300.0 216750.0 ;
      RECT  107700.0 224850.0 106500.0 226050.0 ;
      RECT  107700.0 214950.0 106500.0 216150.0 ;
      RECT  110100.0 218100.0 111300.0 219300.0 ;
      RECT  113100.0 220800.0 114300.0 222000.0 ;
      RECT  112500.0 224250.0 111300.0 225450.0 ;
      RECT  110100.0 215550.0 108900.0 216750.0 ;
      RECT  108900.0 220800.0 110100.0 222000.0 ;
      RECT  114300.0 220800.0 113100.0 222000.0 ;
      RECT  111300.0 218100.0 110100.0 219300.0 ;
      RECT  110100.0 220800.0 108900.0 222000.0 ;
      RECT  116700.0 226950.0 102300.0 227850.0 ;
      RECT  116700.0 213150.0 102300.0 214050.0 ;
      RECT  114900.0 239250.0 113700.0 241650.0 ;
      RECT  114900.0 230550.0 113700.0 226950.0 ;
      RECT  110100.0 230550.0 108900.0 226950.0 ;
      RECT  107700.0 229350.0 106500.0 227400.0 ;
      RECT  107700.0 241200.0 106500.0 239250.0 ;
      RECT  114900.0 230550.0 113700.0 229350.0 ;
      RECT  112500.0 230550.0 111300.0 229350.0 ;
      RECT  112500.0 230550.0 111300.0 229350.0 ;
      RECT  114900.0 230550.0 113700.0 229350.0 ;
      RECT  112500.0 230550.0 111300.0 229350.0 ;
      RECT  110100.0 230550.0 108900.0 229350.0 ;
      RECT  110100.0 230550.0 108900.0 229350.0 ;
      RECT  112500.0 230550.0 111300.0 229350.0 ;
      RECT  114900.0 239250.0 113700.0 238050.0 ;
      RECT  112500.0 239250.0 111300.0 238050.0 ;
      RECT  112500.0 239250.0 111300.0 238050.0 ;
      RECT  114900.0 239250.0 113700.0 238050.0 ;
      RECT  112500.0 239250.0 111300.0 238050.0 ;
      RECT  110100.0 239250.0 108900.0 238050.0 ;
      RECT  110100.0 239250.0 108900.0 238050.0 ;
      RECT  112500.0 239250.0 111300.0 238050.0 ;
      RECT  107700.0 229950.0 106500.0 228750.0 ;
      RECT  107700.0 239850.0 106500.0 238650.0 ;
      RECT  110100.0 236700.0 111300.0 235500.0 ;
      RECT  113100.0 234000.0 114300.0 232800.0 ;
      RECT  112500.0 230550.0 111300.0 229350.0 ;
      RECT  110100.0 239250.0 108900.0 238050.0 ;
      RECT  108900.0 234000.0 110100.0 232800.0 ;
      RECT  114300.0 234000.0 113100.0 232800.0 ;
      RECT  111300.0 236700.0 110100.0 235500.0 ;
      RECT  110100.0 234000.0 108900.0 232800.0 ;
      RECT  116700.0 227850.0 102300.0 226950.0 ;
      RECT  116700.0 241650.0 102300.0 240750.0 ;
      RECT  114900.0 243150.0 113700.0 240750.0 ;
      RECT  114900.0 251850.0 113700.0 255450.0 ;
      RECT  110100.0 251850.0 108900.0 255450.0 ;
      RECT  107700.0 253050.0 106500.0 255000.0 ;
      RECT  107700.0 241200.0 106500.0 243150.0 ;
      RECT  114900.0 251850.0 113700.0 253050.0 ;
      RECT  112500.0 251850.0 111300.0 253050.0 ;
      RECT  112500.0 251850.0 111300.0 253050.0 ;
      RECT  114900.0 251850.0 113700.0 253050.0 ;
      RECT  112500.0 251850.0 111300.0 253050.0 ;
      RECT  110100.0 251850.0 108900.0 253050.0 ;
      RECT  110100.0 251850.0 108900.0 253050.0 ;
      RECT  112500.0 251850.0 111300.0 253050.0 ;
      RECT  114900.0 243150.0 113700.0 244350.0 ;
      RECT  112500.0 243150.0 111300.0 244350.0 ;
      RECT  112500.0 243150.0 111300.0 244350.0 ;
      RECT  114900.0 243150.0 113700.0 244350.0 ;
      RECT  112500.0 243150.0 111300.0 244350.0 ;
      RECT  110100.0 243150.0 108900.0 244350.0 ;
      RECT  110100.0 243150.0 108900.0 244350.0 ;
      RECT  112500.0 243150.0 111300.0 244350.0 ;
      RECT  107700.0 252450.0 106500.0 253650.0 ;
      RECT  107700.0 242550.0 106500.0 243750.0 ;
      RECT  110100.0 245700.0 111300.0 246900.0 ;
      RECT  113100.0 248400.0 114300.0 249600.0 ;
      RECT  112500.0 251850.0 111300.0 253050.0 ;
      RECT  110100.0 243150.0 108900.0 244350.0 ;
      RECT  108900.0 248400.0 110100.0 249600.0 ;
      RECT  114300.0 248400.0 113100.0 249600.0 ;
      RECT  111300.0 245700.0 110100.0 246900.0 ;
      RECT  110100.0 248400.0 108900.0 249600.0 ;
      RECT  116700.0 254550.0 102300.0 255450.0 ;
      RECT  116700.0 240750.0 102300.0 241650.0 ;
      RECT  114900.0 266850.0 113700.0 269250.0 ;
      RECT  114900.0 258150.0 113700.0 254550.0 ;
      RECT  110100.0 258150.0 108900.0 254550.0 ;
      RECT  107700.0 256950.0 106500.0 255000.0 ;
      RECT  107700.0 268800.0 106500.0 266850.0 ;
      RECT  114900.0 258150.0 113700.0 256950.0 ;
      RECT  112500.0 258150.0 111300.0 256950.0 ;
      RECT  112500.0 258150.0 111300.0 256950.0 ;
      RECT  114900.0 258150.0 113700.0 256950.0 ;
      RECT  112500.0 258150.0 111300.0 256950.0 ;
      RECT  110100.0 258150.0 108900.0 256950.0 ;
      RECT  110100.0 258150.0 108900.0 256950.0 ;
      RECT  112500.0 258150.0 111300.0 256950.0 ;
      RECT  114900.0 266850.0 113700.0 265650.0 ;
      RECT  112500.0 266850.0 111300.0 265650.0 ;
      RECT  112500.0 266850.0 111300.0 265650.0 ;
      RECT  114900.0 266850.0 113700.0 265650.0 ;
      RECT  112500.0 266850.0 111300.0 265650.0 ;
      RECT  110100.0 266850.0 108900.0 265650.0 ;
      RECT  110100.0 266850.0 108900.0 265650.0 ;
      RECT  112500.0 266850.0 111300.0 265650.0 ;
      RECT  107700.0 257550.0 106500.0 256350.0 ;
      RECT  107700.0 267450.0 106500.0 266250.0 ;
      RECT  110100.0 264300.0 111300.0 263100.0 ;
      RECT  113100.0 261600.0 114300.0 260400.0 ;
      RECT  112500.0 258150.0 111300.0 256950.0 ;
      RECT  110100.0 266850.0 108900.0 265650.0 ;
      RECT  108900.0 261600.0 110100.0 260400.0 ;
      RECT  114300.0 261600.0 113100.0 260400.0 ;
      RECT  111300.0 264300.0 110100.0 263100.0 ;
      RECT  110100.0 261600.0 108900.0 260400.0 ;
      RECT  116700.0 255450.0 102300.0 254550.0 ;
      RECT  116700.0 269250.0 102300.0 268350.0 ;
      RECT  127650.0 224100.0 128850.0 225300.0 ;
      RECT  146250.0 219600.0 147450.0 220800.0 ;
      RECT  124650.0 237900.0 125850.0 239100.0 ;
      RECT  143250.0 234000.0 144450.0 235200.0 ;
      RECT  146250.0 242700.0 147450.0 243900.0 ;
      RECT  121650.0 242700.0 122850.0 243900.0 ;
      RECT  143250.0 256500.0 144450.0 257700.0 ;
      RECT  118650.0 256500.0 119850.0 257700.0 ;
      RECT  127650.0 220800.0 128850.0 222000.0 ;
      RECT  124650.0 218100.0 125850.0 219300.0 ;
      RECT  121650.0 232800.0 122850.0 234000.0 ;
      RECT  124650.0 235500.0 125850.0 236700.0 ;
      RECT  127650.0 248400.0 128850.0 249600.0 ;
      RECT  118650.0 245700.0 119850.0 246900.0 ;
      RECT  121650.0 260400.0 122850.0 261600.0 ;
      RECT  118650.0 263100.0 119850.0 264300.0 ;
      RECT  96450.0 219750.0 92700.0 220650.0 ;
      RECT  96450.0 234150.0 92700.0 235050.0 ;
      RECT  96450.0 247350.0 92700.0 248250.0 ;
      RECT  96450.0 261750.0 92700.0 262650.0 ;
      RECT  147300.0 226950.0 92700.0 227850.0 ;
      RECT  147300.0 254550.0 92700.0 255450.0 ;
      RECT  147300.0 213150.0 92700.0 214050.0 ;
      RECT  147300.0 240750.0 92700.0 241650.0 ;
      RECT  147300.0 268350.0 92700.0 269250.0 ;
      RECT  138450.0 274950.0 137550.0 275850.0 ;
      RECT  138450.0 279450.0 137550.0 280350.0 ;
      RECT  142650.0 274950.0 138000.0 275850.0 ;
      RECT  138450.0 275400.0 137550.0 279900.0 ;
      RECT  138000.0 279450.0 135450.0 280350.0 ;
      RECT  157050.0 274950.0 146100.0 275850.0 ;
      RECT  138450.0 289350.0 137550.0 290250.0 ;
      RECT  138450.0 293250.0 137550.0 294150.0 ;
      RECT  142650.0 289350.0 138000.0 290250.0 ;
      RECT  138450.0 289800.0 137550.0 293700.0 ;
      RECT  138000.0 293250.0 132450.0 294150.0 ;
      RECT  154050.0 289350.0 146100.0 290250.0 ;
      RECT  138450.0 302550.0 137550.0 303450.0 ;
      RECT  138450.0 307050.0 137550.0 307950.0 ;
      RECT  142650.0 302550.0 138000.0 303450.0 ;
      RECT  138450.0 303000.0 137550.0 307500.0 ;
      RECT  138000.0 307050.0 129450.0 307950.0 ;
      RECT  151050.0 302550.0 146100.0 303450.0 ;
      RECT  157050.0 311850.0 126450.0 312750.0 ;
      RECT  154050.0 325650.0 123450.0 326550.0 ;
      RECT  151050.0 339450.0 120450.0 340350.0 ;
      RECT  135450.0 276900.0 114900.0 277800.0 ;
      RECT  132450.0 274950.0 112500.0 275850.0 ;
      RECT  129450.0 273000.0 110100.0 273900.0 ;
      RECT  126450.0 287400.0 114900.0 288300.0 ;
      RECT  132450.0 289350.0 112500.0 290250.0 ;
      RECT  129450.0 291300.0 110100.0 292200.0 ;
      RECT  135450.0 304500.0 114900.0 305400.0 ;
      RECT  123450.0 302550.0 112500.0 303450.0 ;
      RECT  129450.0 300600.0 110100.0 301500.0 ;
      RECT  126450.0 315000.0 114900.0 315900.0 ;
      RECT  123450.0 316950.0 112500.0 317850.0 ;
      RECT  129450.0 318900.0 110100.0 319800.0 ;
      RECT  135450.0 332100.0 114900.0 333000.0 ;
      RECT  132450.0 330150.0 112500.0 331050.0 ;
      RECT  120450.0 328200.0 110100.0 329100.0 ;
      RECT  126450.0 342600.0 114900.0 343500.0 ;
      RECT  132450.0 344550.0 112500.0 345450.0 ;
      RECT  120450.0 346500.0 110100.0 347400.0 ;
      RECT  135450.0 359700.0 114900.0 360600.0 ;
      RECT  123450.0 357750.0 112500.0 358650.0 ;
      RECT  120450.0 355800.0 110100.0 356700.0 ;
      RECT  126450.0 370200.0 114900.0 371100.0 ;
      RECT  123450.0 372150.0 112500.0 373050.0 ;
      RECT  120450.0 374100.0 110100.0 375000.0 ;
      RECT  104250.0 276900.0 103350.0 277800.0 ;
      RECT  104250.0 274950.0 103350.0 275850.0 ;
      RECT  107700.0 276900.0 103800.0 277800.0 ;
      RECT  104250.0 275400.0 103350.0 277350.0 ;
      RECT  103800.0 274950.0 99900.0 275850.0 ;
      RECT  104250.0 287400.0 103350.0 288300.0 ;
      RECT  104250.0 289350.0 103350.0 290250.0 ;
      RECT  107700.0 287400.0 103800.0 288300.0 ;
      RECT  104250.0 287850.0 103350.0 289800.0 ;
      RECT  103800.0 289350.0 99900.0 290250.0 ;
      RECT  104250.0 304500.0 103350.0 305400.0 ;
      RECT  104250.0 302550.0 103350.0 303450.0 ;
      RECT  107700.0 304500.0 103800.0 305400.0 ;
      RECT  104250.0 303000.0 103350.0 304950.0 ;
      RECT  103800.0 302550.0 99900.0 303450.0 ;
      RECT  104250.0 315000.0 103350.0 315900.0 ;
      RECT  104250.0 316950.0 103350.0 317850.0 ;
      RECT  107700.0 315000.0 103800.0 315900.0 ;
      RECT  104250.0 315450.0 103350.0 317400.0 ;
      RECT  103800.0 316950.0 99900.0 317850.0 ;
      RECT  104250.0 332100.0 103350.0 333000.0 ;
      RECT  104250.0 330150.0 103350.0 331050.0 ;
      RECT  107700.0 332100.0 103800.0 333000.0 ;
      RECT  104250.0 330600.0 103350.0 332550.0 ;
      RECT  103800.0 330150.0 99900.0 331050.0 ;
      RECT  104250.0 342600.0 103350.0 343500.0 ;
      RECT  104250.0 344550.0 103350.0 345450.0 ;
      RECT  107700.0 342600.0 103800.0 343500.0 ;
      RECT  104250.0 343050.0 103350.0 345000.0 ;
      RECT  103800.0 344550.0 99900.0 345450.0 ;
      RECT  104250.0 359700.0 103350.0 360600.0 ;
      RECT  104250.0 357750.0 103350.0 358650.0 ;
      RECT  107700.0 359700.0 103800.0 360600.0 ;
      RECT  104250.0 358200.0 103350.0 360150.0 ;
      RECT  103800.0 357750.0 99900.0 358650.0 ;
      RECT  104250.0 370200.0 103350.0 371100.0 ;
      RECT  104250.0 372150.0 103350.0 373050.0 ;
      RECT  107700.0 370200.0 103800.0 371100.0 ;
      RECT  104250.0 370650.0 103350.0 372600.0 ;
      RECT  103800.0 372150.0 99900.0 373050.0 ;
      RECT  141900.0 280650.0 140700.0 282600.0 ;
      RECT  141900.0 268800.0 140700.0 270750.0 ;
      RECT  146700.0 270150.0 145500.0 268350.0 ;
      RECT  146700.0 279450.0 145500.0 283050.0 ;
      RECT  144000.0 270150.0 143100.0 279450.0 ;
      RECT  146700.0 279450.0 145500.0 280650.0 ;
      RECT  144300.0 279450.0 143100.0 280650.0 ;
      RECT  144300.0 279450.0 143100.0 280650.0 ;
      RECT  146700.0 279450.0 145500.0 280650.0 ;
      RECT  146700.0 270150.0 145500.0 271350.0 ;
      RECT  144300.0 270150.0 143100.0 271350.0 ;
      RECT  144300.0 270150.0 143100.0 271350.0 ;
      RECT  146700.0 270150.0 145500.0 271350.0 ;
      RECT  141900.0 280050.0 140700.0 281250.0 ;
      RECT  141900.0 270150.0 140700.0 271350.0 ;
      RECT  146100.0 274800.0 144900.0 276000.0 ;
      RECT  146100.0 274800.0 144900.0 276000.0 ;
      RECT  143550.0 274950.0 142650.0 275850.0 ;
      RECT  148500.0 282150.0 138900.0 283050.0 ;
      RECT  148500.0 268350.0 138900.0 269250.0 ;
      RECT  141900.0 284550.0 140700.0 282600.0 ;
      RECT  141900.0 296400.0 140700.0 294450.0 ;
      RECT  146700.0 295050.0 145500.0 296850.0 ;
      RECT  146700.0 285750.0 145500.0 282150.0 ;
      RECT  144000.0 295050.0 143100.0 285750.0 ;
      RECT  146700.0 285750.0 145500.0 284550.0 ;
      RECT  144300.0 285750.0 143100.0 284550.0 ;
      RECT  144300.0 285750.0 143100.0 284550.0 ;
      RECT  146700.0 285750.0 145500.0 284550.0 ;
      RECT  146700.0 295050.0 145500.0 293850.0 ;
      RECT  144300.0 295050.0 143100.0 293850.0 ;
      RECT  144300.0 295050.0 143100.0 293850.0 ;
      RECT  146700.0 295050.0 145500.0 293850.0 ;
      RECT  141900.0 285150.0 140700.0 283950.0 ;
      RECT  141900.0 295050.0 140700.0 293850.0 ;
      RECT  146100.0 290400.0 144900.0 289200.0 ;
      RECT  146100.0 290400.0 144900.0 289200.0 ;
      RECT  143550.0 290250.0 142650.0 289350.0 ;
      RECT  148500.0 283050.0 138900.0 282150.0 ;
      RECT  148500.0 296850.0 138900.0 295950.0 ;
      RECT  141900.0 308250.0 140700.0 310200.0 ;
      RECT  141900.0 296400.0 140700.0 298350.0 ;
      RECT  146700.0 297750.0 145500.0 295950.0 ;
      RECT  146700.0 307050.0 145500.0 310650.0 ;
      RECT  144000.0 297750.0 143100.0 307050.0 ;
      RECT  146700.0 307050.0 145500.0 308250.0 ;
      RECT  144300.0 307050.0 143100.0 308250.0 ;
      RECT  144300.0 307050.0 143100.0 308250.0 ;
      RECT  146700.0 307050.0 145500.0 308250.0 ;
      RECT  146700.0 297750.0 145500.0 298950.0 ;
      RECT  144300.0 297750.0 143100.0 298950.0 ;
      RECT  144300.0 297750.0 143100.0 298950.0 ;
      RECT  146700.0 297750.0 145500.0 298950.0 ;
      RECT  141900.0 307650.0 140700.0 308850.0 ;
      RECT  141900.0 297750.0 140700.0 298950.0 ;
      RECT  146100.0 302400.0 144900.0 303600.0 ;
      RECT  146100.0 302400.0 144900.0 303600.0 ;
      RECT  143550.0 302550.0 142650.0 303450.0 ;
      RECT  148500.0 309750.0 138900.0 310650.0 ;
      RECT  148500.0 295950.0 138900.0 296850.0 ;
      RECT  95700.0 280650.0 94500.0 282600.0 ;
      RECT  95700.0 268800.0 94500.0 270750.0 ;
      RECT  100500.0 270150.0 99300.0 268350.0 ;
      RECT  100500.0 279450.0 99300.0 283050.0 ;
      RECT  97800.0 270150.0 96900.0 279450.0 ;
      RECT  100500.0 279450.0 99300.0 280650.0 ;
      RECT  98100.0 279450.0 96900.0 280650.0 ;
      RECT  98100.0 279450.0 96900.0 280650.0 ;
      RECT  100500.0 279450.0 99300.0 280650.0 ;
      RECT  100500.0 270150.0 99300.0 271350.0 ;
      RECT  98100.0 270150.0 96900.0 271350.0 ;
      RECT  98100.0 270150.0 96900.0 271350.0 ;
      RECT  100500.0 270150.0 99300.0 271350.0 ;
      RECT  95700.0 280050.0 94500.0 281250.0 ;
      RECT  95700.0 270150.0 94500.0 271350.0 ;
      RECT  99900.0 274800.0 98700.0 276000.0 ;
      RECT  99900.0 274800.0 98700.0 276000.0 ;
      RECT  97350.0 274950.0 96450.0 275850.0 ;
      RECT  102300.0 282150.0 92700.0 283050.0 ;
      RECT  102300.0 268350.0 92700.0 269250.0 ;
      RECT  95700.0 284550.0 94500.0 282600.0 ;
      RECT  95700.0 296400.0 94500.0 294450.0 ;
      RECT  100500.0 295050.0 99300.0 296850.0 ;
      RECT  100500.0 285750.0 99300.0 282150.0 ;
      RECT  97800.0 295050.0 96900.0 285750.0 ;
      RECT  100500.0 285750.0 99300.0 284550.0 ;
      RECT  98100.0 285750.0 96900.0 284550.0 ;
      RECT  98100.0 285750.0 96900.0 284550.0 ;
      RECT  100500.0 285750.0 99300.0 284550.0 ;
      RECT  100500.0 295050.0 99300.0 293850.0 ;
      RECT  98100.0 295050.0 96900.0 293850.0 ;
      RECT  98100.0 295050.0 96900.0 293850.0 ;
      RECT  100500.0 295050.0 99300.0 293850.0 ;
      RECT  95700.0 285150.0 94500.0 283950.0 ;
      RECT  95700.0 295050.0 94500.0 293850.0 ;
      RECT  99900.0 290400.0 98700.0 289200.0 ;
      RECT  99900.0 290400.0 98700.0 289200.0 ;
      RECT  97350.0 290250.0 96450.0 289350.0 ;
      RECT  102300.0 283050.0 92700.0 282150.0 ;
      RECT  102300.0 296850.0 92700.0 295950.0 ;
      RECT  95700.0 308250.0 94500.0 310200.0 ;
      RECT  95700.0 296400.0 94500.0 298350.0 ;
      RECT  100500.0 297750.0 99300.0 295950.0 ;
      RECT  100500.0 307050.0 99300.0 310650.0 ;
      RECT  97800.0 297750.0 96900.0 307050.0 ;
      RECT  100500.0 307050.0 99300.0 308250.0 ;
      RECT  98100.0 307050.0 96900.0 308250.0 ;
      RECT  98100.0 307050.0 96900.0 308250.0 ;
      RECT  100500.0 307050.0 99300.0 308250.0 ;
      RECT  100500.0 297750.0 99300.0 298950.0 ;
      RECT  98100.0 297750.0 96900.0 298950.0 ;
      RECT  98100.0 297750.0 96900.0 298950.0 ;
      RECT  100500.0 297750.0 99300.0 298950.0 ;
      RECT  95700.0 307650.0 94500.0 308850.0 ;
      RECT  95700.0 297750.0 94500.0 298950.0 ;
      RECT  99900.0 302400.0 98700.0 303600.0 ;
      RECT  99900.0 302400.0 98700.0 303600.0 ;
      RECT  97350.0 302550.0 96450.0 303450.0 ;
      RECT  102300.0 309750.0 92700.0 310650.0 ;
      RECT  102300.0 295950.0 92700.0 296850.0 ;
      RECT  95700.0 312150.0 94500.0 310200.0 ;
      RECT  95700.0 324000.0 94500.0 322050.0 ;
      RECT  100500.0 322650.0 99300.0 324450.0 ;
      RECT  100500.0 313350.0 99300.0 309750.0 ;
      RECT  97800.0 322650.0 96900.0 313350.0 ;
      RECT  100500.0 313350.0 99300.0 312150.0 ;
      RECT  98100.0 313350.0 96900.0 312150.0 ;
      RECT  98100.0 313350.0 96900.0 312150.0 ;
      RECT  100500.0 313350.0 99300.0 312150.0 ;
      RECT  100500.0 322650.0 99300.0 321450.0 ;
      RECT  98100.0 322650.0 96900.0 321450.0 ;
      RECT  98100.0 322650.0 96900.0 321450.0 ;
      RECT  100500.0 322650.0 99300.0 321450.0 ;
      RECT  95700.0 312750.0 94500.0 311550.0 ;
      RECT  95700.0 322650.0 94500.0 321450.0 ;
      RECT  99900.0 318000.0 98700.0 316800.0 ;
      RECT  99900.0 318000.0 98700.0 316800.0 ;
      RECT  97350.0 317850.0 96450.0 316950.0 ;
      RECT  102300.0 310650.0 92700.0 309750.0 ;
      RECT  102300.0 324450.0 92700.0 323550.0 ;
      RECT  95700.0 335850.0 94500.0 337800.0 ;
      RECT  95700.0 324000.0 94500.0 325950.0 ;
      RECT  100500.0 325350.0 99300.0 323550.0 ;
      RECT  100500.0 334650.0 99300.0 338250.0 ;
      RECT  97800.0 325350.0 96900.0 334650.0 ;
      RECT  100500.0 334650.0 99300.0 335850.0 ;
      RECT  98100.0 334650.0 96900.0 335850.0 ;
      RECT  98100.0 334650.0 96900.0 335850.0 ;
      RECT  100500.0 334650.0 99300.0 335850.0 ;
      RECT  100500.0 325350.0 99300.0 326550.0 ;
      RECT  98100.0 325350.0 96900.0 326550.0 ;
      RECT  98100.0 325350.0 96900.0 326550.0 ;
      RECT  100500.0 325350.0 99300.0 326550.0 ;
      RECT  95700.0 335250.0 94500.0 336450.0 ;
      RECT  95700.0 325350.0 94500.0 326550.0 ;
      RECT  99900.0 330000.0 98700.0 331200.0 ;
      RECT  99900.0 330000.0 98700.0 331200.0 ;
      RECT  97350.0 330150.0 96450.0 331050.0 ;
      RECT  102300.0 337350.0 92700.0 338250.0 ;
      RECT  102300.0 323550.0 92700.0 324450.0 ;
      RECT  95700.0 339750.0 94500.0 337800.0 ;
      RECT  95700.0 351600.0 94500.0 349650.0 ;
      RECT  100500.0 350250.0 99300.0 352050.0 ;
      RECT  100500.0 340950.0 99300.0 337350.0 ;
      RECT  97800.0 350250.0 96900.0 340950.0 ;
      RECT  100500.0 340950.0 99300.0 339750.0 ;
      RECT  98100.0 340950.0 96900.0 339750.0 ;
      RECT  98100.0 340950.0 96900.0 339750.0 ;
      RECT  100500.0 340950.0 99300.0 339750.0 ;
      RECT  100500.0 350250.0 99300.0 349050.0 ;
      RECT  98100.0 350250.0 96900.0 349050.0 ;
      RECT  98100.0 350250.0 96900.0 349050.0 ;
      RECT  100500.0 350250.0 99300.0 349050.0 ;
      RECT  95700.0 340350.0 94500.0 339150.0 ;
      RECT  95700.0 350250.0 94500.0 349050.0 ;
      RECT  99900.0 345600.0 98700.0 344400.0 ;
      RECT  99900.0 345600.0 98700.0 344400.0 ;
      RECT  97350.0 345450.0 96450.0 344550.0 ;
      RECT  102300.0 338250.0 92700.0 337350.0 ;
      RECT  102300.0 352050.0 92700.0 351150.0 ;
      RECT  95700.0 363450.0 94500.0 365400.0 ;
      RECT  95700.0 351600.0 94500.0 353550.0 ;
      RECT  100500.0 352950.0 99300.0 351150.0 ;
      RECT  100500.0 362250.0 99300.0 365850.0 ;
      RECT  97800.0 352950.0 96900.0 362250.0 ;
      RECT  100500.0 362250.0 99300.0 363450.0 ;
      RECT  98100.0 362250.0 96900.0 363450.0 ;
      RECT  98100.0 362250.0 96900.0 363450.0 ;
      RECT  100500.0 362250.0 99300.0 363450.0 ;
      RECT  100500.0 352950.0 99300.0 354150.0 ;
      RECT  98100.0 352950.0 96900.0 354150.0 ;
      RECT  98100.0 352950.0 96900.0 354150.0 ;
      RECT  100500.0 352950.0 99300.0 354150.0 ;
      RECT  95700.0 362850.0 94500.0 364050.0 ;
      RECT  95700.0 352950.0 94500.0 354150.0 ;
      RECT  99900.0 357600.0 98700.0 358800.0 ;
      RECT  99900.0 357600.0 98700.0 358800.0 ;
      RECT  97350.0 357750.0 96450.0 358650.0 ;
      RECT  102300.0 364950.0 92700.0 365850.0 ;
      RECT  102300.0 351150.0 92700.0 352050.0 ;
      RECT  95700.0 367350.0 94500.0 365400.0 ;
      RECT  95700.0 379200.0 94500.0 377250.0 ;
      RECT  100500.0 377850.0 99300.0 379650.0 ;
      RECT  100500.0 368550.0 99300.0 364950.0 ;
      RECT  97800.0 377850.0 96900.0 368550.0 ;
      RECT  100500.0 368550.0 99300.0 367350.0 ;
      RECT  98100.0 368550.0 96900.0 367350.0 ;
      RECT  98100.0 368550.0 96900.0 367350.0 ;
      RECT  100500.0 368550.0 99300.0 367350.0 ;
      RECT  100500.0 377850.0 99300.0 376650.0 ;
      RECT  98100.0 377850.0 96900.0 376650.0 ;
      RECT  98100.0 377850.0 96900.0 376650.0 ;
      RECT  100500.0 377850.0 99300.0 376650.0 ;
      RECT  95700.0 367950.0 94500.0 366750.0 ;
      RECT  95700.0 377850.0 94500.0 376650.0 ;
      RECT  99900.0 373200.0 98700.0 372000.0 ;
      RECT  99900.0 373200.0 98700.0 372000.0 ;
      RECT  97350.0 373050.0 96450.0 372150.0 ;
      RECT  102300.0 365850.0 92700.0 364950.0 ;
      RECT  102300.0 379650.0 92700.0 378750.0 ;
      RECT  116100.0 270750.0 114900.0 268350.0 ;
      RECT  116100.0 279450.0 114900.0 283050.0 ;
      RECT  111300.0 279450.0 110100.0 283050.0 ;
      RECT  106500.0 280650.0 105300.0 282600.0 ;
      RECT  106500.0 268800.0 105300.0 270750.0 ;
      RECT  116100.0 279450.0 114900.0 280650.0 ;
      RECT  113700.0 279450.0 112500.0 280650.0 ;
      RECT  113700.0 279450.0 112500.0 280650.0 ;
      RECT  116100.0 279450.0 114900.0 280650.0 ;
      RECT  113700.0 279450.0 112500.0 280650.0 ;
      RECT  111300.0 279450.0 110100.0 280650.0 ;
      RECT  111300.0 279450.0 110100.0 280650.0 ;
      RECT  113700.0 279450.0 112500.0 280650.0 ;
      RECT  111300.0 279450.0 110100.0 280650.0 ;
      RECT  108900.0 279450.0 107700.0 280650.0 ;
      RECT  108900.0 279450.0 107700.0 280650.0 ;
      RECT  111300.0 279450.0 110100.0 280650.0 ;
      RECT  116100.0 270750.0 114900.0 271950.0 ;
      RECT  113700.0 270750.0 112500.0 271950.0 ;
      RECT  113700.0 270750.0 112500.0 271950.0 ;
      RECT  116100.0 270750.0 114900.0 271950.0 ;
      RECT  113700.0 270750.0 112500.0 271950.0 ;
      RECT  111300.0 270750.0 110100.0 271950.0 ;
      RECT  111300.0 270750.0 110100.0 271950.0 ;
      RECT  113700.0 270750.0 112500.0 271950.0 ;
      RECT  111300.0 270750.0 110100.0 271950.0 ;
      RECT  108900.0 270750.0 107700.0 271950.0 ;
      RECT  108900.0 270750.0 107700.0 271950.0 ;
      RECT  111300.0 270750.0 110100.0 271950.0 ;
      RECT  106500.0 280050.0 105300.0 281250.0 ;
      RECT  106500.0 270150.0 105300.0 271350.0 ;
      RECT  108900.0 272850.0 110100.0 274050.0 ;
      RECT  111300.0 274800.0 112500.0 276000.0 ;
      RECT  113700.0 276750.0 114900.0 277950.0 ;
      RECT  113700.0 279450.0 112500.0 280650.0 ;
      RECT  108900.0 279450.0 107700.0 280650.0 ;
      RECT  108900.0 270750.0 107700.0 271950.0 ;
      RECT  108900.0 276750.0 107700.0 277950.0 ;
      RECT  114900.0 276750.0 113700.0 277950.0 ;
      RECT  112500.0 274800.0 111300.0 276000.0 ;
      RECT  110100.0 272850.0 108900.0 274050.0 ;
      RECT  108900.0 276750.0 107700.0 277950.0 ;
      RECT  117900.0 282150.0 102300.0 283050.0 ;
      RECT  117900.0 268350.0 102300.0 269250.0 ;
      RECT  116100.0 294450.0 114900.0 296850.0 ;
      RECT  116100.0 285750.0 114900.0 282150.0 ;
      RECT  111300.0 285750.0 110100.0 282150.0 ;
      RECT  106500.0 284550.0 105300.0 282600.0 ;
      RECT  106500.0 296400.0 105300.0 294450.0 ;
      RECT  116100.0 285750.0 114900.0 284550.0 ;
      RECT  113700.0 285750.0 112500.0 284550.0 ;
      RECT  113700.0 285750.0 112500.0 284550.0 ;
      RECT  116100.0 285750.0 114900.0 284550.0 ;
      RECT  113700.0 285750.0 112500.0 284550.0 ;
      RECT  111300.0 285750.0 110100.0 284550.0 ;
      RECT  111300.0 285750.0 110100.0 284550.0 ;
      RECT  113700.0 285750.0 112500.0 284550.0 ;
      RECT  111300.0 285750.0 110100.0 284550.0 ;
      RECT  108900.0 285750.0 107700.0 284550.0 ;
      RECT  108900.0 285750.0 107700.0 284550.0 ;
      RECT  111300.0 285750.0 110100.0 284550.0 ;
      RECT  116100.0 294450.0 114900.0 293250.0 ;
      RECT  113700.0 294450.0 112500.0 293250.0 ;
      RECT  113700.0 294450.0 112500.0 293250.0 ;
      RECT  116100.0 294450.0 114900.0 293250.0 ;
      RECT  113700.0 294450.0 112500.0 293250.0 ;
      RECT  111300.0 294450.0 110100.0 293250.0 ;
      RECT  111300.0 294450.0 110100.0 293250.0 ;
      RECT  113700.0 294450.0 112500.0 293250.0 ;
      RECT  111300.0 294450.0 110100.0 293250.0 ;
      RECT  108900.0 294450.0 107700.0 293250.0 ;
      RECT  108900.0 294450.0 107700.0 293250.0 ;
      RECT  111300.0 294450.0 110100.0 293250.0 ;
      RECT  106500.0 285150.0 105300.0 283950.0 ;
      RECT  106500.0 295050.0 105300.0 293850.0 ;
      RECT  108900.0 292350.0 110100.0 291150.0 ;
      RECT  111300.0 290400.0 112500.0 289200.0 ;
      RECT  113700.0 288450.0 114900.0 287250.0 ;
      RECT  113700.0 285750.0 112500.0 284550.0 ;
      RECT  108900.0 285750.0 107700.0 284550.0 ;
      RECT  108900.0 294450.0 107700.0 293250.0 ;
      RECT  108900.0 288450.0 107700.0 287250.0 ;
      RECT  114900.0 288450.0 113700.0 287250.0 ;
      RECT  112500.0 290400.0 111300.0 289200.0 ;
      RECT  110100.0 292350.0 108900.0 291150.0 ;
      RECT  108900.0 288450.0 107700.0 287250.0 ;
      RECT  117900.0 283050.0 102300.0 282150.0 ;
      RECT  117900.0 296850.0 102300.0 295950.0 ;
      RECT  116100.0 298350.0 114900.0 295950.0 ;
      RECT  116100.0 307050.0 114900.0 310650.0 ;
      RECT  111300.0 307050.0 110100.0 310650.0 ;
      RECT  106500.0 308250.0 105300.0 310200.0 ;
      RECT  106500.0 296400.0 105300.0 298350.0 ;
      RECT  116100.0 307050.0 114900.0 308250.0 ;
      RECT  113700.0 307050.0 112500.0 308250.0 ;
      RECT  113700.0 307050.0 112500.0 308250.0 ;
      RECT  116100.0 307050.0 114900.0 308250.0 ;
      RECT  113700.0 307050.0 112500.0 308250.0 ;
      RECT  111300.0 307050.0 110100.0 308250.0 ;
      RECT  111300.0 307050.0 110100.0 308250.0 ;
      RECT  113700.0 307050.0 112500.0 308250.0 ;
      RECT  111300.0 307050.0 110100.0 308250.0 ;
      RECT  108900.0 307050.0 107700.0 308250.0 ;
      RECT  108900.0 307050.0 107700.0 308250.0 ;
      RECT  111300.0 307050.0 110100.0 308250.0 ;
      RECT  116100.0 298350.0 114900.0 299550.0 ;
      RECT  113700.0 298350.0 112500.0 299550.0 ;
      RECT  113700.0 298350.0 112500.0 299550.0 ;
      RECT  116100.0 298350.0 114900.0 299550.0 ;
      RECT  113700.0 298350.0 112500.0 299550.0 ;
      RECT  111300.0 298350.0 110100.0 299550.0 ;
      RECT  111300.0 298350.0 110100.0 299550.0 ;
      RECT  113700.0 298350.0 112500.0 299550.0 ;
      RECT  111300.0 298350.0 110100.0 299550.0 ;
      RECT  108900.0 298350.0 107700.0 299550.0 ;
      RECT  108900.0 298350.0 107700.0 299550.0 ;
      RECT  111300.0 298350.0 110100.0 299550.0 ;
      RECT  106500.0 307650.0 105300.0 308850.0 ;
      RECT  106500.0 297750.0 105300.0 298950.0 ;
      RECT  108900.0 300450.0 110100.0 301650.0 ;
      RECT  111300.0 302400.0 112500.0 303600.0 ;
      RECT  113700.0 304350.0 114900.0 305550.0 ;
      RECT  113700.0 307050.0 112500.0 308250.0 ;
      RECT  108900.0 307050.0 107700.0 308250.0 ;
      RECT  108900.0 298350.0 107700.0 299550.0 ;
      RECT  108900.0 304350.0 107700.0 305550.0 ;
      RECT  114900.0 304350.0 113700.0 305550.0 ;
      RECT  112500.0 302400.0 111300.0 303600.0 ;
      RECT  110100.0 300450.0 108900.0 301650.0 ;
      RECT  108900.0 304350.0 107700.0 305550.0 ;
      RECT  117900.0 309750.0 102300.0 310650.0 ;
      RECT  117900.0 295950.0 102300.0 296850.0 ;
      RECT  116100.0 322050.0 114900.0 324450.0 ;
      RECT  116100.0 313350.0 114900.0 309750.0 ;
      RECT  111300.0 313350.0 110100.0 309750.0 ;
      RECT  106500.0 312150.0 105300.0 310200.0 ;
      RECT  106500.0 324000.0 105300.0 322050.0 ;
      RECT  116100.0 313350.0 114900.0 312150.0 ;
      RECT  113700.0 313350.0 112500.0 312150.0 ;
      RECT  113700.0 313350.0 112500.0 312150.0 ;
      RECT  116100.0 313350.0 114900.0 312150.0 ;
      RECT  113700.0 313350.0 112500.0 312150.0 ;
      RECT  111300.0 313350.0 110100.0 312150.0 ;
      RECT  111300.0 313350.0 110100.0 312150.0 ;
      RECT  113700.0 313350.0 112500.0 312150.0 ;
      RECT  111300.0 313350.0 110100.0 312150.0 ;
      RECT  108900.0 313350.0 107700.0 312150.0 ;
      RECT  108900.0 313350.0 107700.0 312150.0 ;
      RECT  111300.0 313350.0 110100.0 312150.0 ;
      RECT  116100.0 322050.0 114900.0 320850.0 ;
      RECT  113700.0 322050.0 112500.0 320850.0 ;
      RECT  113700.0 322050.0 112500.0 320850.0 ;
      RECT  116100.0 322050.0 114900.0 320850.0 ;
      RECT  113700.0 322050.0 112500.0 320850.0 ;
      RECT  111300.0 322050.0 110100.0 320850.0 ;
      RECT  111300.0 322050.0 110100.0 320850.0 ;
      RECT  113700.0 322050.0 112500.0 320850.0 ;
      RECT  111300.0 322050.0 110100.0 320850.0 ;
      RECT  108900.0 322050.0 107700.0 320850.0 ;
      RECT  108900.0 322050.0 107700.0 320850.0 ;
      RECT  111300.0 322050.0 110100.0 320850.0 ;
      RECT  106500.0 312750.0 105300.0 311550.0 ;
      RECT  106500.0 322650.0 105300.0 321450.0 ;
      RECT  108900.0 319950.0 110100.0 318750.0 ;
      RECT  111300.0 318000.0 112500.0 316800.0 ;
      RECT  113700.0 316050.0 114900.0 314850.0 ;
      RECT  113700.0 313350.0 112500.0 312150.0 ;
      RECT  108900.0 313350.0 107700.0 312150.0 ;
      RECT  108900.0 322050.0 107700.0 320850.0 ;
      RECT  108900.0 316050.0 107700.0 314850.0 ;
      RECT  114900.0 316050.0 113700.0 314850.0 ;
      RECT  112500.0 318000.0 111300.0 316800.0 ;
      RECT  110100.0 319950.0 108900.0 318750.0 ;
      RECT  108900.0 316050.0 107700.0 314850.0 ;
      RECT  117900.0 310650.0 102300.0 309750.0 ;
      RECT  117900.0 324450.0 102300.0 323550.0 ;
      RECT  116100.0 325950.0 114900.0 323550.0 ;
      RECT  116100.0 334650.0 114900.0 338250.0 ;
      RECT  111300.0 334650.0 110100.0 338250.0 ;
      RECT  106500.0 335850.0 105300.0 337800.0 ;
      RECT  106500.0 324000.0 105300.0 325950.0 ;
      RECT  116100.0 334650.0 114900.0 335850.0 ;
      RECT  113700.0 334650.0 112500.0 335850.0 ;
      RECT  113700.0 334650.0 112500.0 335850.0 ;
      RECT  116100.0 334650.0 114900.0 335850.0 ;
      RECT  113700.0 334650.0 112500.0 335850.0 ;
      RECT  111300.0 334650.0 110100.0 335850.0 ;
      RECT  111300.0 334650.0 110100.0 335850.0 ;
      RECT  113700.0 334650.0 112500.0 335850.0 ;
      RECT  111300.0 334650.0 110100.0 335850.0 ;
      RECT  108900.0 334650.0 107700.0 335850.0 ;
      RECT  108900.0 334650.0 107700.0 335850.0 ;
      RECT  111300.0 334650.0 110100.0 335850.0 ;
      RECT  116100.0 325950.0 114900.0 327150.0 ;
      RECT  113700.0 325950.0 112500.0 327150.0 ;
      RECT  113700.0 325950.0 112500.0 327150.0 ;
      RECT  116100.0 325950.0 114900.0 327150.0 ;
      RECT  113700.0 325950.0 112500.0 327150.0 ;
      RECT  111300.0 325950.0 110100.0 327150.0 ;
      RECT  111300.0 325950.0 110100.0 327150.0 ;
      RECT  113700.0 325950.0 112500.0 327150.0 ;
      RECT  111300.0 325950.0 110100.0 327150.0 ;
      RECT  108900.0 325950.0 107700.0 327150.0 ;
      RECT  108900.0 325950.0 107700.0 327150.0 ;
      RECT  111300.0 325950.0 110100.0 327150.0 ;
      RECT  106500.0 335250.0 105300.0 336450.0 ;
      RECT  106500.0 325350.0 105300.0 326550.0 ;
      RECT  108900.0 328050.0 110100.0 329250.0 ;
      RECT  111300.0 330000.0 112500.0 331200.0 ;
      RECT  113700.0 331950.0 114900.0 333150.0 ;
      RECT  113700.0 334650.0 112500.0 335850.0 ;
      RECT  108900.0 334650.0 107700.0 335850.0 ;
      RECT  108900.0 325950.0 107700.0 327150.0 ;
      RECT  108900.0 331950.0 107700.0 333150.0 ;
      RECT  114900.0 331950.0 113700.0 333150.0 ;
      RECT  112500.0 330000.0 111300.0 331200.0 ;
      RECT  110100.0 328050.0 108900.0 329250.0 ;
      RECT  108900.0 331950.0 107700.0 333150.0 ;
      RECT  117900.0 337350.0 102300.0 338250.0 ;
      RECT  117900.0 323550.0 102300.0 324450.0 ;
      RECT  116100.0 349650.0 114900.0 352050.0 ;
      RECT  116100.0 340950.0 114900.0 337350.0 ;
      RECT  111300.0 340950.0 110100.0 337350.0 ;
      RECT  106500.0 339750.0 105300.0 337800.0 ;
      RECT  106500.0 351600.0 105300.0 349650.0 ;
      RECT  116100.0 340950.0 114900.0 339750.0 ;
      RECT  113700.0 340950.0 112500.0 339750.0 ;
      RECT  113700.0 340950.0 112500.0 339750.0 ;
      RECT  116100.0 340950.0 114900.0 339750.0 ;
      RECT  113700.0 340950.0 112500.0 339750.0 ;
      RECT  111300.0 340950.0 110100.0 339750.0 ;
      RECT  111300.0 340950.0 110100.0 339750.0 ;
      RECT  113700.0 340950.0 112500.0 339750.0 ;
      RECT  111300.0 340950.0 110100.0 339750.0 ;
      RECT  108900.0 340950.0 107700.0 339750.0 ;
      RECT  108900.0 340950.0 107700.0 339750.0 ;
      RECT  111300.0 340950.0 110100.0 339750.0 ;
      RECT  116100.0 349650.0 114900.0 348450.0 ;
      RECT  113700.0 349650.0 112500.0 348450.0 ;
      RECT  113700.0 349650.0 112500.0 348450.0 ;
      RECT  116100.0 349650.0 114900.0 348450.0 ;
      RECT  113700.0 349650.0 112500.0 348450.0 ;
      RECT  111300.0 349650.0 110100.0 348450.0 ;
      RECT  111300.0 349650.0 110100.0 348450.0 ;
      RECT  113700.0 349650.0 112500.0 348450.0 ;
      RECT  111300.0 349650.0 110100.0 348450.0 ;
      RECT  108900.0 349650.0 107700.0 348450.0 ;
      RECT  108900.0 349650.0 107700.0 348450.0 ;
      RECT  111300.0 349650.0 110100.0 348450.0 ;
      RECT  106500.0 340350.0 105300.0 339150.0 ;
      RECT  106500.0 350250.0 105300.0 349050.0 ;
      RECT  108900.0 347550.0 110100.0 346350.0 ;
      RECT  111300.0 345600.0 112500.0 344400.0 ;
      RECT  113700.0 343650.0 114900.0 342450.0 ;
      RECT  113700.0 340950.0 112500.0 339750.0 ;
      RECT  108900.0 340950.0 107700.0 339750.0 ;
      RECT  108900.0 349650.0 107700.0 348450.0 ;
      RECT  108900.0 343650.0 107700.0 342450.0 ;
      RECT  114900.0 343650.0 113700.0 342450.0 ;
      RECT  112500.0 345600.0 111300.0 344400.0 ;
      RECT  110100.0 347550.0 108900.0 346350.0 ;
      RECT  108900.0 343650.0 107700.0 342450.0 ;
      RECT  117900.0 338250.0 102300.0 337350.0 ;
      RECT  117900.0 352050.0 102300.0 351150.0 ;
      RECT  116100.0 353550.0 114900.0 351150.0 ;
      RECT  116100.0 362250.0 114900.0 365850.0 ;
      RECT  111300.0 362250.0 110100.0 365850.0 ;
      RECT  106500.0 363450.0 105300.0 365400.0 ;
      RECT  106500.0 351600.0 105300.0 353550.0 ;
      RECT  116100.0 362250.0 114900.0 363450.0 ;
      RECT  113700.0 362250.0 112500.0 363450.0 ;
      RECT  113700.0 362250.0 112500.0 363450.0 ;
      RECT  116100.0 362250.0 114900.0 363450.0 ;
      RECT  113700.0 362250.0 112500.0 363450.0 ;
      RECT  111300.0 362250.0 110100.0 363450.0 ;
      RECT  111300.0 362250.0 110100.0 363450.0 ;
      RECT  113700.0 362250.0 112500.0 363450.0 ;
      RECT  111300.0 362250.0 110100.0 363450.0 ;
      RECT  108900.0 362250.0 107700.0 363450.0 ;
      RECT  108900.0 362250.0 107700.0 363450.0 ;
      RECT  111300.0 362250.0 110100.0 363450.0 ;
      RECT  116100.0 353550.0 114900.0 354750.0 ;
      RECT  113700.0 353550.0 112500.0 354750.0 ;
      RECT  113700.0 353550.0 112500.0 354750.0 ;
      RECT  116100.0 353550.0 114900.0 354750.0 ;
      RECT  113700.0 353550.0 112500.0 354750.0 ;
      RECT  111300.0 353550.0 110100.0 354750.0 ;
      RECT  111300.0 353550.0 110100.0 354750.0 ;
      RECT  113700.0 353550.0 112500.0 354750.0 ;
      RECT  111300.0 353550.0 110100.0 354750.0 ;
      RECT  108900.0 353550.0 107700.0 354750.0 ;
      RECT  108900.0 353550.0 107700.0 354750.0 ;
      RECT  111300.0 353550.0 110100.0 354750.0 ;
      RECT  106500.0 362850.0 105300.0 364050.0 ;
      RECT  106500.0 352950.0 105300.0 354150.0 ;
      RECT  108900.0 355650.0 110100.0 356850.0 ;
      RECT  111300.0 357600.0 112500.0 358800.0 ;
      RECT  113700.0 359550.0 114900.0 360750.0 ;
      RECT  113700.0 362250.0 112500.0 363450.0 ;
      RECT  108900.0 362250.0 107700.0 363450.0 ;
      RECT  108900.0 353550.0 107700.0 354750.0 ;
      RECT  108900.0 359550.0 107700.0 360750.0 ;
      RECT  114900.0 359550.0 113700.0 360750.0 ;
      RECT  112500.0 357600.0 111300.0 358800.0 ;
      RECT  110100.0 355650.0 108900.0 356850.0 ;
      RECT  108900.0 359550.0 107700.0 360750.0 ;
      RECT  117900.0 364950.0 102300.0 365850.0 ;
      RECT  117900.0 351150.0 102300.0 352050.0 ;
      RECT  116100.0 377250.0 114900.0 379650.0 ;
      RECT  116100.0 368550.0 114900.0 364950.0 ;
      RECT  111300.0 368550.0 110100.0 364950.0 ;
      RECT  106500.0 367350.0 105300.0 365400.0 ;
      RECT  106500.0 379200.0 105300.0 377250.0 ;
      RECT  116100.0 368550.0 114900.0 367350.0 ;
      RECT  113700.0 368550.0 112500.0 367350.0 ;
      RECT  113700.0 368550.0 112500.0 367350.0 ;
      RECT  116100.0 368550.0 114900.0 367350.0 ;
      RECT  113700.0 368550.0 112500.0 367350.0 ;
      RECT  111300.0 368550.0 110100.0 367350.0 ;
      RECT  111300.0 368550.0 110100.0 367350.0 ;
      RECT  113700.0 368550.0 112500.0 367350.0 ;
      RECT  111300.0 368550.0 110100.0 367350.0 ;
      RECT  108900.0 368550.0 107700.0 367350.0 ;
      RECT  108900.0 368550.0 107700.0 367350.0 ;
      RECT  111300.0 368550.0 110100.0 367350.0 ;
      RECT  116100.0 377250.0 114900.0 376050.0 ;
      RECT  113700.0 377250.0 112500.0 376050.0 ;
      RECT  113700.0 377250.0 112500.0 376050.0 ;
      RECT  116100.0 377250.0 114900.0 376050.0 ;
      RECT  113700.0 377250.0 112500.0 376050.0 ;
      RECT  111300.0 377250.0 110100.0 376050.0 ;
      RECT  111300.0 377250.0 110100.0 376050.0 ;
      RECT  113700.0 377250.0 112500.0 376050.0 ;
      RECT  111300.0 377250.0 110100.0 376050.0 ;
      RECT  108900.0 377250.0 107700.0 376050.0 ;
      RECT  108900.0 377250.0 107700.0 376050.0 ;
      RECT  111300.0 377250.0 110100.0 376050.0 ;
      RECT  106500.0 367950.0 105300.0 366750.0 ;
      RECT  106500.0 377850.0 105300.0 376650.0 ;
      RECT  108900.0 375150.0 110100.0 373950.0 ;
      RECT  111300.0 373200.0 112500.0 372000.0 ;
      RECT  113700.0 371250.0 114900.0 370050.0 ;
      RECT  113700.0 368550.0 112500.0 367350.0 ;
      RECT  108900.0 368550.0 107700.0 367350.0 ;
      RECT  108900.0 377250.0 107700.0 376050.0 ;
      RECT  108900.0 371250.0 107700.0 370050.0 ;
      RECT  114900.0 371250.0 113700.0 370050.0 ;
      RECT  112500.0 373200.0 111300.0 372000.0 ;
      RECT  110100.0 375150.0 108900.0 373950.0 ;
      RECT  108900.0 371250.0 107700.0 370050.0 ;
      RECT  117900.0 365850.0 102300.0 364950.0 ;
      RECT  117900.0 379650.0 102300.0 378750.0 ;
      RECT  134850.0 279300.0 136050.0 280500.0 ;
      RECT  156450.0 274800.0 157650.0 276000.0 ;
      RECT  131850.0 293100.0 133050.0 294300.0 ;
      RECT  153450.0 289200.0 154650.0 290400.0 ;
      RECT  128850.0 306900.0 130050.0 308100.0 ;
      RECT  150450.0 302400.0 151650.0 303600.0 ;
      RECT  156450.0 311700.0 157650.0 312900.0 ;
      RECT  125850.0 311700.0 127050.0 312900.0 ;
      RECT  153450.0 325500.0 154650.0 326700.0 ;
      RECT  122850.0 325500.0 124050.0 326700.0 ;
      RECT  150450.0 339300.0 151650.0 340500.0 ;
      RECT  119850.0 339300.0 121050.0 340500.0 ;
      RECT  134850.0 276750.0 136050.0 277950.0 ;
      RECT  131850.0 274800.0 133050.0 276000.0 ;
      RECT  128850.0 272850.0 130050.0 274050.0 ;
      RECT  125850.0 287250.0 127050.0 288450.0 ;
      RECT  131850.0 289200.0 133050.0 290400.0 ;
      RECT  128850.0 291150.0 130050.0 292350.0 ;
      RECT  134850.0 304350.0 136050.0 305550.0 ;
      RECT  122850.0 302400.0 124050.0 303600.0 ;
      RECT  128850.0 300450.0 130050.0 301650.0 ;
      RECT  125850.0 314850.0 127050.0 316050.0 ;
      RECT  122850.0 316800.0 124050.0 318000.0 ;
      RECT  128850.0 318750.0 130050.0 319950.0 ;
      RECT  134850.0 331950.0 136050.0 333150.0 ;
      RECT  131850.0 330000.0 133050.0 331200.0 ;
      RECT  119850.0 328050.0 121050.0 329250.0 ;
      RECT  125850.0 342450.0 127050.0 343650.0 ;
      RECT  131850.0 344400.0 133050.0 345600.0 ;
      RECT  119850.0 346350.0 121050.0 347550.0 ;
      RECT  134850.0 359550.0 136050.0 360750.0 ;
      RECT  122850.0 357600.0 124050.0 358800.0 ;
      RECT  119850.0 355650.0 121050.0 356850.0 ;
      RECT  125850.0 370050.0 127050.0 371250.0 ;
      RECT  122850.0 372000.0 124050.0 373200.0 ;
      RECT  119850.0 373950.0 121050.0 375150.0 ;
      RECT  96450.0 274950.0 92700.0 275850.0 ;
      RECT  96450.0 289350.0 92700.0 290250.0 ;
      RECT  96450.0 302550.0 92700.0 303450.0 ;
      RECT  96450.0 316950.0 92700.0 317850.0 ;
      RECT  96450.0 330150.0 92700.0 331050.0 ;
      RECT  96450.0 344550.0 92700.0 345450.0 ;
      RECT  96450.0 357750.0 92700.0 358650.0 ;
      RECT  96450.0 372150.0 92700.0 373050.0 ;
      RECT  157500.0 282150.0 92700.0 283050.0 ;
      RECT  157500.0 309750.0 92700.0 310650.0 ;
      RECT  157500.0 337350.0 92700.0 338250.0 ;
      RECT  157500.0 364950.0 92700.0 365850.0 ;
      RECT  157500.0 268350.0 92700.0 269250.0 ;
      RECT  157500.0 295950.0 92700.0 296850.0 ;
      RECT  157500.0 323550.0 92700.0 324450.0 ;
      RECT  157500.0 351150.0 92700.0 352050.0 ;
      RECT  157500.0 378750.0 92700.0 379650.0 ;
      RECT  94500.0 381150.0 95700.0 378750.0 ;
      RECT  94500.0 389850.0 95700.0 393450.0 ;
      RECT  99300.0 389850.0 100500.0 393450.0 ;
      RECT  104100.0 391050.0 105300.0 393000.0 ;
      RECT  104100.0 379200.0 105300.0 381150.0 ;
      RECT  94500.0 389850.0 95700.0 391050.0 ;
      RECT  96900.0 389850.0 98100.0 391050.0 ;
      RECT  96900.0 389850.0 98100.0 391050.0 ;
      RECT  94500.0 389850.0 95700.0 391050.0 ;
      RECT  96900.0 389850.0 98100.0 391050.0 ;
      RECT  99300.0 389850.0 100500.0 391050.0 ;
      RECT  99300.0 389850.0 100500.0 391050.0 ;
      RECT  96900.0 389850.0 98100.0 391050.0 ;
      RECT  99300.0 389850.0 100500.0 391050.0 ;
      RECT  101700.0 389850.0 102900.0 391050.0 ;
      RECT  101700.0 389850.0 102900.0 391050.0 ;
      RECT  99300.0 389850.0 100500.0 391050.0 ;
      RECT  94500.0 381150.0 95700.0 382350.0 ;
      RECT  96900.0 381150.0 98100.0 382350.0 ;
      RECT  96900.0 381150.0 98100.0 382350.0 ;
      RECT  94500.0 381150.0 95700.0 382350.0 ;
      RECT  96900.0 381150.0 98100.0 382350.0 ;
      RECT  99300.0 381150.0 100500.0 382350.0 ;
      RECT  99300.0 381150.0 100500.0 382350.0 ;
      RECT  96900.0 381150.0 98100.0 382350.0 ;
      RECT  99300.0 381150.0 100500.0 382350.0 ;
      RECT  101700.0 381150.0 102900.0 382350.0 ;
      RECT  101700.0 381150.0 102900.0 382350.0 ;
      RECT  99300.0 381150.0 100500.0 382350.0 ;
      RECT  104100.0 390450.0 105300.0 391650.0 ;
      RECT  104100.0 380550.0 105300.0 381750.0 ;
      RECT  101700.0 383250.0 100500.0 384450.0 ;
      RECT  99300.0 385200.0 98100.0 386400.0 ;
      RECT  96900.0 387150.0 95700.0 388350.0 ;
      RECT  96900.0 389850.0 98100.0 391050.0 ;
      RECT  101700.0 389850.0 102900.0 391050.0 ;
      RECT  101700.0 381150.0 102900.0 382350.0 ;
      RECT  101700.0 387150.0 102900.0 388350.0 ;
      RECT  95700.0 387150.0 96900.0 388350.0 ;
      RECT  98100.0 385200.0 99300.0 386400.0 ;
      RECT  100500.0 383250.0 101700.0 384450.0 ;
      RECT  101700.0 387150.0 102900.0 388350.0 ;
      RECT  92700.0 392550.0 108300.0 393450.0 ;
      RECT  92700.0 378750.0 108300.0 379650.0 ;
      RECT  94500.0 404850.0 95700.0 407250.0 ;
      RECT  94500.0 396150.0 95700.0 392550.0 ;
      RECT  99300.0 396150.0 100500.0 392550.0 ;
      RECT  104100.0 394950.0 105300.0 393000.0 ;
      RECT  104100.0 406800.0 105300.0 404850.0 ;
      RECT  94500.0 396150.0 95700.0 394950.0 ;
      RECT  96900.0 396150.0 98100.0 394950.0 ;
      RECT  96900.0 396150.0 98100.0 394950.0 ;
      RECT  94500.0 396150.0 95700.0 394950.0 ;
      RECT  96900.0 396150.0 98100.0 394950.0 ;
      RECT  99300.0 396150.0 100500.0 394950.0 ;
      RECT  99300.0 396150.0 100500.0 394950.0 ;
      RECT  96900.0 396150.0 98100.0 394950.0 ;
      RECT  99300.0 396150.0 100500.0 394950.0 ;
      RECT  101700.0 396150.0 102900.0 394950.0 ;
      RECT  101700.0 396150.0 102900.0 394950.0 ;
      RECT  99300.0 396150.0 100500.0 394950.0 ;
      RECT  94500.0 404850.0 95700.0 403650.0 ;
      RECT  96900.0 404850.0 98100.0 403650.0 ;
      RECT  96900.0 404850.0 98100.0 403650.0 ;
      RECT  94500.0 404850.0 95700.0 403650.0 ;
      RECT  96900.0 404850.0 98100.0 403650.0 ;
      RECT  99300.0 404850.0 100500.0 403650.0 ;
      RECT  99300.0 404850.0 100500.0 403650.0 ;
      RECT  96900.0 404850.0 98100.0 403650.0 ;
      RECT  99300.0 404850.0 100500.0 403650.0 ;
      RECT  101700.0 404850.0 102900.0 403650.0 ;
      RECT  101700.0 404850.0 102900.0 403650.0 ;
      RECT  99300.0 404850.0 100500.0 403650.0 ;
      RECT  104100.0 395550.0 105300.0 394350.0 ;
      RECT  104100.0 405450.0 105300.0 404250.0 ;
      RECT  101700.0 402750.0 100500.0 401550.0 ;
      RECT  99300.0 400800.0 98100.0 399600.0 ;
      RECT  96900.0 398850.0 95700.0 397650.0 ;
      RECT  96900.0 396150.0 98100.0 394950.0 ;
      RECT  101700.0 396150.0 102900.0 394950.0 ;
      RECT  101700.0 404850.0 102900.0 403650.0 ;
      RECT  101700.0 398850.0 102900.0 397650.0 ;
      RECT  95700.0 398850.0 96900.0 397650.0 ;
      RECT  98100.0 400800.0 99300.0 399600.0 ;
      RECT  100500.0 402750.0 101700.0 401550.0 ;
      RECT  101700.0 398850.0 102900.0 397650.0 ;
      RECT  92700.0 393450.0 108300.0 392550.0 ;
      RECT  92700.0 407250.0 108300.0 406350.0 ;
      RECT  94500.0 408750.0 95700.0 406350.0 ;
      RECT  94500.0 417450.0 95700.0 421050.0 ;
      RECT  99300.0 417450.0 100500.0 421050.0 ;
      RECT  104100.0 418650.0 105300.0 420600.0 ;
      RECT  104100.0 406800.0 105300.0 408750.0 ;
      RECT  94500.0 417450.0 95700.0 418650.0 ;
      RECT  96900.0 417450.0 98100.0 418650.0 ;
      RECT  96900.0 417450.0 98100.0 418650.0 ;
      RECT  94500.0 417450.0 95700.0 418650.0 ;
      RECT  96900.0 417450.0 98100.0 418650.0 ;
      RECT  99300.0 417450.0 100500.0 418650.0 ;
      RECT  99300.0 417450.0 100500.0 418650.0 ;
      RECT  96900.0 417450.0 98100.0 418650.0 ;
      RECT  99300.0 417450.0 100500.0 418650.0 ;
      RECT  101700.0 417450.0 102900.0 418650.0 ;
      RECT  101700.0 417450.0 102900.0 418650.0 ;
      RECT  99300.0 417450.0 100500.0 418650.0 ;
      RECT  94500.0 408750.0 95700.0 409950.0 ;
      RECT  96900.0 408750.0 98100.0 409950.0 ;
      RECT  96900.0 408750.0 98100.0 409950.0 ;
      RECT  94500.0 408750.0 95700.0 409950.0 ;
      RECT  96900.0 408750.0 98100.0 409950.0 ;
      RECT  99300.0 408750.0 100500.0 409950.0 ;
      RECT  99300.0 408750.0 100500.0 409950.0 ;
      RECT  96900.0 408750.0 98100.0 409950.0 ;
      RECT  99300.0 408750.0 100500.0 409950.0 ;
      RECT  101700.0 408750.0 102900.0 409950.0 ;
      RECT  101700.0 408750.0 102900.0 409950.0 ;
      RECT  99300.0 408750.0 100500.0 409950.0 ;
      RECT  104100.0 418050.0 105300.0 419250.0 ;
      RECT  104100.0 408150.0 105300.0 409350.0 ;
      RECT  101700.0 410850.0 100500.0 412050.0 ;
      RECT  99300.0 412800.0 98100.0 414000.0 ;
      RECT  96900.0 414750.0 95700.0 415950.0 ;
      RECT  96900.0 417450.0 98100.0 418650.0 ;
      RECT  101700.0 417450.0 102900.0 418650.0 ;
      RECT  101700.0 408750.0 102900.0 409950.0 ;
      RECT  101700.0 414750.0 102900.0 415950.0 ;
      RECT  95700.0 414750.0 96900.0 415950.0 ;
      RECT  98100.0 412800.0 99300.0 414000.0 ;
      RECT  100500.0 410850.0 101700.0 412050.0 ;
      RECT  101700.0 414750.0 102900.0 415950.0 ;
      RECT  92700.0 420150.0 108300.0 421050.0 ;
      RECT  92700.0 406350.0 108300.0 407250.0 ;
      RECT  94500.0 432450.0 95700.0 434850.0 ;
      RECT  94500.0 423750.0 95700.0 420150.0 ;
      RECT  99300.0 423750.0 100500.0 420150.0 ;
      RECT  104100.0 422550.0 105300.0 420600.0 ;
      RECT  104100.0 434400.0 105300.0 432450.0 ;
      RECT  94500.0 423750.0 95700.0 422550.0 ;
      RECT  96900.0 423750.0 98100.0 422550.0 ;
      RECT  96900.0 423750.0 98100.0 422550.0 ;
      RECT  94500.0 423750.0 95700.0 422550.0 ;
      RECT  96900.0 423750.0 98100.0 422550.0 ;
      RECT  99300.0 423750.0 100500.0 422550.0 ;
      RECT  99300.0 423750.0 100500.0 422550.0 ;
      RECT  96900.0 423750.0 98100.0 422550.0 ;
      RECT  99300.0 423750.0 100500.0 422550.0 ;
      RECT  101700.0 423750.0 102900.0 422550.0 ;
      RECT  101700.0 423750.0 102900.0 422550.0 ;
      RECT  99300.0 423750.0 100500.0 422550.0 ;
      RECT  94500.0 432450.0 95700.0 431250.0 ;
      RECT  96900.0 432450.0 98100.0 431250.0 ;
      RECT  96900.0 432450.0 98100.0 431250.0 ;
      RECT  94500.0 432450.0 95700.0 431250.0 ;
      RECT  96900.0 432450.0 98100.0 431250.0 ;
      RECT  99300.0 432450.0 100500.0 431250.0 ;
      RECT  99300.0 432450.0 100500.0 431250.0 ;
      RECT  96900.0 432450.0 98100.0 431250.0 ;
      RECT  99300.0 432450.0 100500.0 431250.0 ;
      RECT  101700.0 432450.0 102900.0 431250.0 ;
      RECT  101700.0 432450.0 102900.0 431250.0 ;
      RECT  99300.0 432450.0 100500.0 431250.0 ;
      RECT  104100.0 423150.0 105300.0 421950.0 ;
      RECT  104100.0 433050.0 105300.0 431850.0 ;
      RECT  101700.0 430350.0 100500.0 429150.0 ;
      RECT  99300.0 428400.0 98100.0 427200.0 ;
      RECT  96900.0 426450.0 95700.0 425250.0 ;
      RECT  96900.0 423750.0 98100.0 422550.0 ;
      RECT  101700.0 423750.0 102900.0 422550.0 ;
      RECT  101700.0 432450.0 102900.0 431250.0 ;
      RECT  101700.0 426450.0 102900.0 425250.0 ;
      RECT  95700.0 426450.0 96900.0 425250.0 ;
      RECT  98100.0 428400.0 99300.0 427200.0 ;
      RECT  100500.0 430350.0 101700.0 429150.0 ;
      RECT  101700.0 426450.0 102900.0 425250.0 ;
      RECT  92700.0 421050.0 108300.0 420150.0 ;
      RECT  92700.0 434850.0 108300.0 433950.0 ;
      RECT  94500.0 436350.0 95700.0 433950.0 ;
      RECT  94500.0 445050.0 95700.0 448650.0 ;
      RECT  99300.0 445050.0 100500.0 448650.0 ;
      RECT  104100.0 446250.0 105300.0 448200.0 ;
      RECT  104100.0 434400.0 105300.0 436350.0 ;
      RECT  94500.0 445050.0 95700.0 446250.0 ;
      RECT  96900.0 445050.0 98100.0 446250.0 ;
      RECT  96900.0 445050.0 98100.0 446250.0 ;
      RECT  94500.0 445050.0 95700.0 446250.0 ;
      RECT  96900.0 445050.0 98100.0 446250.0 ;
      RECT  99300.0 445050.0 100500.0 446250.0 ;
      RECT  99300.0 445050.0 100500.0 446250.0 ;
      RECT  96900.0 445050.0 98100.0 446250.0 ;
      RECT  99300.0 445050.0 100500.0 446250.0 ;
      RECT  101700.0 445050.0 102900.0 446250.0 ;
      RECT  101700.0 445050.0 102900.0 446250.0 ;
      RECT  99300.0 445050.0 100500.0 446250.0 ;
      RECT  94500.0 436350.0 95700.0 437550.0 ;
      RECT  96900.0 436350.0 98100.0 437550.0 ;
      RECT  96900.0 436350.0 98100.0 437550.0 ;
      RECT  94500.0 436350.0 95700.0 437550.0 ;
      RECT  96900.0 436350.0 98100.0 437550.0 ;
      RECT  99300.0 436350.0 100500.0 437550.0 ;
      RECT  99300.0 436350.0 100500.0 437550.0 ;
      RECT  96900.0 436350.0 98100.0 437550.0 ;
      RECT  99300.0 436350.0 100500.0 437550.0 ;
      RECT  101700.0 436350.0 102900.0 437550.0 ;
      RECT  101700.0 436350.0 102900.0 437550.0 ;
      RECT  99300.0 436350.0 100500.0 437550.0 ;
      RECT  104100.0 445650.0 105300.0 446850.0 ;
      RECT  104100.0 435750.0 105300.0 436950.0 ;
      RECT  101700.0 438450.0 100500.0 439650.0 ;
      RECT  99300.0 440400.0 98100.0 441600.0 ;
      RECT  96900.0 442350.0 95700.0 443550.0 ;
      RECT  96900.0 445050.0 98100.0 446250.0 ;
      RECT  101700.0 445050.0 102900.0 446250.0 ;
      RECT  101700.0 436350.0 102900.0 437550.0 ;
      RECT  101700.0 442350.0 102900.0 443550.0 ;
      RECT  95700.0 442350.0 96900.0 443550.0 ;
      RECT  98100.0 440400.0 99300.0 441600.0 ;
      RECT  100500.0 438450.0 101700.0 439650.0 ;
      RECT  101700.0 442350.0 102900.0 443550.0 ;
      RECT  92700.0 447750.0 108300.0 448650.0 ;
      RECT  92700.0 433950.0 108300.0 434850.0 ;
      RECT  94500.0 460050.0 95700.0 462450.0 ;
      RECT  94500.0 451350.0 95700.0 447750.0 ;
      RECT  99300.0 451350.0 100500.0 447750.0 ;
      RECT  104100.0 450150.0 105300.0 448200.0 ;
      RECT  104100.0 462000.0 105300.0 460050.0 ;
      RECT  94500.0 451350.0 95700.0 450150.0 ;
      RECT  96900.0 451350.0 98100.0 450150.0 ;
      RECT  96900.0 451350.0 98100.0 450150.0 ;
      RECT  94500.0 451350.0 95700.0 450150.0 ;
      RECT  96900.0 451350.0 98100.0 450150.0 ;
      RECT  99300.0 451350.0 100500.0 450150.0 ;
      RECT  99300.0 451350.0 100500.0 450150.0 ;
      RECT  96900.0 451350.0 98100.0 450150.0 ;
      RECT  99300.0 451350.0 100500.0 450150.0 ;
      RECT  101700.0 451350.0 102900.0 450150.0 ;
      RECT  101700.0 451350.0 102900.0 450150.0 ;
      RECT  99300.0 451350.0 100500.0 450150.0 ;
      RECT  94500.0 460050.0 95700.0 458850.0 ;
      RECT  96900.0 460050.0 98100.0 458850.0 ;
      RECT  96900.0 460050.0 98100.0 458850.0 ;
      RECT  94500.0 460050.0 95700.0 458850.0 ;
      RECT  96900.0 460050.0 98100.0 458850.0 ;
      RECT  99300.0 460050.0 100500.0 458850.0 ;
      RECT  99300.0 460050.0 100500.0 458850.0 ;
      RECT  96900.0 460050.0 98100.0 458850.0 ;
      RECT  99300.0 460050.0 100500.0 458850.0 ;
      RECT  101700.0 460050.0 102900.0 458850.0 ;
      RECT  101700.0 460050.0 102900.0 458850.0 ;
      RECT  99300.0 460050.0 100500.0 458850.0 ;
      RECT  104100.0 450750.0 105300.0 449550.0 ;
      RECT  104100.0 460650.0 105300.0 459450.0 ;
      RECT  101700.0 457950.0 100500.0 456750.0 ;
      RECT  99300.0 456000.0 98100.0 454800.0 ;
      RECT  96900.0 454050.0 95700.0 452850.0 ;
      RECT  96900.0 451350.0 98100.0 450150.0 ;
      RECT  101700.0 451350.0 102900.0 450150.0 ;
      RECT  101700.0 460050.0 102900.0 458850.0 ;
      RECT  101700.0 454050.0 102900.0 452850.0 ;
      RECT  95700.0 454050.0 96900.0 452850.0 ;
      RECT  98100.0 456000.0 99300.0 454800.0 ;
      RECT  100500.0 457950.0 101700.0 456750.0 ;
      RECT  101700.0 454050.0 102900.0 452850.0 ;
      RECT  92700.0 448650.0 108300.0 447750.0 ;
      RECT  92700.0 462450.0 108300.0 461550.0 ;
      RECT  94500.0 463950.0 95700.0 461550.0 ;
      RECT  94500.0 472650.0 95700.0 476250.0 ;
      RECT  99300.0 472650.0 100500.0 476250.0 ;
      RECT  104100.0 473850.0 105300.0 475800.0 ;
      RECT  104100.0 462000.0 105300.0 463950.0 ;
      RECT  94500.0 472650.0 95700.0 473850.0 ;
      RECT  96900.0 472650.0 98100.0 473850.0 ;
      RECT  96900.0 472650.0 98100.0 473850.0 ;
      RECT  94500.0 472650.0 95700.0 473850.0 ;
      RECT  96900.0 472650.0 98100.0 473850.0 ;
      RECT  99300.0 472650.0 100500.0 473850.0 ;
      RECT  99300.0 472650.0 100500.0 473850.0 ;
      RECT  96900.0 472650.0 98100.0 473850.0 ;
      RECT  99300.0 472650.0 100500.0 473850.0 ;
      RECT  101700.0 472650.0 102900.0 473850.0 ;
      RECT  101700.0 472650.0 102900.0 473850.0 ;
      RECT  99300.0 472650.0 100500.0 473850.0 ;
      RECT  94500.0 463950.0 95700.0 465150.0 ;
      RECT  96900.0 463950.0 98100.0 465150.0 ;
      RECT  96900.0 463950.0 98100.0 465150.0 ;
      RECT  94500.0 463950.0 95700.0 465150.0 ;
      RECT  96900.0 463950.0 98100.0 465150.0 ;
      RECT  99300.0 463950.0 100500.0 465150.0 ;
      RECT  99300.0 463950.0 100500.0 465150.0 ;
      RECT  96900.0 463950.0 98100.0 465150.0 ;
      RECT  99300.0 463950.0 100500.0 465150.0 ;
      RECT  101700.0 463950.0 102900.0 465150.0 ;
      RECT  101700.0 463950.0 102900.0 465150.0 ;
      RECT  99300.0 463950.0 100500.0 465150.0 ;
      RECT  104100.0 473250.0 105300.0 474450.0 ;
      RECT  104100.0 463350.0 105300.0 464550.0 ;
      RECT  101700.0 466050.0 100500.0 467250.0 ;
      RECT  99300.0 468000.0 98100.0 469200.0 ;
      RECT  96900.0 469950.0 95700.0 471150.0 ;
      RECT  96900.0 472650.0 98100.0 473850.0 ;
      RECT  101700.0 472650.0 102900.0 473850.0 ;
      RECT  101700.0 463950.0 102900.0 465150.0 ;
      RECT  101700.0 469950.0 102900.0 471150.0 ;
      RECT  95700.0 469950.0 96900.0 471150.0 ;
      RECT  98100.0 468000.0 99300.0 469200.0 ;
      RECT  100500.0 466050.0 101700.0 467250.0 ;
      RECT  101700.0 469950.0 102900.0 471150.0 ;
      RECT  92700.0 475350.0 108300.0 476250.0 ;
      RECT  92700.0 461550.0 108300.0 462450.0 ;
      RECT  94500.0 487650.0 95700.0 490050.0 ;
      RECT  94500.0 478950.0 95700.0 475350.0 ;
      RECT  99300.0 478950.0 100500.0 475350.0 ;
      RECT  104100.0 477750.0 105300.0 475800.0 ;
      RECT  104100.0 489600.0 105300.0 487650.0 ;
      RECT  94500.0 478950.0 95700.0 477750.0 ;
      RECT  96900.0 478950.0 98100.0 477750.0 ;
      RECT  96900.0 478950.0 98100.0 477750.0 ;
      RECT  94500.0 478950.0 95700.0 477750.0 ;
      RECT  96900.0 478950.0 98100.0 477750.0 ;
      RECT  99300.0 478950.0 100500.0 477750.0 ;
      RECT  99300.0 478950.0 100500.0 477750.0 ;
      RECT  96900.0 478950.0 98100.0 477750.0 ;
      RECT  99300.0 478950.0 100500.0 477750.0 ;
      RECT  101700.0 478950.0 102900.0 477750.0 ;
      RECT  101700.0 478950.0 102900.0 477750.0 ;
      RECT  99300.0 478950.0 100500.0 477750.0 ;
      RECT  94500.0 487650.0 95700.0 486450.0 ;
      RECT  96900.0 487650.0 98100.0 486450.0 ;
      RECT  96900.0 487650.0 98100.0 486450.0 ;
      RECT  94500.0 487650.0 95700.0 486450.0 ;
      RECT  96900.0 487650.0 98100.0 486450.0 ;
      RECT  99300.0 487650.0 100500.0 486450.0 ;
      RECT  99300.0 487650.0 100500.0 486450.0 ;
      RECT  96900.0 487650.0 98100.0 486450.0 ;
      RECT  99300.0 487650.0 100500.0 486450.0 ;
      RECT  101700.0 487650.0 102900.0 486450.0 ;
      RECT  101700.0 487650.0 102900.0 486450.0 ;
      RECT  99300.0 487650.0 100500.0 486450.0 ;
      RECT  104100.0 478350.0 105300.0 477150.0 ;
      RECT  104100.0 488250.0 105300.0 487050.0 ;
      RECT  101700.0 485550.0 100500.0 484350.0 ;
      RECT  99300.0 483600.0 98100.0 482400.0 ;
      RECT  96900.0 481650.0 95700.0 480450.0 ;
      RECT  96900.0 478950.0 98100.0 477750.0 ;
      RECT  101700.0 478950.0 102900.0 477750.0 ;
      RECT  101700.0 487650.0 102900.0 486450.0 ;
      RECT  101700.0 481650.0 102900.0 480450.0 ;
      RECT  95700.0 481650.0 96900.0 480450.0 ;
      RECT  98100.0 483600.0 99300.0 482400.0 ;
      RECT  100500.0 485550.0 101700.0 484350.0 ;
      RECT  101700.0 481650.0 102900.0 480450.0 ;
      RECT  92700.0 476250.0 108300.0 475350.0 ;
      RECT  92700.0 490050.0 108300.0 489150.0 ;
      RECT  94500.0 491550.0 95700.0 489150.0 ;
      RECT  94500.0 500250.0 95700.0 503850.0 ;
      RECT  99300.0 500250.0 100500.0 503850.0 ;
      RECT  104100.0 501450.0 105300.0 503400.0 ;
      RECT  104100.0 489600.0 105300.0 491550.0 ;
      RECT  94500.0 500250.0 95700.0 501450.0 ;
      RECT  96900.0 500250.0 98100.0 501450.0 ;
      RECT  96900.0 500250.0 98100.0 501450.0 ;
      RECT  94500.0 500250.0 95700.0 501450.0 ;
      RECT  96900.0 500250.0 98100.0 501450.0 ;
      RECT  99300.0 500250.0 100500.0 501450.0 ;
      RECT  99300.0 500250.0 100500.0 501450.0 ;
      RECT  96900.0 500250.0 98100.0 501450.0 ;
      RECT  99300.0 500250.0 100500.0 501450.0 ;
      RECT  101700.0 500250.0 102900.0 501450.0 ;
      RECT  101700.0 500250.0 102900.0 501450.0 ;
      RECT  99300.0 500250.0 100500.0 501450.0 ;
      RECT  94500.0 491550.0 95700.0 492750.0 ;
      RECT  96900.0 491550.0 98100.0 492750.0 ;
      RECT  96900.0 491550.0 98100.0 492750.0 ;
      RECT  94500.0 491550.0 95700.0 492750.0 ;
      RECT  96900.0 491550.0 98100.0 492750.0 ;
      RECT  99300.0 491550.0 100500.0 492750.0 ;
      RECT  99300.0 491550.0 100500.0 492750.0 ;
      RECT  96900.0 491550.0 98100.0 492750.0 ;
      RECT  99300.0 491550.0 100500.0 492750.0 ;
      RECT  101700.0 491550.0 102900.0 492750.0 ;
      RECT  101700.0 491550.0 102900.0 492750.0 ;
      RECT  99300.0 491550.0 100500.0 492750.0 ;
      RECT  104100.0 500850.0 105300.0 502050.0 ;
      RECT  104100.0 490950.0 105300.0 492150.0 ;
      RECT  101700.0 493650.0 100500.0 494850.0 ;
      RECT  99300.0 495600.0 98100.0 496800.0 ;
      RECT  96900.0 497550.0 95700.0 498750.0 ;
      RECT  96900.0 500250.0 98100.0 501450.0 ;
      RECT  101700.0 500250.0 102900.0 501450.0 ;
      RECT  101700.0 491550.0 102900.0 492750.0 ;
      RECT  101700.0 497550.0 102900.0 498750.0 ;
      RECT  95700.0 497550.0 96900.0 498750.0 ;
      RECT  98100.0 495600.0 99300.0 496800.0 ;
      RECT  100500.0 493650.0 101700.0 494850.0 ;
      RECT  101700.0 497550.0 102900.0 498750.0 ;
      RECT  92700.0 502950.0 108300.0 503850.0 ;
      RECT  92700.0 489150.0 108300.0 490050.0 ;
      RECT  94500.0 515250.0 95700.0 517650.0 ;
      RECT  94500.0 506550.0 95700.0 502950.0 ;
      RECT  99300.0 506550.0 100500.0 502950.0 ;
      RECT  104100.0 505350.0 105300.0 503400.0 ;
      RECT  104100.0 517200.0 105300.0 515250.0 ;
      RECT  94500.0 506550.0 95700.0 505350.0 ;
      RECT  96900.0 506550.0 98100.0 505350.0 ;
      RECT  96900.0 506550.0 98100.0 505350.0 ;
      RECT  94500.0 506550.0 95700.0 505350.0 ;
      RECT  96900.0 506550.0 98100.0 505350.0 ;
      RECT  99300.0 506550.0 100500.0 505350.0 ;
      RECT  99300.0 506550.0 100500.0 505350.0 ;
      RECT  96900.0 506550.0 98100.0 505350.0 ;
      RECT  99300.0 506550.0 100500.0 505350.0 ;
      RECT  101700.0 506550.0 102900.0 505350.0 ;
      RECT  101700.0 506550.0 102900.0 505350.0 ;
      RECT  99300.0 506550.0 100500.0 505350.0 ;
      RECT  94500.0 515250.0 95700.0 514050.0 ;
      RECT  96900.0 515250.0 98100.0 514050.0 ;
      RECT  96900.0 515250.0 98100.0 514050.0 ;
      RECT  94500.0 515250.0 95700.0 514050.0 ;
      RECT  96900.0 515250.0 98100.0 514050.0 ;
      RECT  99300.0 515250.0 100500.0 514050.0 ;
      RECT  99300.0 515250.0 100500.0 514050.0 ;
      RECT  96900.0 515250.0 98100.0 514050.0 ;
      RECT  99300.0 515250.0 100500.0 514050.0 ;
      RECT  101700.0 515250.0 102900.0 514050.0 ;
      RECT  101700.0 515250.0 102900.0 514050.0 ;
      RECT  99300.0 515250.0 100500.0 514050.0 ;
      RECT  104100.0 505950.0 105300.0 504750.0 ;
      RECT  104100.0 515850.0 105300.0 514650.0 ;
      RECT  101700.0 513150.0 100500.0 511950.0 ;
      RECT  99300.0 511200.0 98100.0 510000.0 ;
      RECT  96900.0 509250.0 95700.0 508050.0 ;
      RECT  96900.0 506550.0 98100.0 505350.0 ;
      RECT  101700.0 506550.0 102900.0 505350.0 ;
      RECT  101700.0 515250.0 102900.0 514050.0 ;
      RECT  101700.0 509250.0 102900.0 508050.0 ;
      RECT  95700.0 509250.0 96900.0 508050.0 ;
      RECT  98100.0 511200.0 99300.0 510000.0 ;
      RECT  100500.0 513150.0 101700.0 511950.0 ;
      RECT  101700.0 509250.0 102900.0 508050.0 ;
      RECT  92700.0 503850.0 108300.0 502950.0 ;
      RECT  92700.0 517650.0 108300.0 516750.0 ;
      RECT  94500.0 519150.0 95700.0 516750.0 ;
      RECT  94500.0 527850.0 95700.0 531450.0 ;
      RECT  99300.0 527850.0 100500.0 531450.0 ;
      RECT  104100.0 529050.0 105300.0 531000.0 ;
      RECT  104100.0 517200.0 105300.0 519150.0 ;
      RECT  94500.0 527850.0 95700.0 529050.0 ;
      RECT  96900.0 527850.0 98100.0 529050.0 ;
      RECT  96900.0 527850.0 98100.0 529050.0 ;
      RECT  94500.0 527850.0 95700.0 529050.0 ;
      RECT  96900.0 527850.0 98100.0 529050.0 ;
      RECT  99300.0 527850.0 100500.0 529050.0 ;
      RECT  99300.0 527850.0 100500.0 529050.0 ;
      RECT  96900.0 527850.0 98100.0 529050.0 ;
      RECT  99300.0 527850.0 100500.0 529050.0 ;
      RECT  101700.0 527850.0 102900.0 529050.0 ;
      RECT  101700.0 527850.0 102900.0 529050.0 ;
      RECT  99300.0 527850.0 100500.0 529050.0 ;
      RECT  94500.0 519150.0 95700.0 520350.0 ;
      RECT  96900.0 519150.0 98100.0 520350.0 ;
      RECT  96900.0 519150.0 98100.0 520350.0 ;
      RECT  94500.0 519150.0 95700.0 520350.0 ;
      RECT  96900.0 519150.0 98100.0 520350.0 ;
      RECT  99300.0 519150.0 100500.0 520350.0 ;
      RECT  99300.0 519150.0 100500.0 520350.0 ;
      RECT  96900.0 519150.0 98100.0 520350.0 ;
      RECT  99300.0 519150.0 100500.0 520350.0 ;
      RECT  101700.0 519150.0 102900.0 520350.0 ;
      RECT  101700.0 519150.0 102900.0 520350.0 ;
      RECT  99300.0 519150.0 100500.0 520350.0 ;
      RECT  104100.0 528450.0 105300.0 529650.0 ;
      RECT  104100.0 518550.0 105300.0 519750.0 ;
      RECT  101700.0 521250.0 100500.0 522450.0 ;
      RECT  99300.0 523200.0 98100.0 524400.0 ;
      RECT  96900.0 525150.0 95700.0 526350.0 ;
      RECT  96900.0 527850.0 98100.0 529050.0 ;
      RECT  101700.0 527850.0 102900.0 529050.0 ;
      RECT  101700.0 519150.0 102900.0 520350.0 ;
      RECT  101700.0 525150.0 102900.0 526350.0 ;
      RECT  95700.0 525150.0 96900.0 526350.0 ;
      RECT  98100.0 523200.0 99300.0 524400.0 ;
      RECT  100500.0 521250.0 101700.0 522450.0 ;
      RECT  101700.0 525150.0 102900.0 526350.0 ;
      RECT  92700.0 530550.0 108300.0 531450.0 ;
      RECT  92700.0 516750.0 108300.0 517650.0 ;
      RECT  94500.0 542850.0 95700.0 545250.0 ;
      RECT  94500.0 534150.0 95700.0 530550.0 ;
      RECT  99300.0 534150.0 100500.0 530550.0 ;
      RECT  104100.0 532950.0 105300.0 531000.0 ;
      RECT  104100.0 544800.0 105300.0 542850.0 ;
      RECT  94500.0 534150.0 95700.0 532950.0 ;
      RECT  96900.0 534150.0 98100.0 532950.0 ;
      RECT  96900.0 534150.0 98100.0 532950.0 ;
      RECT  94500.0 534150.0 95700.0 532950.0 ;
      RECT  96900.0 534150.0 98100.0 532950.0 ;
      RECT  99300.0 534150.0 100500.0 532950.0 ;
      RECT  99300.0 534150.0 100500.0 532950.0 ;
      RECT  96900.0 534150.0 98100.0 532950.0 ;
      RECT  99300.0 534150.0 100500.0 532950.0 ;
      RECT  101700.0 534150.0 102900.0 532950.0 ;
      RECT  101700.0 534150.0 102900.0 532950.0 ;
      RECT  99300.0 534150.0 100500.0 532950.0 ;
      RECT  94500.0 542850.0 95700.0 541650.0 ;
      RECT  96900.0 542850.0 98100.0 541650.0 ;
      RECT  96900.0 542850.0 98100.0 541650.0 ;
      RECT  94500.0 542850.0 95700.0 541650.0 ;
      RECT  96900.0 542850.0 98100.0 541650.0 ;
      RECT  99300.0 542850.0 100500.0 541650.0 ;
      RECT  99300.0 542850.0 100500.0 541650.0 ;
      RECT  96900.0 542850.0 98100.0 541650.0 ;
      RECT  99300.0 542850.0 100500.0 541650.0 ;
      RECT  101700.0 542850.0 102900.0 541650.0 ;
      RECT  101700.0 542850.0 102900.0 541650.0 ;
      RECT  99300.0 542850.0 100500.0 541650.0 ;
      RECT  104100.0 533550.0 105300.0 532350.0 ;
      RECT  104100.0 543450.0 105300.0 542250.0 ;
      RECT  101700.0 540750.0 100500.0 539550.0 ;
      RECT  99300.0 538800.0 98100.0 537600.0 ;
      RECT  96900.0 536850.0 95700.0 535650.0 ;
      RECT  96900.0 534150.0 98100.0 532950.0 ;
      RECT  101700.0 534150.0 102900.0 532950.0 ;
      RECT  101700.0 542850.0 102900.0 541650.0 ;
      RECT  101700.0 536850.0 102900.0 535650.0 ;
      RECT  95700.0 536850.0 96900.0 535650.0 ;
      RECT  98100.0 538800.0 99300.0 537600.0 ;
      RECT  100500.0 540750.0 101700.0 539550.0 ;
      RECT  101700.0 536850.0 102900.0 535650.0 ;
      RECT  92700.0 531450.0 108300.0 530550.0 ;
      RECT  92700.0 545250.0 108300.0 544350.0 ;
      RECT  94500.0 546750.0 95700.0 544350.0 ;
      RECT  94500.0 555450.0 95700.0 559050.0 ;
      RECT  99300.0 555450.0 100500.0 559050.0 ;
      RECT  104100.0 556650.0 105300.0 558600.0 ;
      RECT  104100.0 544800.0 105300.0 546750.0 ;
      RECT  94500.0 555450.0 95700.0 556650.0 ;
      RECT  96900.0 555450.0 98100.0 556650.0 ;
      RECT  96900.0 555450.0 98100.0 556650.0 ;
      RECT  94500.0 555450.0 95700.0 556650.0 ;
      RECT  96900.0 555450.0 98100.0 556650.0 ;
      RECT  99300.0 555450.0 100500.0 556650.0 ;
      RECT  99300.0 555450.0 100500.0 556650.0 ;
      RECT  96900.0 555450.0 98100.0 556650.0 ;
      RECT  99300.0 555450.0 100500.0 556650.0 ;
      RECT  101700.0 555450.0 102900.0 556650.0 ;
      RECT  101700.0 555450.0 102900.0 556650.0 ;
      RECT  99300.0 555450.0 100500.0 556650.0 ;
      RECT  94500.0 546750.0 95700.0 547950.0 ;
      RECT  96900.0 546750.0 98100.0 547950.0 ;
      RECT  96900.0 546750.0 98100.0 547950.0 ;
      RECT  94500.0 546750.0 95700.0 547950.0 ;
      RECT  96900.0 546750.0 98100.0 547950.0 ;
      RECT  99300.0 546750.0 100500.0 547950.0 ;
      RECT  99300.0 546750.0 100500.0 547950.0 ;
      RECT  96900.0 546750.0 98100.0 547950.0 ;
      RECT  99300.0 546750.0 100500.0 547950.0 ;
      RECT  101700.0 546750.0 102900.0 547950.0 ;
      RECT  101700.0 546750.0 102900.0 547950.0 ;
      RECT  99300.0 546750.0 100500.0 547950.0 ;
      RECT  104100.0 556050.0 105300.0 557250.0 ;
      RECT  104100.0 546150.0 105300.0 547350.0 ;
      RECT  101700.0 548850.0 100500.0 550050.0 ;
      RECT  99300.0 550800.0 98100.0 552000.0 ;
      RECT  96900.0 552750.0 95700.0 553950.0 ;
      RECT  96900.0 555450.0 98100.0 556650.0 ;
      RECT  101700.0 555450.0 102900.0 556650.0 ;
      RECT  101700.0 546750.0 102900.0 547950.0 ;
      RECT  101700.0 552750.0 102900.0 553950.0 ;
      RECT  95700.0 552750.0 96900.0 553950.0 ;
      RECT  98100.0 550800.0 99300.0 552000.0 ;
      RECT  100500.0 548850.0 101700.0 550050.0 ;
      RECT  101700.0 552750.0 102900.0 553950.0 ;
      RECT  92700.0 558150.0 108300.0 559050.0 ;
      RECT  92700.0 544350.0 108300.0 545250.0 ;
      RECT  94500.0 570450.0 95700.0 572850.0 ;
      RECT  94500.0 561750.0 95700.0 558150.0 ;
      RECT  99300.0 561750.0 100500.0 558150.0 ;
      RECT  104100.0 560550.0 105300.0 558600.0 ;
      RECT  104100.0 572400.0 105300.0 570450.0 ;
      RECT  94500.0 561750.0 95700.0 560550.0 ;
      RECT  96900.0 561750.0 98100.0 560550.0 ;
      RECT  96900.0 561750.0 98100.0 560550.0 ;
      RECT  94500.0 561750.0 95700.0 560550.0 ;
      RECT  96900.0 561750.0 98100.0 560550.0 ;
      RECT  99300.0 561750.0 100500.0 560550.0 ;
      RECT  99300.0 561750.0 100500.0 560550.0 ;
      RECT  96900.0 561750.0 98100.0 560550.0 ;
      RECT  99300.0 561750.0 100500.0 560550.0 ;
      RECT  101700.0 561750.0 102900.0 560550.0 ;
      RECT  101700.0 561750.0 102900.0 560550.0 ;
      RECT  99300.0 561750.0 100500.0 560550.0 ;
      RECT  94500.0 570450.0 95700.0 569250.0 ;
      RECT  96900.0 570450.0 98100.0 569250.0 ;
      RECT  96900.0 570450.0 98100.0 569250.0 ;
      RECT  94500.0 570450.0 95700.0 569250.0 ;
      RECT  96900.0 570450.0 98100.0 569250.0 ;
      RECT  99300.0 570450.0 100500.0 569250.0 ;
      RECT  99300.0 570450.0 100500.0 569250.0 ;
      RECT  96900.0 570450.0 98100.0 569250.0 ;
      RECT  99300.0 570450.0 100500.0 569250.0 ;
      RECT  101700.0 570450.0 102900.0 569250.0 ;
      RECT  101700.0 570450.0 102900.0 569250.0 ;
      RECT  99300.0 570450.0 100500.0 569250.0 ;
      RECT  104100.0 561150.0 105300.0 559950.0 ;
      RECT  104100.0 571050.0 105300.0 569850.0 ;
      RECT  101700.0 568350.0 100500.0 567150.0 ;
      RECT  99300.0 566400.0 98100.0 565200.0 ;
      RECT  96900.0 564450.0 95700.0 563250.0 ;
      RECT  96900.0 561750.0 98100.0 560550.0 ;
      RECT  101700.0 561750.0 102900.0 560550.0 ;
      RECT  101700.0 570450.0 102900.0 569250.0 ;
      RECT  101700.0 564450.0 102900.0 563250.0 ;
      RECT  95700.0 564450.0 96900.0 563250.0 ;
      RECT  98100.0 566400.0 99300.0 565200.0 ;
      RECT  100500.0 568350.0 101700.0 567150.0 ;
      RECT  101700.0 564450.0 102900.0 563250.0 ;
      RECT  92700.0 559050.0 108300.0 558150.0 ;
      RECT  92700.0 572850.0 108300.0 571950.0 ;
      RECT  94500.0 574350.0 95700.0 571950.0 ;
      RECT  94500.0 583050.0 95700.0 586650.0 ;
      RECT  99300.0 583050.0 100500.0 586650.0 ;
      RECT  104100.0 584250.0 105300.0 586200.0 ;
      RECT  104100.0 572400.0 105300.0 574350.0 ;
      RECT  94500.0 583050.0 95700.0 584250.0 ;
      RECT  96900.0 583050.0 98100.0 584250.0 ;
      RECT  96900.0 583050.0 98100.0 584250.0 ;
      RECT  94500.0 583050.0 95700.0 584250.0 ;
      RECT  96900.0 583050.0 98100.0 584250.0 ;
      RECT  99300.0 583050.0 100500.0 584250.0 ;
      RECT  99300.0 583050.0 100500.0 584250.0 ;
      RECT  96900.0 583050.0 98100.0 584250.0 ;
      RECT  99300.0 583050.0 100500.0 584250.0 ;
      RECT  101700.0 583050.0 102900.0 584250.0 ;
      RECT  101700.0 583050.0 102900.0 584250.0 ;
      RECT  99300.0 583050.0 100500.0 584250.0 ;
      RECT  94500.0 574350.0 95700.0 575550.0 ;
      RECT  96900.0 574350.0 98100.0 575550.0 ;
      RECT  96900.0 574350.0 98100.0 575550.0 ;
      RECT  94500.0 574350.0 95700.0 575550.0 ;
      RECT  96900.0 574350.0 98100.0 575550.0 ;
      RECT  99300.0 574350.0 100500.0 575550.0 ;
      RECT  99300.0 574350.0 100500.0 575550.0 ;
      RECT  96900.0 574350.0 98100.0 575550.0 ;
      RECT  99300.0 574350.0 100500.0 575550.0 ;
      RECT  101700.0 574350.0 102900.0 575550.0 ;
      RECT  101700.0 574350.0 102900.0 575550.0 ;
      RECT  99300.0 574350.0 100500.0 575550.0 ;
      RECT  104100.0 583650.0 105300.0 584850.0 ;
      RECT  104100.0 573750.0 105300.0 574950.0 ;
      RECT  101700.0 576450.0 100500.0 577650.0 ;
      RECT  99300.0 578400.0 98100.0 579600.0 ;
      RECT  96900.0 580350.0 95700.0 581550.0 ;
      RECT  96900.0 583050.0 98100.0 584250.0 ;
      RECT  101700.0 583050.0 102900.0 584250.0 ;
      RECT  101700.0 574350.0 102900.0 575550.0 ;
      RECT  101700.0 580350.0 102900.0 581550.0 ;
      RECT  95700.0 580350.0 96900.0 581550.0 ;
      RECT  98100.0 578400.0 99300.0 579600.0 ;
      RECT  100500.0 576450.0 101700.0 577650.0 ;
      RECT  101700.0 580350.0 102900.0 581550.0 ;
      RECT  92700.0 585750.0 108300.0 586650.0 ;
      RECT  92700.0 571950.0 108300.0 572850.0 ;
      RECT  94500.0 598050.0 95700.0 600450.0 ;
      RECT  94500.0 589350.0 95700.0 585750.0 ;
      RECT  99300.0 589350.0 100500.0 585750.0 ;
      RECT  104100.0 588150.0 105300.0 586200.0 ;
      RECT  104100.0 600000.0 105300.0 598050.0 ;
      RECT  94500.0 589350.0 95700.0 588150.0 ;
      RECT  96900.0 589350.0 98100.0 588150.0 ;
      RECT  96900.0 589350.0 98100.0 588150.0 ;
      RECT  94500.0 589350.0 95700.0 588150.0 ;
      RECT  96900.0 589350.0 98100.0 588150.0 ;
      RECT  99300.0 589350.0 100500.0 588150.0 ;
      RECT  99300.0 589350.0 100500.0 588150.0 ;
      RECT  96900.0 589350.0 98100.0 588150.0 ;
      RECT  99300.0 589350.0 100500.0 588150.0 ;
      RECT  101700.0 589350.0 102900.0 588150.0 ;
      RECT  101700.0 589350.0 102900.0 588150.0 ;
      RECT  99300.0 589350.0 100500.0 588150.0 ;
      RECT  94500.0 598050.0 95700.0 596850.0 ;
      RECT  96900.0 598050.0 98100.0 596850.0 ;
      RECT  96900.0 598050.0 98100.0 596850.0 ;
      RECT  94500.0 598050.0 95700.0 596850.0 ;
      RECT  96900.0 598050.0 98100.0 596850.0 ;
      RECT  99300.0 598050.0 100500.0 596850.0 ;
      RECT  99300.0 598050.0 100500.0 596850.0 ;
      RECT  96900.0 598050.0 98100.0 596850.0 ;
      RECT  99300.0 598050.0 100500.0 596850.0 ;
      RECT  101700.0 598050.0 102900.0 596850.0 ;
      RECT  101700.0 598050.0 102900.0 596850.0 ;
      RECT  99300.0 598050.0 100500.0 596850.0 ;
      RECT  104100.0 588750.0 105300.0 587550.0 ;
      RECT  104100.0 598650.0 105300.0 597450.0 ;
      RECT  101700.0 595950.0 100500.0 594750.0 ;
      RECT  99300.0 594000.0 98100.0 592800.0 ;
      RECT  96900.0 592050.0 95700.0 590850.0 ;
      RECT  96900.0 589350.0 98100.0 588150.0 ;
      RECT  101700.0 589350.0 102900.0 588150.0 ;
      RECT  101700.0 598050.0 102900.0 596850.0 ;
      RECT  101700.0 592050.0 102900.0 590850.0 ;
      RECT  95700.0 592050.0 96900.0 590850.0 ;
      RECT  98100.0 594000.0 99300.0 592800.0 ;
      RECT  100500.0 595950.0 101700.0 594750.0 ;
      RECT  101700.0 592050.0 102900.0 590850.0 ;
      RECT  92700.0 586650.0 108300.0 585750.0 ;
      RECT  92700.0 600450.0 108300.0 599550.0 ;
      RECT  94500.0 601950.0 95700.0 599550.0 ;
      RECT  94500.0 610650.0 95700.0 614250.0 ;
      RECT  99300.0 610650.0 100500.0 614250.0 ;
      RECT  104100.0 611850.0 105300.0 613800.0 ;
      RECT  104100.0 600000.0 105300.0 601950.0 ;
      RECT  94500.0 610650.0 95700.0 611850.0 ;
      RECT  96900.0 610650.0 98100.0 611850.0 ;
      RECT  96900.0 610650.0 98100.0 611850.0 ;
      RECT  94500.0 610650.0 95700.0 611850.0 ;
      RECT  96900.0 610650.0 98100.0 611850.0 ;
      RECT  99300.0 610650.0 100500.0 611850.0 ;
      RECT  99300.0 610650.0 100500.0 611850.0 ;
      RECT  96900.0 610650.0 98100.0 611850.0 ;
      RECT  99300.0 610650.0 100500.0 611850.0 ;
      RECT  101700.0 610650.0 102900.0 611850.0 ;
      RECT  101700.0 610650.0 102900.0 611850.0 ;
      RECT  99300.0 610650.0 100500.0 611850.0 ;
      RECT  94500.0 601950.0 95700.0 603150.0 ;
      RECT  96900.0 601950.0 98100.0 603150.0 ;
      RECT  96900.0 601950.0 98100.0 603150.0 ;
      RECT  94500.0 601950.0 95700.0 603150.0 ;
      RECT  96900.0 601950.0 98100.0 603150.0 ;
      RECT  99300.0 601950.0 100500.0 603150.0 ;
      RECT  99300.0 601950.0 100500.0 603150.0 ;
      RECT  96900.0 601950.0 98100.0 603150.0 ;
      RECT  99300.0 601950.0 100500.0 603150.0 ;
      RECT  101700.0 601950.0 102900.0 603150.0 ;
      RECT  101700.0 601950.0 102900.0 603150.0 ;
      RECT  99300.0 601950.0 100500.0 603150.0 ;
      RECT  104100.0 611250.0 105300.0 612450.0 ;
      RECT  104100.0 601350.0 105300.0 602550.0 ;
      RECT  101700.0 604050.0 100500.0 605250.0 ;
      RECT  99300.0 606000.0 98100.0 607200.0 ;
      RECT  96900.0 607950.0 95700.0 609150.0 ;
      RECT  96900.0 610650.0 98100.0 611850.0 ;
      RECT  101700.0 610650.0 102900.0 611850.0 ;
      RECT  101700.0 601950.0 102900.0 603150.0 ;
      RECT  101700.0 607950.0 102900.0 609150.0 ;
      RECT  95700.0 607950.0 96900.0 609150.0 ;
      RECT  98100.0 606000.0 99300.0 607200.0 ;
      RECT  100500.0 604050.0 101700.0 605250.0 ;
      RECT  101700.0 607950.0 102900.0 609150.0 ;
      RECT  92700.0 613350.0 108300.0 614250.0 ;
      RECT  92700.0 599550.0 108300.0 600450.0 ;
      RECT  94500.0 625650.0 95700.0 628050.0 ;
      RECT  94500.0 616950.0 95700.0 613350.0 ;
      RECT  99300.0 616950.0 100500.0 613350.0 ;
      RECT  104100.0 615750.0 105300.0 613800.0 ;
      RECT  104100.0 627600.0 105300.0 625650.0 ;
      RECT  94500.0 616950.0 95700.0 615750.0 ;
      RECT  96900.0 616950.0 98100.0 615750.0 ;
      RECT  96900.0 616950.0 98100.0 615750.0 ;
      RECT  94500.0 616950.0 95700.0 615750.0 ;
      RECT  96900.0 616950.0 98100.0 615750.0 ;
      RECT  99300.0 616950.0 100500.0 615750.0 ;
      RECT  99300.0 616950.0 100500.0 615750.0 ;
      RECT  96900.0 616950.0 98100.0 615750.0 ;
      RECT  99300.0 616950.0 100500.0 615750.0 ;
      RECT  101700.0 616950.0 102900.0 615750.0 ;
      RECT  101700.0 616950.0 102900.0 615750.0 ;
      RECT  99300.0 616950.0 100500.0 615750.0 ;
      RECT  94500.0 625650.0 95700.0 624450.0 ;
      RECT  96900.0 625650.0 98100.0 624450.0 ;
      RECT  96900.0 625650.0 98100.0 624450.0 ;
      RECT  94500.0 625650.0 95700.0 624450.0 ;
      RECT  96900.0 625650.0 98100.0 624450.0 ;
      RECT  99300.0 625650.0 100500.0 624450.0 ;
      RECT  99300.0 625650.0 100500.0 624450.0 ;
      RECT  96900.0 625650.0 98100.0 624450.0 ;
      RECT  99300.0 625650.0 100500.0 624450.0 ;
      RECT  101700.0 625650.0 102900.0 624450.0 ;
      RECT  101700.0 625650.0 102900.0 624450.0 ;
      RECT  99300.0 625650.0 100500.0 624450.0 ;
      RECT  104100.0 616350.0 105300.0 615150.0 ;
      RECT  104100.0 626250.0 105300.0 625050.0 ;
      RECT  101700.0 623550.0 100500.0 622350.0 ;
      RECT  99300.0 621600.0 98100.0 620400.0 ;
      RECT  96900.0 619650.0 95700.0 618450.0 ;
      RECT  96900.0 616950.0 98100.0 615750.0 ;
      RECT  101700.0 616950.0 102900.0 615750.0 ;
      RECT  101700.0 625650.0 102900.0 624450.0 ;
      RECT  101700.0 619650.0 102900.0 618450.0 ;
      RECT  95700.0 619650.0 96900.0 618450.0 ;
      RECT  98100.0 621600.0 99300.0 620400.0 ;
      RECT  100500.0 623550.0 101700.0 622350.0 ;
      RECT  101700.0 619650.0 102900.0 618450.0 ;
      RECT  92700.0 614250.0 108300.0 613350.0 ;
      RECT  92700.0 628050.0 108300.0 627150.0 ;
      RECT  94500.0 629550.0 95700.0 627150.0 ;
      RECT  94500.0 638250.0 95700.0 641850.0 ;
      RECT  99300.0 638250.0 100500.0 641850.0 ;
      RECT  104100.0 639450.0 105300.0 641400.0 ;
      RECT  104100.0 627600.0 105300.0 629550.0 ;
      RECT  94500.0 638250.0 95700.0 639450.0 ;
      RECT  96900.0 638250.0 98100.0 639450.0 ;
      RECT  96900.0 638250.0 98100.0 639450.0 ;
      RECT  94500.0 638250.0 95700.0 639450.0 ;
      RECT  96900.0 638250.0 98100.0 639450.0 ;
      RECT  99300.0 638250.0 100500.0 639450.0 ;
      RECT  99300.0 638250.0 100500.0 639450.0 ;
      RECT  96900.0 638250.0 98100.0 639450.0 ;
      RECT  99300.0 638250.0 100500.0 639450.0 ;
      RECT  101700.0 638250.0 102900.0 639450.0 ;
      RECT  101700.0 638250.0 102900.0 639450.0 ;
      RECT  99300.0 638250.0 100500.0 639450.0 ;
      RECT  94500.0 629550.0 95700.0 630750.0 ;
      RECT  96900.0 629550.0 98100.0 630750.0 ;
      RECT  96900.0 629550.0 98100.0 630750.0 ;
      RECT  94500.0 629550.0 95700.0 630750.0 ;
      RECT  96900.0 629550.0 98100.0 630750.0 ;
      RECT  99300.0 629550.0 100500.0 630750.0 ;
      RECT  99300.0 629550.0 100500.0 630750.0 ;
      RECT  96900.0 629550.0 98100.0 630750.0 ;
      RECT  99300.0 629550.0 100500.0 630750.0 ;
      RECT  101700.0 629550.0 102900.0 630750.0 ;
      RECT  101700.0 629550.0 102900.0 630750.0 ;
      RECT  99300.0 629550.0 100500.0 630750.0 ;
      RECT  104100.0 638850.0 105300.0 640050.0 ;
      RECT  104100.0 628950.0 105300.0 630150.0 ;
      RECT  101700.0 631650.0 100500.0 632850.0 ;
      RECT  99300.0 633600.0 98100.0 634800.0 ;
      RECT  96900.0 635550.0 95700.0 636750.0 ;
      RECT  96900.0 638250.0 98100.0 639450.0 ;
      RECT  101700.0 638250.0 102900.0 639450.0 ;
      RECT  101700.0 629550.0 102900.0 630750.0 ;
      RECT  101700.0 635550.0 102900.0 636750.0 ;
      RECT  95700.0 635550.0 96900.0 636750.0 ;
      RECT  98100.0 633600.0 99300.0 634800.0 ;
      RECT  100500.0 631650.0 101700.0 632850.0 ;
      RECT  101700.0 635550.0 102900.0 636750.0 ;
      RECT  92700.0 640950.0 108300.0 641850.0 ;
      RECT  92700.0 627150.0 108300.0 628050.0 ;
      RECT  94500.0 653250.0 95700.0 655650.0 ;
      RECT  94500.0 644550.0 95700.0 640950.0 ;
      RECT  99300.0 644550.0 100500.0 640950.0 ;
      RECT  104100.0 643350.0 105300.0 641400.0 ;
      RECT  104100.0 655200.0 105300.0 653250.0 ;
      RECT  94500.0 644550.0 95700.0 643350.0 ;
      RECT  96900.0 644550.0 98100.0 643350.0 ;
      RECT  96900.0 644550.0 98100.0 643350.0 ;
      RECT  94500.0 644550.0 95700.0 643350.0 ;
      RECT  96900.0 644550.0 98100.0 643350.0 ;
      RECT  99300.0 644550.0 100500.0 643350.0 ;
      RECT  99300.0 644550.0 100500.0 643350.0 ;
      RECT  96900.0 644550.0 98100.0 643350.0 ;
      RECT  99300.0 644550.0 100500.0 643350.0 ;
      RECT  101700.0 644550.0 102900.0 643350.0 ;
      RECT  101700.0 644550.0 102900.0 643350.0 ;
      RECT  99300.0 644550.0 100500.0 643350.0 ;
      RECT  94500.0 653250.0 95700.0 652050.0 ;
      RECT  96900.0 653250.0 98100.0 652050.0 ;
      RECT  96900.0 653250.0 98100.0 652050.0 ;
      RECT  94500.0 653250.0 95700.0 652050.0 ;
      RECT  96900.0 653250.0 98100.0 652050.0 ;
      RECT  99300.0 653250.0 100500.0 652050.0 ;
      RECT  99300.0 653250.0 100500.0 652050.0 ;
      RECT  96900.0 653250.0 98100.0 652050.0 ;
      RECT  99300.0 653250.0 100500.0 652050.0 ;
      RECT  101700.0 653250.0 102900.0 652050.0 ;
      RECT  101700.0 653250.0 102900.0 652050.0 ;
      RECT  99300.0 653250.0 100500.0 652050.0 ;
      RECT  104100.0 643950.0 105300.0 642750.0 ;
      RECT  104100.0 653850.0 105300.0 652650.0 ;
      RECT  101700.0 651150.0 100500.0 649950.0 ;
      RECT  99300.0 649200.0 98100.0 648000.0 ;
      RECT  96900.0 647250.0 95700.0 646050.0 ;
      RECT  96900.0 644550.0 98100.0 643350.0 ;
      RECT  101700.0 644550.0 102900.0 643350.0 ;
      RECT  101700.0 653250.0 102900.0 652050.0 ;
      RECT  101700.0 647250.0 102900.0 646050.0 ;
      RECT  95700.0 647250.0 96900.0 646050.0 ;
      RECT  98100.0 649200.0 99300.0 648000.0 ;
      RECT  100500.0 651150.0 101700.0 649950.0 ;
      RECT  101700.0 647250.0 102900.0 646050.0 ;
      RECT  92700.0 641850.0 108300.0 640950.0 ;
      RECT  92700.0 655650.0 108300.0 654750.0 ;
      RECT  94500.0 657150.0 95700.0 654750.0 ;
      RECT  94500.0 665850.0 95700.0 669450.0 ;
      RECT  99300.0 665850.0 100500.0 669450.0 ;
      RECT  104100.0 667050.0 105300.0 669000.0 ;
      RECT  104100.0 655200.0 105300.0 657150.0 ;
      RECT  94500.0 665850.0 95700.0 667050.0 ;
      RECT  96900.0 665850.0 98100.0 667050.0 ;
      RECT  96900.0 665850.0 98100.0 667050.0 ;
      RECT  94500.0 665850.0 95700.0 667050.0 ;
      RECT  96900.0 665850.0 98100.0 667050.0 ;
      RECT  99300.0 665850.0 100500.0 667050.0 ;
      RECT  99300.0 665850.0 100500.0 667050.0 ;
      RECT  96900.0 665850.0 98100.0 667050.0 ;
      RECT  99300.0 665850.0 100500.0 667050.0 ;
      RECT  101700.0 665850.0 102900.0 667050.0 ;
      RECT  101700.0 665850.0 102900.0 667050.0 ;
      RECT  99300.0 665850.0 100500.0 667050.0 ;
      RECT  94500.0 657150.0 95700.0 658350.0 ;
      RECT  96900.0 657150.0 98100.0 658350.0 ;
      RECT  96900.0 657150.0 98100.0 658350.0 ;
      RECT  94500.0 657150.0 95700.0 658350.0 ;
      RECT  96900.0 657150.0 98100.0 658350.0 ;
      RECT  99300.0 657150.0 100500.0 658350.0 ;
      RECT  99300.0 657150.0 100500.0 658350.0 ;
      RECT  96900.0 657150.0 98100.0 658350.0 ;
      RECT  99300.0 657150.0 100500.0 658350.0 ;
      RECT  101700.0 657150.0 102900.0 658350.0 ;
      RECT  101700.0 657150.0 102900.0 658350.0 ;
      RECT  99300.0 657150.0 100500.0 658350.0 ;
      RECT  104100.0 666450.0 105300.0 667650.0 ;
      RECT  104100.0 656550.0 105300.0 657750.0 ;
      RECT  101700.0 659250.0 100500.0 660450.0 ;
      RECT  99300.0 661200.0 98100.0 662400.0 ;
      RECT  96900.0 663150.0 95700.0 664350.0 ;
      RECT  96900.0 665850.0 98100.0 667050.0 ;
      RECT  101700.0 665850.0 102900.0 667050.0 ;
      RECT  101700.0 657150.0 102900.0 658350.0 ;
      RECT  101700.0 663150.0 102900.0 664350.0 ;
      RECT  95700.0 663150.0 96900.0 664350.0 ;
      RECT  98100.0 661200.0 99300.0 662400.0 ;
      RECT  100500.0 659250.0 101700.0 660450.0 ;
      RECT  101700.0 663150.0 102900.0 664350.0 ;
      RECT  92700.0 668550.0 108300.0 669450.0 ;
      RECT  92700.0 654750.0 108300.0 655650.0 ;
      RECT  94500.0 680850.0 95700.0 683250.0 ;
      RECT  94500.0 672150.0 95700.0 668550.0 ;
      RECT  99300.0 672150.0 100500.0 668550.0 ;
      RECT  104100.0 670950.0 105300.0 669000.0 ;
      RECT  104100.0 682800.0 105300.0 680850.0 ;
      RECT  94500.0 672150.0 95700.0 670950.0 ;
      RECT  96900.0 672150.0 98100.0 670950.0 ;
      RECT  96900.0 672150.0 98100.0 670950.0 ;
      RECT  94500.0 672150.0 95700.0 670950.0 ;
      RECT  96900.0 672150.0 98100.0 670950.0 ;
      RECT  99300.0 672150.0 100500.0 670950.0 ;
      RECT  99300.0 672150.0 100500.0 670950.0 ;
      RECT  96900.0 672150.0 98100.0 670950.0 ;
      RECT  99300.0 672150.0 100500.0 670950.0 ;
      RECT  101700.0 672150.0 102900.0 670950.0 ;
      RECT  101700.0 672150.0 102900.0 670950.0 ;
      RECT  99300.0 672150.0 100500.0 670950.0 ;
      RECT  94500.0 680850.0 95700.0 679650.0 ;
      RECT  96900.0 680850.0 98100.0 679650.0 ;
      RECT  96900.0 680850.0 98100.0 679650.0 ;
      RECT  94500.0 680850.0 95700.0 679650.0 ;
      RECT  96900.0 680850.0 98100.0 679650.0 ;
      RECT  99300.0 680850.0 100500.0 679650.0 ;
      RECT  99300.0 680850.0 100500.0 679650.0 ;
      RECT  96900.0 680850.0 98100.0 679650.0 ;
      RECT  99300.0 680850.0 100500.0 679650.0 ;
      RECT  101700.0 680850.0 102900.0 679650.0 ;
      RECT  101700.0 680850.0 102900.0 679650.0 ;
      RECT  99300.0 680850.0 100500.0 679650.0 ;
      RECT  104100.0 671550.0 105300.0 670350.0 ;
      RECT  104100.0 681450.0 105300.0 680250.0 ;
      RECT  101700.0 678750.0 100500.0 677550.0 ;
      RECT  99300.0 676800.0 98100.0 675600.0 ;
      RECT  96900.0 674850.0 95700.0 673650.0 ;
      RECT  96900.0 672150.0 98100.0 670950.0 ;
      RECT  101700.0 672150.0 102900.0 670950.0 ;
      RECT  101700.0 680850.0 102900.0 679650.0 ;
      RECT  101700.0 674850.0 102900.0 673650.0 ;
      RECT  95700.0 674850.0 96900.0 673650.0 ;
      RECT  98100.0 676800.0 99300.0 675600.0 ;
      RECT  100500.0 678750.0 101700.0 677550.0 ;
      RECT  101700.0 674850.0 102900.0 673650.0 ;
      RECT  92700.0 669450.0 108300.0 668550.0 ;
      RECT  92700.0 683250.0 108300.0 682350.0 ;
      RECT  94500.0 684750.0 95700.0 682350.0 ;
      RECT  94500.0 693450.0 95700.0 697050.0 ;
      RECT  99300.0 693450.0 100500.0 697050.0 ;
      RECT  104100.0 694650.0 105300.0 696600.0 ;
      RECT  104100.0 682800.0 105300.0 684750.0 ;
      RECT  94500.0 693450.0 95700.0 694650.0 ;
      RECT  96900.0 693450.0 98100.0 694650.0 ;
      RECT  96900.0 693450.0 98100.0 694650.0 ;
      RECT  94500.0 693450.0 95700.0 694650.0 ;
      RECT  96900.0 693450.0 98100.0 694650.0 ;
      RECT  99300.0 693450.0 100500.0 694650.0 ;
      RECT  99300.0 693450.0 100500.0 694650.0 ;
      RECT  96900.0 693450.0 98100.0 694650.0 ;
      RECT  99300.0 693450.0 100500.0 694650.0 ;
      RECT  101700.0 693450.0 102900.0 694650.0 ;
      RECT  101700.0 693450.0 102900.0 694650.0 ;
      RECT  99300.0 693450.0 100500.0 694650.0 ;
      RECT  94500.0 684750.0 95700.0 685950.0 ;
      RECT  96900.0 684750.0 98100.0 685950.0 ;
      RECT  96900.0 684750.0 98100.0 685950.0 ;
      RECT  94500.0 684750.0 95700.0 685950.0 ;
      RECT  96900.0 684750.0 98100.0 685950.0 ;
      RECT  99300.0 684750.0 100500.0 685950.0 ;
      RECT  99300.0 684750.0 100500.0 685950.0 ;
      RECT  96900.0 684750.0 98100.0 685950.0 ;
      RECT  99300.0 684750.0 100500.0 685950.0 ;
      RECT  101700.0 684750.0 102900.0 685950.0 ;
      RECT  101700.0 684750.0 102900.0 685950.0 ;
      RECT  99300.0 684750.0 100500.0 685950.0 ;
      RECT  104100.0 694050.0 105300.0 695250.0 ;
      RECT  104100.0 684150.0 105300.0 685350.0 ;
      RECT  101700.0 686850.0 100500.0 688050.0 ;
      RECT  99300.0 688800.0 98100.0 690000.0 ;
      RECT  96900.0 690750.0 95700.0 691950.0 ;
      RECT  96900.0 693450.0 98100.0 694650.0 ;
      RECT  101700.0 693450.0 102900.0 694650.0 ;
      RECT  101700.0 684750.0 102900.0 685950.0 ;
      RECT  101700.0 690750.0 102900.0 691950.0 ;
      RECT  95700.0 690750.0 96900.0 691950.0 ;
      RECT  98100.0 688800.0 99300.0 690000.0 ;
      RECT  100500.0 686850.0 101700.0 688050.0 ;
      RECT  101700.0 690750.0 102900.0 691950.0 ;
      RECT  92700.0 696150.0 108300.0 697050.0 ;
      RECT  92700.0 682350.0 108300.0 683250.0 ;
      RECT  94500.0 708450.0 95700.0 710850.0 ;
      RECT  94500.0 699750.0 95700.0 696150.0 ;
      RECT  99300.0 699750.0 100500.0 696150.0 ;
      RECT  104100.0 698550.0 105300.0 696600.0 ;
      RECT  104100.0 710400.0 105300.0 708450.0 ;
      RECT  94500.0 699750.0 95700.0 698550.0 ;
      RECT  96900.0 699750.0 98100.0 698550.0 ;
      RECT  96900.0 699750.0 98100.0 698550.0 ;
      RECT  94500.0 699750.0 95700.0 698550.0 ;
      RECT  96900.0 699750.0 98100.0 698550.0 ;
      RECT  99300.0 699750.0 100500.0 698550.0 ;
      RECT  99300.0 699750.0 100500.0 698550.0 ;
      RECT  96900.0 699750.0 98100.0 698550.0 ;
      RECT  99300.0 699750.0 100500.0 698550.0 ;
      RECT  101700.0 699750.0 102900.0 698550.0 ;
      RECT  101700.0 699750.0 102900.0 698550.0 ;
      RECT  99300.0 699750.0 100500.0 698550.0 ;
      RECT  94500.0 708450.0 95700.0 707250.0 ;
      RECT  96900.0 708450.0 98100.0 707250.0 ;
      RECT  96900.0 708450.0 98100.0 707250.0 ;
      RECT  94500.0 708450.0 95700.0 707250.0 ;
      RECT  96900.0 708450.0 98100.0 707250.0 ;
      RECT  99300.0 708450.0 100500.0 707250.0 ;
      RECT  99300.0 708450.0 100500.0 707250.0 ;
      RECT  96900.0 708450.0 98100.0 707250.0 ;
      RECT  99300.0 708450.0 100500.0 707250.0 ;
      RECT  101700.0 708450.0 102900.0 707250.0 ;
      RECT  101700.0 708450.0 102900.0 707250.0 ;
      RECT  99300.0 708450.0 100500.0 707250.0 ;
      RECT  104100.0 699150.0 105300.0 697950.0 ;
      RECT  104100.0 709050.0 105300.0 707850.0 ;
      RECT  101700.0 706350.0 100500.0 705150.0 ;
      RECT  99300.0 704400.0 98100.0 703200.0 ;
      RECT  96900.0 702450.0 95700.0 701250.0 ;
      RECT  96900.0 699750.0 98100.0 698550.0 ;
      RECT  101700.0 699750.0 102900.0 698550.0 ;
      RECT  101700.0 708450.0 102900.0 707250.0 ;
      RECT  101700.0 702450.0 102900.0 701250.0 ;
      RECT  95700.0 702450.0 96900.0 701250.0 ;
      RECT  98100.0 704400.0 99300.0 703200.0 ;
      RECT  100500.0 706350.0 101700.0 705150.0 ;
      RECT  101700.0 702450.0 102900.0 701250.0 ;
      RECT  92700.0 697050.0 108300.0 696150.0 ;
      RECT  92700.0 710850.0 108300.0 709950.0 ;
      RECT  94500.0 712350.0 95700.0 709950.0 ;
      RECT  94500.0 721050.0 95700.0 724650.0 ;
      RECT  99300.0 721050.0 100500.0 724650.0 ;
      RECT  104100.0 722250.0 105300.0 724200.0 ;
      RECT  104100.0 710400.0 105300.0 712350.0 ;
      RECT  94500.0 721050.0 95700.0 722250.0 ;
      RECT  96900.0 721050.0 98100.0 722250.0 ;
      RECT  96900.0 721050.0 98100.0 722250.0 ;
      RECT  94500.0 721050.0 95700.0 722250.0 ;
      RECT  96900.0 721050.0 98100.0 722250.0 ;
      RECT  99300.0 721050.0 100500.0 722250.0 ;
      RECT  99300.0 721050.0 100500.0 722250.0 ;
      RECT  96900.0 721050.0 98100.0 722250.0 ;
      RECT  99300.0 721050.0 100500.0 722250.0 ;
      RECT  101700.0 721050.0 102900.0 722250.0 ;
      RECT  101700.0 721050.0 102900.0 722250.0 ;
      RECT  99300.0 721050.0 100500.0 722250.0 ;
      RECT  94500.0 712350.0 95700.0 713550.0 ;
      RECT  96900.0 712350.0 98100.0 713550.0 ;
      RECT  96900.0 712350.0 98100.0 713550.0 ;
      RECT  94500.0 712350.0 95700.0 713550.0 ;
      RECT  96900.0 712350.0 98100.0 713550.0 ;
      RECT  99300.0 712350.0 100500.0 713550.0 ;
      RECT  99300.0 712350.0 100500.0 713550.0 ;
      RECT  96900.0 712350.0 98100.0 713550.0 ;
      RECT  99300.0 712350.0 100500.0 713550.0 ;
      RECT  101700.0 712350.0 102900.0 713550.0 ;
      RECT  101700.0 712350.0 102900.0 713550.0 ;
      RECT  99300.0 712350.0 100500.0 713550.0 ;
      RECT  104100.0 721650.0 105300.0 722850.0 ;
      RECT  104100.0 711750.0 105300.0 712950.0 ;
      RECT  101700.0 714450.0 100500.0 715650.0 ;
      RECT  99300.0 716400.0 98100.0 717600.0 ;
      RECT  96900.0 718350.0 95700.0 719550.0 ;
      RECT  96900.0 721050.0 98100.0 722250.0 ;
      RECT  101700.0 721050.0 102900.0 722250.0 ;
      RECT  101700.0 712350.0 102900.0 713550.0 ;
      RECT  101700.0 718350.0 102900.0 719550.0 ;
      RECT  95700.0 718350.0 96900.0 719550.0 ;
      RECT  98100.0 716400.0 99300.0 717600.0 ;
      RECT  100500.0 714450.0 101700.0 715650.0 ;
      RECT  101700.0 718350.0 102900.0 719550.0 ;
      RECT  92700.0 723750.0 108300.0 724650.0 ;
      RECT  92700.0 709950.0 108300.0 710850.0 ;
      RECT  94500.0 736050.0 95700.0 738450.0 ;
      RECT  94500.0 727350.0 95700.0 723750.0 ;
      RECT  99300.0 727350.0 100500.0 723750.0 ;
      RECT  104100.0 726150.0 105300.0 724200.0 ;
      RECT  104100.0 738000.0 105300.0 736050.0 ;
      RECT  94500.0 727350.0 95700.0 726150.0 ;
      RECT  96900.0 727350.0 98100.0 726150.0 ;
      RECT  96900.0 727350.0 98100.0 726150.0 ;
      RECT  94500.0 727350.0 95700.0 726150.0 ;
      RECT  96900.0 727350.0 98100.0 726150.0 ;
      RECT  99300.0 727350.0 100500.0 726150.0 ;
      RECT  99300.0 727350.0 100500.0 726150.0 ;
      RECT  96900.0 727350.0 98100.0 726150.0 ;
      RECT  99300.0 727350.0 100500.0 726150.0 ;
      RECT  101700.0 727350.0 102900.0 726150.0 ;
      RECT  101700.0 727350.0 102900.0 726150.0 ;
      RECT  99300.0 727350.0 100500.0 726150.0 ;
      RECT  94500.0 736050.0 95700.0 734850.0 ;
      RECT  96900.0 736050.0 98100.0 734850.0 ;
      RECT  96900.0 736050.0 98100.0 734850.0 ;
      RECT  94500.0 736050.0 95700.0 734850.0 ;
      RECT  96900.0 736050.0 98100.0 734850.0 ;
      RECT  99300.0 736050.0 100500.0 734850.0 ;
      RECT  99300.0 736050.0 100500.0 734850.0 ;
      RECT  96900.0 736050.0 98100.0 734850.0 ;
      RECT  99300.0 736050.0 100500.0 734850.0 ;
      RECT  101700.0 736050.0 102900.0 734850.0 ;
      RECT  101700.0 736050.0 102900.0 734850.0 ;
      RECT  99300.0 736050.0 100500.0 734850.0 ;
      RECT  104100.0 726750.0 105300.0 725550.0 ;
      RECT  104100.0 736650.0 105300.0 735450.0 ;
      RECT  101700.0 733950.0 100500.0 732750.0 ;
      RECT  99300.0 732000.0 98100.0 730800.0 ;
      RECT  96900.0 730050.0 95700.0 728850.0 ;
      RECT  96900.0 727350.0 98100.0 726150.0 ;
      RECT  101700.0 727350.0 102900.0 726150.0 ;
      RECT  101700.0 736050.0 102900.0 734850.0 ;
      RECT  101700.0 730050.0 102900.0 728850.0 ;
      RECT  95700.0 730050.0 96900.0 728850.0 ;
      RECT  98100.0 732000.0 99300.0 730800.0 ;
      RECT  100500.0 733950.0 101700.0 732750.0 ;
      RECT  101700.0 730050.0 102900.0 728850.0 ;
      RECT  92700.0 724650.0 108300.0 723750.0 ;
      RECT  92700.0 738450.0 108300.0 737550.0 ;
      RECT  94500.0 739950.0 95700.0 737550.0 ;
      RECT  94500.0 748650.0 95700.0 752250.0 ;
      RECT  99300.0 748650.0 100500.0 752250.0 ;
      RECT  104100.0 749850.0 105300.0 751800.0 ;
      RECT  104100.0 738000.0 105300.0 739950.0 ;
      RECT  94500.0 748650.0 95700.0 749850.0 ;
      RECT  96900.0 748650.0 98100.0 749850.0 ;
      RECT  96900.0 748650.0 98100.0 749850.0 ;
      RECT  94500.0 748650.0 95700.0 749850.0 ;
      RECT  96900.0 748650.0 98100.0 749850.0 ;
      RECT  99300.0 748650.0 100500.0 749850.0 ;
      RECT  99300.0 748650.0 100500.0 749850.0 ;
      RECT  96900.0 748650.0 98100.0 749850.0 ;
      RECT  99300.0 748650.0 100500.0 749850.0 ;
      RECT  101700.0 748650.0 102900.0 749850.0 ;
      RECT  101700.0 748650.0 102900.0 749850.0 ;
      RECT  99300.0 748650.0 100500.0 749850.0 ;
      RECT  94500.0 739950.0 95700.0 741150.0 ;
      RECT  96900.0 739950.0 98100.0 741150.0 ;
      RECT  96900.0 739950.0 98100.0 741150.0 ;
      RECT  94500.0 739950.0 95700.0 741150.0 ;
      RECT  96900.0 739950.0 98100.0 741150.0 ;
      RECT  99300.0 739950.0 100500.0 741150.0 ;
      RECT  99300.0 739950.0 100500.0 741150.0 ;
      RECT  96900.0 739950.0 98100.0 741150.0 ;
      RECT  99300.0 739950.0 100500.0 741150.0 ;
      RECT  101700.0 739950.0 102900.0 741150.0 ;
      RECT  101700.0 739950.0 102900.0 741150.0 ;
      RECT  99300.0 739950.0 100500.0 741150.0 ;
      RECT  104100.0 749250.0 105300.0 750450.0 ;
      RECT  104100.0 739350.0 105300.0 740550.0 ;
      RECT  101700.0 742050.0 100500.0 743250.0 ;
      RECT  99300.0 744000.0 98100.0 745200.0 ;
      RECT  96900.0 745950.0 95700.0 747150.0 ;
      RECT  96900.0 748650.0 98100.0 749850.0 ;
      RECT  101700.0 748650.0 102900.0 749850.0 ;
      RECT  101700.0 739950.0 102900.0 741150.0 ;
      RECT  101700.0 745950.0 102900.0 747150.0 ;
      RECT  95700.0 745950.0 96900.0 747150.0 ;
      RECT  98100.0 744000.0 99300.0 745200.0 ;
      RECT  100500.0 742050.0 101700.0 743250.0 ;
      RECT  101700.0 745950.0 102900.0 747150.0 ;
      RECT  92700.0 751350.0 108300.0 752250.0 ;
      RECT  92700.0 737550.0 108300.0 738450.0 ;
      RECT  94500.0 763650.0 95700.0 766050.0 ;
      RECT  94500.0 754950.0 95700.0 751350.0 ;
      RECT  99300.0 754950.0 100500.0 751350.0 ;
      RECT  104100.0 753750.0 105300.0 751800.0 ;
      RECT  104100.0 765600.0 105300.0 763650.0 ;
      RECT  94500.0 754950.0 95700.0 753750.0 ;
      RECT  96900.0 754950.0 98100.0 753750.0 ;
      RECT  96900.0 754950.0 98100.0 753750.0 ;
      RECT  94500.0 754950.0 95700.0 753750.0 ;
      RECT  96900.0 754950.0 98100.0 753750.0 ;
      RECT  99300.0 754950.0 100500.0 753750.0 ;
      RECT  99300.0 754950.0 100500.0 753750.0 ;
      RECT  96900.0 754950.0 98100.0 753750.0 ;
      RECT  99300.0 754950.0 100500.0 753750.0 ;
      RECT  101700.0 754950.0 102900.0 753750.0 ;
      RECT  101700.0 754950.0 102900.0 753750.0 ;
      RECT  99300.0 754950.0 100500.0 753750.0 ;
      RECT  94500.0 763650.0 95700.0 762450.0 ;
      RECT  96900.0 763650.0 98100.0 762450.0 ;
      RECT  96900.0 763650.0 98100.0 762450.0 ;
      RECT  94500.0 763650.0 95700.0 762450.0 ;
      RECT  96900.0 763650.0 98100.0 762450.0 ;
      RECT  99300.0 763650.0 100500.0 762450.0 ;
      RECT  99300.0 763650.0 100500.0 762450.0 ;
      RECT  96900.0 763650.0 98100.0 762450.0 ;
      RECT  99300.0 763650.0 100500.0 762450.0 ;
      RECT  101700.0 763650.0 102900.0 762450.0 ;
      RECT  101700.0 763650.0 102900.0 762450.0 ;
      RECT  99300.0 763650.0 100500.0 762450.0 ;
      RECT  104100.0 754350.0 105300.0 753150.0 ;
      RECT  104100.0 764250.0 105300.0 763050.0 ;
      RECT  101700.0 761550.0 100500.0 760350.0 ;
      RECT  99300.0 759600.0 98100.0 758400.0 ;
      RECT  96900.0 757650.0 95700.0 756450.0 ;
      RECT  96900.0 754950.0 98100.0 753750.0 ;
      RECT  101700.0 754950.0 102900.0 753750.0 ;
      RECT  101700.0 763650.0 102900.0 762450.0 ;
      RECT  101700.0 757650.0 102900.0 756450.0 ;
      RECT  95700.0 757650.0 96900.0 756450.0 ;
      RECT  98100.0 759600.0 99300.0 758400.0 ;
      RECT  100500.0 761550.0 101700.0 760350.0 ;
      RECT  101700.0 757650.0 102900.0 756450.0 ;
      RECT  92700.0 752250.0 108300.0 751350.0 ;
      RECT  92700.0 766050.0 108300.0 765150.0 ;
      RECT  94500.0 767550.0 95700.0 765150.0 ;
      RECT  94500.0 776250.0 95700.0 779850.0 ;
      RECT  99300.0 776250.0 100500.0 779850.0 ;
      RECT  104100.0 777450.0 105300.0 779400.0 ;
      RECT  104100.0 765600.0 105300.0 767550.0 ;
      RECT  94500.0 776250.0 95700.0 777450.0 ;
      RECT  96900.0 776250.0 98100.0 777450.0 ;
      RECT  96900.0 776250.0 98100.0 777450.0 ;
      RECT  94500.0 776250.0 95700.0 777450.0 ;
      RECT  96900.0 776250.0 98100.0 777450.0 ;
      RECT  99300.0 776250.0 100500.0 777450.0 ;
      RECT  99300.0 776250.0 100500.0 777450.0 ;
      RECT  96900.0 776250.0 98100.0 777450.0 ;
      RECT  99300.0 776250.0 100500.0 777450.0 ;
      RECT  101700.0 776250.0 102900.0 777450.0 ;
      RECT  101700.0 776250.0 102900.0 777450.0 ;
      RECT  99300.0 776250.0 100500.0 777450.0 ;
      RECT  94500.0 767550.0 95700.0 768750.0 ;
      RECT  96900.0 767550.0 98100.0 768750.0 ;
      RECT  96900.0 767550.0 98100.0 768750.0 ;
      RECT  94500.0 767550.0 95700.0 768750.0 ;
      RECT  96900.0 767550.0 98100.0 768750.0 ;
      RECT  99300.0 767550.0 100500.0 768750.0 ;
      RECT  99300.0 767550.0 100500.0 768750.0 ;
      RECT  96900.0 767550.0 98100.0 768750.0 ;
      RECT  99300.0 767550.0 100500.0 768750.0 ;
      RECT  101700.0 767550.0 102900.0 768750.0 ;
      RECT  101700.0 767550.0 102900.0 768750.0 ;
      RECT  99300.0 767550.0 100500.0 768750.0 ;
      RECT  104100.0 776850.0 105300.0 778050.0 ;
      RECT  104100.0 766950.0 105300.0 768150.0 ;
      RECT  101700.0 769650.0 100500.0 770850.0 ;
      RECT  99300.0 771600.0 98100.0 772800.0 ;
      RECT  96900.0 773550.0 95700.0 774750.0 ;
      RECT  96900.0 776250.0 98100.0 777450.0 ;
      RECT  101700.0 776250.0 102900.0 777450.0 ;
      RECT  101700.0 767550.0 102900.0 768750.0 ;
      RECT  101700.0 773550.0 102900.0 774750.0 ;
      RECT  95700.0 773550.0 96900.0 774750.0 ;
      RECT  98100.0 771600.0 99300.0 772800.0 ;
      RECT  100500.0 769650.0 101700.0 770850.0 ;
      RECT  101700.0 773550.0 102900.0 774750.0 ;
      RECT  92700.0 778950.0 108300.0 779850.0 ;
      RECT  92700.0 765150.0 108300.0 766050.0 ;
      RECT  94500.0 791250.0 95700.0 793650.0 ;
      RECT  94500.0 782550.0 95700.0 778950.0 ;
      RECT  99300.0 782550.0 100500.0 778950.0 ;
      RECT  104100.0 781350.0 105300.0 779400.0 ;
      RECT  104100.0 793200.0 105300.0 791250.0 ;
      RECT  94500.0 782550.0 95700.0 781350.0 ;
      RECT  96900.0 782550.0 98100.0 781350.0 ;
      RECT  96900.0 782550.0 98100.0 781350.0 ;
      RECT  94500.0 782550.0 95700.0 781350.0 ;
      RECT  96900.0 782550.0 98100.0 781350.0 ;
      RECT  99300.0 782550.0 100500.0 781350.0 ;
      RECT  99300.0 782550.0 100500.0 781350.0 ;
      RECT  96900.0 782550.0 98100.0 781350.0 ;
      RECT  99300.0 782550.0 100500.0 781350.0 ;
      RECT  101700.0 782550.0 102900.0 781350.0 ;
      RECT  101700.0 782550.0 102900.0 781350.0 ;
      RECT  99300.0 782550.0 100500.0 781350.0 ;
      RECT  94500.0 791250.0 95700.0 790050.0 ;
      RECT  96900.0 791250.0 98100.0 790050.0 ;
      RECT  96900.0 791250.0 98100.0 790050.0 ;
      RECT  94500.0 791250.0 95700.0 790050.0 ;
      RECT  96900.0 791250.0 98100.0 790050.0 ;
      RECT  99300.0 791250.0 100500.0 790050.0 ;
      RECT  99300.0 791250.0 100500.0 790050.0 ;
      RECT  96900.0 791250.0 98100.0 790050.0 ;
      RECT  99300.0 791250.0 100500.0 790050.0 ;
      RECT  101700.0 791250.0 102900.0 790050.0 ;
      RECT  101700.0 791250.0 102900.0 790050.0 ;
      RECT  99300.0 791250.0 100500.0 790050.0 ;
      RECT  104100.0 781950.0 105300.0 780750.0 ;
      RECT  104100.0 791850.0 105300.0 790650.0 ;
      RECT  101700.0 789150.0 100500.0 787950.0 ;
      RECT  99300.0 787200.0 98100.0 786000.0 ;
      RECT  96900.0 785250.0 95700.0 784050.0 ;
      RECT  96900.0 782550.0 98100.0 781350.0 ;
      RECT  101700.0 782550.0 102900.0 781350.0 ;
      RECT  101700.0 791250.0 102900.0 790050.0 ;
      RECT  101700.0 785250.0 102900.0 784050.0 ;
      RECT  95700.0 785250.0 96900.0 784050.0 ;
      RECT  98100.0 787200.0 99300.0 786000.0 ;
      RECT  100500.0 789150.0 101700.0 787950.0 ;
      RECT  101700.0 785250.0 102900.0 784050.0 ;
      RECT  92700.0 779850.0 108300.0 778950.0 ;
      RECT  92700.0 793650.0 108300.0 792750.0 ;
      RECT  94500.0 795150.0 95700.0 792750.0 ;
      RECT  94500.0 803850.0 95700.0 807450.0 ;
      RECT  99300.0 803850.0 100500.0 807450.0 ;
      RECT  104100.0 805050.0 105300.0 807000.0 ;
      RECT  104100.0 793200.0 105300.0 795150.0 ;
      RECT  94500.0 803850.0 95700.0 805050.0 ;
      RECT  96900.0 803850.0 98100.0 805050.0 ;
      RECT  96900.0 803850.0 98100.0 805050.0 ;
      RECT  94500.0 803850.0 95700.0 805050.0 ;
      RECT  96900.0 803850.0 98100.0 805050.0 ;
      RECT  99300.0 803850.0 100500.0 805050.0 ;
      RECT  99300.0 803850.0 100500.0 805050.0 ;
      RECT  96900.0 803850.0 98100.0 805050.0 ;
      RECT  99300.0 803850.0 100500.0 805050.0 ;
      RECT  101700.0 803850.0 102900.0 805050.0 ;
      RECT  101700.0 803850.0 102900.0 805050.0 ;
      RECT  99300.0 803850.0 100500.0 805050.0 ;
      RECT  94500.0 795150.0 95700.0 796350.0 ;
      RECT  96900.0 795150.0 98100.0 796350.0 ;
      RECT  96900.0 795150.0 98100.0 796350.0 ;
      RECT  94500.0 795150.0 95700.0 796350.0 ;
      RECT  96900.0 795150.0 98100.0 796350.0 ;
      RECT  99300.0 795150.0 100500.0 796350.0 ;
      RECT  99300.0 795150.0 100500.0 796350.0 ;
      RECT  96900.0 795150.0 98100.0 796350.0 ;
      RECT  99300.0 795150.0 100500.0 796350.0 ;
      RECT  101700.0 795150.0 102900.0 796350.0 ;
      RECT  101700.0 795150.0 102900.0 796350.0 ;
      RECT  99300.0 795150.0 100500.0 796350.0 ;
      RECT  104100.0 804450.0 105300.0 805650.0 ;
      RECT  104100.0 794550.0 105300.0 795750.0 ;
      RECT  101700.0 797250.0 100500.0 798450.0 ;
      RECT  99300.0 799200.0 98100.0 800400.0 ;
      RECT  96900.0 801150.0 95700.0 802350.0 ;
      RECT  96900.0 803850.0 98100.0 805050.0 ;
      RECT  101700.0 803850.0 102900.0 805050.0 ;
      RECT  101700.0 795150.0 102900.0 796350.0 ;
      RECT  101700.0 801150.0 102900.0 802350.0 ;
      RECT  95700.0 801150.0 96900.0 802350.0 ;
      RECT  98100.0 799200.0 99300.0 800400.0 ;
      RECT  100500.0 797250.0 101700.0 798450.0 ;
      RECT  101700.0 801150.0 102900.0 802350.0 ;
      RECT  92700.0 806550.0 108300.0 807450.0 ;
      RECT  92700.0 792750.0 108300.0 793650.0 ;
      RECT  94500.0 818850.0 95700.0 821250.0 ;
      RECT  94500.0 810150.0 95700.0 806550.0 ;
      RECT  99300.0 810150.0 100500.0 806550.0 ;
      RECT  104100.0 808950.0 105300.0 807000.0 ;
      RECT  104100.0 820800.0 105300.0 818850.0 ;
      RECT  94500.0 810150.0 95700.0 808950.0 ;
      RECT  96900.0 810150.0 98100.0 808950.0 ;
      RECT  96900.0 810150.0 98100.0 808950.0 ;
      RECT  94500.0 810150.0 95700.0 808950.0 ;
      RECT  96900.0 810150.0 98100.0 808950.0 ;
      RECT  99300.0 810150.0 100500.0 808950.0 ;
      RECT  99300.0 810150.0 100500.0 808950.0 ;
      RECT  96900.0 810150.0 98100.0 808950.0 ;
      RECT  99300.0 810150.0 100500.0 808950.0 ;
      RECT  101700.0 810150.0 102900.0 808950.0 ;
      RECT  101700.0 810150.0 102900.0 808950.0 ;
      RECT  99300.0 810150.0 100500.0 808950.0 ;
      RECT  94500.0 818850.0 95700.0 817650.0 ;
      RECT  96900.0 818850.0 98100.0 817650.0 ;
      RECT  96900.0 818850.0 98100.0 817650.0 ;
      RECT  94500.0 818850.0 95700.0 817650.0 ;
      RECT  96900.0 818850.0 98100.0 817650.0 ;
      RECT  99300.0 818850.0 100500.0 817650.0 ;
      RECT  99300.0 818850.0 100500.0 817650.0 ;
      RECT  96900.0 818850.0 98100.0 817650.0 ;
      RECT  99300.0 818850.0 100500.0 817650.0 ;
      RECT  101700.0 818850.0 102900.0 817650.0 ;
      RECT  101700.0 818850.0 102900.0 817650.0 ;
      RECT  99300.0 818850.0 100500.0 817650.0 ;
      RECT  104100.0 809550.0 105300.0 808350.0 ;
      RECT  104100.0 819450.0 105300.0 818250.0 ;
      RECT  101700.0 816750.0 100500.0 815550.0 ;
      RECT  99300.0 814800.0 98100.0 813600.0 ;
      RECT  96900.0 812850.0 95700.0 811650.0 ;
      RECT  96900.0 810150.0 98100.0 808950.0 ;
      RECT  101700.0 810150.0 102900.0 808950.0 ;
      RECT  101700.0 818850.0 102900.0 817650.0 ;
      RECT  101700.0 812850.0 102900.0 811650.0 ;
      RECT  95700.0 812850.0 96900.0 811650.0 ;
      RECT  98100.0 814800.0 99300.0 813600.0 ;
      RECT  100500.0 816750.0 101700.0 815550.0 ;
      RECT  101700.0 812850.0 102900.0 811650.0 ;
      RECT  92700.0 807450.0 108300.0 806550.0 ;
      RECT  92700.0 821250.0 108300.0 820350.0 ;
      RECT  94500.0 822750.0 95700.0 820350.0 ;
      RECT  94500.0 831450.0 95700.0 835050.0 ;
      RECT  99300.0 831450.0 100500.0 835050.0 ;
      RECT  104100.0 832650.0 105300.0 834600.0 ;
      RECT  104100.0 820800.0 105300.0 822750.0 ;
      RECT  94500.0 831450.0 95700.0 832650.0 ;
      RECT  96900.0 831450.0 98100.0 832650.0 ;
      RECT  96900.0 831450.0 98100.0 832650.0 ;
      RECT  94500.0 831450.0 95700.0 832650.0 ;
      RECT  96900.0 831450.0 98100.0 832650.0 ;
      RECT  99300.0 831450.0 100500.0 832650.0 ;
      RECT  99300.0 831450.0 100500.0 832650.0 ;
      RECT  96900.0 831450.0 98100.0 832650.0 ;
      RECT  99300.0 831450.0 100500.0 832650.0 ;
      RECT  101700.0 831450.0 102900.0 832650.0 ;
      RECT  101700.0 831450.0 102900.0 832650.0 ;
      RECT  99300.0 831450.0 100500.0 832650.0 ;
      RECT  94500.0 822750.0 95700.0 823950.0 ;
      RECT  96900.0 822750.0 98100.0 823950.0 ;
      RECT  96900.0 822750.0 98100.0 823950.0 ;
      RECT  94500.0 822750.0 95700.0 823950.0 ;
      RECT  96900.0 822750.0 98100.0 823950.0 ;
      RECT  99300.0 822750.0 100500.0 823950.0 ;
      RECT  99300.0 822750.0 100500.0 823950.0 ;
      RECT  96900.0 822750.0 98100.0 823950.0 ;
      RECT  99300.0 822750.0 100500.0 823950.0 ;
      RECT  101700.0 822750.0 102900.0 823950.0 ;
      RECT  101700.0 822750.0 102900.0 823950.0 ;
      RECT  99300.0 822750.0 100500.0 823950.0 ;
      RECT  104100.0 832050.0 105300.0 833250.0 ;
      RECT  104100.0 822150.0 105300.0 823350.0 ;
      RECT  101700.0 824850.0 100500.0 826050.0 ;
      RECT  99300.0 826800.0 98100.0 828000.0 ;
      RECT  96900.0 828750.0 95700.0 829950.0 ;
      RECT  96900.0 831450.0 98100.0 832650.0 ;
      RECT  101700.0 831450.0 102900.0 832650.0 ;
      RECT  101700.0 822750.0 102900.0 823950.0 ;
      RECT  101700.0 828750.0 102900.0 829950.0 ;
      RECT  95700.0 828750.0 96900.0 829950.0 ;
      RECT  98100.0 826800.0 99300.0 828000.0 ;
      RECT  100500.0 824850.0 101700.0 826050.0 ;
      RECT  101700.0 828750.0 102900.0 829950.0 ;
      RECT  92700.0 834150.0 108300.0 835050.0 ;
      RECT  92700.0 820350.0 108300.0 821250.0 ;
      RECT  94500.0 846450.0 95700.0 848850.0 ;
      RECT  94500.0 837750.0 95700.0 834150.0 ;
      RECT  99300.0 837750.0 100500.0 834150.0 ;
      RECT  104100.0 836550.0 105300.0 834600.0 ;
      RECT  104100.0 848400.0 105300.0 846450.0 ;
      RECT  94500.0 837750.0 95700.0 836550.0 ;
      RECT  96900.0 837750.0 98100.0 836550.0 ;
      RECT  96900.0 837750.0 98100.0 836550.0 ;
      RECT  94500.0 837750.0 95700.0 836550.0 ;
      RECT  96900.0 837750.0 98100.0 836550.0 ;
      RECT  99300.0 837750.0 100500.0 836550.0 ;
      RECT  99300.0 837750.0 100500.0 836550.0 ;
      RECT  96900.0 837750.0 98100.0 836550.0 ;
      RECT  99300.0 837750.0 100500.0 836550.0 ;
      RECT  101700.0 837750.0 102900.0 836550.0 ;
      RECT  101700.0 837750.0 102900.0 836550.0 ;
      RECT  99300.0 837750.0 100500.0 836550.0 ;
      RECT  94500.0 846450.0 95700.0 845250.0 ;
      RECT  96900.0 846450.0 98100.0 845250.0 ;
      RECT  96900.0 846450.0 98100.0 845250.0 ;
      RECT  94500.0 846450.0 95700.0 845250.0 ;
      RECT  96900.0 846450.0 98100.0 845250.0 ;
      RECT  99300.0 846450.0 100500.0 845250.0 ;
      RECT  99300.0 846450.0 100500.0 845250.0 ;
      RECT  96900.0 846450.0 98100.0 845250.0 ;
      RECT  99300.0 846450.0 100500.0 845250.0 ;
      RECT  101700.0 846450.0 102900.0 845250.0 ;
      RECT  101700.0 846450.0 102900.0 845250.0 ;
      RECT  99300.0 846450.0 100500.0 845250.0 ;
      RECT  104100.0 837150.0 105300.0 835950.0 ;
      RECT  104100.0 847050.0 105300.0 845850.0 ;
      RECT  101700.0 844350.0 100500.0 843150.0 ;
      RECT  99300.0 842400.0 98100.0 841200.0 ;
      RECT  96900.0 840450.0 95700.0 839250.0 ;
      RECT  96900.0 837750.0 98100.0 836550.0 ;
      RECT  101700.0 837750.0 102900.0 836550.0 ;
      RECT  101700.0 846450.0 102900.0 845250.0 ;
      RECT  101700.0 840450.0 102900.0 839250.0 ;
      RECT  95700.0 840450.0 96900.0 839250.0 ;
      RECT  98100.0 842400.0 99300.0 841200.0 ;
      RECT  100500.0 844350.0 101700.0 843150.0 ;
      RECT  101700.0 840450.0 102900.0 839250.0 ;
      RECT  92700.0 835050.0 108300.0 834150.0 ;
      RECT  92700.0 848850.0 108300.0 847950.0 ;
      RECT  94500.0 850350.0 95700.0 847950.0 ;
      RECT  94500.0 859050.0 95700.0 862650.0 ;
      RECT  99300.0 859050.0 100500.0 862650.0 ;
      RECT  104100.0 860250.0 105300.0 862200.0 ;
      RECT  104100.0 848400.0 105300.0 850350.0 ;
      RECT  94500.0 859050.0 95700.0 860250.0 ;
      RECT  96900.0 859050.0 98100.0 860250.0 ;
      RECT  96900.0 859050.0 98100.0 860250.0 ;
      RECT  94500.0 859050.0 95700.0 860250.0 ;
      RECT  96900.0 859050.0 98100.0 860250.0 ;
      RECT  99300.0 859050.0 100500.0 860250.0 ;
      RECT  99300.0 859050.0 100500.0 860250.0 ;
      RECT  96900.0 859050.0 98100.0 860250.0 ;
      RECT  99300.0 859050.0 100500.0 860250.0 ;
      RECT  101700.0 859050.0 102900.0 860250.0 ;
      RECT  101700.0 859050.0 102900.0 860250.0 ;
      RECT  99300.0 859050.0 100500.0 860250.0 ;
      RECT  94500.0 850350.0 95700.0 851550.0 ;
      RECT  96900.0 850350.0 98100.0 851550.0 ;
      RECT  96900.0 850350.0 98100.0 851550.0 ;
      RECT  94500.0 850350.0 95700.0 851550.0 ;
      RECT  96900.0 850350.0 98100.0 851550.0 ;
      RECT  99300.0 850350.0 100500.0 851550.0 ;
      RECT  99300.0 850350.0 100500.0 851550.0 ;
      RECT  96900.0 850350.0 98100.0 851550.0 ;
      RECT  99300.0 850350.0 100500.0 851550.0 ;
      RECT  101700.0 850350.0 102900.0 851550.0 ;
      RECT  101700.0 850350.0 102900.0 851550.0 ;
      RECT  99300.0 850350.0 100500.0 851550.0 ;
      RECT  104100.0 859650.0 105300.0 860850.0 ;
      RECT  104100.0 849750.0 105300.0 850950.0 ;
      RECT  101700.0 852450.0 100500.0 853650.0 ;
      RECT  99300.0 854400.0 98100.0 855600.0 ;
      RECT  96900.0 856350.0 95700.0 857550.0 ;
      RECT  96900.0 859050.0 98100.0 860250.0 ;
      RECT  101700.0 859050.0 102900.0 860250.0 ;
      RECT  101700.0 850350.0 102900.0 851550.0 ;
      RECT  101700.0 856350.0 102900.0 857550.0 ;
      RECT  95700.0 856350.0 96900.0 857550.0 ;
      RECT  98100.0 854400.0 99300.0 855600.0 ;
      RECT  100500.0 852450.0 101700.0 853650.0 ;
      RECT  101700.0 856350.0 102900.0 857550.0 ;
      RECT  92700.0 861750.0 108300.0 862650.0 ;
      RECT  92700.0 847950.0 108300.0 848850.0 ;
      RECT  94500.0 874050.0 95700.0 876450.0 ;
      RECT  94500.0 865350.0 95700.0 861750.0 ;
      RECT  99300.0 865350.0 100500.0 861750.0 ;
      RECT  104100.0 864150.0 105300.0 862200.0 ;
      RECT  104100.0 876000.0 105300.0 874050.0 ;
      RECT  94500.0 865350.0 95700.0 864150.0 ;
      RECT  96900.0 865350.0 98100.0 864150.0 ;
      RECT  96900.0 865350.0 98100.0 864150.0 ;
      RECT  94500.0 865350.0 95700.0 864150.0 ;
      RECT  96900.0 865350.0 98100.0 864150.0 ;
      RECT  99300.0 865350.0 100500.0 864150.0 ;
      RECT  99300.0 865350.0 100500.0 864150.0 ;
      RECT  96900.0 865350.0 98100.0 864150.0 ;
      RECT  99300.0 865350.0 100500.0 864150.0 ;
      RECT  101700.0 865350.0 102900.0 864150.0 ;
      RECT  101700.0 865350.0 102900.0 864150.0 ;
      RECT  99300.0 865350.0 100500.0 864150.0 ;
      RECT  94500.0 874050.0 95700.0 872850.0 ;
      RECT  96900.0 874050.0 98100.0 872850.0 ;
      RECT  96900.0 874050.0 98100.0 872850.0 ;
      RECT  94500.0 874050.0 95700.0 872850.0 ;
      RECT  96900.0 874050.0 98100.0 872850.0 ;
      RECT  99300.0 874050.0 100500.0 872850.0 ;
      RECT  99300.0 874050.0 100500.0 872850.0 ;
      RECT  96900.0 874050.0 98100.0 872850.0 ;
      RECT  99300.0 874050.0 100500.0 872850.0 ;
      RECT  101700.0 874050.0 102900.0 872850.0 ;
      RECT  101700.0 874050.0 102900.0 872850.0 ;
      RECT  99300.0 874050.0 100500.0 872850.0 ;
      RECT  104100.0 864750.0 105300.0 863550.0 ;
      RECT  104100.0 874650.0 105300.0 873450.0 ;
      RECT  101700.0 871950.0 100500.0 870750.0 ;
      RECT  99300.0 870000.0 98100.0 868800.0 ;
      RECT  96900.0 868050.0 95700.0 866850.0 ;
      RECT  96900.0 865350.0 98100.0 864150.0 ;
      RECT  101700.0 865350.0 102900.0 864150.0 ;
      RECT  101700.0 874050.0 102900.0 872850.0 ;
      RECT  101700.0 868050.0 102900.0 866850.0 ;
      RECT  95700.0 868050.0 96900.0 866850.0 ;
      RECT  98100.0 870000.0 99300.0 868800.0 ;
      RECT  100500.0 871950.0 101700.0 870750.0 ;
      RECT  101700.0 868050.0 102900.0 866850.0 ;
      RECT  92700.0 862650.0 108300.0 861750.0 ;
      RECT  92700.0 876450.0 108300.0 875550.0 ;
      RECT  94500.0 877950.0 95700.0 875550.0 ;
      RECT  94500.0 886650.0 95700.0 890250.0 ;
      RECT  99300.0 886650.0 100500.0 890250.0 ;
      RECT  104100.0 887850.0 105300.0 889800.0 ;
      RECT  104100.0 876000.0 105300.0 877950.0 ;
      RECT  94500.0 886650.0 95700.0 887850.0 ;
      RECT  96900.0 886650.0 98100.0 887850.0 ;
      RECT  96900.0 886650.0 98100.0 887850.0 ;
      RECT  94500.0 886650.0 95700.0 887850.0 ;
      RECT  96900.0 886650.0 98100.0 887850.0 ;
      RECT  99300.0 886650.0 100500.0 887850.0 ;
      RECT  99300.0 886650.0 100500.0 887850.0 ;
      RECT  96900.0 886650.0 98100.0 887850.0 ;
      RECT  99300.0 886650.0 100500.0 887850.0 ;
      RECT  101700.0 886650.0 102900.0 887850.0 ;
      RECT  101700.0 886650.0 102900.0 887850.0 ;
      RECT  99300.0 886650.0 100500.0 887850.0 ;
      RECT  94500.0 877950.0 95700.0 879150.0 ;
      RECT  96900.0 877950.0 98100.0 879150.0 ;
      RECT  96900.0 877950.0 98100.0 879150.0 ;
      RECT  94500.0 877950.0 95700.0 879150.0 ;
      RECT  96900.0 877950.0 98100.0 879150.0 ;
      RECT  99300.0 877950.0 100500.0 879150.0 ;
      RECT  99300.0 877950.0 100500.0 879150.0 ;
      RECT  96900.0 877950.0 98100.0 879150.0 ;
      RECT  99300.0 877950.0 100500.0 879150.0 ;
      RECT  101700.0 877950.0 102900.0 879150.0 ;
      RECT  101700.0 877950.0 102900.0 879150.0 ;
      RECT  99300.0 877950.0 100500.0 879150.0 ;
      RECT  104100.0 887250.0 105300.0 888450.0 ;
      RECT  104100.0 877350.0 105300.0 878550.0 ;
      RECT  101700.0 880050.0 100500.0 881250.0 ;
      RECT  99300.0 882000.0 98100.0 883200.0 ;
      RECT  96900.0 883950.0 95700.0 885150.0 ;
      RECT  96900.0 886650.0 98100.0 887850.0 ;
      RECT  101700.0 886650.0 102900.0 887850.0 ;
      RECT  101700.0 877950.0 102900.0 879150.0 ;
      RECT  101700.0 883950.0 102900.0 885150.0 ;
      RECT  95700.0 883950.0 96900.0 885150.0 ;
      RECT  98100.0 882000.0 99300.0 883200.0 ;
      RECT  100500.0 880050.0 101700.0 881250.0 ;
      RECT  101700.0 883950.0 102900.0 885150.0 ;
      RECT  92700.0 889350.0 108300.0 890250.0 ;
      RECT  92700.0 875550.0 108300.0 876450.0 ;
      RECT  94500.0 901650.0 95700.0 904050.0 ;
      RECT  94500.0 892950.0 95700.0 889350.0 ;
      RECT  99300.0 892950.0 100500.0 889350.0 ;
      RECT  104100.0 891750.0 105300.0 889800.0 ;
      RECT  104100.0 903600.0 105300.0 901650.0 ;
      RECT  94500.0 892950.0 95700.0 891750.0 ;
      RECT  96900.0 892950.0 98100.0 891750.0 ;
      RECT  96900.0 892950.0 98100.0 891750.0 ;
      RECT  94500.0 892950.0 95700.0 891750.0 ;
      RECT  96900.0 892950.0 98100.0 891750.0 ;
      RECT  99300.0 892950.0 100500.0 891750.0 ;
      RECT  99300.0 892950.0 100500.0 891750.0 ;
      RECT  96900.0 892950.0 98100.0 891750.0 ;
      RECT  99300.0 892950.0 100500.0 891750.0 ;
      RECT  101700.0 892950.0 102900.0 891750.0 ;
      RECT  101700.0 892950.0 102900.0 891750.0 ;
      RECT  99300.0 892950.0 100500.0 891750.0 ;
      RECT  94500.0 901650.0 95700.0 900450.0 ;
      RECT  96900.0 901650.0 98100.0 900450.0 ;
      RECT  96900.0 901650.0 98100.0 900450.0 ;
      RECT  94500.0 901650.0 95700.0 900450.0 ;
      RECT  96900.0 901650.0 98100.0 900450.0 ;
      RECT  99300.0 901650.0 100500.0 900450.0 ;
      RECT  99300.0 901650.0 100500.0 900450.0 ;
      RECT  96900.0 901650.0 98100.0 900450.0 ;
      RECT  99300.0 901650.0 100500.0 900450.0 ;
      RECT  101700.0 901650.0 102900.0 900450.0 ;
      RECT  101700.0 901650.0 102900.0 900450.0 ;
      RECT  99300.0 901650.0 100500.0 900450.0 ;
      RECT  104100.0 892350.0 105300.0 891150.0 ;
      RECT  104100.0 902250.0 105300.0 901050.0 ;
      RECT  101700.0 899550.0 100500.0 898350.0 ;
      RECT  99300.0 897600.0 98100.0 896400.0 ;
      RECT  96900.0 895650.0 95700.0 894450.0 ;
      RECT  96900.0 892950.0 98100.0 891750.0 ;
      RECT  101700.0 892950.0 102900.0 891750.0 ;
      RECT  101700.0 901650.0 102900.0 900450.0 ;
      RECT  101700.0 895650.0 102900.0 894450.0 ;
      RECT  95700.0 895650.0 96900.0 894450.0 ;
      RECT  98100.0 897600.0 99300.0 896400.0 ;
      RECT  100500.0 899550.0 101700.0 898350.0 ;
      RECT  101700.0 895650.0 102900.0 894450.0 ;
      RECT  92700.0 890250.0 108300.0 889350.0 ;
      RECT  92700.0 904050.0 108300.0 903150.0 ;
      RECT  94500.0 905550.0 95700.0 903150.0 ;
      RECT  94500.0 914250.0 95700.0 917850.0 ;
      RECT  99300.0 914250.0 100500.0 917850.0 ;
      RECT  104100.0 915450.0 105300.0 917400.0 ;
      RECT  104100.0 903600.0 105300.0 905550.0 ;
      RECT  94500.0 914250.0 95700.0 915450.0 ;
      RECT  96900.0 914250.0 98100.0 915450.0 ;
      RECT  96900.0 914250.0 98100.0 915450.0 ;
      RECT  94500.0 914250.0 95700.0 915450.0 ;
      RECT  96900.0 914250.0 98100.0 915450.0 ;
      RECT  99300.0 914250.0 100500.0 915450.0 ;
      RECT  99300.0 914250.0 100500.0 915450.0 ;
      RECT  96900.0 914250.0 98100.0 915450.0 ;
      RECT  99300.0 914250.0 100500.0 915450.0 ;
      RECT  101700.0 914250.0 102900.0 915450.0 ;
      RECT  101700.0 914250.0 102900.0 915450.0 ;
      RECT  99300.0 914250.0 100500.0 915450.0 ;
      RECT  94500.0 905550.0 95700.0 906750.0 ;
      RECT  96900.0 905550.0 98100.0 906750.0 ;
      RECT  96900.0 905550.0 98100.0 906750.0 ;
      RECT  94500.0 905550.0 95700.0 906750.0 ;
      RECT  96900.0 905550.0 98100.0 906750.0 ;
      RECT  99300.0 905550.0 100500.0 906750.0 ;
      RECT  99300.0 905550.0 100500.0 906750.0 ;
      RECT  96900.0 905550.0 98100.0 906750.0 ;
      RECT  99300.0 905550.0 100500.0 906750.0 ;
      RECT  101700.0 905550.0 102900.0 906750.0 ;
      RECT  101700.0 905550.0 102900.0 906750.0 ;
      RECT  99300.0 905550.0 100500.0 906750.0 ;
      RECT  104100.0 914850.0 105300.0 916050.0 ;
      RECT  104100.0 904950.0 105300.0 906150.0 ;
      RECT  101700.0 907650.0 100500.0 908850.0 ;
      RECT  99300.0 909600.0 98100.0 910800.0 ;
      RECT  96900.0 911550.0 95700.0 912750.0 ;
      RECT  96900.0 914250.0 98100.0 915450.0 ;
      RECT  101700.0 914250.0 102900.0 915450.0 ;
      RECT  101700.0 905550.0 102900.0 906750.0 ;
      RECT  101700.0 911550.0 102900.0 912750.0 ;
      RECT  95700.0 911550.0 96900.0 912750.0 ;
      RECT  98100.0 909600.0 99300.0 910800.0 ;
      RECT  100500.0 907650.0 101700.0 908850.0 ;
      RECT  101700.0 911550.0 102900.0 912750.0 ;
      RECT  92700.0 916950.0 108300.0 917850.0 ;
      RECT  92700.0 903150.0 108300.0 904050.0 ;
      RECT  94500.0 929250.0 95700.0 931650.0 ;
      RECT  94500.0 920550.0 95700.0 916950.0 ;
      RECT  99300.0 920550.0 100500.0 916950.0 ;
      RECT  104100.0 919350.0 105300.0 917400.0 ;
      RECT  104100.0 931200.0 105300.0 929250.0 ;
      RECT  94500.0 920550.0 95700.0 919350.0 ;
      RECT  96900.0 920550.0 98100.0 919350.0 ;
      RECT  96900.0 920550.0 98100.0 919350.0 ;
      RECT  94500.0 920550.0 95700.0 919350.0 ;
      RECT  96900.0 920550.0 98100.0 919350.0 ;
      RECT  99300.0 920550.0 100500.0 919350.0 ;
      RECT  99300.0 920550.0 100500.0 919350.0 ;
      RECT  96900.0 920550.0 98100.0 919350.0 ;
      RECT  99300.0 920550.0 100500.0 919350.0 ;
      RECT  101700.0 920550.0 102900.0 919350.0 ;
      RECT  101700.0 920550.0 102900.0 919350.0 ;
      RECT  99300.0 920550.0 100500.0 919350.0 ;
      RECT  94500.0 929250.0 95700.0 928050.0 ;
      RECT  96900.0 929250.0 98100.0 928050.0 ;
      RECT  96900.0 929250.0 98100.0 928050.0 ;
      RECT  94500.0 929250.0 95700.0 928050.0 ;
      RECT  96900.0 929250.0 98100.0 928050.0 ;
      RECT  99300.0 929250.0 100500.0 928050.0 ;
      RECT  99300.0 929250.0 100500.0 928050.0 ;
      RECT  96900.0 929250.0 98100.0 928050.0 ;
      RECT  99300.0 929250.0 100500.0 928050.0 ;
      RECT  101700.0 929250.0 102900.0 928050.0 ;
      RECT  101700.0 929250.0 102900.0 928050.0 ;
      RECT  99300.0 929250.0 100500.0 928050.0 ;
      RECT  104100.0 919950.0 105300.0 918750.0 ;
      RECT  104100.0 929850.0 105300.0 928650.0 ;
      RECT  101700.0 927150.0 100500.0 925950.0 ;
      RECT  99300.0 925200.0 98100.0 924000.0 ;
      RECT  96900.0 923250.0 95700.0 922050.0 ;
      RECT  96900.0 920550.0 98100.0 919350.0 ;
      RECT  101700.0 920550.0 102900.0 919350.0 ;
      RECT  101700.0 929250.0 102900.0 928050.0 ;
      RECT  101700.0 923250.0 102900.0 922050.0 ;
      RECT  95700.0 923250.0 96900.0 922050.0 ;
      RECT  98100.0 925200.0 99300.0 924000.0 ;
      RECT  100500.0 927150.0 101700.0 925950.0 ;
      RECT  101700.0 923250.0 102900.0 922050.0 ;
      RECT  92700.0 917850.0 108300.0 916950.0 ;
      RECT  92700.0 931650.0 108300.0 930750.0 ;
      RECT  94500.0 933150.0 95700.0 930750.0 ;
      RECT  94500.0 941850.0 95700.0 945450.0 ;
      RECT  99300.0 941850.0 100500.0 945450.0 ;
      RECT  104100.0 943050.0 105300.0 945000.0 ;
      RECT  104100.0 931200.0 105300.0 933150.0 ;
      RECT  94500.0 941850.0 95700.0 943050.0 ;
      RECT  96900.0 941850.0 98100.0 943050.0 ;
      RECT  96900.0 941850.0 98100.0 943050.0 ;
      RECT  94500.0 941850.0 95700.0 943050.0 ;
      RECT  96900.0 941850.0 98100.0 943050.0 ;
      RECT  99300.0 941850.0 100500.0 943050.0 ;
      RECT  99300.0 941850.0 100500.0 943050.0 ;
      RECT  96900.0 941850.0 98100.0 943050.0 ;
      RECT  99300.0 941850.0 100500.0 943050.0 ;
      RECT  101700.0 941850.0 102900.0 943050.0 ;
      RECT  101700.0 941850.0 102900.0 943050.0 ;
      RECT  99300.0 941850.0 100500.0 943050.0 ;
      RECT  94500.0 933150.0 95700.0 934350.0 ;
      RECT  96900.0 933150.0 98100.0 934350.0 ;
      RECT  96900.0 933150.0 98100.0 934350.0 ;
      RECT  94500.0 933150.0 95700.0 934350.0 ;
      RECT  96900.0 933150.0 98100.0 934350.0 ;
      RECT  99300.0 933150.0 100500.0 934350.0 ;
      RECT  99300.0 933150.0 100500.0 934350.0 ;
      RECT  96900.0 933150.0 98100.0 934350.0 ;
      RECT  99300.0 933150.0 100500.0 934350.0 ;
      RECT  101700.0 933150.0 102900.0 934350.0 ;
      RECT  101700.0 933150.0 102900.0 934350.0 ;
      RECT  99300.0 933150.0 100500.0 934350.0 ;
      RECT  104100.0 942450.0 105300.0 943650.0 ;
      RECT  104100.0 932550.0 105300.0 933750.0 ;
      RECT  101700.0 935250.0 100500.0 936450.0 ;
      RECT  99300.0 937200.0 98100.0 938400.0 ;
      RECT  96900.0 939150.0 95700.0 940350.0 ;
      RECT  96900.0 941850.0 98100.0 943050.0 ;
      RECT  101700.0 941850.0 102900.0 943050.0 ;
      RECT  101700.0 933150.0 102900.0 934350.0 ;
      RECT  101700.0 939150.0 102900.0 940350.0 ;
      RECT  95700.0 939150.0 96900.0 940350.0 ;
      RECT  98100.0 937200.0 99300.0 938400.0 ;
      RECT  100500.0 935250.0 101700.0 936450.0 ;
      RECT  101700.0 939150.0 102900.0 940350.0 ;
      RECT  92700.0 944550.0 108300.0 945450.0 ;
      RECT  92700.0 930750.0 108300.0 931650.0 ;
      RECT  94500.0 956850.0 95700.0 959250.0 ;
      RECT  94500.0 948150.0 95700.0 944550.0 ;
      RECT  99300.0 948150.0 100500.0 944550.0 ;
      RECT  104100.0 946950.0 105300.0 945000.0 ;
      RECT  104100.0 958800.0 105300.0 956850.0 ;
      RECT  94500.0 948150.0 95700.0 946950.0 ;
      RECT  96900.0 948150.0 98100.0 946950.0 ;
      RECT  96900.0 948150.0 98100.0 946950.0 ;
      RECT  94500.0 948150.0 95700.0 946950.0 ;
      RECT  96900.0 948150.0 98100.0 946950.0 ;
      RECT  99300.0 948150.0 100500.0 946950.0 ;
      RECT  99300.0 948150.0 100500.0 946950.0 ;
      RECT  96900.0 948150.0 98100.0 946950.0 ;
      RECT  99300.0 948150.0 100500.0 946950.0 ;
      RECT  101700.0 948150.0 102900.0 946950.0 ;
      RECT  101700.0 948150.0 102900.0 946950.0 ;
      RECT  99300.0 948150.0 100500.0 946950.0 ;
      RECT  94500.0 956850.0 95700.0 955650.0 ;
      RECT  96900.0 956850.0 98100.0 955650.0 ;
      RECT  96900.0 956850.0 98100.0 955650.0 ;
      RECT  94500.0 956850.0 95700.0 955650.0 ;
      RECT  96900.0 956850.0 98100.0 955650.0 ;
      RECT  99300.0 956850.0 100500.0 955650.0 ;
      RECT  99300.0 956850.0 100500.0 955650.0 ;
      RECT  96900.0 956850.0 98100.0 955650.0 ;
      RECT  99300.0 956850.0 100500.0 955650.0 ;
      RECT  101700.0 956850.0 102900.0 955650.0 ;
      RECT  101700.0 956850.0 102900.0 955650.0 ;
      RECT  99300.0 956850.0 100500.0 955650.0 ;
      RECT  104100.0 947550.0 105300.0 946350.0 ;
      RECT  104100.0 957450.0 105300.0 956250.0 ;
      RECT  101700.0 954750.0 100500.0 953550.0 ;
      RECT  99300.0 952800.0 98100.0 951600.0 ;
      RECT  96900.0 950850.0 95700.0 949650.0 ;
      RECT  96900.0 948150.0 98100.0 946950.0 ;
      RECT  101700.0 948150.0 102900.0 946950.0 ;
      RECT  101700.0 956850.0 102900.0 955650.0 ;
      RECT  101700.0 950850.0 102900.0 949650.0 ;
      RECT  95700.0 950850.0 96900.0 949650.0 ;
      RECT  98100.0 952800.0 99300.0 951600.0 ;
      RECT  100500.0 954750.0 101700.0 953550.0 ;
      RECT  101700.0 950850.0 102900.0 949650.0 ;
      RECT  92700.0 945450.0 108300.0 944550.0 ;
      RECT  92700.0 959250.0 108300.0 958350.0 ;
      RECT  94500.0 960750.0 95700.0 958350.0 ;
      RECT  94500.0 969450.0 95700.0 973050.0 ;
      RECT  99300.0 969450.0 100500.0 973050.0 ;
      RECT  104100.0 970650.0 105300.0 972600.0 ;
      RECT  104100.0 958800.0 105300.0 960750.0 ;
      RECT  94500.0 969450.0 95700.0 970650.0 ;
      RECT  96900.0 969450.0 98100.0 970650.0 ;
      RECT  96900.0 969450.0 98100.0 970650.0 ;
      RECT  94500.0 969450.0 95700.0 970650.0 ;
      RECT  96900.0 969450.0 98100.0 970650.0 ;
      RECT  99300.0 969450.0 100500.0 970650.0 ;
      RECT  99300.0 969450.0 100500.0 970650.0 ;
      RECT  96900.0 969450.0 98100.0 970650.0 ;
      RECT  99300.0 969450.0 100500.0 970650.0 ;
      RECT  101700.0 969450.0 102900.0 970650.0 ;
      RECT  101700.0 969450.0 102900.0 970650.0 ;
      RECT  99300.0 969450.0 100500.0 970650.0 ;
      RECT  94500.0 960750.0 95700.0 961950.0 ;
      RECT  96900.0 960750.0 98100.0 961950.0 ;
      RECT  96900.0 960750.0 98100.0 961950.0 ;
      RECT  94500.0 960750.0 95700.0 961950.0 ;
      RECT  96900.0 960750.0 98100.0 961950.0 ;
      RECT  99300.0 960750.0 100500.0 961950.0 ;
      RECT  99300.0 960750.0 100500.0 961950.0 ;
      RECT  96900.0 960750.0 98100.0 961950.0 ;
      RECT  99300.0 960750.0 100500.0 961950.0 ;
      RECT  101700.0 960750.0 102900.0 961950.0 ;
      RECT  101700.0 960750.0 102900.0 961950.0 ;
      RECT  99300.0 960750.0 100500.0 961950.0 ;
      RECT  104100.0 970050.0 105300.0 971250.0 ;
      RECT  104100.0 960150.0 105300.0 961350.0 ;
      RECT  101700.0 962850.0 100500.0 964050.0 ;
      RECT  99300.0 964800.0 98100.0 966000.0 ;
      RECT  96900.0 966750.0 95700.0 967950.0 ;
      RECT  96900.0 969450.0 98100.0 970650.0 ;
      RECT  101700.0 969450.0 102900.0 970650.0 ;
      RECT  101700.0 960750.0 102900.0 961950.0 ;
      RECT  101700.0 966750.0 102900.0 967950.0 ;
      RECT  95700.0 966750.0 96900.0 967950.0 ;
      RECT  98100.0 964800.0 99300.0 966000.0 ;
      RECT  100500.0 962850.0 101700.0 964050.0 ;
      RECT  101700.0 966750.0 102900.0 967950.0 ;
      RECT  92700.0 972150.0 108300.0 973050.0 ;
      RECT  92700.0 958350.0 108300.0 959250.0 ;
      RECT  94500.0 984450.0 95700.0 986850.0 ;
      RECT  94500.0 975750.0 95700.0 972150.0 ;
      RECT  99300.0 975750.0 100500.0 972150.0 ;
      RECT  104100.0 974550.0 105300.0 972600.0 ;
      RECT  104100.0 986400.0 105300.0 984450.0 ;
      RECT  94500.0 975750.0 95700.0 974550.0 ;
      RECT  96900.0 975750.0 98100.0 974550.0 ;
      RECT  96900.0 975750.0 98100.0 974550.0 ;
      RECT  94500.0 975750.0 95700.0 974550.0 ;
      RECT  96900.0 975750.0 98100.0 974550.0 ;
      RECT  99300.0 975750.0 100500.0 974550.0 ;
      RECT  99300.0 975750.0 100500.0 974550.0 ;
      RECT  96900.0 975750.0 98100.0 974550.0 ;
      RECT  99300.0 975750.0 100500.0 974550.0 ;
      RECT  101700.0 975750.0 102900.0 974550.0 ;
      RECT  101700.0 975750.0 102900.0 974550.0 ;
      RECT  99300.0 975750.0 100500.0 974550.0 ;
      RECT  94500.0 984450.0 95700.0 983250.0 ;
      RECT  96900.0 984450.0 98100.0 983250.0 ;
      RECT  96900.0 984450.0 98100.0 983250.0 ;
      RECT  94500.0 984450.0 95700.0 983250.0 ;
      RECT  96900.0 984450.0 98100.0 983250.0 ;
      RECT  99300.0 984450.0 100500.0 983250.0 ;
      RECT  99300.0 984450.0 100500.0 983250.0 ;
      RECT  96900.0 984450.0 98100.0 983250.0 ;
      RECT  99300.0 984450.0 100500.0 983250.0 ;
      RECT  101700.0 984450.0 102900.0 983250.0 ;
      RECT  101700.0 984450.0 102900.0 983250.0 ;
      RECT  99300.0 984450.0 100500.0 983250.0 ;
      RECT  104100.0 975150.0 105300.0 973950.0 ;
      RECT  104100.0 985050.0 105300.0 983850.0 ;
      RECT  101700.0 982350.0 100500.0 981150.0 ;
      RECT  99300.0 980400.0 98100.0 979200.0 ;
      RECT  96900.0 978450.0 95700.0 977250.0 ;
      RECT  96900.0 975750.0 98100.0 974550.0 ;
      RECT  101700.0 975750.0 102900.0 974550.0 ;
      RECT  101700.0 984450.0 102900.0 983250.0 ;
      RECT  101700.0 978450.0 102900.0 977250.0 ;
      RECT  95700.0 978450.0 96900.0 977250.0 ;
      RECT  98100.0 980400.0 99300.0 979200.0 ;
      RECT  100500.0 982350.0 101700.0 981150.0 ;
      RECT  101700.0 978450.0 102900.0 977250.0 ;
      RECT  92700.0 973050.0 108300.0 972150.0 ;
      RECT  92700.0 986850.0 108300.0 985950.0 ;
      RECT  94500.0 988350.0 95700.0 985950.0 ;
      RECT  94500.0 997050.0 95700.0 1000650.0 ;
      RECT  99300.0 997050.0 100500.0 1000650.0 ;
      RECT  104100.0 998250.0 105300.0 1000200.0 ;
      RECT  104100.0 986400.0 105300.0 988350.0 ;
      RECT  94500.0 997050.0 95700.0 998250.0 ;
      RECT  96900.0 997050.0 98100.0 998250.0 ;
      RECT  96900.0 997050.0 98100.0 998250.0 ;
      RECT  94500.0 997050.0 95700.0 998250.0 ;
      RECT  96900.0 997050.0 98100.0 998250.0 ;
      RECT  99300.0 997050.0 100500.0 998250.0 ;
      RECT  99300.0 997050.0 100500.0 998250.0 ;
      RECT  96900.0 997050.0 98100.0 998250.0 ;
      RECT  99300.0 997050.0 100500.0 998250.0 ;
      RECT  101700.0 997050.0 102900.0 998250.0 ;
      RECT  101700.0 997050.0 102900.0 998250.0 ;
      RECT  99300.0 997050.0 100500.0 998250.0 ;
      RECT  94500.0 988350.0 95700.0 989550.0 ;
      RECT  96900.0 988350.0 98100.0 989550.0 ;
      RECT  96900.0 988350.0 98100.0 989550.0 ;
      RECT  94500.0 988350.0 95700.0 989550.0 ;
      RECT  96900.0 988350.0 98100.0 989550.0 ;
      RECT  99300.0 988350.0 100500.0 989550.0 ;
      RECT  99300.0 988350.0 100500.0 989550.0 ;
      RECT  96900.0 988350.0 98100.0 989550.0 ;
      RECT  99300.0 988350.0 100500.0 989550.0 ;
      RECT  101700.0 988350.0 102900.0 989550.0 ;
      RECT  101700.0 988350.0 102900.0 989550.0 ;
      RECT  99300.0 988350.0 100500.0 989550.0 ;
      RECT  104100.0 997650.0 105300.0 998850.0 ;
      RECT  104100.0 987750.0 105300.0 988950.0 ;
      RECT  101700.0 990450.0 100500.0 991650.0 ;
      RECT  99300.0 992400.0 98100.0 993600.0 ;
      RECT  96900.0 994350.0 95700.0 995550.0 ;
      RECT  96900.0 997050.0 98100.0 998250.0 ;
      RECT  101700.0 997050.0 102900.0 998250.0 ;
      RECT  101700.0 988350.0 102900.0 989550.0 ;
      RECT  101700.0 994350.0 102900.0 995550.0 ;
      RECT  95700.0 994350.0 96900.0 995550.0 ;
      RECT  98100.0 992400.0 99300.0 993600.0 ;
      RECT  100500.0 990450.0 101700.0 991650.0 ;
      RECT  101700.0 994350.0 102900.0 995550.0 ;
      RECT  92700.0 999750.0 108300.0 1000650.0 ;
      RECT  92700.0 985950.0 108300.0 986850.0 ;
      RECT  94500.0 1012050.0 95700.0 1014450.0 ;
      RECT  94500.0 1003350.0 95700.0 999750.0 ;
      RECT  99300.0 1003350.0 100500.0 999750.0 ;
      RECT  104100.0 1002150.0 105300.0 1000200.0 ;
      RECT  104100.0 1014000.0 105300.0 1012050.0 ;
      RECT  94500.0 1003350.0 95700.0 1002150.0 ;
      RECT  96900.0 1003350.0 98100.0 1002150.0 ;
      RECT  96900.0 1003350.0 98100.0 1002150.0 ;
      RECT  94500.0 1003350.0 95700.0 1002150.0 ;
      RECT  96900.0 1003350.0 98100.0 1002150.0 ;
      RECT  99300.0 1003350.0 100500.0 1002150.0 ;
      RECT  99300.0 1003350.0 100500.0 1002150.0 ;
      RECT  96900.0 1003350.0 98100.0 1002150.0 ;
      RECT  99300.0 1003350.0 100500.0 1002150.0 ;
      RECT  101700.0 1003350.0 102900.0 1002150.0 ;
      RECT  101700.0 1003350.0 102900.0 1002150.0 ;
      RECT  99300.0 1003350.0 100500.0 1002150.0 ;
      RECT  94500.0 1012050.0 95700.0 1010850.0 ;
      RECT  96900.0 1012050.0 98100.0 1010850.0 ;
      RECT  96900.0 1012050.0 98100.0 1010850.0 ;
      RECT  94500.0 1012050.0 95700.0 1010850.0 ;
      RECT  96900.0 1012050.0 98100.0 1010850.0 ;
      RECT  99300.0 1012050.0 100500.0 1010850.0 ;
      RECT  99300.0 1012050.0 100500.0 1010850.0 ;
      RECT  96900.0 1012050.0 98100.0 1010850.0 ;
      RECT  99300.0 1012050.0 100500.0 1010850.0 ;
      RECT  101700.0 1012050.0 102900.0 1010850.0 ;
      RECT  101700.0 1012050.0 102900.0 1010850.0 ;
      RECT  99300.0 1012050.0 100500.0 1010850.0 ;
      RECT  104100.0 1002750.0 105300.0 1001550.0 ;
      RECT  104100.0 1012650.0 105300.0 1011450.0 ;
      RECT  101700.0 1009950.0 100500.0 1008750.0 ;
      RECT  99300.0 1008000.0 98100.0 1006800.0 ;
      RECT  96900.0 1006050.0 95700.0 1004850.0 ;
      RECT  96900.0 1003350.0 98100.0 1002150.0 ;
      RECT  101700.0 1003350.0 102900.0 1002150.0 ;
      RECT  101700.0 1012050.0 102900.0 1010850.0 ;
      RECT  101700.0 1006050.0 102900.0 1004850.0 ;
      RECT  95700.0 1006050.0 96900.0 1004850.0 ;
      RECT  98100.0 1008000.0 99300.0 1006800.0 ;
      RECT  100500.0 1009950.0 101700.0 1008750.0 ;
      RECT  101700.0 1006050.0 102900.0 1004850.0 ;
      RECT  92700.0 1000650.0 108300.0 999750.0 ;
      RECT  92700.0 1014450.0 108300.0 1013550.0 ;
      RECT  94500.0 1015950.0 95700.0 1013550.0 ;
      RECT  94500.0 1024650.0 95700.0 1028250.0 ;
      RECT  99300.0 1024650.0 100500.0 1028250.0 ;
      RECT  104100.0 1025850.0 105300.0 1027800.0 ;
      RECT  104100.0 1014000.0 105300.0 1015950.0 ;
      RECT  94500.0 1024650.0 95700.0 1025850.0 ;
      RECT  96900.0 1024650.0 98100.0 1025850.0 ;
      RECT  96900.0 1024650.0 98100.0 1025850.0 ;
      RECT  94500.0 1024650.0 95700.0 1025850.0 ;
      RECT  96900.0 1024650.0 98100.0 1025850.0 ;
      RECT  99300.0 1024650.0 100500.0 1025850.0 ;
      RECT  99300.0 1024650.0 100500.0 1025850.0 ;
      RECT  96900.0 1024650.0 98100.0 1025850.0 ;
      RECT  99300.0 1024650.0 100500.0 1025850.0 ;
      RECT  101700.0 1024650.0 102900.0 1025850.0 ;
      RECT  101700.0 1024650.0 102900.0 1025850.0 ;
      RECT  99300.0 1024650.0 100500.0 1025850.0 ;
      RECT  94500.0 1015950.0 95700.0 1017150.0 ;
      RECT  96900.0 1015950.0 98100.0 1017150.0 ;
      RECT  96900.0 1015950.0 98100.0 1017150.0 ;
      RECT  94500.0 1015950.0 95700.0 1017150.0 ;
      RECT  96900.0 1015950.0 98100.0 1017150.0 ;
      RECT  99300.0 1015950.0 100500.0 1017150.0 ;
      RECT  99300.0 1015950.0 100500.0 1017150.0 ;
      RECT  96900.0 1015950.0 98100.0 1017150.0 ;
      RECT  99300.0 1015950.0 100500.0 1017150.0 ;
      RECT  101700.0 1015950.0 102900.0 1017150.0 ;
      RECT  101700.0 1015950.0 102900.0 1017150.0 ;
      RECT  99300.0 1015950.0 100500.0 1017150.0 ;
      RECT  104100.0 1025250.0 105300.0 1026450.0 ;
      RECT  104100.0 1015350.0 105300.0 1016550.0 ;
      RECT  101700.0 1018050.0 100500.0 1019250.0 ;
      RECT  99300.0 1020000.0 98100.0 1021200.0 ;
      RECT  96900.0 1021950.0 95700.0 1023150.0 ;
      RECT  96900.0 1024650.0 98100.0 1025850.0 ;
      RECT  101700.0 1024650.0 102900.0 1025850.0 ;
      RECT  101700.0 1015950.0 102900.0 1017150.0 ;
      RECT  101700.0 1021950.0 102900.0 1023150.0 ;
      RECT  95700.0 1021950.0 96900.0 1023150.0 ;
      RECT  98100.0 1020000.0 99300.0 1021200.0 ;
      RECT  100500.0 1018050.0 101700.0 1019250.0 ;
      RECT  101700.0 1021950.0 102900.0 1023150.0 ;
      RECT  92700.0 1027350.0 108300.0 1028250.0 ;
      RECT  92700.0 1013550.0 108300.0 1014450.0 ;
      RECT  94500.0 1039650.0 95700.0 1042050.0 ;
      RECT  94500.0 1030950.0 95700.0 1027350.0 ;
      RECT  99300.0 1030950.0 100500.0 1027350.0 ;
      RECT  104100.0 1029750.0 105300.0 1027800.0 ;
      RECT  104100.0 1041600.0 105300.0 1039650.0 ;
      RECT  94500.0 1030950.0 95700.0 1029750.0 ;
      RECT  96900.0 1030950.0 98100.0 1029750.0 ;
      RECT  96900.0 1030950.0 98100.0 1029750.0 ;
      RECT  94500.0 1030950.0 95700.0 1029750.0 ;
      RECT  96900.0 1030950.0 98100.0 1029750.0 ;
      RECT  99300.0 1030950.0 100500.0 1029750.0 ;
      RECT  99300.0 1030950.0 100500.0 1029750.0 ;
      RECT  96900.0 1030950.0 98100.0 1029750.0 ;
      RECT  99300.0 1030950.0 100500.0 1029750.0 ;
      RECT  101700.0 1030950.0 102900.0 1029750.0 ;
      RECT  101700.0 1030950.0 102900.0 1029750.0 ;
      RECT  99300.0 1030950.0 100500.0 1029750.0 ;
      RECT  94500.0 1039650.0 95700.0 1038450.0 ;
      RECT  96900.0 1039650.0 98100.0 1038450.0 ;
      RECT  96900.0 1039650.0 98100.0 1038450.0 ;
      RECT  94500.0 1039650.0 95700.0 1038450.0 ;
      RECT  96900.0 1039650.0 98100.0 1038450.0 ;
      RECT  99300.0 1039650.0 100500.0 1038450.0 ;
      RECT  99300.0 1039650.0 100500.0 1038450.0 ;
      RECT  96900.0 1039650.0 98100.0 1038450.0 ;
      RECT  99300.0 1039650.0 100500.0 1038450.0 ;
      RECT  101700.0 1039650.0 102900.0 1038450.0 ;
      RECT  101700.0 1039650.0 102900.0 1038450.0 ;
      RECT  99300.0 1039650.0 100500.0 1038450.0 ;
      RECT  104100.0 1030350.0 105300.0 1029150.0 ;
      RECT  104100.0 1040250.0 105300.0 1039050.0 ;
      RECT  101700.0 1037550.0 100500.0 1036350.0 ;
      RECT  99300.0 1035600.0 98100.0 1034400.0 ;
      RECT  96900.0 1033650.0 95700.0 1032450.0 ;
      RECT  96900.0 1030950.0 98100.0 1029750.0 ;
      RECT  101700.0 1030950.0 102900.0 1029750.0 ;
      RECT  101700.0 1039650.0 102900.0 1038450.0 ;
      RECT  101700.0 1033650.0 102900.0 1032450.0 ;
      RECT  95700.0 1033650.0 96900.0 1032450.0 ;
      RECT  98100.0 1035600.0 99300.0 1034400.0 ;
      RECT  100500.0 1037550.0 101700.0 1036350.0 ;
      RECT  101700.0 1033650.0 102900.0 1032450.0 ;
      RECT  92700.0 1028250.0 108300.0 1027350.0 ;
      RECT  92700.0 1042050.0 108300.0 1041150.0 ;
      RECT  94500.0 1043550.0 95700.0 1041150.0 ;
      RECT  94500.0 1052250.0 95700.0 1055850.0 ;
      RECT  99300.0 1052250.0 100500.0 1055850.0 ;
      RECT  104100.0 1053450.0 105300.0 1055400.0 ;
      RECT  104100.0 1041600.0 105300.0 1043550.0 ;
      RECT  94500.0 1052250.0 95700.0 1053450.0 ;
      RECT  96900.0 1052250.0 98100.0 1053450.0 ;
      RECT  96900.0 1052250.0 98100.0 1053450.0 ;
      RECT  94500.0 1052250.0 95700.0 1053450.0 ;
      RECT  96900.0 1052250.0 98100.0 1053450.0 ;
      RECT  99300.0 1052250.0 100500.0 1053450.0 ;
      RECT  99300.0 1052250.0 100500.0 1053450.0 ;
      RECT  96900.0 1052250.0 98100.0 1053450.0 ;
      RECT  99300.0 1052250.0 100500.0 1053450.0 ;
      RECT  101700.0 1052250.0 102900.0 1053450.0 ;
      RECT  101700.0 1052250.0 102900.0 1053450.0 ;
      RECT  99300.0 1052250.0 100500.0 1053450.0 ;
      RECT  94500.0 1043550.0 95700.0 1044750.0 ;
      RECT  96900.0 1043550.0 98100.0 1044750.0 ;
      RECT  96900.0 1043550.0 98100.0 1044750.0 ;
      RECT  94500.0 1043550.0 95700.0 1044750.0 ;
      RECT  96900.0 1043550.0 98100.0 1044750.0 ;
      RECT  99300.0 1043550.0 100500.0 1044750.0 ;
      RECT  99300.0 1043550.0 100500.0 1044750.0 ;
      RECT  96900.0 1043550.0 98100.0 1044750.0 ;
      RECT  99300.0 1043550.0 100500.0 1044750.0 ;
      RECT  101700.0 1043550.0 102900.0 1044750.0 ;
      RECT  101700.0 1043550.0 102900.0 1044750.0 ;
      RECT  99300.0 1043550.0 100500.0 1044750.0 ;
      RECT  104100.0 1052850.0 105300.0 1054050.0 ;
      RECT  104100.0 1042950.0 105300.0 1044150.0 ;
      RECT  101700.0 1045650.0 100500.0 1046850.0 ;
      RECT  99300.0 1047600.0 98100.0 1048800.0 ;
      RECT  96900.0 1049550.0 95700.0 1050750.0 ;
      RECT  96900.0 1052250.0 98100.0 1053450.0 ;
      RECT  101700.0 1052250.0 102900.0 1053450.0 ;
      RECT  101700.0 1043550.0 102900.0 1044750.0 ;
      RECT  101700.0 1049550.0 102900.0 1050750.0 ;
      RECT  95700.0 1049550.0 96900.0 1050750.0 ;
      RECT  98100.0 1047600.0 99300.0 1048800.0 ;
      RECT  100500.0 1045650.0 101700.0 1046850.0 ;
      RECT  101700.0 1049550.0 102900.0 1050750.0 ;
      RECT  92700.0 1054950.0 108300.0 1055850.0 ;
      RECT  92700.0 1041150.0 108300.0 1042050.0 ;
      RECT  94500.0 1067250.0 95700.0 1069650.0 ;
      RECT  94500.0 1058550.0 95700.0 1054950.0 ;
      RECT  99300.0 1058550.0 100500.0 1054950.0 ;
      RECT  104100.0 1057350.0 105300.0 1055400.0 ;
      RECT  104100.0 1069200.0 105300.0 1067250.0 ;
      RECT  94500.0 1058550.0 95700.0 1057350.0 ;
      RECT  96900.0 1058550.0 98100.0 1057350.0 ;
      RECT  96900.0 1058550.0 98100.0 1057350.0 ;
      RECT  94500.0 1058550.0 95700.0 1057350.0 ;
      RECT  96900.0 1058550.0 98100.0 1057350.0 ;
      RECT  99300.0 1058550.0 100500.0 1057350.0 ;
      RECT  99300.0 1058550.0 100500.0 1057350.0 ;
      RECT  96900.0 1058550.0 98100.0 1057350.0 ;
      RECT  99300.0 1058550.0 100500.0 1057350.0 ;
      RECT  101700.0 1058550.0 102900.0 1057350.0 ;
      RECT  101700.0 1058550.0 102900.0 1057350.0 ;
      RECT  99300.0 1058550.0 100500.0 1057350.0 ;
      RECT  94500.0 1067250.0 95700.0 1066050.0 ;
      RECT  96900.0 1067250.0 98100.0 1066050.0 ;
      RECT  96900.0 1067250.0 98100.0 1066050.0 ;
      RECT  94500.0 1067250.0 95700.0 1066050.0 ;
      RECT  96900.0 1067250.0 98100.0 1066050.0 ;
      RECT  99300.0 1067250.0 100500.0 1066050.0 ;
      RECT  99300.0 1067250.0 100500.0 1066050.0 ;
      RECT  96900.0 1067250.0 98100.0 1066050.0 ;
      RECT  99300.0 1067250.0 100500.0 1066050.0 ;
      RECT  101700.0 1067250.0 102900.0 1066050.0 ;
      RECT  101700.0 1067250.0 102900.0 1066050.0 ;
      RECT  99300.0 1067250.0 100500.0 1066050.0 ;
      RECT  104100.0 1057950.0 105300.0 1056750.0 ;
      RECT  104100.0 1067850.0 105300.0 1066650.0 ;
      RECT  101700.0 1065150.0 100500.0 1063950.0 ;
      RECT  99300.0 1063200.0 98100.0 1062000.0 ;
      RECT  96900.0 1061250.0 95700.0 1060050.0 ;
      RECT  96900.0 1058550.0 98100.0 1057350.0 ;
      RECT  101700.0 1058550.0 102900.0 1057350.0 ;
      RECT  101700.0 1067250.0 102900.0 1066050.0 ;
      RECT  101700.0 1061250.0 102900.0 1060050.0 ;
      RECT  95700.0 1061250.0 96900.0 1060050.0 ;
      RECT  98100.0 1063200.0 99300.0 1062000.0 ;
      RECT  100500.0 1065150.0 101700.0 1063950.0 ;
      RECT  101700.0 1061250.0 102900.0 1060050.0 ;
      RECT  92700.0 1055850.0 108300.0 1054950.0 ;
      RECT  92700.0 1069650.0 108300.0 1068750.0 ;
      RECT  94500.0 1071150.0 95700.0 1068750.0 ;
      RECT  94500.0 1079850.0 95700.0 1083450.0 ;
      RECT  99300.0 1079850.0 100500.0 1083450.0 ;
      RECT  104100.0 1081050.0 105300.0 1083000.0 ;
      RECT  104100.0 1069200.0 105300.0 1071150.0 ;
      RECT  94500.0 1079850.0 95700.0 1081050.0 ;
      RECT  96900.0 1079850.0 98100.0 1081050.0 ;
      RECT  96900.0 1079850.0 98100.0 1081050.0 ;
      RECT  94500.0 1079850.0 95700.0 1081050.0 ;
      RECT  96900.0 1079850.0 98100.0 1081050.0 ;
      RECT  99300.0 1079850.0 100500.0 1081050.0 ;
      RECT  99300.0 1079850.0 100500.0 1081050.0 ;
      RECT  96900.0 1079850.0 98100.0 1081050.0 ;
      RECT  99300.0 1079850.0 100500.0 1081050.0 ;
      RECT  101700.0 1079850.0 102900.0 1081050.0 ;
      RECT  101700.0 1079850.0 102900.0 1081050.0 ;
      RECT  99300.0 1079850.0 100500.0 1081050.0 ;
      RECT  94500.0 1071150.0 95700.0 1072350.0 ;
      RECT  96900.0 1071150.0 98100.0 1072350.0 ;
      RECT  96900.0 1071150.0 98100.0 1072350.0 ;
      RECT  94500.0 1071150.0 95700.0 1072350.0 ;
      RECT  96900.0 1071150.0 98100.0 1072350.0 ;
      RECT  99300.0 1071150.0 100500.0 1072350.0 ;
      RECT  99300.0 1071150.0 100500.0 1072350.0 ;
      RECT  96900.0 1071150.0 98100.0 1072350.0 ;
      RECT  99300.0 1071150.0 100500.0 1072350.0 ;
      RECT  101700.0 1071150.0 102900.0 1072350.0 ;
      RECT  101700.0 1071150.0 102900.0 1072350.0 ;
      RECT  99300.0 1071150.0 100500.0 1072350.0 ;
      RECT  104100.0 1080450.0 105300.0 1081650.0 ;
      RECT  104100.0 1070550.0 105300.0 1071750.0 ;
      RECT  101700.0 1073250.0 100500.0 1074450.0 ;
      RECT  99300.0 1075200.0 98100.0 1076400.0 ;
      RECT  96900.0 1077150.0 95700.0 1078350.0 ;
      RECT  96900.0 1079850.0 98100.0 1081050.0 ;
      RECT  101700.0 1079850.0 102900.0 1081050.0 ;
      RECT  101700.0 1071150.0 102900.0 1072350.0 ;
      RECT  101700.0 1077150.0 102900.0 1078350.0 ;
      RECT  95700.0 1077150.0 96900.0 1078350.0 ;
      RECT  98100.0 1075200.0 99300.0 1076400.0 ;
      RECT  100500.0 1073250.0 101700.0 1074450.0 ;
      RECT  101700.0 1077150.0 102900.0 1078350.0 ;
      RECT  92700.0 1082550.0 108300.0 1083450.0 ;
      RECT  92700.0 1068750.0 108300.0 1069650.0 ;
      RECT  94500.0 1094850.0 95700.0 1097250.0 ;
      RECT  94500.0 1086150.0 95700.0 1082550.0 ;
      RECT  99300.0 1086150.0 100500.0 1082550.0 ;
      RECT  104100.0 1084950.0 105300.0 1083000.0 ;
      RECT  104100.0 1096800.0 105300.0 1094850.0 ;
      RECT  94500.0 1086150.0 95700.0 1084950.0 ;
      RECT  96900.0 1086150.0 98100.0 1084950.0 ;
      RECT  96900.0 1086150.0 98100.0 1084950.0 ;
      RECT  94500.0 1086150.0 95700.0 1084950.0 ;
      RECT  96900.0 1086150.0 98100.0 1084950.0 ;
      RECT  99300.0 1086150.0 100500.0 1084950.0 ;
      RECT  99300.0 1086150.0 100500.0 1084950.0 ;
      RECT  96900.0 1086150.0 98100.0 1084950.0 ;
      RECT  99300.0 1086150.0 100500.0 1084950.0 ;
      RECT  101700.0 1086150.0 102900.0 1084950.0 ;
      RECT  101700.0 1086150.0 102900.0 1084950.0 ;
      RECT  99300.0 1086150.0 100500.0 1084950.0 ;
      RECT  94500.0 1094850.0 95700.0 1093650.0 ;
      RECT  96900.0 1094850.0 98100.0 1093650.0 ;
      RECT  96900.0 1094850.0 98100.0 1093650.0 ;
      RECT  94500.0 1094850.0 95700.0 1093650.0 ;
      RECT  96900.0 1094850.0 98100.0 1093650.0 ;
      RECT  99300.0 1094850.0 100500.0 1093650.0 ;
      RECT  99300.0 1094850.0 100500.0 1093650.0 ;
      RECT  96900.0 1094850.0 98100.0 1093650.0 ;
      RECT  99300.0 1094850.0 100500.0 1093650.0 ;
      RECT  101700.0 1094850.0 102900.0 1093650.0 ;
      RECT  101700.0 1094850.0 102900.0 1093650.0 ;
      RECT  99300.0 1094850.0 100500.0 1093650.0 ;
      RECT  104100.0 1085550.0 105300.0 1084350.0 ;
      RECT  104100.0 1095450.0 105300.0 1094250.0 ;
      RECT  101700.0 1092750.0 100500.0 1091550.0 ;
      RECT  99300.0 1090800.0 98100.0 1089600.0 ;
      RECT  96900.0 1088850.0 95700.0 1087650.0 ;
      RECT  96900.0 1086150.0 98100.0 1084950.0 ;
      RECT  101700.0 1086150.0 102900.0 1084950.0 ;
      RECT  101700.0 1094850.0 102900.0 1093650.0 ;
      RECT  101700.0 1088850.0 102900.0 1087650.0 ;
      RECT  95700.0 1088850.0 96900.0 1087650.0 ;
      RECT  98100.0 1090800.0 99300.0 1089600.0 ;
      RECT  100500.0 1092750.0 101700.0 1091550.0 ;
      RECT  101700.0 1088850.0 102900.0 1087650.0 ;
      RECT  92700.0 1083450.0 108300.0 1082550.0 ;
      RECT  92700.0 1097250.0 108300.0 1096350.0 ;
      RECT  94500.0 1098750.0 95700.0 1096350.0 ;
      RECT  94500.0 1107450.0 95700.0 1111050.0 ;
      RECT  99300.0 1107450.0 100500.0 1111050.0 ;
      RECT  104100.0 1108650.0 105300.0 1110600.0 ;
      RECT  104100.0 1096800.0 105300.0 1098750.0 ;
      RECT  94500.0 1107450.0 95700.0 1108650.0 ;
      RECT  96900.0 1107450.0 98100.0 1108650.0 ;
      RECT  96900.0 1107450.0 98100.0 1108650.0 ;
      RECT  94500.0 1107450.0 95700.0 1108650.0 ;
      RECT  96900.0 1107450.0 98100.0 1108650.0 ;
      RECT  99300.0 1107450.0 100500.0 1108650.0 ;
      RECT  99300.0 1107450.0 100500.0 1108650.0 ;
      RECT  96900.0 1107450.0 98100.0 1108650.0 ;
      RECT  99300.0 1107450.0 100500.0 1108650.0 ;
      RECT  101700.0 1107450.0 102900.0 1108650.0 ;
      RECT  101700.0 1107450.0 102900.0 1108650.0 ;
      RECT  99300.0 1107450.0 100500.0 1108650.0 ;
      RECT  94500.0 1098750.0 95700.0 1099950.0 ;
      RECT  96900.0 1098750.0 98100.0 1099950.0 ;
      RECT  96900.0 1098750.0 98100.0 1099950.0 ;
      RECT  94500.0 1098750.0 95700.0 1099950.0 ;
      RECT  96900.0 1098750.0 98100.0 1099950.0 ;
      RECT  99300.0 1098750.0 100500.0 1099950.0 ;
      RECT  99300.0 1098750.0 100500.0 1099950.0 ;
      RECT  96900.0 1098750.0 98100.0 1099950.0 ;
      RECT  99300.0 1098750.0 100500.0 1099950.0 ;
      RECT  101700.0 1098750.0 102900.0 1099950.0 ;
      RECT  101700.0 1098750.0 102900.0 1099950.0 ;
      RECT  99300.0 1098750.0 100500.0 1099950.0 ;
      RECT  104100.0 1108050.0 105300.0 1109250.0 ;
      RECT  104100.0 1098150.0 105300.0 1099350.0 ;
      RECT  101700.0 1100850.0 100500.0 1102050.0 ;
      RECT  99300.0 1102800.0 98100.0 1104000.0 ;
      RECT  96900.0 1104750.0 95700.0 1105950.0 ;
      RECT  96900.0 1107450.0 98100.0 1108650.0 ;
      RECT  101700.0 1107450.0 102900.0 1108650.0 ;
      RECT  101700.0 1098750.0 102900.0 1099950.0 ;
      RECT  101700.0 1104750.0 102900.0 1105950.0 ;
      RECT  95700.0 1104750.0 96900.0 1105950.0 ;
      RECT  98100.0 1102800.0 99300.0 1104000.0 ;
      RECT  100500.0 1100850.0 101700.0 1102050.0 ;
      RECT  101700.0 1104750.0 102900.0 1105950.0 ;
      RECT  92700.0 1110150.0 108300.0 1111050.0 ;
      RECT  92700.0 1096350.0 108300.0 1097250.0 ;
      RECT  94500.0 1122450.0 95700.0 1124850.0 ;
      RECT  94500.0 1113750.0 95700.0 1110150.0 ;
      RECT  99300.0 1113750.0 100500.0 1110150.0 ;
      RECT  104100.0 1112550.0 105300.0 1110600.0 ;
      RECT  104100.0 1124400.0 105300.0 1122450.0 ;
      RECT  94500.0 1113750.0 95700.0 1112550.0 ;
      RECT  96900.0 1113750.0 98100.0 1112550.0 ;
      RECT  96900.0 1113750.0 98100.0 1112550.0 ;
      RECT  94500.0 1113750.0 95700.0 1112550.0 ;
      RECT  96900.0 1113750.0 98100.0 1112550.0 ;
      RECT  99300.0 1113750.0 100500.0 1112550.0 ;
      RECT  99300.0 1113750.0 100500.0 1112550.0 ;
      RECT  96900.0 1113750.0 98100.0 1112550.0 ;
      RECT  99300.0 1113750.0 100500.0 1112550.0 ;
      RECT  101700.0 1113750.0 102900.0 1112550.0 ;
      RECT  101700.0 1113750.0 102900.0 1112550.0 ;
      RECT  99300.0 1113750.0 100500.0 1112550.0 ;
      RECT  94500.0 1122450.0 95700.0 1121250.0 ;
      RECT  96900.0 1122450.0 98100.0 1121250.0 ;
      RECT  96900.0 1122450.0 98100.0 1121250.0 ;
      RECT  94500.0 1122450.0 95700.0 1121250.0 ;
      RECT  96900.0 1122450.0 98100.0 1121250.0 ;
      RECT  99300.0 1122450.0 100500.0 1121250.0 ;
      RECT  99300.0 1122450.0 100500.0 1121250.0 ;
      RECT  96900.0 1122450.0 98100.0 1121250.0 ;
      RECT  99300.0 1122450.0 100500.0 1121250.0 ;
      RECT  101700.0 1122450.0 102900.0 1121250.0 ;
      RECT  101700.0 1122450.0 102900.0 1121250.0 ;
      RECT  99300.0 1122450.0 100500.0 1121250.0 ;
      RECT  104100.0 1113150.0 105300.0 1111950.0 ;
      RECT  104100.0 1123050.0 105300.0 1121850.0 ;
      RECT  101700.0 1120350.0 100500.0 1119150.0 ;
      RECT  99300.0 1118400.0 98100.0 1117200.0 ;
      RECT  96900.0 1116450.0 95700.0 1115250.0 ;
      RECT  96900.0 1113750.0 98100.0 1112550.0 ;
      RECT  101700.0 1113750.0 102900.0 1112550.0 ;
      RECT  101700.0 1122450.0 102900.0 1121250.0 ;
      RECT  101700.0 1116450.0 102900.0 1115250.0 ;
      RECT  95700.0 1116450.0 96900.0 1115250.0 ;
      RECT  98100.0 1118400.0 99300.0 1117200.0 ;
      RECT  100500.0 1120350.0 101700.0 1119150.0 ;
      RECT  101700.0 1116450.0 102900.0 1115250.0 ;
      RECT  92700.0 1111050.0 108300.0 1110150.0 ;
      RECT  92700.0 1124850.0 108300.0 1123950.0 ;
      RECT  94500.0 1126350.0 95700.0 1123950.0 ;
      RECT  94500.0 1135050.0 95700.0 1138650.0 ;
      RECT  99300.0 1135050.0 100500.0 1138650.0 ;
      RECT  104100.0 1136250.0 105300.0 1138200.0 ;
      RECT  104100.0 1124400.0 105300.0 1126350.0 ;
      RECT  94500.0 1135050.0 95700.0 1136250.0 ;
      RECT  96900.0 1135050.0 98100.0 1136250.0 ;
      RECT  96900.0 1135050.0 98100.0 1136250.0 ;
      RECT  94500.0 1135050.0 95700.0 1136250.0 ;
      RECT  96900.0 1135050.0 98100.0 1136250.0 ;
      RECT  99300.0 1135050.0 100500.0 1136250.0 ;
      RECT  99300.0 1135050.0 100500.0 1136250.0 ;
      RECT  96900.0 1135050.0 98100.0 1136250.0 ;
      RECT  99300.0 1135050.0 100500.0 1136250.0 ;
      RECT  101700.0 1135050.0 102900.0 1136250.0 ;
      RECT  101700.0 1135050.0 102900.0 1136250.0 ;
      RECT  99300.0 1135050.0 100500.0 1136250.0 ;
      RECT  94500.0 1126350.0 95700.0 1127550.0 ;
      RECT  96900.0 1126350.0 98100.0 1127550.0 ;
      RECT  96900.0 1126350.0 98100.0 1127550.0 ;
      RECT  94500.0 1126350.0 95700.0 1127550.0 ;
      RECT  96900.0 1126350.0 98100.0 1127550.0 ;
      RECT  99300.0 1126350.0 100500.0 1127550.0 ;
      RECT  99300.0 1126350.0 100500.0 1127550.0 ;
      RECT  96900.0 1126350.0 98100.0 1127550.0 ;
      RECT  99300.0 1126350.0 100500.0 1127550.0 ;
      RECT  101700.0 1126350.0 102900.0 1127550.0 ;
      RECT  101700.0 1126350.0 102900.0 1127550.0 ;
      RECT  99300.0 1126350.0 100500.0 1127550.0 ;
      RECT  104100.0 1135650.0 105300.0 1136850.0 ;
      RECT  104100.0 1125750.0 105300.0 1126950.0 ;
      RECT  101700.0 1128450.0 100500.0 1129650.0 ;
      RECT  99300.0 1130400.0 98100.0 1131600.0 ;
      RECT  96900.0 1132350.0 95700.0 1133550.0 ;
      RECT  96900.0 1135050.0 98100.0 1136250.0 ;
      RECT  101700.0 1135050.0 102900.0 1136250.0 ;
      RECT  101700.0 1126350.0 102900.0 1127550.0 ;
      RECT  101700.0 1132350.0 102900.0 1133550.0 ;
      RECT  95700.0 1132350.0 96900.0 1133550.0 ;
      RECT  98100.0 1130400.0 99300.0 1131600.0 ;
      RECT  100500.0 1128450.0 101700.0 1129650.0 ;
      RECT  101700.0 1132350.0 102900.0 1133550.0 ;
      RECT  92700.0 1137750.0 108300.0 1138650.0 ;
      RECT  92700.0 1123950.0 108300.0 1124850.0 ;
      RECT  94500.0 1150050.0 95700.0 1152450.0 ;
      RECT  94500.0 1141350.0 95700.0 1137750.0 ;
      RECT  99300.0 1141350.0 100500.0 1137750.0 ;
      RECT  104100.0 1140150.0 105300.0 1138200.0 ;
      RECT  104100.0 1152000.0 105300.0 1150050.0 ;
      RECT  94500.0 1141350.0 95700.0 1140150.0 ;
      RECT  96900.0 1141350.0 98100.0 1140150.0 ;
      RECT  96900.0 1141350.0 98100.0 1140150.0 ;
      RECT  94500.0 1141350.0 95700.0 1140150.0 ;
      RECT  96900.0 1141350.0 98100.0 1140150.0 ;
      RECT  99300.0 1141350.0 100500.0 1140150.0 ;
      RECT  99300.0 1141350.0 100500.0 1140150.0 ;
      RECT  96900.0 1141350.0 98100.0 1140150.0 ;
      RECT  99300.0 1141350.0 100500.0 1140150.0 ;
      RECT  101700.0 1141350.0 102900.0 1140150.0 ;
      RECT  101700.0 1141350.0 102900.0 1140150.0 ;
      RECT  99300.0 1141350.0 100500.0 1140150.0 ;
      RECT  94500.0 1150050.0 95700.0 1148850.0 ;
      RECT  96900.0 1150050.0 98100.0 1148850.0 ;
      RECT  96900.0 1150050.0 98100.0 1148850.0 ;
      RECT  94500.0 1150050.0 95700.0 1148850.0 ;
      RECT  96900.0 1150050.0 98100.0 1148850.0 ;
      RECT  99300.0 1150050.0 100500.0 1148850.0 ;
      RECT  99300.0 1150050.0 100500.0 1148850.0 ;
      RECT  96900.0 1150050.0 98100.0 1148850.0 ;
      RECT  99300.0 1150050.0 100500.0 1148850.0 ;
      RECT  101700.0 1150050.0 102900.0 1148850.0 ;
      RECT  101700.0 1150050.0 102900.0 1148850.0 ;
      RECT  99300.0 1150050.0 100500.0 1148850.0 ;
      RECT  104100.0 1140750.0 105300.0 1139550.0 ;
      RECT  104100.0 1150650.0 105300.0 1149450.0 ;
      RECT  101700.0 1147950.0 100500.0 1146750.0 ;
      RECT  99300.0 1146000.0 98100.0 1144800.0 ;
      RECT  96900.0 1144050.0 95700.0 1142850.0 ;
      RECT  96900.0 1141350.0 98100.0 1140150.0 ;
      RECT  101700.0 1141350.0 102900.0 1140150.0 ;
      RECT  101700.0 1150050.0 102900.0 1148850.0 ;
      RECT  101700.0 1144050.0 102900.0 1142850.0 ;
      RECT  95700.0 1144050.0 96900.0 1142850.0 ;
      RECT  98100.0 1146000.0 99300.0 1144800.0 ;
      RECT  100500.0 1147950.0 101700.0 1146750.0 ;
      RECT  101700.0 1144050.0 102900.0 1142850.0 ;
      RECT  92700.0 1138650.0 108300.0 1137750.0 ;
      RECT  92700.0 1152450.0 108300.0 1151550.0 ;
      RECT  94500.0 1153950.0 95700.0 1151550.0 ;
      RECT  94500.0 1162650.0 95700.0 1166250.0 ;
      RECT  99300.0 1162650.0 100500.0 1166250.0 ;
      RECT  104100.0 1163850.0 105300.0 1165800.0 ;
      RECT  104100.0 1152000.0 105300.0 1153950.0 ;
      RECT  94500.0 1162650.0 95700.0 1163850.0 ;
      RECT  96900.0 1162650.0 98100.0 1163850.0 ;
      RECT  96900.0 1162650.0 98100.0 1163850.0 ;
      RECT  94500.0 1162650.0 95700.0 1163850.0 ;
      RECT  96900.0 1162650.0 98100.0 1163850.0 ;
      RECT  99300.0 1162650.0 100500.0 1163850.0 ;
      RECT  99300.0 1162650.0 100500.0 1163850.0 ;
      RECT  96900.0 1162650.0 98100.0 1163850.0 ;
      RECT  99300.0 1162650.0 100500.0 1163850.0 ;
      RECT  101700.0 1162650.0 102900.0 1163850.0 ;
      RECT  101700.0 1162650.0 102900.0 1163850.0 ;
      RECT  99300.0 1162650.0 100500.0 1163850.0 ;
      RECT  94500.0 1153950.0 95700.0 1155150.0 ;
      RECT  96900.0 1153950.0 98100.0 1155150.0 ;
      RECT  96900.0 1153950.0 98100.0 1155150.0 ;
      RECT  94500.0 1153950.0 95700.0 1155150.0 ;
      RECT  96900.0 1153950.0 98100.0 1155150.0 ;
      RECT  99300.0 1153950.0 100500.0 1155150.0 ;
      RECT  99300.0 1153950.0 100500.0 1155150.0 ;
      RECT  96900.0 1153950.0 98100.0 1155150.0 ;
      RECT  99300.0 1153950.0 100500.0 1155150.0 ;
      RECT  101700.0 1153950.0 102900.0 1155150.0 ;
      RECT  101700.0 1153950.0 102900.0 1155150.0 ;
      RECT  99300.0 1153950.0 100500.0 1155150.0 ;
      RECT  104100.0 1163250.0 105300.0 1164450.0 ;
      RECT  104100.0 1153350.0 105300.0 1154550.0 ;
      RECT  101700.0 1156050.0 100500.0 1157250.0 ;
      RECT  99300.0 1158000.0 98100.0 1159200.0 ;
      RECT  96900.0 1159950.0 95700.0 1161150.0 ;
      RECT  96900.0 1162650.0 98100.0 1163850.0 ;
      RECT  101700.0 1162650.0 102900.0 1163850.0 ;
      RECT  101700.0 1153950.0 102900.0 1155150.0 ;
      RECT  101700.0 1159950.0 102900.0 1161150.0 ;
      RECT  95700.0 1159950.0 96900.0 1161150.0 ;
      RECT  98100.0 1158000.0 99300.0 1159200.0 ;
      RECT  100500.0 1156050.0 101700.0 1157250.0 ;
      RECT  101700.0 1159950.0 102900.0 1161150.0 ;
      RECT  92700.0 1165350.0 108300.0 1166250.0 ;
      RECT  92700.0 1151550.0 108300.0 1152450.0 ;
      RECT  94500.0 1177650.0 95700.0 1180050.0 ;
      RECT  94500.0 1168950.0 95700.0 1165350.0 ;
      RECT  99300.0 1168950.0 100500.0 1165350.0 ;
      RECT  104100.0 1167750.0 105300.0 1165800.0 ;
      RECT  104100.0 1179600.0 105300.0 1177650.0 ;
      RECT  94500.0 1168950.0 95700.0 1167750.0 ;
      RECT  96900.0 1168950.0 98100.0 1167750.0 ;
      RECT  96900.0 1168950.0 98100.0 1167750.0 ;
      RECT  94500.0 1168950.0 95700.0 1167750.0 ;
      RECT  96900.0 1168950.0 98100.0 1167750.0 ;
      RECT  99300.0 1168950.0 100500.0 1167750.0 ;
      RECT  99300.0 1168950.0 100500.0 1167750.0 ;
      RECT  96900.0 1168950.0 98100.0 1167750.0 ;
      RECT  99300.0 1168950.0 100500.0 1167750.0 ;
      RECT  101700.0 1168950.0 102900.0 1167750.0 ;
      RECT  101700.0 1168950.0 102900.0 1167750.0 ;
      RECT  99300.0 1168950.0 100500.0 1167750.0 ;
      RECT  94500.0 1177650.0 95700.0 1176450.0 ;
      RECT  96900.0 1177650.0 98100.0 1176450.0 ;
      RECT  96900.0 1177650.0 98100.0 1176450.0 ;
      RECT  94500.0 1177650.0 95700.0 1176450.0 ;
      RECT  96900.0 1177650.0 98100.0 1176450.0 ;
      RECT  99300.0 1177650.0 100500.0 1176450.0 ;
      RECT  99300.0 1177650.0 100500.0 1176450.0 ;
      RECT  96900.0 1177650.0 98100.0 1176450.0 ;
      RECT  99300.0 1177650.0 100500.0 1176450.0 ;
      RECT  101700.0 1177650.0 102900.0 1176450.0 ;
      RECT  101700.0 1177650.0 102900.0 1176450.0 ;
      RECT  99300.0 1177650.0 100500.0 1176450.0 ;
      RECT  104100.0 1168350.0 105300.0 1167150.0 ;
      RECT  104100.0 1178250.0 105300.0 1177050.0 ;
      RECT  101700.0 1175550.0 100500.0 1174350.0 ;
      RECT  99300.0 1173600.0 98100.0 1172400.0 ;
      RECT  96900.0 1171650.0 95700.0 1170450.0 ;
      RECT  96900.0 1168950.0 98100.0 1167750.0 ;
      RECT  101700.0 1168950.0 102900.0 1167750.0 ;
      RECT  101700.0 1177650.0 102900.0 1176450.0 ;
      RECT  101700.0 1171650.0 102900.0 1170450.0 ;
      RECT  95700.0 1171650.0 96900.0 1170450.0 ;
      RECT  98100.0 1173600.0 99300.0 1172400.0 ;
      RECT  100500.0 1175550.0 101700.0 1174350.0 ;
      RECT  101700.0 1171650.0 102900.0 1170450.0 ;
      RECT  92700.0 1166250.0 108300.0 1165350.0 ;
      RECT  92700.0 1180050.0 108300.0 1179150.0 ;
      RECT  94500.0 1181550.0 95700.0 1179150.0 ;
      RECT  94500.0 1190250.0 95700.0 1193850.0 ;
      RECT  99300.0 1190250.0 100500.0 1193850.0 ;
      RECT  104100.0 1191450.0 105300.0 1193400.0 ;
      RECT  104100.0 1179600.0 105300.0 1181550.0 ;
      RECT  94500.0 1190250.0 95700.0 1191450.0 ;
      RECT  96900.0 1190250.0 98100.0 1191450.0 ;
      RECT  96900.0 1190250.0 98100.0 1191450.0 ;
      RECT  94500.0 1190250.0 95700.0 1191450.0 ;
      RECT  96900.0 1190250.0 98100.0 1191450.0 ;
      RECT  99300.0 1190250.0 100500.0 1191450.0 ;
      RECT  99300.0 1190250.0 100500.0 1191450.0 ;
      RECT  96900.0 1190250.0 98100.0 1191450.0 ;
      RECT  99300.0 1190250.0 100500.0 1191450.0 ;
      RECT  101700.0 1190250.0 102900.0 1191450.0 ;
      RECT  101700.0 1190250.0 102900.0 1191450.0 ;
      RECT  99300.0 1190250.0 100500.0 1191450.0 ;
      RECT  94500.0 1181550.0 95700.0 1182750.0 ;
      RECT  96900.0 1181550.0 98100.0 1182750.0 ;
      RECT  96900.0 1181550.0 98100.0 1182750.0 ;
      RECT  94500.0 1181550.0 95700.0 1182750.0 ;
      RECT  96900.0 1181550.0 98100.0 1182750.0 ;
      RECT  99300.0 1181550.0 100500.0 1182750.0 ;
      RECT  99300.0 1181550.0 100500.0 1182750.0 ;
      RECT  96900.0 1181550.0 98100.0 1182750.0 ;
      RECT  99300.0 1181550.0 100500.0 1182750.0 ;
      RECT  101700.0 1181550.0 102900.0 1182750.0 ;
      RECT  101700.0 1181550.0 102900.0 1182750.0 ;
      RECT  99300.0 1181550.0 100500.0 1182750.0 ;
      RECT  104100.0 1190850.0 105300.0 1192050.0 ;
      RECT  104100.0 1180950.0 105300.0 1182150.0 ;
      RECT  101700.0 1183650.0 100500.0 1184850.0 ;
      RECT  99300.0 1185600.0 98100.0 1186800.0 ;
      RECT  96900.0 1187550.0 95700.0 1188750.0 ;
      RECT  96900.0 1190250.0 98100.0 1191450.0 ;
      RECT  101700.0 1190250.0 102900.0 1191450.0 ;
      RECT  101700.0 1181550.0 102900.0 1182750.0 ;
      RECT  101700.0 1187550.0 102900.0 1188750.0 ;
      RECT  95700.0 1187550.0 96900.0 1188750.0 ;
      RECT  98100.0 1185600.0 99300.0 1186800.0 ;
      RECT  100500.0 1183650.0 101700.0 1184850.0 ;
      RECT  101700.0 1187550.0 102900.0 1188750.0 ;
      RECT  92700.0 1192950.0 108300.0 1193850.0 ;
      RECT  92700.0 1179150.0 108300.0 1180050.0 ;
      RECT  94500.0 1205250.0 95700.0 1207650.0 ;
      RECT  94500.0 1196550.0 95700.0 1192950.0 ;
      RECT  99300.0 1196550.0 100500.0 1192950.0 ;
      RECT  104100.0 1195350.0 105300.0 1193400.0 ;
      RECT  104100.0 1207200.0 105300.0 1205250.0 ;
      RECT  94500.0 1196550.0 95700.0 1195350.0 ;
      RECT  96900.0 1196550.0 98100.0 1195350.0 ;
      RECT  96900.0 1196550.0 98100.0 1195350.0 ;
      RECT  94500.0 1196550.0 95700.0 1195350.0 ;
      RECT  96900.0 1196550.0 98100.0 1195350.0 ;
      RECT  99300.0 1196550.0 100500.0 1195350.0 ;
      RECT  99300.0 1196550.0 100500.0 1195350.0 ;
      RECT  96900.0 1196550.0 98100.0 1195350.0 ;
      RECT  99300.0 1196550.0 100500.0 1195350.0 ;
      RECT  101700.0 1196550.0 102900.0 1195350.0 ;
      RECT  101700.0 1196550.0 102900.0 1195350.0 ;
      RECT  99300.0 1196550.0 100500.0 1195350.0 ;
      RECT  94500.0 1205250.0 95700.0 1204050.0 ;
      RECT  96900.0 1205250.0 98100.0 1204050.0 ;
      RECT  96900.0 1205250.0 98100.0 1204050.0 ;
      RECT  94500.0 1205250.0 95700.0 1204050.0 ;
      RECT  96900.0 1205250.0 98100.0 1204050.0 ;
      RECT  99300.0 1205250.0 100500.0 1204050.0 ;
      RECT  99300.0 1205250.0 100500.0 1204050.0 ;
      RECT  96900.0 1205250.0 98100.0 1204050.0 ;
      RECT  99300.0 1205250.0 100500.0 1204050.0 ;
      RECT  101700.0 1205250.0 102900.0 1204050.0 ;
      RECT  101700.0 1205250.0 102900.0 1204050.0 ;
      RECT  99300.0 1205250.0 100500.0 1204050.0 ;
      RECT  104100.0 1195950.0 105300.0 1194750.0 ;
      RECT  104100.0 1205850.0 105300.0 1204650.0 ;
      RECT  101700.0 1203150.0 100500.0 1201950.0 ;
      RECT  99300.0 1201200.0 98100.0 1200000.0 ;
      RECT  96900.0 1199250.0 95700.0 1198050.0 ;
      RECT  96900.0 1196550.0 98100.0 1195350.0 ;
      RECT  101700.0 1196550.0 102900.0 1195350.0 ;
      RECT  101700.0 1205250.0 102900.0 1204050.0 ;
      RECT  101700.0 1199250.0 102900.0 1198050.0 ;
      RECT  95700.0 1199250.0 96900.0 1198050.0 ;
      RECT  98100.0 1201200.0 99300.0 1200000.0 ;
      RECT  100500.0 1203150.0 101700.0 1201950.0 ;
      RECT  101700.0 1199250.0 102900.0 1198050.0 ;
      RECT  92700.0 1193850.0 108300.0 1192950.0 ;
      RECT  92700.0 1207650.0 108300.0 1206750.0 ;
      RECT  94500.0 1209150.0 95700.0 1206750.0 ;
      RECT  94500.0 1217850.0 95700.0 1221450.0 ;
      RECT  99300.0 1217850.0 100500.0 1221450.0 ;
      RECT  104100.0 1219050.0 105300.0 1221000.0 ;
      RECT  104100.0 1207200.0 105300.0 1209150.0 ;
      RECT  94500.0 1217850.0 95700.0 1219050.0 ;
      RECT  96900.0 1217850.0 98100.0 1219050.0 ;
      RECT  96900.0 1217850.0 98100.0 1219050.0 ;
      RECT  94500.0 1217850.0 95700.0 1219050.0 ;
      RECT  96900.0 1217850.0 98100.0 1219050.0 ;
      RECT  99300.0 1217850.0 100500.0 1219050.0 ;
      RECT  99300.0 1217850.0 100500.0 1219050.0 ;
      RECT  96900.0 1217850.0 98100.0 1219050.0 ;
      RECT  99300.0 1217850.0 100500.0 1219050.0 ;
      RECT  101700.0 1217850.0 102900.0 1219050.0 ;
      RECT  101700.0 1217850.0 102900.0 1219050.0 ;
      RECT  99300.0 1217850.0 100500.0 1219050.0 ;
      RECT  94500.0 1209150.0 95700.0 1210350.0 ;
      RECT  96900.0 1209150.0 98100.0 1210350.0 ;
      RECT  96900.0 1209150.0 98100.0 1210350.0 ;
      RECT  94500.0 1209150.0 95700.0 1210350.0 ;
      RECT  96900.0 1209150.0 98100.0 1210350.0 ;
      RECT  99300.0 1209150.0 100500.0 1210350.0 ;
      RECT  99300.0 1209150.0 100500.0 1210350.0 ;
      RECT  96900.0 1209150.0 98100.0 1210350.0 ;
      RECT  99300.0 1209150.0 100500.0 1210350.0 ;
      RECT  101700.0 1209150.0 102900.0 1210350.0 ;
      RECT  101700.0 1209150.0 102900.0 1210350.0 ;
      RECT  99300.0 1209150.0 100500.0 1210350.0 ;
      RECT  104100.0 1218450.0 105300.0 1219650.0 ;
      RECT  104100.0 1208550.0 105300.0 1209750.0 ;
      RECT  101700.0 1211250.0 100500.0 1212450.0 ;
      RECT  99300.0 1213200.0 98100.0 1214400.0 ;
      RECT  96900.0 1215150.0 95700.0 1216350.0 ;
      RECT  96900.0 1217850.0 98100.0 1219050.0 ;
      RECT  101700.0 1217850.0 102900.0 1219050.0 ;
      RECT  101700.0 1209150.0 102900.0 1210350.0 ;
      RECT  101700.0 1215150.0 102900.0 1216350.0 ;
      RECT  95700.0 1215150.0 96900.0 1216350.0 ;
      RECT  98100.0 1213200.0 99300.0 1214400.0 ;
      RECT  100500.0 1211250.0 101700.0 1212450.0 ;
      RECT  101700.0 1215150.0 102900.0 1216350.0 ;
      RECT  92700.0 1220550.0 108300.0 1221450.0 ;
      RECT  92700.0 1206750.0 108300.0 1207650.0 ;
      RECT  94500.0 1232850.0 95700.0 1235250.0 ;
      RECT  94500.0 1224150.0 95700.0 1220550.0 ;
      RECT  99300.0 1224150.0 100500.0 1220550.0 ;
      RECT  104100.0 1222950.0 105300.0 1221000.0 ;
      RECT  104100.0 1234800.0 105300.0 1232850.0 ;
      RECT  94500.0 1224150.0 95700.0 1222950.0 ;
      RECT  96900.0 1224150.0 98100.0 1222950.0 ;
      RECT  96900.0 1224150.0 98100.0 1222950.0 ;
      RECT  94500.0 1224150.0 95700.0 1222950.0 ;
      RECT  96900.0 1224150.0 98100.0 1222950.0 ;
      RECT  99300.0 1224150.0 100500.0 1222950.0 ;
      RECT  99300.0 1224150.0 100500.0 1222950.0 ;
      RECT  96900.0 1224150.0 98100.0 1222950.0 ;
      RECT  99300.0 1224150.0 100500.0 1222950.0 ;
      RECT  101700.0 1224150.0 102900.0 1222950.0 ;
      RECT  101700.0 1224150.0 102900.0 1222950.0 ;
      RECT  99300.0 1224150.0 100500.0 1222950.0 ;
      RECT  94500.0 1232850.0 95700.0 1231650.0 ;
      RECT  96900.0 1232850.0 98100.0 1231650.0 ;
      RECT  96900.0 1232850.0 98100.0 1231650.0 ;
      RECT  94500.0 1232850.0 95700.0 1231650.0 ;
      RECT  96900.0 1232850.0 98100.0 1231650.0 ;
      RECT  99300.0 1232850.0 100500.0 1231650.0 ;
      RECT  99300.0 1232850.0 100500.0 1231650.0 ;
      RECT  96900.0 1232850.0 98100.0 1231650.0 ;
      RECT  99300.0 1232850.0 100500.0 1231650.0 ;
      RECT  101700.0 1232850.0 102900.0 1231650.0 ;
      RECT  101700.0 1232850.0 102900.0 1231650.0 ;
      RECT  99300.0 1232850.0 100500.0 1231650.0 ;
      RECT  104100.0 1223550.0 105300.0 1222350.0 ;
      RECT  104100.0 1233450.0 105300.0 1232250.0 ;
      RECT  101700.0 1230750.0 100500.0 1229550.0 ;
      RECT  99300.0 1228800.0 98100.0 1227600.0 ;
      RECT  96900.0 1226850.0 95700.0 1225650.0 ;
      RECT  96900.0 1224150.0 98100.0 1222950.0 ;
      RECT  101700.0 1224150.0 102900.0 1222950.0 ;
      RECT  101700.0 1232850.0 102900.0 1231650.0 ;
      RECT  101700.0 1226850.0 102900.0 1225650.0 ;
      RECT  95700.0 1226850.0 96900.0 1225650.0 ;
      RECT  98100.0 1228800.0 99300.0 1227600.0 ;
      RECT  100500.0 1230750.0 101700.0 1229550.0 ;
      RECT  101700.0 1226850.0 102900.0 1225650.0 ;
      RECT  92700.0 1221450.0 108300.0 1220550.0 ;
      RECT  92700.0 1235250.0 108300.0 1234350.0 ;
      RECT  94500.0 1236750.0 95700.0 1234350.0 ;
      RECT  94500.0 1245450.0 95700.0 1249050.0 ;
      RECT  99300.0 1245450.0 100500.0 1249050.0 ;
      RECT  104100.0 1246650.0 105300.0 1248600.0 ;
      RECT  104100.0 1234800.0 105300.0 1236750.0 ;
      RECT  94500.0 1245450.0 95700.0 1246650.0 ;
      RECT  96900.0 1245450.0 98100.0 1246650.0 ;
      RECT  96900.0 1245450.0 98100.0 1246650.0 ;
      RECT  94500.0 1245450.0 95700.0 1246650.0 ;
      RECT  96900.0 1245450.0 98100.0 1246650.0 ;
      RECT  99300.0 1245450.0 100500.0 1246650.0 ;
      RECT  99300.0 1245450.0 100500.0 1246650.0 ;
      RECT  96900.0 1245450.0 98100.0 1246650.0 ;
      RECT  99300.0 1245450.0 100500.0 1246650.0 ;
      RECT  101700.0 1245450.0 102900.0 1246650.0 ;
      RECT  101700.0 1245450.0 102900.0 1246650.0 ;
      RECT  99300.0 1245450.0 100500.0 1246650.0 ;
      RECT  94500.0 1236750.0 95700.0 1237950.0 ;
      RECT  96900.0 1236750.0 98100.0 1237950.0 ;
      RECT  96900.0 1236750.0 98100.0 1237950.0 ;
      RECT  94500.0 1236750.0 95700.0 1237950.0 ;
      RECT  96900.0 1236750.0 98100.0 1237950.0 ;
      RECT  99300.0 1236750.0 100500.0 1237950.0 ;
      RECT  99300.0 1236750.0 100500.0 1237950.0 ;
      RECT  96900.0 1236750.0 98100.0 1237950.0 ;
      RECT  99300.0 1236750.0 100500.0 1237950.0 ;
      RECT  101700.0 1236750.0 102900.0 1237950.0 ;
      RECT  101700.0 1236750.0 102900.0 1237950.0 ;
      RECT  99300.0 1236750.0 100500.0 1237950.0 ;
      RECT  104100.0 1246050.0 105300.0 1247250.0 ;
      RECT  104100.0 1236150.0 105300.0 1237350.0 ;
      RECT  101700.0 1238850.0 100500.0 1240050.0 ;
      RECT  99300.0 1240800.0 98100.0 1242000.0 ;
      RECT  96900.0 1242750.0 95700.0 1243950.0 ;
      RECT  96900.0 1245450.0 98100.0 1246650.0 ;
      RECT  101700.0 1245450.0 102900.0 1246650.0 ;
      RECT  101700.0 1236750.0 102900.0 1237950.0 ;
      RECT  101700.0 1242750.0 102900.0 1243950.0 ;
      RECT  95700.0 1242750.0 96900.0 1243950.0 ;
      RECT  98100.0 1240800.0 99300.0 1242000.0 ;
      RECT  100500.0 1238850.0 101700.0 1240050.0 ;
      RECT  101700.0 1242750.0 102900.0 1243950.0 ;
      RECT  92700.0 1248150.0 108300.0 1249050.0 ;
      RECT  92700.0 1234350.0 108300.0 1235250.0 ;
      RECT  94500.0 1260450.0 95700.0 1262850.0 ;
      RECT  94500.0 1251750.0 95700.0 1248150.0 ;
      RECT  99300.0 1251750.0 100500.0 1248150.0 ;
      RECT  104100.0 1250550.0 105300.0 1248600.0 ;
      RECT  104100.0 1262400.0 105300.0 1260450.0 ;
      RECT  94500.0 1251750.0 95700.0 1250550.0 ;
      RECT  96900.0 1251750.0 98100.0 1250550.0 ;
      RECT  96900.0 1251750.0 98100.0 1250550.0 ;
      RECT  94500.0 1251750.0 95700.0 1250550.0 ;
      RECT  96900.0 1251750.0 98100.0 1250550.0 ;
      RECT  99300.0 1251750.0 100500.0 1250550.0 ;
      RECT  99300.0 1251750.0 100500.0 1250550.0 ;
      RECT  96900.0 1251750.0 98100.0 1250550.0 ;
      RECT  99300.0 1251750.0 100500.0 1250550.0 ;
      RECT  101700.0 1251750.0 102900.0 1250550.0 ;
      RECT  101700.0 1251750.0 102900.0 1250550.0 ;
      RECT  99300.0 1251750.0 100500.0 1250550.0 ;
      RECT  94500.0 1260450.0 95700.0 1259250.0 ;
      RECT  96900.0 1260450.0 98100.0 1259250.0 ;
      RECT  96900.0 1260450.0 98100.0 1259250.0 ;
      RECT  94500.0 1260450.0 95700.0 1259250.0 ;
      RECT  96900.0 1260450.0 98100.0 1259250.0 ;
      RECT  99300.0 1260450.0 100500.0 1259250.0 ;
      RECT  99300.0 1260450.0 100500.0 1259250.0 ;
      RECT  96900.0 1260450.0 98100.0 1259250.0 ;
      RECT  99300.0 1260450.0 100500.0 1259250.0 ;
      RECT  101700.0 1260450.0 102900.0 1259250.0 ;
      RECT  101700.0 1260450.0 102900.0 1259250.0 ;
      RECT  99300.0 1260450.0 100500.0 1259250.0 ;
      RECT  104100.0 1251150.0 105300.0 1249950.0 ;
      RECT  104100.0 1261050.0 105300.0 1259850.0 ;
      RECT  101700.0 1258350.0 100500.0 1257150.0 ;
      RECT  99300.0 1256400.0 98100.0 1255200.0 ;
      RECT  96900.0 1254450.0 95700.0 1253250.0 ;
      RECT  96900.0 1251750.0 98100.0 1250550.0 ;
      RECT  101700.0 1251750.0 102900.0 1250550.0 ;
      RECT  101700.0 1260450.0 102900.0 1259250.0 ;
      RECT  101700.0 1254450.0 102900.0 1253250.0 ;
      RECT  95700.0 1254450.0 96900.0 1253250.0 ;
      RECT  98100.0 1256400.0 99300.0 1255200.0 ;
      RECT  100500.0 1258350.0 101700.0 1257150.0 ;
      RECT  101700.0 1254450.0 102900.0 1253250.0 ;
      RECT  92700.0 1249050.0 108300.0 1248150.0 ;
      RECT  92700.0 1262850.0 108300.0 1261950.0 ;
      RECT  94500.0 1264350.0 95700.0 1261950.0 ;
      RECT  94500.0 1273050.0 95700.0 1276650.0 ;
      RECT  99300.0 1273050.0 100500.0 1276650.0 ;
      RECT  104100.0 1274250.0 105300.0 1276200.0 ;
      RECT  104100.0 1262400.0 105300.0 1264350.0 ;
      RECT  94500.0 1273050.0 95700.0 1274250.0 ;
      RECT  96900.0 1273050.0 98100.0 1274250.0 ;
      RECT  96900.0 1273050.0 98100.0 1274250.0 ;
      RECT  94500.0 1273050.0 95700.0 1274250.0 ;
      RECT  96900.0 1273050.0 98100.0 1274250.0 ;
      RECT  99300.0 1273050.0 100500.0 1274250.0 ;
      RECT  99300.0 1273050.0 100500.0 1274250.0 ;
      RECT  96900.0 1273050.0 98100.0 1274250.0 ;
      RECT  99300.0 1273050.0 100500.0 1274250.0 ;
      RECT  101700.0 1273050.0 102900.0 1274250.0 ;
      RECT  101700.0 1273050.0 102900.0 1274250.0 ;
      RECT  99300.0 1273050.0 100500.0 1274250.0 ;
      RECT  94500.0 1264350.0 95700.0 1265550.0 ;
      RECT  96900.0 1264350.0 98100.0 1265550.0 ;
      RECT  96900.0 1264350.0 98100.0 1265550.0 ;
      RECT  94500.0 1264350.0 95700.0 1265550.0 ;
      RECT  96900.0 1264350.0 98100.0 1265550.0 ;
      RECT  99300.0 1264350.0 100500.0 1265550.0 ;
      RECT  99300.0 1264350.0 100500.0 1265550.0 ;
      RECT  96900.0 1264350.0 98100.0 1265550.0 ;
      RECT  99300.0 1264350.0 100500.0 1265550.0 ;
      RECT  101700.0 1264350.0 102900.0 1265550.0 ;
      RECT  101700.0 1264350.0 102900.0 1265550.0 ;
      RECT  99300.0 1264350.0 100500.0 1265550.0 ;
      RECT  104100.0 1273650.0 105300.0 1274850.0 ;
      RECT  104100.0 1263750.0 105300.0 1264950.0 ;
      RECT  101700.0 1266450.0 100500.0 1267650.0 ;
      RECT  99300.0 1268400.0 98100.0 1269600.0 ;
      RECT  96900.0 1270350.0 95700.0 1271550.0 ;
      RECT  96900.0 1273050.0 98100.0 1274250.0 ;
      RECT  101700.0 1273050.0 102900.0 1274250.0 ;
      RECT  101700.0 1264350.0 102900.0 1265550.0 ;
      RECT  101700.0 1270350.0 102900.0 1271550.0 ;
      RECT  95700.0 1270350.0 96900.0 1271550.0 ;
      RECT  98100.0 1268400.0 99300.0 1269600.0 ;
      RECT  100500.0 1266450.0 101700.0 1267650.0 ;
      RECT  101700.0 1270350.0 102900.0 1271550.0 ;
      RECT  92700.0 1275750.0 108300.0 1276650.0 ;
      RECT  92700.0 1261950.0 108300.0 1262850.0 ;
      RECT  94500.0 1288050.0 95700.0 1290450.0 ;
      RECT  94500.0 1279350.0 95700.0 1275750.0 ;
      RECT  99300.0 1279350.0 100500.0 1275750.0 ;
      RECT  104100.0 1278150.0 105300.0 1276200.0 ;
      RECT  104100.0 1290000.0 105300.0 1288050.0 ;
      RECT  94500.0 1279350.0 95700.0 1278150.0 ;
      RECT  96900.0 1279350.0 98100.0 1278150.0 ;
      RECT  96900.0 1279350.0 98100.0 1278150.0 ;
      RECT  94500.0 1279350.0 95700.0 1278150.0 ;
      RECT  96900.0 1279350.0 98100.0 1278150.0 ;
      RECT  99300.0 1279350.0 100500.0 1278150.0 ;
      RECT  99300.0 1279350.0 100500.0 1278150.0 ;
      RECT  96900.0 1279350.0 98100.0 1278150.0 ;
      RECT  99300.0 1279350.0 100500.0 1278150.0 ;
      RECT  101700.0 1279350.0 102900.0 1278150.0 ;
      RECT  101700.0 1279350.0 102900.0 1278150.0 ;
      RECT  99300.0 1279350.0 100500.0 1278150.0 ;
      RECT  94500.0 1288050.0 95700.0 1286850.0 ;
      RECT  96900.0 1288050.0 98100.0 1286850.0 ;
      RECT  96900.0 1288050.0 98100.0 1286850.0 ;
      RECT  94500.0 1288050.0 95700.0 1286850.0 ;
      RECT  96900.0 1288050.0 98100.0 1286850.0 ;
      RECT  99300.0 1288050.0 100500.0 1286850.0 ;
      RECT  99300.0 1288050.0 100500.0 1286850.0 ;
      RECT  96900.0 1288050.0 98100.0 1286850.0 ;
      RECT  99300.0 1288050.0 100500.0 1286850.0 ;
      RECT  101700.0 1288050.0 102900.0 1286850.0 ;
      RECT  101700.0 1288050.0 102900.0 1286850.0 ;
      RECT  99300.0 1288050.0 100500.0 1286850.0 ;
      RECT  104100.0 1278750.0 105300.0 1277550.0 ;
      RECT  104100.0 1288650.0 105300.0 1287450.0 ;
      RECT  101700.0 1285950.0 100500.0 1284750.0 ;
      RECT  99300.0 1284000.0 98100.0 1282800.0 ;
      RECT  96900.0 1282050.0 95700.0 1280850.0 ;
      RECT  96900.0 1279350.0 98100.0 1278150.0 ;
      RECT  101700.0 1279350.0 102900.0 1278150.0 ;
      RECT  101700.0 1288050.0 102900.0 1286850.0 ;
      RECT  101700.0 1282050.0 102900.0 1280850.0 ;
      RECT  95700.0 1282050.0 96900.0 1280850.0 ;
      RECT  98100.0 1284000.0 99300.0 1282800.0 ;
      RECT  100500.0 1285950.0 101700.0 1284750.0 ;
      RECT  101700.0 1282050.0 102900.0 1280850.0 ;
      RECT  92700.0 1276650.0 108300.0 1275750.0 ;
      RECT  92700.0 1290450.0 108300.0 1289550.0 ;
      RECT  94500.0 1291950.0 95700.0 1289550.0 ;
      RECT  94500.0 1300650.0 95700.0 1304250.0 ;
      RECT  99300.0 1300650.0 100500.0 1304250.0 ;
      RECT  104100.0 1301850.0 105300.0 1303800.0 ;
      RECT  104100.0 1290000.0 105300.0 1291950.0 ;
      RECT  94500.0 1300650.0 95700.0 1301850.0 ;
      RECT  96900.0 1300650.0 98100.0 1301850.0 ;
      RECT  96900.0 1300650.0 98100.0 1301850.0 ;
      RECT  94500.0 1300650.0 95700.0 1301850.0 ;
      RECT  96900.0 1300650.0 98100.0 1301850.0 ;
      RECT  99300.0 1300650.0 100500.0 1301850.0 ;
      RECT  99300.0 1300650.0 100500.0 1301850.0 ;
      RECT  96900.0 1300650.0 98100.0 1301850.0 ;
      RECT  99300.0 1300650.0 100500.0 1301850.0 ;
      RECT  101700.0 1300650.0 102900.0 1301850.0 ;
      RECT  101700.0 1300650.0 102900.0 1301850.0 ;
      RECT  99300.0 1300650.0 100500.0 1301850.0 ;
      RECT  94500.0 1291950.0 95700.0 1293150.0 ;
      RECT  96900.0 1291950.0 98100.0 1293150.0 ;
      RECT  96900.0 1291950.0 98100.0 1293150.0 ;
      RECT  94500.0 1291950.0 95700.0 1293150.0 ;
      RECT  96900.0 1291950.0 98100.0 1293150.0 ;
      RECT  99300.0 1291950.0 100500.0 1293150.0 ;
      RECT  99300.0 1291950.0 100500.0 1293150.0 ;
      RECT  96900.0 1291950.0 98100.0 1293150.0 ;
      RECT  99300.0 1291950.0 100500.0 1293150.0 ;
      RECT  101700.0 1291950.0 102900.0 1293150.0 ;
      RECT  101700.0 1291950.0 102900.0 1293150.0 ;
      RECT  99300.0 1291950.0 100500.0 1293150.0 ;
      RECT  104100.0 1301250.0 105300.0 1302450.0 ;
      RECT  104100.0 1291350.0 105300.0 1292550.0 ;
      RECT  101700.0 1294050.0 100500.0 1295250.0 ;
      RECT  99300.0 1296000.0 98100.0 1297200.0 ;
      RECT  96900.0 1297950.0 95700.0 1299150.0 ;
      RECT  96900.0 1300650.0 98100.0 1301850.0 ;
      RECT  101700.0 1300650.0 102900.0 1301850.0 ;
      RECT  101700.0 1291950.0 102900.0 1293150.0 ;
      RECT  101700.0 1297950.0 102900.0 1299150.0 ;
      RECT  95700.0 1297950.0 96900.0 1299150.0 ;
      RECT  98100.0 1296000.0 99300.0 1297200.0 ;
      RECT  100500.0 1294050.0 101700.0 1295250.0 ;
      RECT  101700.0 1297950.0 102900.0 1299150.0 ;
      RECT  92700.0 1303350.0 108300.0 1304250.0 ;
      RECT  92700.0 1289550.0 108300.0 1290450.0 ;
      RECT  94500.0 1315650.0 95700.0 1318050.0 ;
      RECT  94500.0 1306950.0 95700.0 1303350.0 ;
      RECT  99300.0 1306950.0 100500.0 1303350.0 ;
      RECT  104100.0 1305750.0 105300.0 1303800.0 ;
      RECT  104100.0 1317600.0 105300.0 1315650.0 ;
      RECT  94500.0 1306950.0 95700.0 1305750.0 ;
      RECT  96900.0 1306950.0 98100.0 1305750.0 ;
      RECT  96900.0 1306950.0 98100.0 1305750.0 ;
      RECT  94500.0 1306950.0 95700.0 1305750.0 ;
      RECT  96900.0 1306950.0 98100.0 1305750.0 ;
      RECT  99300.0 1306950.0 100500.0 1305750.0 ;
      RECT  99300.0 1306950.0 100500.0 1305750.0 ;
      RECT  96900.0 1306950.0 98100.0 1305750.0 ;
      RECT  99300.0 1306950.0 100500.0 1305750.0 ;
      RECT  101700.0 1306950.0 102900.0 1305750.0 ;
      RECT  101700.0 1306950.0 102900.0 1305750.0 ;
      RECT  99300.0 1306950.0 100500.0 1305750.0 ;
      RECT  94500.0 1315650.0 95700.0 1314450.0 ;
      RECT  96900.0 1315650.0 98100.0 1314450.0 ;
      RECT  96900.0 1315650.0 98100.0 1314450.0 ;
      RECT  94500.0 1315650.0 95700.0 1314450.0 ;
      RECT  96900.0 1315650.0 98100.0 1314450.0 ;
      RECT  99300.0 1315650.0 100500.0 1314450.0 ;
      RECT  99300.0 1315650.0 100500.0 1314450.0 ;
      RECT  96900.0 1315650.0 98100.0 1314450.0 ;
      RECT  99300.0 1315650.0 100500.0 1314450.0 ;
      RECT  101700.0 1315650.0 102900.0 1314450.0 ;
      RECT  101700.0 1315650.0 102900.0 1314450.0 ;
      RECT  99300.0 1315650.0 100500.0 1314450.0 ;
      RECT  104100.0 1306350.0 105300.0 1305150.0 ;
      RECT  104100.0 1316250.0 105300.0 1315050.0 ;
      RECT  101700.0 1313550.0 100500.0 1312350.0 ;
      RECT  99300.0 1311600.0 98100.0 1310400.0 ;
      RECT  96900.0 1309650.0 95700.0 1308450.0 ;
      RECT  96900.0 1306950.0 98100.0 1305750.0 ;
      RECT  101700.0 1306950.0 102900.0 1305750.0 ;
      RECT  101700.0 1315650.0 102900.0 1314450.0 ;
      RECT  101700.0 1309650.0 102900.0 1308450.0 ;
      RECT  95700.0 1309650.0 96900.0 1308450.0 ;
      RECT  98100.0 1311600.0 99300.0 1310400.0 ;
      RECT  100500.0 1313550.0 101700.0 1312350.0 ;
      RECT  101700.0 1309650.0 102900.0 1308450.0 ;
      RECT  92700.0 1304250.0 108300.0 1303350.0 ;
      RECT  92700.0 1318050.0 108300.0 1317150.0 ;
      RECT  94500.0 1319550.0 95700.0 1317150.0 ;
      RECT  94500.0 1328250.0 95700.0 1331850.0 ;
      RECT  99300.0 1328250.0 100500.0 1331850.0 ;
      RECT  104100.0 1329450.0 105300.0 1331400.0 ;
      RECT  104100.0 1317600.0 105300.0 1319550.0 ;
      RECT  94500.0 1328250.0 95700.0 1329450.0 ;
      RECT  96900.0 1328250.0 98100.0 1329450.0 ;
      RECT  96900.0 1328250.0 98100.0 1329450.0 ;
      RECT  94500.0 1328250.0 95700.0 1329450.0 ;
      RECT  96900.0 1328250.0 98100.0 1329450.0 ;
      RECT  99300.0 1328250.0 100500.0 1329450.0 ;
      RECT  99300.0 1328250.0 100500.0 1329450.0 ;
      RECT  96900.0 1328250.0 98100.0 1329450.0 ;
      RECT  99300.0 1328250.0 100500.0 1329450.0 ;
      RECT  101700.0 1328250.0 102900.0 1329450.0 ;
      RECT  101700.0 1328250.0 102900.0 1329450.0 ;
      RECT  99300.0 1328250.0 100500.0 1329450.0 ;
      RECT  94500.0 1319550.0 95700.0 1320750.0 ;
      RECT  96900.0 1319550.0 98100.0 1320750.0 ;
      RECT  96900.0 1319550.0 98100.0 1320750.0 ;
      RECT  94500.0 1319550.0 95700.0 1320750.0 ;
      RECT  96900.0 1319550.0 98100.0 1320750.0 ;
      RECT  99300.0 1319550.0 100500.0 1320750.0 ;
      RECT  99300.0 1319550.0 100500.0 1320750.0 ;
      RECT  96900.0 1319550.0 98100.0 1320750.0 ;
      RECT  99300.0 1319550.0 100500.0 1320750.0 ;
      RECT  101700.0 1319550.0 102900.0 1320750.0 ;
      RECT  101700.0 1319550.0 102900.0 1320750.0 ;
      RECT  99300.0 1319550.0 100500.0 1320750.0 ;
      RECT  104100.0 1328850.0 105300.0 1330050.0 ;
      RECT  104100.0 1318950.0 105300.0 1320150.0 ;
      RECT  101700.0 1321650.0 100500.0 1322850.0 ;
      RECT  99300.0 1323600.0 98100.0 1324800.0 ;
      RECT  96900.0 1325550.0 95700.0 1326750.0 ;
      RECT  96900.0 1328250.0 98100.0 1329450.0 ;
      RECT  101700.0 1328250.0 102900.0 1329450.0 ;
      RECT  101700.0 1319550.0 102900.0 1320750.0 ;
      RECT  101700.0 1325550.0 102900.0 1326750.0 ;
      RECT  95700.0 1325550.0 96900.0 1326750.0 ;
      RECT  98100.0 1323600.0 99300.0 1324800.0 ;
      RECT  100500.0 1321650.0 101700.0 1322850.0 ;
      RECT  101700.0 1325550.0 102900.0 1326750.0 ;
      RECT  92700.0 1330950.0 108300.0 1331850.0 ;
      RECT  92700.0 1317150.0 108300.0 1318050.0 ;
      RECT  94500.0 1343250.0 95700.0 1345650.0 ;
      RECT  94500.0 1334550.0 95700.0 1330950.0 ;
      RECT  99300.0 1334550.0 100500.0 1330950.0 ;
      RECT  104100.0 1333350.0 105300.0 1331400.0 ;
      RECT  104100.0 1345200.0 105300.0 1343250.0 ;
      RECT  94500.0 1334550.0 95700.0 1333350.0 ;
      RECT  96900.0 1334550.0 98100.0 1333350.0 ;
      RECT  96900.0 1334550.0 98100.0 1333350.0 ;
      RECT  94500.0 1334550.0 95700.0 1333350.0 ;
      RECT  96900.0 1334550.0 98100.0 1333350.0 ;
      RECT  99300.0 1334550.0 100500.0 1333350.0 ;
      RECT  99300.0 1334550.0 100500.0 1333350.0 ;
      RECT  96900.0 1334550.0 98100.0 1333350.0 ;
      RECT  99300.0 1334550.0 100500.0 1333350.0 ;
      RECT  101700.0 1334550.0 102900.0 1333350.0 ;
      RECT  101700.0 1334550.0 102900.0 1333350.0 ;
      RECT  99300.0 1334550.0 100500.0 1333350.0 ;
      RECT  94500.0 1343250.0 95700.0 1342050.0 ;
      RECT  96900.0 1343250.0 98100.0 1342050.0 ;
      RECT  96900.0 1343250.0 98100.0 1342050.0 ;
      RECT  94500.0 1343250.0 95700.0 1342050.0 ;
      RECT  96900.0 1343250.0 98100.0 1342050.0 ;
      RECT  99300.0 1343250.0 100500.0 1342050.0 ;
      RECT  99300.0 1343250.0 100500.0 1342050.0 ;
      RECT  96900.0 1343250.0 98100.0 1342050.0 ;
      RECT  99300.0 1343250.0 100500.0 1342050.0 ;
      RECT  101700.0 1343250.0 102900.0 1342050.0 ;
      RECT  101700.0 1343250.0 102900.0 1342050.0 ;
      RECT  99300.0 1343250.0 100500.0 1342050.0 ;
      RECT  104100.0 1333950.0 105300.0 1332750.0 ;
      RECT  104100.0 1343850.0 105300.0 1342650.0 ;
      RECT  101700.0 1341150.0 100500.0 1339950.0 ;
      RECT  99300.0 1339200.0 98100.0 1338000.0 ;
      RECT  96900.0 1337250.0 95700.0 1336050.0 ;
      RECT  96900.0 1334550.0 98100.0 1333350.0 ;
      RECT  101700.0 1334550.0 102900.0 1333350.0 ;
      RECT  101700.0 1343250.0 102900.0 1342050.0 ;
      RECT  101700.0 1337250.0 102900.0 1336050.0 ;
      RECT  95700.0 1337250.0 96900.0 1336050.0 ;
      RECT  98100.0 1339200.0 99300.0 1338000.0 ;
      RECT  100500.0 1341150.0 101700.0 1339950.0 ;
      RECT  101700.0 1337250.0 102900.0 1336050.0 ;
      RECT  92700.0 1331850.0 108300.0 1330950.0 ;
      RECT  92700.0 1345650.0 108300.0 1344750.0 ;
      RECT  94500.0 1347150.0 95700.0 1344750.0 ;
      RECT  94500.0 1355850.0 95700.0 1359450.0 ;
      RECT  99300.0 1355850.0 100500.0 1359450.0 ;
      RECT  104100.0 1357050.0 105300.0 1359000.0 ;
      RECT  104100.0 1345200.0 105300.0 1347150.0 ;
      RECT  94500.0 1355850.0 95700.0 1357050.0 ;
      RECT  96900.0 1355850.0 98100.0 1357050.0 ;
      RECT  96900.0 1355850.0 98100.0 1357050.0 ;
      RECT  94500.0 1355850.0 95700.0 1357050.0 ;
      RECT  96900.0 1355850.0 98100.0 1357050.0 ;
      RECT  99300.0 1355850.0 100500.0 1357050.0 ;
      RECT  99300.0 1355850.0 100500.0 1357050.0 ;
      RECT  96900.0 1355850.0 98100.0 1357050.0 ;
      RECT  99300.0 1355850.0 100500.0 1357050.0 ;
      RECT  101700.0 1355850.0 102900.0 1357050.0 ;
      RECT  101700.0 1355850.0 102900.0 1357050.0 ;
      RECT  99300.0 1355850.0 100500.0 1357050.0 ;
      RECT  94500.0 1347150.0 95700.0 1348350.0 ;
      RECT  96900.0 1347150.0 98100.0 1348350.0 ;
      RECT  96900.0 1347150.0 98100.0 1348350.0 ;
      RECT  94500.0 1347150.0 95700.0 1348350.0 ;
      RECT  96900.0 1347150.0 98100.0 1348350.0 ;
      RECT  99300.0 1347150.0 100500.0 1348350.0 ;
      RECT  99300.0 1347150.0 100500.0 1348350.0 ;
      RECT  96900.0 1347150.0 98100.0 1348350.0 ;
      RECT  99300.0 1347150.0 100500.0 1348350.0 ;
      RECT  101700.0 1347150.0 102900.0 1348350.0 ;
      RECT  101700.0 1347150.0 102900.0 1348350.0 ;
      RECT  99300.0 1347150.0 100500.0 1348350.0 ;
      RECT  104100.0 1356450.0 105300.0 1357650.0 ;
      RECT  104100.0 1346550.0 105300.0 1347750.0 ;
      RECT  101700.0 1349250.0 100500.0 1350450.0 ;
      RECT  99300.0 1351200.0 98100.0 1352400.0 ;
      RECT  96900.0 1353150.0 95700.0 1354350.0 ;
      RECT  96900.0 1355850.0 98100.0 1357050.0 ;
      RECT  101700.0 1355850.0 102900.0 1357050.0 ;
      RECT  101700.0 1347150.0 102900.0 1348350.0 ;
      RECT  101700.0 1353150.0 102900.0 1354350.0 ;
      RECT  95700.0 1353150.0 96900.0 1354350.0 ;
      RECT  98100.0 1351200.0 99300.0 1352400.0 ;
      RECT  100500.0 1349250.0 101700.0 1350450.0 ;
      RECT  101700.0 1353150.0 102900.0 1354350.0 ;
      RECT  92700.0 1358550.0 108300.0 1359450.0 ;
      RECT  92700.0 1344750.0 108300.0 1345650.0 ;
      RECT  94500.0 1370850.0 95700.0 1373250.0 ;
      RECT  94500.0 1362150.0 95700.0 1358550.0 ;
      RECT  99300.0 1362150.0 100500.0 1358550.0 ;
      RECT  104100.0 1360950.0 105300.0 1359000.0 ;
      RECT  104100.0 1372800.0 105300.0 1370850.0 ;
      RECT  94500.0 1362150.0 95700.0 1360950.0 ;
      RECT  96900.0 1362150.0 98100.0 1360950.0 ;
      RECT  96900.0 1362150.0 98100.0 1360950.0 ;
      RECT  94500.0 1362150.0 95700.0 1360950.0 ;
      RECT  96900.0 1362150.0 98100.0 1360950.0 ;
      RECT  99300.0 1362150.0 100500.0 1360950.0 ;
      RECT  99300.0 1362150.0 100500.0 1360950.0 ;
      RECT  96900.0 1362150.0 98100.0 1360950.0 ;
      RECT  99300.0 1362150.0 100500.0 1360950.0 ;
      RECT  101700.0 1362150.0 102900.0 1360950.0 ;
      RECT  101700.0 1362150.0 102900.0 1360950.0 ;
      RECT  99300.0 1362150.0 100500.0 1360950.0 ;
      RECT  94500.0 1370850.0 95700.0 1369650.0 ;
      RECT  96900.0 1370850.0 98100.0 1369650.0 ;
      RECT  96900.0 1370850.0 98100.0 1369650.0 ;
      RECT  94500.0 1370850.0 95700.0 1369650.0 ;
      RECT  96900.0 1370850.0 98100.0 1369650.0 ;
      RECT  99300.0 1370850.0 100500.0 1369650.0 ;
      RECT  99300.0 1370850.0 100500.0 1369650.0 ;
      RECT  96900.0 1370850.0 98100.0 1369650.0 ;
      RECT  99300.0 1370850.0 100500.0 1369650.0 ;
      RECT  101700.0 1370850.0 102900.0 1369650.0 ;
      RECT  101700.0 1370850.0 102900.0 1369650.0 ;
      RECT  99300.0 1370850.0 100500.0 1369650.0 ;
      RECT  104100.0 1361550.0 105300.0 1360350.0 ;
      RECT  104100.0 1371450.0 105300.0 1370250.0 ;
      RECT  101700.0 1368750.0 100500.0 1367550.0 ;
      RECT  99300.0 1366800.0 98100.0 1365600.0 ;
      RECT  96900.0 1364850.0 95700.0 1363650.0 ;
      RECT  96900.0 1362150.0 98100.0 1360950.0 ;
      RECT  101700.0 1362150.0 102900.0 1360950.0 ;
      RECT  101700.0 1370850.0 102900.0 1369650.0 ;
      RECT  101700.0 1364850.0 102900.0 1363650.0 ;
      RECT  95700.0 1364850.0 96900.0 1363650.0 ;
      RECT  98100.0 1366800.0 99300.0 1365600.0 ;
      RECT  100500.0 1368750.0 101700.0 1367550.0 ;
      RECT  101700.0 1364850.0 102900.0 1363650.0 ;
      RECT  92700.0 1359450.0 108300.0 1358550.0 ;
      RECT  92700.0 1373250.0 108300.0 1372350.0 ;
      RECT  94500.0 1374750.0 95700.0 1372350.0 ;
      RECT  94500.0 1383450.0 95700.0 1387050.0 ;
      RECT  99300.0 1383450.0 100500.0 1387050.0 ;
      RECT  104100.0 1384650.0 105300.0 1386600.0 ;
      RECT  104100.0 1372800.0 105300.0 1374750.0 ;
      RECT  94500.0 1383450.0 95700.0 1384650.0 ;
      RECT  96900.0 1383450.0 98100.0 1384650.0 ;
      RECT  96900.0 1383450.0 98100.0 1384650.0 ;
      RECT  94500.0 1383450.0 95700.0 1384650.0 ;
      RECT  96900.0 1383450.0 98100.0 1384650.0 ;
      RECT  99300.0 1383450.0 100500.0 1384650.0 ;
      RECT  99300.0 1383450.0 100500.0 1384650.0 ;
      RECT  96900.0 1383450.0 98100.0 1384650.0 ;
      RECT  99300.0 1383450.0 100500.0 1384650.0 ;
      RECT  101700.0 1383450.0 102900.0 1384650.0 ;
      RECT  101700.0 1383450.0 102900.0 1384650.0 ;
      RECT  99300.0 1383450.0 100500.0 1384650.0 ;
      RECT  94500.0 1374750.0 95700.0 1375950.0 ;
      RECT  96900.0 1374750.0 98100.0 1375950.0 ;
      RECT  96900.0 1374750.0 98100.0 1375950.0 ;
      RECT  94500.0 1374750.0 95700.0 1375950.0 ;
      RECT  96900.0 1374750.0 98100.0 1375950.0 ;
      RECT  99300.0 1374750.0 100500.0 1375950.0 ;
      RECT  99300.0 1374750.0 100500.0 1375950.0 ;
      RECT  96900.0 1374750.0 98100.0 1375950.0 ;
      RECT  99300.0 1374750.0 100500.0 1375950.0 ;
      RECT  101700.0 1374750.0 102900.0 1375950.0 ;
      RECT  101700.0 1374750.0 102900.0 1375950.0 ;
      RECT  99300.0 1374750.0 100500.0 1375950.0 ;
      RECT  104100.0 1384050.0 105300.0 1385250.0 ;
      RECT  104100.0 1374150.0 105300.0 1375350.0 ;
      RECT  101700.0 1376850.0 100500.0 1378050.0 ;
      RECT  99300.0 1378800.0 98100.0 1380000.0 ;
      RECT  96900.0 1380750.0 95700.0 1381950.0 ;
      RECT  96900.0 1383450.0 98100.0 1384650.0 ;
      RECT  101700.0 1383450.0 102900.0 1384650.0 ;
      RECT  101700.0 1374750.0 102900.0 1375950.0 ;
      RECT  101700.0 1380750.0 102900.0 1381950.0 ;
      RECT  95700.0 1380750.0 96900.0 1381950.0 ;
      RECT  98100.0 1378800.0 99300.0 1380000.0 ;
      RECT  100500.0 1376850.0 101700.0 1378050.0 ;
      RECT  101700.0 1380750.0 102900.0 1381950.0 ;
      RECT  92700.0 1386150.0 108300.0 1387050.0 ;
      RECT  92700.0 1372350.0 108300.0 1373250.0 ;
      RECT  94500.0 1398450.0 95700.0 1400850.0 ;
      RECT  94500.0 1389750.0 95700.0 1386150.0 ;
      RECT  99300.0 1389750.0 100500.0 1386150.0 ;
      RECT  104100.0 1388550.0 105300.0 1386600.0 ;
      RECT  104100.0 1400400.0 105300.0 1398450.0 ;
      RECT  94500.0 1389750.0 95700.0 1388550.0 ;
      RECT  96900.0 1389750.0 98100.0 1388550.0 ;
      RECT  96900.0 1389750.0 98100.0 1388550.0 ;
      RECT  94500.0 1389750.0 95700.0 1388550.0 ;
      RECT  96900.0 1389750.0 98100.0 1388550.0 ;
      RECT  99300.0 1389750.0 100500.0 1388550.0 ;
      RECT  99300.0 1389750.0 100500.0 1388550.0 ;
      RECT  96900.0 1389750.0 98100.0 1388550.0 ;
      RECT  99300.0 1389750.0 100500.0 1388550.0 ;
      RECT  101700.0 1389750.0 102900.0 1388550.0 ;
      RECT  101700.0 1389750.0 102900.0 1388550.0 ;
      RECT  99300.0 1389750.0 100500.0 1388550.0 ;
      RECT  94500.0 1398450.0 95700.0 1397250.0 ;
      RECT  96900.0 1398450.0 98100.0 1397250.0 ;
      RECT  96900.0 1398450.0 98100.0 1397250.0 ;
      RECT  94500.0 1398450.0 95700.0 1397250.0 ;
      RECT  96900.0 1398450.0 98100.0 1397250.0 ;
      RECT  99300.0 1398450.0 100500.0 1397250.0 ;
      RECT  99300.0 1398450.0 100500.0 1397250.0 ;
      RECT  96900.0 1398450.0 98100.0 1397250.0 ;
      RECT  99300.0 1398450.0 100500.0 1397250.0 ;
      RECT  101700.0 1398450.0 102900.0 1397250.0 ;
      RECT  101700.0 1398450.0 102900.0 1397250.0 ;
      RECT  99300.0 1398450.0 100500.0 1397250.0 ;
      RECT  104100.0 1389150.0 105300.0 1387950.0 ;
      RECT  104100.0 1399050.0 105300.0 1397850.0 ;
      RECT  101700.0 1396350.0 100500.0 1395150.0 ;
      RECT  99300.0 1394400.0 98100.0 1393200.0 ;
      RECT  96900.0 1392450.0 95700.0 1391250.0 ;
      RECT  96900.0 1389750.0 98100.0 1388550.0 ;
      RECT  101700.0 1389750.0 102900.0 1388550.0 ;
      RECT  101700.0 1398450.0 102900.0 1397250.0 ;
      RECT  101700.0 1392450.0 102900.0 1391250.0 ;
      RECT  95700.0 1392450.0 96900.0 1391250.0 ;
      RECT  98100.0 1394400.0 99300.0 1393200.0 ;
      RECT  100500.0 1396350.0 101700.0 1395150.0 ;
      RECT  101700.0 1392450.0 102900.0 1391250.0 ;
      RECT  92700.0 1387050.0 108300.0 1386150.0 ;
      RECT  92700.0 1400850.0 108300.0 1399950.0 ;
      RECT  94500.0 1402350.0 95700.0 1399950.0 ;
      RECT  94500.0 1411050.0 95700.0 1414650.0 ;
      RECT  99300.0 1411050.0 100500.0 1414650.0 ;
      RECT  104100.0 1412250.0 105300.0 1414200.0 ;
      RECT  104100.0 1400400.0 105300.0 1402350.0 ;
      RECT  94500.0 1411050.0 95700.0 1412250.0 ;
      RECT  96900.0 1411050.0 98100.0 1412250.0 ;
      RECT  96900.0 1411050.0 98100.0 1412250.0 ;
      RECT  94500.0 1411050.0 95700.0 1412250.0 ;
      RECT  96900.0 1411050.0 98100.0 1412250.0 ;
      RECT  99300.0 1411050.0 100500.0 1412250.0 ;
      RECT  99300.0 1411050.0 100500.0 1412250.0 ;
      RECT  96900.0 1411050.0 98100.0 1412250.0 ;
      RECT  99300.0 1411050.0 100500.0 1412250.0 ;
      RECT  101700.0 1411050.0 102900.0 1412250.0 ;
      RECT  101700.0 1411050.0 102900.0 1412250.0 ;
      RECT  99300.0 1411050.0 100500.0 1412250.0 ;
      RECT  94500.0 1402350.0 95700.0 1403550.0 ;
      RECT  96900.0 1402350.0 98100.0 1403550.0 ;
      RECT  96900.0 1402350.0 98100.0 1403550.0 ;
      RECT  94500.0 1402350.0 95700.0 1403550.0 ;
      RECT  96900.0 1402350.0 98100.0 1403550.0 ;
      RECT  99300.0 1402350.0 100500.0 1403550.0 ;
      RECT  99300.0 1402350.0 100500.0 1403550.0 ;
      RECT  96900.0 1402350.0 98100.0 1403550.0 ;
      RECT  99300.0 1402350.0 100500.0 1403550.0 ;
      RECT  101700.0 1402350.0 102900.0 1403550.0 ;
      RECT  101700.0 1402350.0 102900.0 1403550.0 ;
      RECT  99300.0 1402350.0 100500.0 1403550.0 ;
      RECT  104100.0 1411650.0 105300.0 1412850.0 ;
      RECT  104100.0 1401750.0 105300.0 1402950.0 ;
      RECT  101700.0 1404450.0 100500.0 1405650.0 ;
      RECT  99300.0 1406400.0 98100.0 1407600.0 ;
      RECT  96900.0 1408350.0 95700.0 1409550.0 ;
      RECT  96900.0 1411050.0 98100.0 1412250.0 ;
      RECT  101700.0 1411050.0 102900.0 1412250.0 ;
      RECT  101700.0 1402350.0 102900.0 1403550.0 ;
      RECT  101700.0 1408350.0 102900.0 1409550.0 ;
      RECT  95700.0 1408350.0 96900.0 1409550.0 ;
      RECT  98100.0 1406400.0 99300.0 1407600.0 ;
      RECT  100500.0 1404450.0 101700.0 1405650.0 ;
      RECT  101700.0 1408350.0 102900.0 1409550.0 ;
      RECT  92700.0 1413750.0 108300.0 1414650.0 ;
      RECT  92700.0 1399950.0 108300.0 1400850.0 ;
      RECT  94500.0 1426050.0 95700.0 1428450.0 ;
      RECT  94500.0 1417350.0 95700.0 1413750.0 ;
      RECT  99300.0 1417350.0 100500.0 1413750.0 ;
      RECT  104100.0 1416150.0 105300.0 1414200.0 ;
      RECT  104100.0 1428000.0 105300.0 1426050.0 ;
      RECT  94500.0 1417350.0 95700.0 1416150.0 ;
      RECT  96900.0 1417350.0 98100.0 1416150.0 ;
      RECT  96900.0 1417350.0 98100.0 1416150.0 ;
      RECT  94500.0 1417350.0 95700.0 1416150.0 ;
      RECT  96900.0 1417350.0 98100.0 1416150.0 ;
      RECT  99300.0 1417350.0 100500.0 1416150.0 ;
      RECT  99300.0 1417350.0 100500.0 1416150.0 ;
      RECT  96900.0 1417350.0 98100.0 1416150.0 ;
      RECT  99300.0 1417350.0 100500.0 1416150.0 ;
      RECT  101700.0 1417350.0 102900.0 1416150.0 ;
      RECT  101700.0 1417350.0 102900.0 1416150.0 ;
      RECT  99300.0 1417350.0 100500.0 1416150.0 ;
      RECT  94500.0 1426050.0 95700.0 1424850.0 ;
      RECT  96900.0 1426050.0 98100.0 1424850.0 ;
      RECT  96900.0 1426050.0 98100.0 1424850.0 ;
      RECT  94500.0 1426050.0 95700.0 1424850.0 ;
      RECT  96900.0 1426050.0 98100.0 1424850.0 ;
      RECT  99300.0 1426050.0 100500.0 1424850.0 ;
      RECT  99300.0 1426050.0 100500.0 1424850.0 ;
      RECT  96900.0 1426050.0 98100.0 1424850.0 ;
      RECT  99300.0 1426050.0 100500.0 1424850.0 ;
      RECT  101700.0 1426050.0 102900.0 1424850.0 ;
      RECT  101700.0 1426050.0 102900.0 1424850.0 ;
      RECT  99300.0 1426050.0 100500.0 1424850.0 ;
      RECT  104100.0 1416750.0 105300.0 1415550.0 ;
      RECT  104100.0 1426650.0 105300.0 1425450.0 ;
      RECT  101700.0 1423950.0 100500.0 1422750.0 ;
      RECT  99300.0 1422000.0 98100.0 1420800.0 ;
      RECT  96900.0 1420050.0 95700.0 1418850.0 ;
      RECT  96900.0 1417350.0 98100.0 1416150.0 ;
      RECT  101700.0 1417350.0 102900.0 1416150.0 ;
      RECT  101700.0 1426050.0 102900.0 1424850.0 ;
      RECT  101700.0 1420050.0 102900.0 1418850.0 ;
      RECT  95700.0 1420050.0 96900.0 1418850.0 ;
      RECT  98100.0 1422000.0 99300.0 1420800.0 ;
      RECT  100500.0 1423950.0 101700.0 1422750.0 ;
      RECT  101700.0 1420050.0 102900.0 1418850.0 ;
      RECT  92700.0 1414650.0 108300.0 1413750.0 ;
      RECT  92700.0 1428450.0 108300.0 1427550.0 ;
      RECT  94500.0 1429950.0 95700.0 1427550.0 ;
      RECT  94500.0 1438650.0 95700.0 1442250.0 ;
      RECT  99300.0 1438650.0 100500.0 1442250.0 ;
      RECT  104100.0 1439850.0 105300.0 1441800.0 ;
      RECT  104100.0 1428000.0 105300.0 1429950.0 ;
      RECT  94500.0 1438650.0 95700.0 1439850.0 ;
      RECT  96900.0 1438650.0 98100.0 1439850.0 ;
      RECT  96900.0 1438650.0 98100.0 1439850.0 ;
      RECT  94500.0 1438650.0 95700.0 1439850.0 ;
      RECT  96900.0 1438650.0 98100.0 1439850.0 ;
      RECT  99300.0 1438650.0 100500.0 1439850.0 ;
      RECT  99300.0 1438650.0 100500.0 1439850.0 ;
      RECT  96900.0 1438650.0 98100.0 1439850.0 ;
      RECT  99300.0 1438650.0 100500.0 1439850.0 ;
      RECT  101700.0 1438650.0 102900.0 1439850.0 ;
      RECT  101700.0 1438650.0 102900.0 1439850.0 ;
      RECT  99300.0 1438650.0 100500.0 1439850.0 ;
      RECT  94500.0 1429950.0 95700.0 1431150.0 ;
      RECT  96900.0 1429950.0 98100.0 1431150.0 ;
      RECT  96900.0 1429950.0 98100.0 1431150.0 ;
      RECT  94500.0 1429950.0 95700.0 1431150.0 ;
      RECT  96900.0 1429950.0 98100.0 1431150.0 ;
      RECT  99300.0 1429950.0 100500.0 1431150.0 ;
      RECT  99300.0 1429950.0 100500.0 1431150.0 ;
      RECT  96900.0 1429950.0 98100.0 1431150.0 ;
      RECT  99300.0 1429950.0 100500.0 1431150.0 ;
      RECT  101700.0 1429950.0 102900.0 1431150.0 ;
      RECT  101700.0 1429950.0 102900.0 1431150.0 ;
      RECT  99300.0 1429950.0 100500.0 1431150.0 ;
      RECT  104100.0 1439250.0 105300.0 1440450.0 ;
      RECT  104100.0 1429350.0 105300.0 1430550.0 ;
      RECT  101700.0 1432050.0 100500.0 1433250.0 ;
      RECT  99300.0 1434000.0 98100.0 1435200.0 ;
      RECT  96900.0 1435950.0 95700.0 1437150.0 ;
      RECT  96900.0 1438650.0 98100.0 1439850.0 ;
      RECT  101700.0 1438650.0 102900.0 1439850.0 ;
      RECT  101700.0 1429950.0 102900.0 1431150.0 ;
      RECT  101700.0 1435950.0 102900.0 1437150.0 ;
      RECT  95700.0 1435950.0 96900.0 1437150.0 ;
      RECT  98100.0 1434000.0 99300.0 1435200.0 ;
      RECT  100500.0 1432050.0 101700.0 1433250.0 ;
      RECT  101700.0 1435950.0 102900.0 1437150.0 ;
      RECT  92700.0 1441350.0 108300.0 1442250.0 ;
      RECT  92700.0 1427550.0 108300.0 1428450.0 ;
      RECT  94500.0 1453650.0 95700.0 1456050.0 ;
      RECT  94500.0 1444950.0 95700.0 1441350.0 ;
      RECT  99300.0 1444950.0 100500.0 1441350.0 ;
      RECT  104100.0 1443750.0 105300.0 1441800.0 ;
      RECT  104100.0 1455600.0 105300.0 1453650.0 ;
      RECT  94500.0 1444950.0 95700.0 1443750.0 ;
      RECT  96900.0 1444950.0 98100.0 1443750.0 ;
      RECT  96900.0 1444950.0 98100.0 1443750.0 ;
      RECT  94500.0 1444950.0 95700.0 1443750.0 ;
      RECT  96900.0 1444950.0 98100.0 1443750.0 ;
      RECT  99300.0 1444950.0 100500.0 1443750.0 ;
      RECT  99300.0 1444950.0 100500.0 1443750.0 ;
      RECT  96900.0 1444950.0 98100.0 1443750.0 ;
      RECT  99300.0 1444950.0 100500.0 1443750.0 ;
      RECT  101700.0 1444950.0 102900.0 1443750.0 ;
      RECT  101700.0 1444950.0 102900.0 1443750.0 ;
      RECT  99300.0 1444950.0 100500.0 1443750.0 ;
      RECT  94500.0 1453650.0 95700.0 1452450.0 ;
      RECT  96900.0 1453650.0 98100.0 1452450.0 ;
      RECT  96900.0 1453650.0 98100.0 1452450.0 ;
      RECT  94500.0 1453650.0 95700.0 1452450.0 ;
      RECT  96900.0 1453650.0 98100.0 1452450.0 ;
      RECT  99300.0 1453650.0 100500.0 1452450.0 ;
      RECT  99300.0 1453650.0 100500.0 1452450.0 ;
      RECT  96900.0 1453650.0 98100.0 1452450.0 ;
      RECT  99300.0 1453650.0 100500.0 1452450.0 ;
      RECT  101700.0 1453650.0 102900.0 1452450.0 ;
      RECT  101700.0 1453650.0 102900.0 1452450.0 ;
      RECT  99300.0 1453650.0 100500.0 1452450.0 ;
      RECT  104100.0 1444350.0 105300.0 1443150.0 ;
      RECT  104100.0 1454250.0 105300.0 1453050.0 ;
      RECT  101700.0 1451550.0 100500.0 1450350.0 ;
      RECT  99300.0 1449600.0 98100.0 1448400.0 ;
      RECT  96900.0 1447650.0 95700.0 1446450.0 ;
      RECT  96900.0 1444950.0 98100.0 1443750.0 ;
      RECT  101700.0 1444950.0 102900.0 1443750.0 ;
      RECT  101700.0 1453650.0 102900.0 1452450.0 ;
      RECT  101700.0 1447650.0 102900.0 1446450.0 ;
      RECT  95700.0 1447650.0 96900.0 1446450.0 ;
      RECT  98100.0 1449600.0 99300.0 1448400.0 ;
      RECT  100500.0 1451550.0 101700.0 1450350.0 ;
      RECT  101700.0 1447650.0 102900.0 1446450.0 ;
      RECT  92700.0 1442250.0 108300.0 1441350.0 ;
      RECT  92700.0 1456050.0 108300.0 1455150.0 ;
      RECT  94500.0 1457550.0 95700.0 1455150.0 ;
      RECT  94500.0 1466250.0 95700.0 1469850.0 ;
      RECT  99300.0 1466250.0 100500.0 1469850.0 ;
      RECT  104100.0 1467450.0 105300.0 1469400.0 ;
      RECT  104100.0 1455600.0 105300.0 1457550.0 ;
      RECT  94500.0 1466250.0 95700.0 1467450.0 ;
      RECT  96900.0 1466250.0 98100.0 1467450.0 ;
      RECT  96900.0 1466250.0 98100.0 1467450.0 ;
      RECT  94500.0 1466250.0 95700.0 1467450.0 ;
      RECT  96900.0 1466250.0 98100.0 1467450.0 ;
      RECT  99300.0 1466250.0 100500.0 1467450.0 ;
      RECT  99300.0 1466250.0 100500.0 1467450.0 ;
      RECT  96900.0 1466250.0 98100.0 1467450.0 ;
      RECT  99300.0 1466250.0 100500.0 1467450.0 ;
      RECT  101700.0 1466250.0 102900.0 1467450.0 ;
      RECT  101700.0 1466250.0 102900.0 1467450.0 ;
      RECT  99300.0 1466250.0 100500.0 1467450.0 ;
      RECT  94500.0 1457550.0 95700.0 1458750.0 ;
      RECT  96900.0 1457550.0 98100.0 1458750.0 ;
      RECT  96900.0 1457550.0 98100.0 1458750.0 ;
      RECT  94500.0 1457550.0 95700.0 1458750.0 ;
      RECT  96900.0 1457550.0 98100.0 1458750.0 ;
      RECT  99300.0 1457550.0 100500.0 1458750.0 ;
      RECT  99300.0 1457550.0 100500.0 1458750.0 ;
      RECT  96900.0 1457550.0 98100.0 1458750.0 ;
      RECT  99300.0 1457550.0 100500.0 1458750.0 ;
      RECT  101700.0 1457550.0 102900.0 1458750.0 ;
      RECT  101700.0 1457550.0 102900.0 1458750.0 ;
      RECT  99300.0 1457550.0 100500.0 1458750.0 ;
      RECT  104100.0 1466850.0 105300.0 1468050.0 ;
      RECT  104100.0 1456950.0 105300.0 1458150.0 ;
      RECT  101700.0 1459650.0 100500.0 1460850.0 ;
      RECT  99300.0 1461600.0 98100.0 1462800.0 ;
      RECT  96900.0 1463550.0 95700.0 1464750.0 ;
      RECT  96900.0 1466250.0 98100.0 1467450.0 ;
      RECT  101700.0 1466250.0 102900.0 1467450.0 ;
      RECT  101700.0 1457550.0 102900.0 1458750.0 ;
      RECT  101700.0 1463550.0 102900.0 1464750.0 ;
      RECT  95700.0 1463550.0 96900.0 1464750.0 ;
      RECT  98100.0 1461600.0 99300.0 1462800.0 ;
      RECT  100500.0 1459650.0 101700.0 1460850.0 ;
      RECT  101700.0 1463550.0 102900.0 1464750.0 ;
      RECT  92700.0 1468950.0 108300.0 1469850.0 ;
      RECT  92700.0 1455150.0 108300.0 1456050.0 ;
      RECT  94500.0 1481250.0 95700.0 1483650.0 ;
      RECT  94500.0 1472550.0 95700.0 1468950.0 ;
      RECT  99300.0 1472550.0 100500.0 1468950.0 ;
      RECT  104100.0 1471350.0 105300.0 1469400.0 ;
      RECT  104100.0 1483200.0 105300.0 1481250.0 ;
      RECT  94500.0 1472550.0 95700.0 1471350.0 ;
      RECT  96900.0 1472550.0 98100.0 1471350.0 ;
      RECT  96900.0 1472550.0 98100.0 1471350.0 ;
      RECT  94500.0 1472550.0 95700.0 1471350.0 ;
      RECT  96900.0 1472550.0 98100.0 1471350.0 ;
      RECT  99300.0 1472550.0 100500.0 1471350.0 ;
      RECT  99300.0 1472550.0 100500.0 1471350.0 ;
      RECT  96900.0 1472550.0 98100.0 1471350.0 ;
      RECT  99300.0 1472550.0 100500.0 1471350.0 ;
      RECT  101700.0 1472550.0 102900.0 1471350.0 ;
      RECT  101700.0 1472550.0 102900.0 1471350.0 ;
      RECT  99300.0 1472550.0 100500.0 1471350.0 ;
      RECT  94500.0 1481250.0 95700.0 1480050.0 ;
      RECT  96900.0 1481250.0 98100.0 1480050.0 ;
      RECT  96900.0 1481250.0 98100.0 1480050.0 ;
      RECT  94500.0 1481250.0 95700.0 1480050.0 ;
      RECT  96900.0 1481250.0 98100.0 1480050.0 ;
      RECT  99300.0 1481250.0 100500.0 1480050.0 ;
      RECT  99300.0 1481250.0 100500.0 1480050.0 ;
      RECT  96900.0 1481250.0 98100.0 1480050.0 ;
      RECT  99300.0 1481250.0 100500.0 1480050.0 ;
      RECT  101700.0 1481250.0 102900.0 1480050.0 ;
      RECT  101700.0 1481250.0 102900.0 1480050.0 ;
      RECT  99300.0 1481250.0 100500.0 1480050.0 ;
      RECT  104100.0 1471950.0 105300.0 1470750.0 ;
      RECT  104100.0 1481850.0 105300.0 1480650.0 ;
      RECT  101700.0 1479150.0 100500.0 1477950.0 ;
      RECT  99300.0 1477200.0 98100.0 1476000.0 ;
      RECT  96900.0 1475250.0 95700.0 1474050.0 ;
      RECT  96900.0 1472550.0 98100.0 1471350.0 ;
      RECT  101700.0 1472550.0 102900.0 1471350.0 ;
      RECT  101700.0 1481250.0 102900.0 1480050.0 ;
      RECT  101700.0 1475250.0 102900.0 1474050.0 ;
      RECT  95700.0 1475250.0 96900.0 1474050.0 ;
      RECT  98100.0 1477200.0 99300.0 1476000.0 ;
      RECT  100500.0 1479150.0 101700.0 1477950.0 ;
      RECT  101700.0 1475250.0 102900.0 1474050.0 ;
      RECT  92700.0 1469850.0 108300.0 1468950.0 ;
      RECT  92700.0 1483650.0 108300.0 1482750.0 ;
      RECT  94500.0 1485150.0 95700.0 1482750.0 ;
      RECT  94500.0 1493850.0 95700.0 1497450.0 ;
      RECT  99300.0 1493850.0 100500.0 1497450.0 ;
      RECT  104100.0 1495050.0 105300.0 1497000.0 ;
      RECT  104100.0 1483200.0 105300.0 1485150.0 ;
      RECT  94500.0 1493850.0 95700.0 1495050.0 ;
      RECT  96900.0 1493850.0 98100.0 1495050.0 ;
      RECT  96900.0 1493850.0 98100.0 1495050.0 ;
      RECT  94500.0 1493850.0 95700.0 1495050.0 ;
      RECT  96900.0 1493850.0 98100.0 1495050.0 ;
      RECT  99300.0 1493850.0 100500.0 1495050.0 ;
      RECT  99300.0 1493850.0 100500.0 1495050.0 ;
      RECT  96900.0 1493850.0 98100.0 1495050.0 ;
      RECT  99300.0 1493850.0 100500.0 1495050.0 ;
      RECT  101700.0 1493850.0 102900.0 1495050.0 ;
      RECT  101700.0 1493850.0 102900.0 1495050.0 ;
      RECT  99300.0 1493850.0 100500.0 1495050.0 ;
      RECT  94500.0 1485150.0 95700.0 1486350.0 ;
      RECT  96900.0 1485150.0 98100.0 1486350.0 ;
      RECT  96900.0 1485150.0 98100.0 1486350.0 ;
      RECT  94500.0 1485150.0 95700.0 1486350.0 ;
      RECT  96900.0 1485150.0 98100.0 1486350.0 ;
      RECT  99300.0 1485150.0 100500.0 1486350.0 ;
      RECT  99300.0 1485150.0 100500.0 1486350.0 ;
      RECT  96900.0 1485150.0 98100.0 1486350.0 ;
      RECT  99300.0 1485150.0 100500.0 1486350.0 ;
      RECT  101700.0 1485150.0 102900.0 1486350.0 ;
      RECT  101700.0 1485150.0 102900.0 1486350.0 ;
      RECT  99300.0 1485150.0 100500.0 1486350.0 ;
      RECT  104100.0 1494450.0 105300.0 1495650.0 ;
      RECT  104100.0 1484550.0 105300.0 1485750.0 ;
      RECT  101700.0 1487250.0 100500.0 1488450.0 ;
      RECT  99300.0 1489200.0 98100.0 1490400.0 ;
      RECT  96900.0 1491150.0 95700.0 1492350.0 ;
      RECT  96900.0 1493850.0 98100.0 1495050.0 ;
      RECT  101700.0 1493850.0 102900.0 1495050.0 ;
      RECT  101700.0 1485150.0 102900.0 1486350.0 ;
      RECT  101700.0 1491150.0 102900.0 1492350.0 ;
      RECT  95700.0 1491150.0 96900.0 1492350.0 ;
      RECT  98100.0 1489200.0 99300.0 1490400.0 ;
      RECT  100500.0 1487250.0 101700.0 1488450.0 ;
      RECT  101700.0 1491150.0 102900.0 1492350.0 ;
      RECT  92700.0 1496550.0 108300.0 1497450.0 ;
      RECT  92700.0 1482750.0 108300.0 1483650.0 ;
      RECT  94500.0 1508850.0 95700.0 1511250.0 ;
      RECT  94500.0 1500150.0 95700.0 1496550.0 ;
      RECT  99300.0 1500150.0 100500.0 1496550.0 ;
      RECT  104100.0 1498950.0 105300.0 1497000.0 ;
      RECT  104100.0 1510800.0 105300.0 1508850.0 ;
      RECT  94500.0 1500150.0 95700.0 1498950.0 ;
      RECT  96900.0 1500150.0 98100.0 1498950.0 ;
      RECT  96900.0 1500150.0 98100.0 1498950.0 ;
      RECT  94500.0 1500150.0 95700.0 1498950.0 ;
      RECT  96900.0 1500150.0 98100.0 1498950.0 ;
      RECT  99300.0 1500150.0 100500.0 1498950.0 ;
      RECT  99300.0 1500150.0 100500.0 1498950.0 ;
      RECT  96900.0 1500150.0 98100.0 1498950.0 ;
      RECT  99300.0 1500150.0 100500.0 1498950.0 ;
      RECT  101700.0 1500150.0 102900.0 1498950.0 ;
      RECT  101700.0 1500150.0 102900.0 1498950.0 ;
      RECT  99300.0 1500150.0 100500.0 1498950.0 ;
      RECT  94500.0 1508850.0 95700.0 1507650.0 ;
      RECT  96900.0 1508850.0 98100.0 1507650.0 ;
      RECT  96900.0 1508850.0 98100.0 1507650.0 ;
      RECT  94500.0 1508850.0 95700.0 1507650.0 ;
      RECT  96900.0 1508850.0 98100.0 1507650.0 ;
      RECT  99300.0 1508850.0 100500.0 1507650.0 ;
      RECT  99300.0 1508850.0 100500.0 1507650.0 ;
      RECT  96900.0 1508850.0 98100.0 1507650.0 ;
      RECT  99300.0 1508850.0 100500.0 1507650.0 ;
      RECT  101700.0 1508850.0 102900.0 1507650.0 ;
      RECT  101700.0 1508850.0 102900.0 1507650.0 ;
      RECT  99300.0 1508850.0 100500.0 1507650.0 ;
      RECT  104100.0 1499550.0 105300.0 1498350.0 ;
      RECT  104100.0 1509450.0 105300.0 1508250.0 ;
      RECT  101700.0 1506750.0 100500.0 1505550.0 ;
      RECT  99300.0 1504800.0 98100.0 1503600.0 ;
      RECT  96900.0 1502850.0 95700.0 1501650.0 ;
      RECT  96900.0 1500150.0 98100.0 1498950.0 ;
      RECT  101700.0 1500150.0 102900.0 1498950.0 ;
      RECT  101700.0 1508850.0 102900.0 1507650.0 ;
      RECT  101700.0 1502850.0 102900.0 1501650.0 ;
      RECT  95700.0 1502850.0 96900.0 1501650.0 ;
      RECT  98100.0 1504800.0 99300.0 1503600.0 ;
      RECT  100500.0 1506750.0 101700.0 1505550.0 ;
      RECT  101700.0 1502850.0 102900.0 1501650.0 ;
      RECT  92700.0 1497450.0 108300.0 1496550.0 ;
      RECT  92700.0 1511250.0 108300.0 1510350.0 ;
      RECT  94500.0 1512750.0 95700.0 1510350.0 ;
      RECT  94500.0 1521450.0 95700.0 1525050.0 ;
      RECT  99300.0 1521450.0 100500.0 1525050.0 ;
      RECT  104100.0 1522650.0 105300.0 1524600.0 ;
      RECT  104100.0 1510800.0 105300.0 1512750.0 ;
      RECT  94500.0 1521450.0 95700.0 1522650.0 ;
      RECT  96900.0 1521450.0 98100.0 1522650.0 ;
      RECT  96900.0 1521450.0 98100.0 1522650.0 ;
      RECT  94500.0 1521450.0 95700.0 1522650.0 ;
      RECT  96900.0 1521450.0 98100.0 1522650.0 ;
      RECT  99300.0 1521450.0 100500.0 1522650.0 ;
      RECT  99300.0 1521450.0 100500.0 1522650.0 ;
      RECT  96900.0 1521450.0 98100.0 1522650.0 ;
      RECT  99300.0 1521450.0 100500.0 1522650.0 ;
      RECT  101700.0 1521450.0 102900.0 1522650.0 ;
      RECT  101700.0 1521450.0 102900.0 1522650.0 ;
      RECT  99300.0 1521450.0 100500.0 1522650.0 ;
      RECT  94500.0 1512750.0 95700.0 1513950.0 ;
      RECT  96900.0 1512750.0 98100.0 1513950.0 ;
      RECT  96900.0 1512750.0 98100.0 1513950.0 ;
      RECT  94500.0 1512750.0 95700.0 1513950.0 ;
      RECT  96900.0 1512750.0 98100.0 1513950.0 ;
      RECT  99300.0 1512750.0 100500.0 1513950.0 ;
      RECT  99300.0 1512750.0 100500.0 1513950.0 ;
      RECT  96900.0 1512750.0 98100.0 1513950.0 ;
      RECT  99300.0 1512750.0 100500.0 1513950.0 ;
      RECT  101700.0 1512750.0 102900.0 1513950.0 ;
      RECT  101700.0 1512750.0 102900.0 1513950.0 ;
      RECT  99300.0 1512750.0 100500.0 1513950.0 ;
      RECT  104100.0 1522050.0 105300.0 1523250.0 ;
      RECT  104100.0 1512150.0 105300.0 1513350.0 ;
      RECT  101700.0 1514850.0 100500.0 1516050.0 ;
      RECT  99300.0 1516800.0 98100.0 1518000.0 ;
      RECT  96900.0 1518750.0 95700.0 1519950.0 ;
      RECT  96900.0 1521450.0 98100.0 1522650.0 ;
      RECT  101700.0 1521450.0 102900.0 1522650.0 ;
      RECT  101700.0 1512750.0 102900.0 1513950.0 ;
      RECT  101700.0 1518750.0 102900.0 1519950.0 ;
      RECT  95700.0 1518750.0 96900.0 1519950.0 ;
      RECT  98100.0 1516800.0 99300.0 1518000.0 ;
      RECT  100500.0 1514850.0 101700.0 1516050.0 ;
      RECT  101700.0 1518750.0 102900.0 1519950.0 ;
      RECT  92700.0 1524150.0 108300.0 1525050.0 ;
      RECT  92700.0 1510350.0 108300.0 1511250.0 ;
      RECT  94500.0 1536450.0 95700.0 1538850.0 ;
      RECT  94500.0 1527750.0 95700.0 1524150.0 ;
      RECT  99300.0 1527750.0 100500.0 1524150.0 ;
      RECT  104100.0 1526550.0 105300.0 1524600.0 ;
      RECT  104100.0 1538400.0 105300.0 1536450.0 ;
      RECT  94500.0 1527750.0 95700.0 1526550.0 ;
      RECT  96900.0 1527750.0 98100.0 1526550.0 ;
      RECT  96900.0 1527750.0 98100.0 1526550.0 ;
      RECT  94500.0 1527750.0 95700.0 1526550.0 ;
      RECT  96900.0 1527750.0 98100.0 1526550.0 ;
      RECT  99300.0 1527750.0 100500.0 1526550.0 ;
      RECT  99300.0 1527750.0 100500.0 1526550.0 ;
      RECT  96900.0 1527750.0 98100.0 1526550.0 ;
      RECT  99300.0 1527750.0 100500.0 1526550.0 ;
      RECT  101700.0 1527750.0 102900.0 1526550.0 ;
      RECT  101700.0 1527750.0 102900.0 1526550.0 ;
      RECT  99300.0 1527750.0 100500.0 1526550.0 ;
      RECT  94500.0 1536450.0 95700.0 1535250.0 ;
      RECT  96900.0 1536450.0 98100.0 1535250.0 ;
      RECT  96900.0 1536450.0 98100.0 1535250.0 ;
      RECT  94500.0 1536450.0 95700.0 1535250.0 ;
      RECT  96900.0 1536450.0 98100.0 1535250.0 ;
      RECT  99300.0 1536450.0 100500.0 1535250.0 ;
      RECT  99300.0 1536450.0 100500.0 1535250.0 ;
      RECT  96900.0 1536450.0 98100.0 1535250.0 ;
      RECT  99300.0 1536450.0 100500.0 1535250.0 ;
      RECT  101700.0 1536450.0 102900.0 1535250.0 ;
      RECT  101700.0 1536450.0 102900.0 1535250.0 ;
      RECT  99300.0 1536450.0 100500.0 1535250.0 ;
      RECT  104100.0 1527150.0 105300.0 1525950.0 ;
      RECT  104100.0 1537050.0 105300.0 1535850.0 ;
      RECT  101700.0 1534350.0 100500.0 1533150.0 ;
      RECT  99300.0 1532400.0 98100.0 1531200.0 ;
      RECT  96900.0 1530450.0 95700.0 1529250.0 ;
      RECT  96900.0 1527750.0 98100.0 1526550.0 ;
      RECT  101700.0 1527750.0 102900.0 1526550.0 ;
      RECT  101700.0 1536450.0 102900.0 1535250.0 ;
      RECT  101700.0 1530450.0 102900.0 1529250.0 ;
      RECT  95700.0 1530450.0 96900.0 1529250.0 ;
      RECT  98100.0 1532400.0 99300.0 1531200.0 ;
      RECT  100500.0 1534350.0 101700.0 1533150.0 ;
      RECT  101700.0 1530450.0 102900.0 1529250.0 ;
      RECT  92700.0 1525050.0 108300.0 1524150.0 ;
      RECT  92700.0 1538850.0 108300.0 1537950.0 ;
      RECT  94500.0 1540350.0 95700.0 1537950.0 ;
      RECT  94500.0 1549050.0 95700.0 1552650.0 ;
      RECT  99300.0 1549050.0 100500.0 1552650.0 ;
      RECT  104100.0 1550250.0 105300.0 1552200.0 ;
      RECT  104100.0 1538400.0 105300.0 1540350.0 ;
      RECT  94500.0 1549050.0 95700.0 1550250.0 ;
      RECT  96900.0 1549050.0 98100.0 1550250.0 ;
      RECT  96900.0 1549050.0 98100.0 1550250.0 ;
      RECT  94500.0 1549050.0 95700.0 1550250.0 ;
      RECT  96900.0 1549050.0 98100.0 1550250.0 ;
      RECT  99300.0 1549050.0 100500.0 1550250.0 ;
      RECT  99300.0 1549050.0 100500.0 1550250.0 ;
      RECT  96900.0 1549050.0 98100.0 1550250.0 ;
      RECT  99300.0 1549050.0 100500.0 1550250.0 ;
      RECT  101700.0 1549050.0 102900.0 1550250.0 ;
      RECT  101700.0 1549050.0 102900.0 1550250.0 ;
      RECT  99300.0 1549050.0 100500.0 1550250.0 ;
      RECT  94500.0 1540350.0 95700.0 1541550.0 ;
      RECT  96900.0 1540350.0 98100.0 1541550.0 ;
      RECT  96900.0 1540350.0 98100.0 1541550.0 ;
      RECT  94500.0 1540350.0 95700.0 1541550.0 ;
      RECT  96900.0 1540350.0 98100.0 1541550.0 ;
      RECT  99300.0 1540350.0 100500.0 1541550.0 ;
      RECT  99300.0 1540350.0 100500.0 1541550.0 ;
      RECT  96900.0 1540350.0 98100.0 1541550.0 ;
      RECT  99300.0 1540350.0 100500.0 1541550.0 ;
      RECT  101700.0 1540350.0 102900.0 1541550.0 ;
      RECT  101700.0 1540350.0 102900.0 1541550.0 ;
      RECT  99300.0 1540350.0 100500.0 1541550.0 ;
      RECT  104100.0 1549650.0 105300.0 1550850.0 ;
      RECT  104100.0 1539750.0 105300.0 1540950.0 ;
      RECT  101700.0 1542450.0 100500.0 1543650.0 ;
      RECT  99300.0 1544400.0 98100.0 1545600.0 ;
      RECT  96900.0 1546350.0 95700.0 1547550.0 ;
      RECT  96900.0 1549050.0 98100.0 1550250.0 ;
      RECT  101700.0 1549050.0 102900.0 1550250.0 ;
      RECT  101700.0 1540350.0 102900.0 1541550.0 ;
      RECT  101700.0 1546350.0 102900.0 1547550.0 ;
      RECT  95700.0 1546350.0 96900.0 1547550.0 ;
      RECT  98100.0 1544400.0 99300.0 1545600.0 ;
      RECT  100500.0 1542450.0 101700.0 1543650.0 ;
      RECT  101700.0 1546350.0 102900.0 1547550.0 ;
      RECT  92700.0 1551750.0 108300.0 1552650.0 ;
      RECT  92700.0 1537950.0 108300.0 1538850.0 ;
      RECT  94500.0 1564050.0 95700.0 1566450.0 ;
      RECT  94500.0 1555350.0 95700.0 1551750.0 ;
      RECT  99300.0 1555350.0 100500.0 1551750.0 ;
      RECT  104100.0 1554150.0 105300.0 1552200.0 ;
      RECT  104100.0 1566000.0 105300.0 1564050.0 ;
      RECT  94500.0 1555350.0 95700.0 1554150.0 ;
      RECT  96900.0 1555350.0 98100.0 1554150.0 ;
      RECT  96900.0 1555350.0 98100.0 1554150.0 ;
      RECT  94500.0 1555350.0 95700.0 1554150.0 ;
      RECT  96900.0 1555350.0 98100.0 1554150.0 ;
      RECT  99300.0 1555350.0 100500.0 1554150.0 ;
      RECT  99300.0 1555350.0 100500.0 1554150.0 ;
      RECT  96900.0 1555350.0 98100.0 1554150.0 ;
      RECT  99300.0 1555350.0 100500.0 1554150.0 ;
      RECT  101700.0 1555350.0 102900.0 1554150.0 ;
      RECT  101700.0 1555350.0 102900.0 1554150.0 ;
      RECT  99300.0 1555350.0 100500.0 1554150.0 ;
      RECT  94500.0 1564050.0 95700.0 1562850.0 ;
      RECT  96900.0 1564050.0 98100.0 1562850.0 ;
      RECT  96900.0 1564050.0 98100.0 1562850.0 ;
      RECT  94500.0 1564050.0 95700.0 1562850.0 ;
      RECT  96900.0 1564050.0 98100.0 1562850.0 ;
      RECT  99300.0 1564050.0 100500.0 1562850.0 ;
      RECT  99300.0 1564050.0 100500.0 1562850.0 ;
      RECT  96900.0 1564050.0 98100.0 1562850.0 ;
      RECT  99300.0 1564050.0 100500.0 1562850.0 ;
      RECT  101700.0 1564050.0 102900.0 1562850.0 ;
      RECT  101700.0 1564050.0 102900.0 1562850.0 ;
      RECT  99300.0 1564050.0 100500.0 1562850.0 ;
      RECT  104100.0 1554750.0 105300.0 1553550.0 ;
      RECT  104100.0 1564650.0 105300.0 1563450.0 ;
      RECT  101700.0 1561950.0 100500.0 1560750.0 ;
      RECT  99300.0 1560000.0 98100.0 1558800.0 ;
      RECT  96900.0 1558050.0 95700.0 1556850.0 ;
      RECT  96900.0 1555350.0 98100.0 1554150.0 ;
      RECT  101700.0 1555350.0 102900.0 1554150.0 ;
      RECT  101700.0 1564050.0 102900.0 1562850.0 ;
      RECT  101700.0 1558050.0 102900.0 1556850.0 ;
      RECT  95700.0 1558050.0 96900.0 1556850.0 ;
      RECT  98100.0 1560000.0 99300.0 1558800.0 ;
      RECT  100500.0 1561950.0 101700.0 1560750.0 ;
      RECT  101700.0 1558050.0 102900.0 1556850.0 ;
      RECT  92700.0 1552650.0 108300.0 1551750.0 ;
      RECT  92700.0 1566450.0 108300.0 1565550.0 ;
      RECT  94500.0 1567950.0 95700.0 1565550.0 ;
      RECT  94500.0 1576650.0 95700.0 1580250.0 ;
      RECT  99300.0 1576650.0 100500.0 1580250.0 ;
      RECT  104100.0 1577850.0 105300.0 1579800.0 ;
      RECT  104100.0 1566000.0 105300.0 1567950.0 ;
      RECT  94500.0 1576650.0 95700.0 1577850.0 ;
      RECT  96900.0 1576650.0 98100.0 1577850.0 ;
      RECT  96900.0 1576650.0 98100.0 1577850.0 ;
      RECT  94500.0 1576650.0 95700.0 1577850.0 ;
      RECT  96900.0 1576650.0 98100.0 1577850.0 ;
      RECT  99300.0 1576650.0 100500.0 1577850.0 ;
      RECT  99300.0 1576650.0 100500.0 1577850.0 ;
      RECT  96900.0 1576650.0 98100.0 1577850.0 ;
      RECT  99300.0 1576650.0 100500.0 1577850.0 ;
      RECT  101700.0 1576650.0 102900.0 1577850.0 ;
      RECT  101700.0 1576650.0 102900.0 1577850.0 ;
      RECT  99300.0 1576650.0 100500.0 1577850.0 ;
      RECT  94500.0 1567950.0 95700.0 1569150.0 ;
      RECT  96900.0 1567950.0 98100.0 1569150.0 ;
      RECT  96900.0 1567950.0 98100.0 1569150.0 ;
      RECT  94500.0 1567950.0 95700.0 1569150.0 ;
      RECT  96900.0 1567950.0 98100.0 1569150.0 ;
      RECT  99300.0 1567950.0 100500.0 1569150.0 ;
      RECT  99300.0 1567950.0 100500.0 1569150.0 ;
      RECT  96900.0 1567950.0 98100.0 1569150.0 ;
      RECT  99300.0 1567950.0 100500.0 1569150.0 ;
      RECT  101700.0 1567950.0 102900.0 1569150.0 ;
      RECT  101700.0 1567950.0 102900.0 1569150.0 ;
      RECT  99300.0 1567950.0 100500.0 1569150.0 ;
      RECT  104100.0 1577250.0 105300.0 1578450.0 ;
      RECT  104100.0 1567350.0 105300.0 1568550.0 ;
      RECT  101700.0 1570050.0 100500.0 1571250.0 ;
      RECT  99300.0 1572000.0 98100.0 1573200.0 ;
      RECT  96900.0 1573950.0 95700.0 1575150.0 ;
      RECT  96900.0 1576650.0 98100.0 1577850.0 ;
      RECT  101700.0 1576650.0 102900.0 1577850.0 ;
      RECT  101700.0 1567950.0 102900.0 1569150.0 ;
      RECT  101700.0 1573950.0 102900.0 1575150.0 ;
      RECT  95700.0 1573950.0 96900.0 1575150.0 ;
      RECT  98100.0 1572000.0 99300.0 1573200.0 ;
      RECT  100500.0 1570050.0 101700.0 1571250.0 ;
      RECT  101700.0 1573950.0 102900.0 1575150.0 ;
      RECT  92700.0 1579350.0 108300.0 1580250.0 ;
      RECT  92700.0 1565550.0 108300.0 1566450.0 ;
      RECT  94500.0 1591650.0 95700.0 1594050.0 ;
      RECT  94500.0 1582950.0 95700.0 1579350.0 ;
      RECT  99300.0 1582950.0 100500.0 1579350.0 ;
      RECT  104100.0 1581750.0 105300.0 1579800.0 ;
      RECT  104100.0 1593600.0 105300.0 1591650.0 ;
      RECT  94500.0 1582950.0 95700.0 1581750.0 ;
      RECT  96900.0 1582950.0 98100.0 1581750.0 ;
      RECT  96900.0 1582950.0 98100.0 1581750.0 ;
      RECT  94500.0 1582950.0 95700.0 1581750.0 ;
      RECT  96900.0 1582950.0 98100.0 1581750.0 ;
      RECT  99300.0 1582950.0 100500.0 1581750.0 ;
      RECT  99300.0 1582950.0 100500.0 1581750.0 ;
      RECT  96900.0 1582950.0 98100.0 1581750.0 ;
      RECT  99300.0 1582950.0 100500.0 1581750.0 ;
      RECT  101700.0 1582950.0 102900.0 1581750.0 ;
      RECT  101700.0 1582950.0 102900.0 1581750.0 ;
      RECT  99300.0 1582950.0 100500.0 1581750.0 ;
      RECT  94500.0 1591650.0 95700.0 1590450.0 ;
      RECT  96900.0 1591650.0 98100.0 1590450.0 ;
      RECT  96900.0 1591650.0 98100.0 1590450.0 ;
      RECT  94500.0 1591650.0 95700.0 1590450.0 ;
      RECT  96900.0 1591650.0 98100.0 1590450.0 ;
      RECT  99300.0 1591650.0 100500.0 1590450.0 ;
      RECT  99300.0 1591650.0 100500.0 1590450.0 ;
      RECT  96900.0 1591650.0 98100.0 1590450.0 ;
      RECT  99300.0 1591650.0 100500.0 1590450.0 ;
      RECT  101700.0 1591650.0 102900.0 1590450.0 ;
      RECT  101700.0 1591650.0 102900.0 1590450.0 ;
      RECT  99300.0 1591650.0 100500.0 1590450.0 ;
      RECT  104100.0 1582350.0 105300.0 1581150.0 ;
      RECT  104100.0 1592250.0 105300.0 1591050.0 ;
      RECT  101700.0 1589550.0 100500.0 1588350.0 ;
      RECT  99300.0 1587600.0 98100.0 1586400.0 ;
      RECT  96900.0 1585650.0 95700.0 1584450.0 ;
      RECT  96900.0 1582950.0 98100.0 1581750.0 ;
      RECT  101700.0 1582950.0 102900.0 1581750.0 ;
      RECT  101700.0 1591650.0 102900.0 1590450.0 ;
      RECT  101700.0 1585650.0 102900.0 1584450.0 ;
      RECT  95700.0 1585650.0 96900.0 1584450.0 ;
      RECT  98100.0 1587600.0 99300.0 1586400.0 ;
      RECT  100500.0 1589550.0 101700.0 1588350.0 ;
      RECT  101700.0 1585650.0 102900.0 1584450.0 ;
      RECT  92700.0 1580250.0 108300.0 1579350.0 ;
      RECT  92700.0 1594050.0 108300.0 1593150.0 ;
      RECT  94500.0 1595550.0 95700.0 1593150.0 ;
      RECT  94500.0 1604250.0 95700.0 1607850.0 ;
      RECT  99300.0 1604250.0 100500.0 1607850.0 ;
      RECT  104100.0 1605450.0 105300.0 1607400.0 ;
      RECT  104100.0 1593600.0 105300.0 1595550.0 ;
      RECT  94500.0 1604250.0 95700.0 1605450.0 ;
      RECT  96900.0 1604250.0 98100.0 1605450.0 ;
      RECT  96900.0 1604250.0 98100.0 1605450.0 ;
      RECT  94500.0 1604250.0 95700.0 1605450.0 ;
      RECT  96900.0 1604250.0 98100.0 1605450.0 ;
      RECT  99300.0 1604250.0 100500.0 1605450.0 ;
      RECT  99300.0 1604250.0 100500.0 1605450.0 ;
      RECT  96900.0 1604250.0 98100.0 1605450.0 ;
      RECT  99300.0 1604250.0 100500.0 1605450.0 ;
      RECT  101700.0 1604250.0 102900.0 1605450.0 ;
      RECT  101700.0 1604250.0 102900.0 1605450.0 ;
      RECT  99300.0 1604250.0 100500.0 1605450.0 ;
      RECT  94500.0 1595550.0 95700.0 1596750.0 ;
      RECT  96900.0 1595550.0 98100.0 1596750.0 ;
      RECT  96900.0 1595550.0 98100.0 1596750.0 ;
      RECT  94500.0 1595550.0 95700.0 1596750.0 ;
      RECT  96900.0 1595550.0 98100.0 1596750.0 ;
      RECT  99300.0 1595550.0 100500.0 1596750.0 ;
      RECT  99300.0 1595550.0 100500.0 1596750.0 ;
      RECT  96900.0 1595550.0 98100.0 1596750.0 ;
      RECT  99300.0 1595550.0 100500.0 1596750.0 ;
      RECT  101700.0 1595550.0 102900.0 1596750.0 ;
      RECT  101700.0 1595550.0 102900.0 1596750.0 ;
      RECT  99300.0 1595550.0 100500.0 1596750.0 ;
      RECT  104100.0 1604850.0 105300.0 1606050.0 ;
      RECT  104100.0 1594950.0 105300.0 1596150.0 ;
      RECT  101700.0 1597650.0 100500.0 1598850.0 ;
      RECT  99300.0 1599600.0 98100.0 1600800.0 ;
      RECT  96900.0 1601550.0 95700.0 1602750.0 ;
      RECT  96900.0 1604250.0 98100.0 1605450.0 ;
      RECT  101700.0 1604250.0 102900.0 1605450.0 ;
      RECT  101700.0 1595550.0 102900.0 1596750.0 ;
      RECT  101700.0 1601550.0 102900.0 1602750.0 ;
      RECT  95700.0 1601550.0 96900.0 1602750.0 ;
      RECT  98100.0 1599600.0 99300.0 1600800.0 ;
      RECT  100500.0 1597650.0 101700.0 1598850.0 ;
      RECT  101700.0 1601550.0 102900.0 1602750.0 ;
      RECT  92700.0 1606950.0 108300.0 1607850.0 ;
      RECT  92700.0 1593150.0 108300.0 1594050.0 ;
      RECT  94500.0 1619250.0 95700.0 1621650.0 ;
      RECT  94500.0 1610550.0 95700.0 1606950.0 ;
      RECT  99300.0 1610550.0 100500.0 1606950.0 ;
      RECT  104100.0 1609350.0 105300.0 1607400.0 ;
      RECT  104100.0 1621200.0 105300.0 1619250.0 ;
      RECT  94500.0 1610550.0 95700.0 1609350.0 ;
      RECT  96900.0 1610550.0 98100.0 1609350.0 ;
      RECT  96900.0 1610550.0 98100.0 1609350.0 ;
      RECT  94500.0 1610550.0 95700.0 1609350.0 ;
      RECT  96900.0 1610550.0 98100.0 1609350.0 ;
      RECT  99300.0 1610550.0 100500.0 1609350.0 ;
      RECT  99300.0 1610550.0 100500.0 1609350.0 ;
      RECT  96900.0 1610550.0 98100.0 1609350.0 ;
      RECT  99300.0 1610550.0 100500.0 1609350.0 ;
      RECT  101700.0 1610550.0 102900.0 1609350.0 ;
      RECT  101700.0 1610550.0 102900.0 1609350.0 ;
      RECT  99300.0 1610550.0 100500.0 1609350.0 ;
      RECT  94500.0 1619250.0 95700.0 1618050.0 ;
      RECT  96900.0 1619250.0 98100.0 1618050.0 ;
      RECT  96900.0 1619250.0 98100.0 1618050.0 ;
      RECT  94500.0 1619250.0 95700.0 1618050.0 ;
      RECT  96900.0 1619250.0 98100.0 1618050.0 ;
      RECT  99300.0 1619250.0 100500.0 1618050.0 ;
      RECT  99300.0 1619250.0 100500.0 1618050.0 ;
      RECT  96900.0 1619250.0 98100.0 1618050.0 ;
      RECT  99300.0 1619250.0 100500.0 1618050.0 ;
      RECT  101700.0 1619250.0 102900.0 1618050.0 ;
      RECT  101700.0 1619250.0 102900.0 1618050.0 ;
      RECT  99300.0 1619250.0 100500.0 1618050.0 ;
      RECT  104100.0 1609950.0 105300.0 1608750.0 ;
      RECT  104100.0 1619850.0 105300.0 1618650.0 ;
      RECT  101700.0 1617150.0 100500.0 1615950.0 ;
      RECT  99300.0 1615200.0 98100.0 1614000.0 ;
      RECT  96900.0 1613250.0 95700.0 1612050.0 ;
      RECT  96900.0 1610550.0 98100.0 1609350.0 ;
      RECT  101700.0 1610550.0 102900.0 1609350.0 ;
      RECT  101700.0 1619250.0 102900.0 1618050.0 ;
      RECT  101700.0 1613250.0 102900.0 1612050.0 ;
      RECT  95700.0 1613250.0 96900.0 1612050.0 ;
      RECT  98100.0 1615200.0 99300.0 1614000.0 ;
      RECT  100500.0 1617150.0 101700.0 1615950.0 ;
      RECT  101700.0 1613250.0 102900.0 1612050.0 ;
      RECT  92700.0 1607850.0 108300.0 1606950.0 ;
      RECT  92700.0 1621650.0 108300.0 1620750.0 ;
      RECT  94500.0 1623150.0 95700.0 1620750.0 ;
      RECT  94500.0 1631850.0 95700.0 1635450.0 ;
      RECT  99300.0 1631850.0 100500.0 1635450.0 ;
      RECT  104100.0 1633050.0 105300.0 1635000.0 ;
      RECT  104100.0 1621200.0 105300.0 1623150.0 ;
      RECT  94500.0 1631850.0 95700.0 1633050.0 ;
      RECT  96900.0 1631850.0 98100.0 1633050.0 ;
      RECT  96900.0 1631850.0 98100.0 1633050.0 ;
      RECT  94500.0 1631850.0 95700.0 1633050.0 ;
      RECT  96900.0 1631850.0 98100.0 1633050.0 ;
      RECT  99300.0 1631850.0 100500.0 1633050.0 ;
      RECT  99300.0 1631850.0 100500.0 1633050.0 ;
      RECT  96900.0 1631850.0 98100.0 1633050.0 ;
      RECT  99300.0 1631850.0 100500.0 1633050.0 ;
      RECT  101700.0 1631850.0 102900.0 1633050.0 ;
      RECT  101700.0 1631850.0 102900.0 1633050.0 ;
      RECT  99300.0 1631850.0 100500.0 1633050.0 ;
      RECT  94500.0 1623150.0 95700.0 1624350.0 ;
      RECT  96900.0 1623150.0 98100.0 1624350.0 ;
      RECT  96900.0 1623150.0 98100.0 1624350.0 ;
      RECT  94500.0 1623150.0 95700.0 1624350.0 ;
      RECT  96900.0 1623150.0 98100.0 1624350.0 ;
      RECT  99300.0 1623150.0 100500.0 1624350.0 ;
      RECT  99300.0 1623150.0 100500.0 1624350.0 ;
      RECT  96900.0 1623150.0 98100.0 1624350.0 ;
      RECT  99300.0 1623150.0 100500.0 1624350.0 ;
      RECT  101700.0 1623150.0 102900.0 1624350.0 ;
      RECT  101700.0 1623150.0 102900.0 1624350.0 ;
      RECT  99300.0 1623150.0 100500.0 1624350.0 ;
      RECT  104100.0 1632450.0 105300.0 1633650.0 ;
      RECT  104100.0 1622550.0 105300.0 1623750.0 ;
      RECT  101700.0 1625250.0 100500.0 1626450.0 ;
      RECT  99300.0 1627200.0 98100.0 1628400.0 ;
      RECT  96900.0 1629150.0 95700.0 1630350.0 ;
      RECT  96900.0 1631850.0 98100.0 1633050.0 ;
      RECT  101700.0 1631850.0 102900.0 1633050.0 ;
      RECT  101700.0 1623150.0 102900.0 1624350.0 ;
      RECT  101700.0 1629150.0 102900.0 1630350.0 ;
      RECT  95700.0 1629150.0 96900.0 1630350.0 ;
      RECT  98100.0 1627200.0 99300.0 1628400.0 ;
      RECT  100500.0 1625250.0 101700.0 1626450.0 ;
      RECT  101700.0 1629150.0 102900.0 1630350.0 ;
      RECT  92700.0 1634550.0 108300.0 1635450.0 ;
      RECT  92700.0 1620750.0 108300.0 1621650.0 ;
      RECT  94500.0 1646850.0 95700.0 1649250.0 ;
      RECT  94500.0 1638150.0 95700.0 1634550.0 ;
      RECT  99300.0 1638150.0 100500.0 1634550.0 ;
      RECT  104100.0 1636950.0 105300.0 1635000.0 ;
      RECT  104100.0 1648800.0 105300.0 1646850.0 ;
      RECT  94500.0 1638150.0 95700.0 1636950.0 ;
      RECT  96900.0 1638150.0 98100.0 1636950.0 ;
      RECT  96900.0 1638150.0 98100.0 1636950.0 ;
      RECT  94500.0 1638150.0 95700.0 1636950.0 ;
      RECT  96900.0 1638150.0 98100.0 1636950.0 ;
      RECT  99300.0 1638150.0 100500.0 1636950.0 ;
      RECT  99300.0 1638150.0 100500.0 1636950.0 ;
      RECT  96900.0 1638150.0 98100.0 1636950.0 ;
      RECT  99300.0 1638150.0 100500.0 1636950.0 ;
      RECT  101700.0 1638150.0 102900.0 1636950.0 ;
      RECT  101700.0 1638150.0 102900.0 1636950.0 ;
      RECT  99300.0 1638150.0 100500.0 1636950.0 ;
      RECT  94500.0 1646850.0 95700.0 1645650.0 ;
      RECT  96900.0 1646850.0 98100.0 1645650.0 ;
      RECT  96900.0 1646850.0 98100.0 1645650.0 ;
      RECT  94500.0 1646850.0 95700.0 1645650.0 ;
      RECT  96900.0 1646850.0 98100.0 1645650.0 ;
      RECT  99300.0 1646850.0 100500.0 1645650.0 ;
      RECT  99300.0 1646850.0 100500.0 1645650.0 ;
      RECT  96900.0 1646850.0 98100.0 1645650.0 ;
      RECT  99300.0 1646850.0 100500.0 1645650.0 ;
      RECT  101700.0 1646850.0 102900.0 1645650.0 ;
      RECT  101700.0 1646850.0 102900.0 1645650.0 ;
      RECT  99300.0 1646850.0 100500.0 1645650.0 ;
      RECT  104100.0 1637550.0 105300.0 1636350.0 ;
      RECT  104100.0 1647450.0 105300.0 1646250.0 ;
      RECT  101700.0 1644750.0 100500.0 1643550.0 ;
      RECT  99300.0 1642800.0 98100.0 1641600.0 ;
      RECT  96900.0 1640850.0 95700.0 1639650.0 ;
      RECT  96900.0 1638150.0 98100.0 1636950.0 ;
      RECT  101700.0 1638150.0 102900.0 1636950.0 ;
      RECT  101700.0 1646850.0 102900.0 1645650.0 ;
      RECT  101700.0 1640850.0 102900.0 1639650.0 ;
      RECT  95700.0 1640850.0 96900.0 1639650.0 ;
      RECT  98100.0 1642800.0 99300.0 1641600.0 ;
      RECT  100500.0 1644750.0 101700.0 1643550.0 ;
      RECT  101700.0 1640850.0 102900.0 1639650.0 ;
      RECT  92700.0 1635450.0 108300.0 1634550.0 ;
      RECT  92700.0 1649250.0 108300.0 1648350.0 ;
      RECT  94500.0 1650750.0 95700.0 1648350.0 ;
      RECT  94500.0 1659450.0 95700.0 1663050.0 ;
      RECT  99300.0 1659450.0 100500.0 1663050.0 ;
      RECT  104100.0 1660650.0 105300.0 1662600.0 ;
      RECT  104100.0 1648800.0 105300.0 1650750.0 ;
      RECT  94500.0 1659450.0 95700.0 1660650.0 ;
      RECT  96900.0 1659450.0 98100.0 1660650.0 ;
      RECT  96900.0 1659450.0 98100.0 1660650.0 ;
      RECT  94500.0 1659450.0 95700.0 1660650.0 ;
      RECT  96900.0 1659450.0 98100.0 1660650.0 ;
      RECT  99300.0 1659450.0 100500.0 1660650.0 ;
      RECT  99300.0 1659450.0 100500.0 1660650.0 ;
      RECT  96900.0 1659450.0 98100.0 1660650.0 ;
      RECT  99300.0 1659450.0 100500.0 1660650.0 ;
      RECT  101700.0 1659450.0 102900.0 1660650.0 ;
      RECT  101700.0 1659450.0 102900.0 1660650.0 ;
      RECT  99300.0 1659450.0 100500.0 1660650.0 ;
      RECT  94500.0 1650750.0 95700.0 1651950.0 ;
      RECT  96900.0 1650750.0 98100.0 1651950.0 ;
      RECT  96900.0 1650750.0 98100.0 1651950.0 ;
      RECT  94500.0 1650750.0 95700.0 1651950.0 ;
      RECT  96900.0 1650750.0 98100.0 1651950.0 ;
      RECT  99300.0 1650750.0 100500.0 1651950.0 ;
      RECT  99300.0 1650750.0 100500.0 1651950.0 ;
      RECT  96900.0 1650750.0 98100.0 1651950.0 ;
      RECT  99300.0 1650750.0 100500.0 1651950.0 ;
      RECT  101700.0 1650750.0 102900.0 1651950.0 ;
      RECT  101700.0 1650750.0 102900.0 1651950.0 ;
      RECT  99300.0 1650750.0 100500.0 1651950.0 ;
      RECT  104100.0 1660050.0 105300.0 1661250.0 ;
      RECT  104100.0 1650150.0 105300.0 1651350.0 ;
      RECT  101700.0 1652850.0 100500.0 1654050.0 ;
      RECT  99300.0 1654800.0 98100.0 1656000.0 ;
      RECT  96900.0 1656750.0 95700.0 1657950.0 ;
      RECT  96900.0 1659450.0 98100.0 1660650.0 ;
      RECT  101700.0 1659450.0 102900.0 1660650.0 ;
      RECT  101700.0 1650750.0 102900.0 1651950.0 ;
      RECT  101700.0 1656750.0 102900.0 1657950.0 ;
      RECT  95700.0 1656750.0 96900.0 1657950.0 ;
      RECT  98100.0 1654800.0 99300.0 1656000.0 ;
      RECT  100500.0 1652850.0 101700.0 1654050.0 ;
      RECT  101700.0 1656750.0 102900.0 1657950.0 ;
      RECT  92700.0 1662150.0 108300.0 1663050.0 ;
      RECT  92700.0 1648350.0 108300.0 1649250.0 ;
      RECT  94500.0 1674450.0 95700.0 1676850.0 ;
      RECT  94500.0 1665750.0 95700.0 1662150.0 ;
      RECT  99300.0 1665750.0 100500.0 1662150.0 ;
      RECT  104100.0 1664550.0 105300.0 1662600.0 ;
      RECT  104100.0 1676400.0 105300.0 1674450.0 ;
      RECT  94500.0 1665750.0 95700.0 1664550.0 ;
      RECT  96900.0 1665750.0 98100.0 1664550.0 ;
      RECT  96900.0 1665750.0 98100.0 1664550.0 ;
      RECT  94500.0 1665750.0 95700.0 1664550.0 ;
      RECT  96900.0 1665750.0 98100.0 1664550.0 ;
      RECT  99300.0 1665750.0 100500.0 1664550.0 ;
      RECT  99300.0 1665750.0 100500.0 1664550.0 ;
      RECT  96900.0 1665750.0 98100.0 1664550.0 ;
      RECT  99300.0 1665750.0 100500.0 1664550.0 ;
      RECT  101700.0 1665750.0 102900.0 1664550.0 ;
      RECT  101700.0 1665750.0 102900.0 1664550.0 ;
      RECT  99300.0 1665750.0 100500.0 1664550.0 ;
      RECT  94500.0 1674450.0 95700.0 1673250.0 ;
      RECT  96900.0 1674450.0 98100.0 1673250.0 ;
      RECT  96900.0 1674450.0 98100.0 1673250.0 ;
      RECT  94500.0 1674450.0 95700.0 1673250.0 ;
      RECT  96900.0 1674450.0 98100.0 1673250.0 ;
      RECT  99300.0 1674450.0 100500.0 1673250.0 ;
      RECT  99300.0 1674450.0 100500.0 1673250.0 ;
      RECT  96900.0 1674450.0 98100.0 1673250.0 ;
      RECT  99300.0 1674450.0 100500.0 1673250.0 ;
      RECT  101700.0 1674450.0 102900.0 1673250.0 ;
      RECT  101700.0 1674450.0 102900.0 1673250.0 ;
      RECT  99300.0 1674450.0 100500.0 1673250.0 ;
      RECT  104100.0 1665150.0 105300.0 1663950.0 ;
      RECT  104100.0 1675050.0 105300.0 1673850.0 ;
      RECT  101700.0 1672350.0 100500.0 1671150.0 ;
      RECT  99300.0 1670400.0 98100.0 1669200.0 ;
      RECT  96900.0 1668450.0 95700.0 1667250.0 ;
      RECT  96900.0 1665750.0 98100.0 1664550.0 ;
      RECT  101700.0 1665750.0 102900.0 1664550.0 ;
      RECT  101700.0 1674450.0 102900.0 1673250.0 ;
      RECT  101700.0 1668450.0 102900.0 1667250.0 ;
      RECT  95700.0 1668450.0 96900.0 1667250.0 ;
      RECT  98100.0 1670400.0 99300.0 1669200.0 ;
      RECT  100500.0 1672350.0 101700.0 1671150.0 ;
      RECT  101700.0 1668450.0 102900.0 1667250.0 ;
      RECT  92700.0 1663050.0 108300.0 1662150.0 ;
      RECT  92700.0 1676850.0 108300.0 1675950.0 ;
      RECT  94500.0 1678350.0 95700.0 1675950.0 ;
      RECT  94500.0 1687050.0 95700.0 1690650.0 ;
      RECT  99300.0 1687050.0 100500.0 1690650.0 ;
      RECT  104100.0 1688250.0 105300.0 1690200.0 ;
      RECT  104100.0 1676400.0 105300.0 1678350.0 ;
      RECT  94500.0 1687050.0 95700.0 1688250.0 ;
      RECT  96900.0 1687050.0 98100.0 1688250.0 ;
      RECT  96900.0 1687050.0 98100.0 1688250.0 ;
      RECT  94500.0 1687050.0 95700.0 1688250.0 ;
      RECT  96900.0 1687050.0 98100.0 1688250.0 ;
      RECT  99300.0 1687050.0 100500.0 1688250.0 ;
      RECT  99300.0 1687050.0 100500.0 1688250.0 ;
      RECT  96900.0 1687050.0 98100.0 1688250.0 ;
      RECT  99300.0 1687050.0 100500.0 1688250.0 ;
      RECT  101700.0 1687050.0 102900.0 1688250.0 ;
      RECT  101700.0 1687050.0 102900.0 1688250.0 ;
      RECT  99300.0 1687050.0 100500.0 1688250.0 ;
      RECT  94500.0 1678350.0 95700.0 1679550.0 ;
      RECT  96900.0 1678350.0 98100.0 1679550.0 ;
      RECT  96900.0 1678350.0 98100.0 1679550.0 ;
      RECT  94500.0 1678350.0 95700.0 1679550.0 ;
      RECT  96900.0 1678350.0 98100.0 1679550.0 ;
      RECT  99300.0 1678350.0 100500.0 1679550.0 ;
      RECT  99300.0 1678350.0 100500.0 1679550.0 ;
      RECT  96900.0 1678350.0 98100.0 1679550.0 ;
      RECT  99300.0 1678350.0 100500.0 1679550.0 ;
      RECT  101700.0 1678350.0 102900.0 1679550.0 ;
      RECT  101700.0 1678350.0 102900.0 1679550.0 ;
      RECT  99300.0 1678350.0 100500.0 1679550.0 ;
      RECT  104100.0 1687650.0 105300.0 1688850.0 ;
      RECT  104100.0 1677750.0 105300.0 1678950.0 ;
      RECT  101700.0 1680450.0 100500.0 1681650.0 ;
      RECT  99300.0 1682400.0 98100.0 1683600.0 ;
      RECT  96900.0 1684350.0 95700.0 1685550.0 ;
      RECT  96900.0 1687050.0 98100.0 1688250.0 ;
      RECT  101700.0 1687050.0 102900.0 1688250.0 ;
      RECT  101700.0 1678350.0 102900.0 1679550.0 ;
      RECT  101700.0 1684350.0 102900.0 1685550.0 ;
      RECT  95700.0 1684350.0 96900.0 1685550.0 ;
      RECT  98100.0 1682400.0 99300.0 1683600.0 ;
      RECT  100500.0 1680450.0 101700.0 1681650.0 ;
      RECT  101700.0 1684350.0 102900.0 1685550.0 ;
      RECT  92700.0 1689750.0 108300.0 1690650.0 ;
      RECT  92700.0 1675950.0 108300.0 1676850.0 ;
      RECT  94500.0 1702050.0 95700.0 1704450.0 ;
      RECT  94500.0 1693350.0 95700.0 1689750.0 ;
      RECT  99300.0 1693350.0 100500.0 1689750.0 ;
      RECT  104100.0 1692150.0 105300.0 1690200.0 ;
      RECT  104100.0 1704000.0 105300.0 1702050.0 ;
      RECT  94500.0 1693350.0 95700.0 1692150.0 ;
      RECT  96900.0 1693350.0 98100.0 1692150.0 ;
      RECT  96900.0 1693350.0 98100.0 1692150.0 ;
      RECT  94500.0 1693350.0 95700.0 1692150.0 ;
      RECT  96900.0 1693350.0 98100.0 1692150.0 ;
      RECT  99300.0 1693350.0 100500.0 1692150.0 ;
      RECT  99300.0 1693350.0 100500.0 1692150.0 ;
      RECT  96900.0 1693350.0 98100.0 1692150.0 ;
      RECT  99300.0 1693350.0 100500.0 1692150.0 ;
      RECT  101700.0 1693350.0 102900.0 1692150.0 ;
      RECT  101700.0 1693350.0 102900.0 1692150.0 ;
      RECT  99300.0 1693350.0 100500.0 1692150.0 ;
      RECT  94500.0 1702050.0 95700.0 1700850.0 ;
      RECT  96900.0 1702050.0 98100.0 1700850.0 ;
      RECT  96900.0 1702050.0 98100.0 1700850.0 ;
      RECT  94500.0 1702050.0 95700.0 1700850.0 ;
      RECT  96900.0 1702050.0 98100.0 1700850.0 ;
      RECT  99300.0 1702050.0 100500.0 1700850.0 ;
      RECT  99300.0 1702050.0 100500.0 1700850.0 ;
      RECT  96900.0 1702050.0 98100.0 1700850.0 ;
      RECT  99300.0 1702050.0 100500.0 1700850.0 ;
      RECT  101700.0 1702050.0 102900.0 1700850.0 ;
      RECT  101700.0 1702050.0 102900.0 1700850.0 ;
      RECT  99300.0 1702050.0 100500.0 1700850.0 ;
      RECT  104100.0 1692750.0 105300.0 1691550.0 ;
      RECT  104100.0 1702650.0 105300.0 1701450.0 ;
      RECT  101700.0 1699950.0 100500.0 1698750.0 ;
      RECT  99300.0 1698000.0 98100.0 1696800.0 ;
      RECT  96900.0 1696050.0 95700.0 1694850.0 ;
      RECT  96900.0 1693350.0 98100.0 1692150.0 ;
      RECT  101700.0 1693350.0 102900.0 1692150.0 ;
      RECT  101700.0 1702050.0 102900.0 1700850.0 ;
      RECT  101700.0 1696050.0 102900.0 1694850.0 ;
      RECT  95700.0 1696050.0 96900.0 1694850.0 ;
      RECT  98100.0 1698000.0 99300.0 1696800.0 ;
      RECT  100500.0 1699950.0 101700.0 1698750.0 ;
      RECT  101700.0 1696050.0 102900.0 1694850.0 ;
      RECT  92700.0 1690650.0 108300.0 1689750.0 ;
      RECT  92700.0 1704450.0 108300.0 1703550.0 ;
      RECT  94500.0 1705950.0 95700.0 1703550.0 ;
      RECT  94500.0 1714650.0 95700.0 1718250.0 ;
      RECT  99300.0 1714650.0 100500.0 1718250.0 ;
      RECT  104100.0 1715850.0 105300.0 1717800.0 ;
      RECT  104100.0 1704000.0 105300.0 1705950.0 ;
      RECT  94500.0 1714650.0 95700.0 1715850.0 ;
      RECT  96900.0 1714650.0 98100.0 1715850.0 ;
      RECT  96900.0 1714650.0 98100.0 1715850.0 ;
      RECT  94500.0 1714650.0 95700.0 1715850.0 ;
      RECT  96900.0 1714650.0 98100.0 1715850.0 ;
      RECT  99300.0 1714650.0 100500.0 1715850.0 ;
      RECT  99300.0 1714650.0 100500.0 1715850.0 ;
      RECT  96900.0 1714650.0 98100.0 1715850.0 ;
      RECT  99300.0 1714650.0 100500.0 1715850.0 ;
      RECT  101700.0 1714650.0 102900.0 1715850.0 ;
      RECT  101700.0 1714650.0 102900.0 1715850.0 ;
      RECT  99300.0 1714650.0 100500.0 1715850.0 ;
      RECT  94500.0 1705950.0 95700.0 1707150.0 ;
      RECT  96900.0 1705950.0 98100.0 1707150.0 ;
      RECT  96900.0 1705950.0 98100.0 1707150.0 ;
      RECT  94500.0 1705950.0 95700.0 1707150.0 ;
      RECT  96900.0 1705950.0 98100.0 1707150.0 ;
      RECT  99300.0 1705950.0 100500.0 1707150.0 ;
      RECT  99300.0 1705950.0 100500.0 1707150.0 ;
      RECT  96900.0 1705950.0 98100.0 1707150.0 ;
      RECT  99300.0 1705950.0 100500.0 1707150.0 ;
      RECT  101700.0 1705950.0 102900.0 1707150.0 ;
      RECT  101700.0 1705950.0 102900.0 1707150.0 ;
      RECT  99300.0 1705950.0 100500.0 1707150.0 ;
      RECT  104100.0 1715250.0 105300.0 1716450.0 ;
      RECT  104100.0 1705350.0 105300.0 1706550.0 ;
      RECT  101700.0 1708050.0 100500.0 1709250.0 ;
      RECT  99300.0 1710000.0 98100.0 1711200.0 ;
      RECT  96900.0 1711950.0 95700.0 1713150.0 ;
      RECT  96900.0 1714650.0 98100.0 1715850.0 ;
      RECT  101700.0 1714650.0 102900.0 1715850.0 ;
      RECT  101700.0 1705950.0 102900.0 1707150.0 ;
      RECT  101700.0 1711950.0 102900.0 1713150.0 ;
      RECT  95700.0 1711950.0 96900.0 1713150.0 ;
      RECT  98100.0 1710000.0 99300.0 1711200.0 ;
      RECT  100500.0 1708050.0 101700.0 1709250.0 ;
      RECT  101700.0 1711950.0 102900.0 1713150.0 ;
      RECT  92700.0 1717350.0 108300.0 1718250.0 ;
      RECT  92700.0 1703550.0 108300.0 1704450.0 ;
      RECT  94500.0 1729650.0 95700.0 1732050.0 ;
      RECT  94500.0 1720950.0 95700.0 1717350.0 ;
      RECT  99300.0 1720950.0 100500.0 1717350.0 ;
      RECT  104100.0 1719750.0 105300.0 1717800.0 ;
      RECT  104100.0 1731600.0 105300.0 1729650.0 ;
      RECT  94500.0 1720950.0 95700.0 1719750.0 ;
      RECT  96900.0 1720950.0 98100.0 1719750.0 ;
      RECT  96900.0 1720950.0 98100.0 1719750.0 ;
      RECT  94500.0 1720950.0 95700.0 1719750.0 ;
      RECT  96900.0 1720950.0 98100.0 1719750.0 ;
      RECT  99300.0 1720950.0 100500.0 1719750.0 ;
      RECT  99300.0 1720950.0 100500.0 1719750.0 ;
      RECT  96900.0 1720950.0 98100.0 1719750.0 ;
      RECT  99300.0 1720950.0 100500.0 1719750.0 ;
      RECT  101700.0 1720950.0 102900.0 1719750.0 ;
      RECT  101700.0 1720950.0 102900.0 1719750.0 ;
      RECT  99300.0 1720950.0 100500.0 1719750.0 ;
      RECT  94500.0 1729650.0 95700.0 1728450.0 ;
      RECT  96900.0 1729650.0 98100.0 1728450.0 ;
      RECT  96900.0 1729650.0 98100.0 1728450.0 ;
      RECT  94500.0 1729650.0 95700.0 1728450.0 ;
      RECT  96900.0 1729650.0 98100.0 1728450.0 ;
      RECT  99300.0 1729650.0 100500.0 1728450.0 ;
      RECT  99300.0 1729650.0 100500.0 1728450.0 ;
      RECT  96900.0 1729650.0 98100.0 1728450.0 ;
      RECT  99300.0 1729650.0 100500.0 1728450.0 ;
      RECT  101700.0 1729650.0 102900.0 1728450.0 ;
      RECT  101700.0 1729650.0 102900.0 1728450.0 ;
      RECT  99300.0 1729650.0 100500.0 1728450.0 ;
      RECT  104100.0 1720350.0 105300.0 1719150.0 ;
      RECT  104100.0 1730250.0 105300.0 1729050.0 ;
      RECT  101700.0 1727550.0 100500.0 1726350.0 ;
      RECT  99300.0 1725600.0 98100.0 1724400.0 ;
      RECT  96900.0 1723650.0 95700.0 1722450.0 ;
      RECT  96900.0 1720950.0 98100.0 1719750.0 ;
      RECT  101700.0 1720950.0 102900.0 1719750.0 ;
      RECT  101700.0 1729650.0 102900.0 1728450.0 ;
      RECT  101700.0 1723650.0 102900.0 1722450.0 ;
      RECT  95700.0 1723650.0 96900.0 1722450.0 ;
      RECT  98100.0 1725600.0 99300.0 1724400.0 ;
      RECT  100500.0 1727550.0 101700.0 1726350.0 ;
      RECT  101700.0 1723650.0 102900.0 1722450.0 ;
      RECT  92700.0 1718250.0 108300.0 1717350.0 ;
      RECT  92700.0 1732050.0 108300.0 1731150.0 ;
      RECT  94500.0 1733550.0 95700.0 1731150.0 ;
      RECT  94500.0 1742250.0 95700.0 1745850.0 ;
      RECT  99300.0 1742250.0 100500.0 1745850.0 ;
      RECT  104100.0 1743450.0 105300.0 1745400.0 ;
      RECT  104100.0 1731600.0 105300.0 1733550.0 ;
      RECT  94500.0 1742250.0 95700.0 1743450.0 ;
      RECT  96900.0 1742250.0 98100.0 1743450.0 ;
      RECT  96900.0 1742250.0 98100.0 1743450.0 ;
      RECT  94500.0 1742250.0 95700.0 1743450.0 ;
      RECT  96900.0 1742250.0 98100.0 1743450.0 ;
      RECT  99300.0 1742250.0 100500.0 1743450.0 ;
      RECT  99300.0 1742250.0 100500.0 1743450.0 ;
      RECT  96900.0 1742250.0 98100.0 1743450.0 ;
      RECT  99300.0 1742250.0 100500.0 1743450.0 ;
      RECT  101700.0 1742250.0 102900.0 1743450.0 ;
      RECT  101700.0 1742250.0 102900.0 1743450.0 ;
      RECT  99300.0 1742250.0 100500.0 1743450.0 ;
      RECT  94500.0 1733550.0 95700.0 1734750.0 ;
      RECT  96900.0 1733550.0 98100.0 1734750.0 ;
      RECT  96900.0 1733550.0 98100.0 1734750.0 ;
      RECT  94500.0 1733550.0 95700.0 1734750.0 ;
      RECT  96900.0 1733550.0 98100.0 1734750.0 ;
      RECT  99300.0 1733550.0 100500.0 1734750.0 ;
      RECT  99300.0 1733550.0 100500.0 1734750.0 ;
      RECT  96900.0 1733550.0 98100.0 1734750.0 ;
      RECT  99300.0 1733550.0 100500.0 1734750.0 ;
      RECT  101700.0 1733550.0 102900.0 1734750.0 ;
      RECT  101700.0 1733550.0 102900.0 1734750.0 ;
      RECT  99300.0 1733550.0 100500.0 1734750.0 ;
      RECT  104100.0 1742850.0 105300.0 1744050.0 ;
      RECT  104100.0 1732950.0 105300.0 1734150.0 ;
      RECT  101700.0 1735650.0 100500.0 1736850.0 ;
      RECT  99300.0 1737600.0 98100.0 1738800.0 ;
      RECT  96900.0 1739550.0 95700.0 1740750.0 ;
      RECT  96900.0 1742250.0 98100.0 1743450.0 ;
      RECT  101700.0 1742250.0 102900.0 1743450.0 ;
      RECT  101700.0 1733550.0 102900.0 1734750.0 ;
      RECT  101700.0 1739550.0 102900.0 1740750.0 ;
      RECT  95700.0 1739550.0 96900.0 1740750.0 ;
      RECT  98100.0 1737600.0 99300.0 1738800.0 ;
      RECT  100500.0 1735650.0 101700.0 1736850.0 ;
      RECT  101700.0 1739550.0 102900.0 1740750.0 ;
      RECT  92700.0 1744950.0 108300.0 1745850.0 ;
      RECT  92700.0 1731150.0 108300.0 1732050.0 ;
      RECT  94500.0 1757250.0 95700.0 1759650.0 ;
      RECT  94500.0 1748550.0 95700.0 1744950.0 ;
      RECT  99300.0 1748550.0 100500.0 1744950.0 ;
      RECT  104100.0 1747350.0 105300.0 1745400.0 ;
      RECT  104100.0 1759200.0 105300.0 1757250.0 ;
      RECT  94500.0 1748550.0 95700.0 1747350.0 ;
      RECT  96900.0 1748550.0 98100.0 1747350.0 ;
      RECT  96900.0 1748550.0 98100.0 1747350.0 ;
      RECT  94500.0 1748550.0 95700.0 1747350.0 ;
      RECT  96900.0 1748550.0 98100.0 1747350.0 ;
      RECT  99300.0 1748550.0 100500.0 1747350.0 ;
      RECT  99300.0 1748550.0 100500.0 1747350.0 ;
      RECT  96900.0 1748550.0 98100.0 1747350.0 ;
      RECT  99300.0 1748550.0 100500.0 1747350.0 ;
      RECT  101700.0 1748550.0 102900.0 1747350.0 ;
      RECT  101700.0 1748550.0 102900.0 1747350.0 ;
      RECT  99300.0 1748550.0 100500.0 1747350.0 ;
      RECT  94500.0 1757250.0 95700.0 1756050.0 ;
      RECT  96900.0 1757250.0 98100.0 1756050.0 ;
      RECT  96900.0 1757250.0 98100.0 1756050.0 ;
      RECT  94500.0 1757250.0 95700.0 1756050.0 ;
      RECT  96900.0 1757250.0 98100.0 1756050.0 ;
      RECT  99300.0 1757250.0 100500.0 1756050.0 ;
      RECT  99300.0 1757250.0 100500.0 1756050.0 ;
      RECT  96900.0 1757250.0 98100.0 1756050.0 ;
      RECT  99300.0 1757250.0 100500.0 1756050.0 ;
      RECT  101700.0 1757250.0 102900.0 1756050.0 ;
      RECT  101700.0 1757250.0 102900.0 1756050.0 ;
      RECT  99300.0 1757250.0 100500.0 1756050.0 ;
      RECT  104100.0 1747950.0 105300.0 1746750.0 ;
      RECT  104100.0 1757850.0 105300.0 1756650.0 ;
      RECT  101700.0 1755150.0 100500.0 1753950.0 ;
      RECT  99300.0 1753200.0 98100.0 1752000.0 ;
      RECT  96900.0 1751250.0 95700.0 1750050.0 ;
      RECT  96900.0 1748550.0 98100.0 1747350.0 ;
      RECT  101700.0 1748550.0 102900.0 1747350.0 ;
      RECT  101700.0 1757250.0 102900.0 1756050.0 ;
      RECT  101700.0 1751250.0 102900.0 1750050.0 ;
      RECT  95700.0 1751250.0 96900.0 1750050.0 ;
      RECT  98100.0 1753200.0 99300.0 1752000.0 ;
      RECT  100500.0 1755150.0 101700.0 1753950.0 ;
      RECT  101700.0 1751250.0 102900.0 1750050.0 ;
      RECT  92700.0 1745850.0 108300.0 1744950.0 ;
      RECT  92700.0 1759650.0 108300.0 1758750.0 ;
      RECT  94500.0 1761150.0 95700.0 1758750.0 ;
      RECT  94500.0 1769850.0 95700.0 1773450.0 ;
      RECT  99300.0 1769850.0 100500.0 1773450.0 ;
      RECT  104100.0 1771050.0 105300.0 1773000.0 ;
      RECT  104100.0 1759200.0 105300.0 1761150.0 ;
      RECT  94500.0 1769850.0 95700.0 1771050.0 ;
      RECT  96900.0 1769850.0 98100.0 1771050.0 ;
      RECT  96900.0 1769850.0 98100.0 1771050.0 ;
      RECT  94500.0 1769850.0 95700.0 1771050.0 ;
      RECT  96900.0 1769850.0 98100.0 1771050.0 ;
      RECT  99300.0 1769850.0 100500.0 1771050.0 ;
      RECT  99300.0 1769850.0 100500.0 1771050.0 ;
      RECT  96900.0 1769850.0 98100.0 1771050.0 ;
      RECT  99300.0 1769850.0 100500.0 1771050.0 ;
      RECT  101700.0 1769850.0 102900.0 1771050.0 ;
      RECT  101700.0 1769850.0 102900.0 1771050.0 ;
      RECT  99300.0 1769850.0 100500.0 1771050.0 ;
      RECT  94500.0 1761150.0 95700.0 1762350.0 ;
      RECT  96900.0 1761150.0 98100.0 1762350.0 ;
      RECT  96900.0 1761150.0 98100.0 1762350.0 ;
      RECT  94500.0 1761150.0 95700.0 1762350.0 ;
      RECT  96900.0 1761150.0 98100.0 1762350.0 ;
      RECT  99300.0 1761150.0 100500.0 1762350.0 ;
      RECT  99300.0 1761150.0 100500.0 1762350.0 ;
      RECT  96900.0 1761150.0 98100.0 1762350.0 ;
      RECT  99300.0 1761150.0 100500.0 1762350.0 ;
      RECT  101700.0 1761150.0 102900.0 1762350.0 ;
      RECT  101700.0 1761150.0 102900.0 1762350.0 ;
      RECT  99300.0 1761150.0 100500.0 1762350.0 ;
      RECT  104100.0 1770450.0 105300.0 1771650.0 ;
      RECT  104100.0 1760550.0 105300.0 1761750.0 ;
      RECT  101700.0 1763250.0 100500.0 1764450.0 ;
      RECT  99300.0 1765200.0 98100.0 1766400.0 ;
      RECT  96900.0 1767150.0 95700.0 1768350.0 ;
      RECT  96900.0 1769850.0 98100.0 1771050.0 ;
      RECT  101700.0 1769850.0 102900.0 1771050.0 ;
      RECT  101700.0 1761150.0 102900.0 1762350.0 ;
      RECT  101700.0 1767150.0 102900.0 1768350.0 ;
      RECT  95700.0 1767150.0 96900.0 1768350.0 ;
      RECT  98100.0 1765200.0 99300.0 1766400.0 ;
      RECT  100500.0 1763250.0 101700.0 1764450.0 ;
      RECT  101700.0 1767150.0 102900.0 1768350.0 ;
      RECT  92700.0 1772550.0 108300.0 1773450.0 ;
      RECT  92700.0 1758750.0 108300.0 1759650.0 ;
      RECT  94500.0 1784850.0 95700.0 1787250.0 ;
      RECT  94500.0 1776150.0 95700.0 1772550.0 ;
      RECT  99300.0 1776150.0 100500.0 1772550.0 ;
      RECT  104100.0 1774950.0 105300.0 1773000.0 ;
      RECT  104100.0 1786800.0 105300.0 1784850.0 ;
      RECT  94500.0 1776150.0 95700.0 1774950.0 ;
      RECT  96900.0 1776150.0 98100.0 1774950.0 ;
      RECT  96900.0 1776150.0 98100.0 1774950.0 ;
      RECT  94500.0 1776150.0 95700.0 1774950.0 ;
      RECT  96900.0 1776150.0 98100.0 1774950.0 ;
      RECT  99300.0 1776150.0 100500.0 1774950.0 ;
      RECT  99300.0 1776150.0 100500.0 1774950.0 ;
      RECT  96900.0 1776150.0 98100.0 1774950.0 ;
      RECT  99300.0 1776150.0 100500.0 1774950.0 ;
      RECT  101700.0 1776150.0 102900.0 1774950.0 ;
      RECT  101700.0 1776150.0 102900.0 1774950.0 ;
      RECT  99300.0 1776150.0 100500.0 1774950.0 ;
      RECT  94500.0 1784850.0 95700.0 1783650.0 ;
      RECT  96900.0 1784850.0 98100.0 1783650.0 ;
      RECT  96900.0 1784850.0 98100.0 1783650.0 ;
      RECT  94500.0 1784850.0 95700.0 1783650.0 ;
      RECT  96900.0 1784850.0 98100.0 1783650.0 ;
      RECT  99300.0 1784850.0 100500.0 1783650.0 ;
      RECT  99300.0 1784850.0 100500.0 1783650.0 ;
      RECT  96900.0 1784850.0 98100.0 1783650.0 ;
      RECT  99300.0 1784850.0 100500.0 1783650.0 ;
      RECT  101700.0 1784850.0 102900.0 1783650.0 ;
      RECT  101700.0 1784850.0 102900.0 1783650.0 ;
      RECT  99300.0 1784850.0 100500.0 1783650.0 ;
      RECT  104100.0 1775550.0 105300.0 1774350.0 ;
      RECT  104100.0 1785450.0 105300.0 1784250.0 ;
      RECT  101700.0 1782750.0 100500.0 1781550.0 ;
      RECT  99300.0 1780800.0 98100.0 1779600.0 ;
      RECT  96900.0 1778850.0 95700.0 1777650.0 ;
      RECT  96900.0 1776150.0 98100.0 1774950.0 ;
      RECT  101700.0 1776150.0 102900.0 1774950.0 ;
      RECT  101700.0 1784850.0 102900.0 1783650.0 ;
      RECT  101700.0 1778850.0 102900.0 1777650.0 ;
      RECT  95700.0 1778850.0 96900.0 1777650.0 ;
      RECT  98100.0 1780800.0 99300.0 1779600.0 ;
      RECT  100500.0 1782750.0 101700.0 1781550.0 ;
      RECT  101700.0 1778850.0 102900.0 1777650.0 ;
      RECT  92700.0 1773450.0 108300.0 1772550.0 ;
      RECT  92700.0 1787250.0 108300.0 1786350.0 ;
      RECT  94500.0 1788750.0 95700.0 1786350.0 ;
      RECT  94500.0 1797450.0 95700.0 1801050.0 ;
      RECT  99300.0 1797450.0 100500.0 1801050.0 ;
      RECT  104100.0 1798650.0 105300.0 1800600.0 ;
      RECT  104100.0 1786800.0 105300.0 1788750.0 ;
      RECT  94500.0 1797450.0 95700.0 1798650.0 ;
      RECT  96900.0 1797450.0 98100.0 1798650.0 ;
      RECT  96900.0 1797450.0 98100.0 1798650.0 ;
      RECT  94500.0 1797450.0 95700.0 1798650.0 ;
      RECT  96900.0 1797450.0 98100.0 1798650.0 ;
      RECT  99300.0 1797450.0 100500.0 1798650.0 ;
      RECT  99300.0 1797450.0 100500.0 1798650.0 ;
      RECT  96900.0 1797450.0 98100.0 1798650.0 ;
      RECT  99300.0 1797450.0 100500.0 1798650.0 ;
      RECT  101700.0 1797450.0 102900.0 1798650.0 ;
      RECT  101700.0 1797450.0 102900.0 1798650.0 ;
      RECT  99300.0 1797450.0 100500.0 1798650.0 ;
      RECT  94500.0 1788750.0 95700.0 1789950.0 ;
      RECT  96900.0 1788750.0 98100.0 1789950.0 ;
      RECT  96900.0 1788750.0 98100.0 1789950.0 ;
      RECT  94500.0 1788750.0 95700.0 1789950.0 ;
      RECT  96900.0 1788750.0 98100.0 1789950.0 ;
      RECT  99300.0 1788750.0 100500.0 1789950.0 ;
      RECT  99300.0 1788750.0 100500.0 1789950.0 ;
      RECT  96900.0 1788750.0 98100.0 1789950.0 ;
      RECT  99300.0 1788750.0 100500.0 1789950.0 ;
      RECT  101700.0 1788750.0 102900.0 1789950.0 ;
      RECT  101700.0 1788750.0 102900.0 1789950.0 ;
      RECT  99300.0 1788750.0 100500.0 1789950.0 ;
      RECT  104100.0 1798050.0 105300.0 1799250.0 ;
      RECT  104100.0 1788150.0 105300.0 1789350.0 ;
      RECT  101700.0 1790850.0 100500.0 1792050.0 ;
      RECT  99300.0 1792800.0 98100.0 1794000.0 ;
      RECT  96900.0 1794750.0 95700.0 1795950.0 ;
      RECT  96900.0 1797450.0 98100.0 1798650.0 ;
      RECT  101700.0 1797450.0 102900.0 1798650.0 ;
      RECT  101700.0 1788750.0 102900.0 1789950.0 ;
      RECT  101700.0 1794750.0 102900.0 1795950.0 ;
      RECT  95700.0 1794750.0 96900.0 1795950.0 ;
      RECT  98100.0 1792800.0 99300.0 1794000.0 ;
      RECT  100500.0 1790850.0 101700.0 1792050.0 ;
      RECT  101700.0 1794750.0 102900.0 1795950.0 ;
      RECT  92700.0 1800150.0 108300.0 1801050.0 ;
      RECT  92700.0 1786350.0 108300.0 1787250.0 ;
      RECT  94500.0 1812450.0 95700.0 1814850.0 ;
      RECT  94500.0 1803750.0 95700.0 1800150.0 ;
      RECT  99300.0 1803750.0 100500.0 1800150.0 ;
      RECT  104100.0 1802550.0 105300.0 1800600.0 ;
      RECT  104100.0 1814400.0 105300.0 1812450.0 ;
      RECT  94500.0 1803750.0 95700.0 1802550.0 ;
      RECT  96900.0 1803750.0 98100.0 1802550.0 ;
      RECT  96900.0 1803750.0 98100.0 1802550.0 ;
      RECT  94500.0 1803750.0 95700.0 1802550.0 ;
      RECT  96900.0 1803750.0 98100.0 1802550.0 ;
      RECT  99300.0 1803750.0 100500.0 1802550.0 ;
      RECT  99300.0 1803750.0 100500.0 1802550.0 ;
      RECT  96900.0 1803750.0 98100.0 1802550.0 ;
      RECT  99300.0 1803750.0 100500.0 1802550.0 ;
      RECT  101700.0 1803750.0 102900.0 1802550.0 ;
      RECT  101700.0 1803750.0 102900.0 1802550.0 ;
      RECT  99300.0 1803750.0 100500.0 1802550.0 ;
      RECT  94500.0 1812450.0 95700.0 1811250.0 ;
      RECT  96900.0 1812450.0 98100.0 1811250.0 ;
      RECT  96900.0 1812450.0 98100.0 1811250.0 ;
      RECT  94500.0 1812450.0 95700.0 1811250.0 ;
      RECT  96900.0 1812450.0 98100.0 1811250.0 ;
      RECT  99300.0 1812450.0 100500.0 1811250.0 ;
      RECT  99300.0 1812450.0 100500.0 1811250.0 ;
      RECT  96900.0 1812450.0 98100.0 1811250.0 ;
      RECT  99300.0 1812450.0 100500.0 1811250.0 ;
      RECT  101700.0 1812450.0 102900.0 1811250.0 ;
      RECT  101700.0 1812450.0 102900.0 1811250.0 ;
      RECT  99300.0 1812450.0 100500.0 1811250.0 ;
      RECT  104100.0 1803150.0 105300.0 1801950.0 ;
      RECT  104100.0 1813050.0 105300.0 1811850.0 ;
      RECT  101700.0 1810350.0 100500.0 1809150.0 ;
      RECT  99300.0 1808400.0 98100.0 1807200.0 ;
      RECT  96900.0 1806450.0 95700.0 1805250.0 ;
      RECT  96900.0 1803750.0 98100.0 1802550.0 ;
      RECT  101700.0 1803750.0 102900.0 1802550.0 ;
      RECT  101700.0 1812450.0 102900.0 1811250.0 ;
      RECT  101700.0 1806450.0 102900.0 1805250.0 ;
      RECT  95700.0 1806450.0 96900.0 1805250.0 ;
      RECT  98100.0 1808400.0 99300.0 1807200.0 ;
      RECT  100500.0 1810350.0 101700.0 1809150.0 ;
      RECT  101700.0 1806450.0 102900.0 1805250.0 ;
      RECT  92700.0 1801050.0 108300.0 1800150.0 ;
      RECT  92700.0 1814850.0 108300.0 1813950.0 ;
      RECT  94500.0 1816350.0 95700.0 1813950.0 ;
      RECT  94500.0 1825050.0 95700.0 1828650.0 ;
      RECT  99300.0 1825050.0 100500.0 1828650.0 ;
      RECT  104100.0 1826250.0 105300.0 1828200.0 ;
      RECT  104100.0 1814400.0 105300.0 1816350.0 ;
      RECT  94500.0 1825050.0 95700.0 1826250.0 ;
      RECT  96900.0 1825050.0 98100.0 1826250.0 ;
      RECT  96900.0 1825050.0 98100.0 1826250.0 ;
      RECT  94500.0 1825050.0 95700.0 1826250.0 ;
      RECT  96900.0 1825050.0 98100.0 1826250.0 ;
      RECT  99300.0 1825050.0 100500.0 1826250.0 ;
      RECT  99300.0 1825050.0 100500.0 1826250.0 ;
      RECT  96900.0 1825050.0 98100.0 1826250.0 ;
      RECT  99300.0 1825050.0 100500.0 1826250.0 ;
      RECT  101700.0 1825050.0 102900.0 1826250.0 ;
      RECT  101700.0 1825050.0 102900.0 1826250.0 ;
      RECT  99300.0 1825050.0 100500.0 1826250.0 ;
      RECT  94500.0 1816350.0 95700.0 1817550.0 ;
      RECT  96900.0 1816350.0 98100.0 1817550.0 ;
      RECT  96900.0 1816350.0 98100.0 1817550.0 ;
      RECT  94500.0 1816350.0 95700.0 1817550.0 ;
      RECT  96900.0 1816350.0 98100.0 1817550.0 ;
      RECT  99300.0 1816350.0 100500.0 1817550.0 ;
      RECT  99300.0 1816350.0 100500.0 1817550.0 ;
      RECT  96900.0 1816350.0 98100.0 1817550.0 ;
      RECT  99300.0 1816350.0 100500.0 1817550.0 ;
      RECT  101700.0 1816350.0 102900.0 1817550.0 ;
      RECT  101700.0 1816350.0 102900.0 1817550.0 ;
      RECT  99300.0 1816350.0 100500.0 1817550.0 ;
      RECT  104100.0 1825650.0 105300.0 1826850.0 ;
      RECT  104100.0 1815750.0 105300.0 1816950.0 ;
      RECT  101700.0 1818450.0 100500.0 1819650.0 ;
      RECT  99300.0 1820400.0 98100.0 1821600.0 ;
      RECT  96900.0 1822350.0 95700.0 1823550.0 ;
      RECT  96900.0 1825050.0 98100.0 1826250.0 ;
      RECT  101700.0 1825050.0 102900.0 1826250.0 ;
      RECT  101700.0 1816350.0 102900.0 1817550.0 ;
      RECT  101700.0 1822350.0 102900.0 1823550.0 ;
      RECT  95700.0 1822350.0 96900.0 1823550.0 ;
      RECT  98100.0 1820400.0 99300.0 1821600.0 ;
      RECT  100500.0 1818450.0 101700.0 1819650.0 ;
      RECT  101700.0 1822350.0 102900.0 1823550.0 ;
      RECT  92700.0 1827750.0 108300.0 1828650.0 ;
      RECT  92700.0 1813950.0 108300.0 1814850.0 ;
      RECT  94500.0 1840050.0 95700.0 1842450.0 ;
      RECT  94500.0 1831350.0 95700.0 1827750.0 ;
      RECT  99300.0 1831350.0 100500.0 1827750.0 ;
      RECT  104100.0 1830150.0 105300.0 1828200.0 ;
      RECT  104100.0 1842000.0 105300.0 1840050.0 ;
      RECT  94500.0 1831350.0 95700.0 1830150.0 ;
      RECT  96900.0 1831350.0 98100.0 1830150.0 ;
      RECT  96900.0 1831350.0 98100.0 1830150.0 ;
      RECT  94500.0 1831350.0 95700.0 1830150.0 ;
      RECT  96900.0 1831350.0 98100.0 1830150.0 ;
      RECT  99300.0 1831350.0 100500.0 1830150.0 ;
      RECT  99300.0 1831350.0 100500.0 1830150.0 ;
      RECT  96900.0 1831350.0 98100.0 1830150.0 ;
      RECT  99300.0 1831350.0 100500.0 1830150.0 ;
      RECT  101700.0 1831350.0 102900.0 1830150.0 ;
      RECT  101700.0 1831350.0 102900.0 1830150.0 ;
      RECT  99300.0 1831350.0 100500.0 1830150.0 ;
      RECT  94500.0 1840050.0 95700.0 1838850.0 ;
      RECT  96900.0 1840050.0 98100.0 1838850.0 ;
      RECT  96900.0 1840050.0 98100.0 1838850.0 ;
      RECT  94500.0 1840050.0 95700.0 1838850.0 ;
      RECT  96900.0 1840050.0 98100.0 1838850.0 ;
      RECT  99300.0 1840050.0 100500.0 1838850.0 ;
      RECT  99300.0 1840050.0 100500.0 1838850.0 ;
      RECT  96900.0 1840050.0 98100.0 1838850.0 ;
      RECT  99300.0 1840050.0 100500.0 1838850.0 ;
      RECT  101700.0 1840050.0 102900.0 1838850.0 ;
      RECT  101700.0 1840050.0 102900.0 1838850.0 ;
      RECT  99300.0 1840050.0 100500.0 1838850.0 ;
      RECT  104100.0 1830750.0 105300.0 1829550.0 ;
      RECT  104100.0 1840650.0 105300.0 1839450.0 ;
      RECT  101700.0 1837950.0 100500.0 1836750.0 ;
      RECT  99300.0 1836000.0 98100.0 1834800.0 ;
      RECT  96900.0 1834050.0 95700.0 1832850.0 ;
      RECT  96900.0 1831350.0 98100.0 1830150.0 ;
      RECT  101700.0 1831350.0 102900.0 1830150.0 ;
      RECT  101700.0 1840050.0 102900.0 1838850.0 ;
      RECT  101700.0 1834050.0 102900.0 1832850.0 ;
      RECT  95700.0 1834050.0 96900.0 1832850.0 ;
      RECT  98100.0 1836000.0 99300.0 1834800.0 ;
      RECT  100500.0 1837950.0 101700.0 1836750.0 ;
      RECT  101700.0 1834050.0 102900.0 1832850.0 ;
      RECT  92700.0 1828650.0 108300.0 1827750.0 ;
      RECT  92700.0 1842450.0 108300.0 1841550.0 ;
      RECT  94500.0 1843950.0 95700.0 1841550.0 ;
      RECT  94500.0 1852650.0 95700.0 1856250.0 ;
      RECT  99300.0 1852650.0 100500.0 1856250.0 ;
      RECT  104100.0 1853850.0 105300.0 1855800.0 ;
      RECT  104100.0 1842000.0 105300.0 1843950.0 ;
      RECT  94500.0 1852650.0 95700.0 1853850.0 ;
      RECT  96900.0 1852650.0 98100.0 1853850.0 ;
      RECT  96900.0 1852650.0 98100.0 1853850.0 ;
      RECT  94500.0 1852650.0 95700.0 1853850.0 ;
      RECT  96900.0 1852650.0 98100.0 1853850.0 ;
      RECT  99300.0 1852650.0 100500.0 1853850.0 ;
      RECT  99300.0 1852650.0 100500.0 1853850.0 ;
      RECT  96900.0 1852650.0 98100.0 1853850.0 ;
      RECT  99300.0 1852650.0 100500.0 1853850.0 ;
      RECT  101700.0 1852650.0 102900.0 1853850.0 ;
      RECT  101700.0 1852650.0 102900.0 1853850.0 ;
      RECT  99300.0 1852650.0 100500.0 1853850.0 ;
      RECT  94500.0 1843950.0 95700.0 1845150.0 ;
      RECT  96900.0 1843950.0 98100.0 1845150.0 ;
      RECT  96900.0 1843950.0 98100.0 1845150.0 ;
      RECT  94500.0 1843950.0 95700.0 1845150.0 ;
      RECT  96900.0 1843950.0 98100.0 1845150.0 ;
      RECT  99300.0 1843950.0 100500.0 1845150.0 ;
      RECT  99300.0 1843950.0 100500.0 1845150.0 ;
      RECT  96900.0 1843950.0 98100.0 1845150.0 ;
      RECT  99300.0 1843950.0 100500.0 1845150.0 ;
      RECT  101700.0 1843950.0 102900.0 1845150.0 ;
      RECT  101700.0 1843950.0 102900.0 1845150.0 ;
      RECT  99300.0 1843950.0 100500.0 1845150.0 ;
      RECT  104100.0 1853250.0 105300.0 1854450.0 ;
      RECT  104100.0 1843350.0 105300.0 1844550.0 ;
      RECT  101700.0 1846050.0 100500.0 1847250.0 ;
      RECT  99300.0 1848000.0 98100.0 1849200.0 ;
      RECT  96900.0 1849950.0 95700.0 1851150.0 ;
      RECT  96900.0 1852650.0 98100.0 1853850.0 ;
      RECT  101700.0 1852650.0 102900.0 1853850.0 ;
      RECT  101700.0 1843950.0 102900.0 1845150.0 ;
      RECT  101700.0 1849950.0 102900.0 1851150.0 ;
      RECT  95700.0 1849950.0 96900.0 1851150.0 ;
      RECT  98100.0 1848000.0 99300.0 1849200.0 ;
      RECT  100500.0 1846050.0 101700.0 1847250.0 ;
      RECT  101700.0 1849950.0 102900.0 1851150.0 ;
      RECT  92700.0 1855350.0 108300.0 1856250.0 ;
      RECT  92700.0 1841550.0 108300.0 1842450.0 ;
      RECT  94500.0 1867650.0 95700.0 1870050.0 ;
      RECT  94500.0 1858950.0 95700.0 1855350.0 ;
      RECT  99300.0 1858950.0 100500.0 1855350.0 ;
      RECT  104100.0 1857750.0 105300.0 1855800.0 ;
      RECT  104100.0 1869600.0 105300.0 1867650.0 ;
      RECT  94500.0 1858950.0 95700.0 1857750.0 ;
      RECT  96900.0 1858950.0 98100.0 1857750.0 ;
      RECT  96900.0 1858950.0 98100.0 1857750.0 ;
      RECT  94500.0 1858950.0 95700.0 1857750.0 ;
      RECT  96900.0 1858950.0 98100.0 1857750.0 ;
      RECT  99300.0 1858950.0 100500.0 1857750.0 ;
      RECT  99300.0 1858950.0 100500.0 1857750.0 ;
      RECT  96900.0 1858950.0 98100.0 1857750.0 ;
      RECT  99300.0 1858950.0 100500.0 1857750.0 ;
      RECT  101700.0 1858950.0 102900.0 1857750.0 ;
      RECT  101700.0 1858950.0 102900.0 1857750.0 ;
      RECT  99300.0 1858950.0 100500.0 1857750.0 ;
      RECT  94500.0 1867650.0 95700.0 1866450.0 ;
      RECT  96900.0 1867650.0 98100.0 1866450.0 ;
      RECT  96900.0 1867650.0 98100.0 1866450.0 ;
      RECT  94500.0 1867650.0 95700.0 1866450.0 ;
      RECT  96900.0 1867650.0 98100.0 1866450.0 ;
      RECT  99300.0 1867650.0 100500.0 1866450.0 ;
      RECT  99300.0 1867650.0 100500.0 1866450.0 ;
      RECT  96900.0 1867650.0 98100.0 1866450.0 ;
      RECT  99300.0 1867650.0 100500.0 1866450.0 ;
      RECT  101700.0 1867650.0 102900.0 1866450.0 ;
      RECT  101700.0 1867650.0 102900.0 1866450.0 ;
      RECT  99300.0 1867650.0 100500.0 1866450.0 ;
      RECT  104100.0 1858350.0 105300.0 1857150.0 ;
      RECT  104100.0 1868250.0 105300.0 1867050.0 ;
      RECT  101700.0 1865550.0 100500.0 1864350.0 ;
      RECT  99300.0 1863600.0 98100.0 1862400.0 ;
      RECT  96900.0 1861650.0 95700.0 1860450.0 ;
      RECT  96900.0 1858950.0 98100.0 1857750.0 ;
      RECT  101700.0 1858950.0 102900.0 1857750.0 ;
      RECT  101700.0 1867650.0 102900.0 1866450.0 ;
      RECT  101700.0 1861650.0 102900.0 1860450.0 ;
      RECT  95700.0 1861650.0 96900.0 1860450.0 ;
      RECT  98100.0 1863600.0 99300.0 1862400.0 ;
      RECT  100500.0 1865550.0 101700.0 1864350.0 ;
      RECT  101700.0 1861650.0 102900.0 1860450.0 ;
      RECT  92700.0 1856250.0 108300.0 1855350.0 ;
      RECT  92700.0 1870050.0 108300.0 1869150.0 ;
      RECT  94500.0 1871550.0 95700.0 1869150.0 ;
      RECT  94500.0 1880250.0 95700.0 1883850.0 ;
      RECT  99300.0 1880250.0 100500.0 1883850.0 ;
      RECT  104100.0 1881450.0 105300.0 1883400.0 ;
      RECT  104100.0 1869600.0 105300.0 1871550.0 ;
      RECT  94500.0 1880250.0 95700.0 1881450.0 ;
      RECT  96900.0 1880250.0 98100.0 1881450.0 ;
      RECT  96900.0 1880250.0 98100.0 1881450.0 ;
      RECT  94500.0 1880250.0 95700.0 1881450.0 ;
      RECT  96900.0 1880250.0 98100.0 1881450.0 ;
      RECT  99300.0 1880250.0 100500.0 1881450.0 ;
      RECT  99300.0 1880250.0 100500.0 1881450.0 ;
      RECT  96900.0 1880250.0 98100.0 1881450.0 ;
      RECT  99300.0 1880250.0 100500.0 1881450.0 ;
      RECT  101700.0 1880250.0 102900.0 1881450.0 ;
      RECT  101700.0 1880250.0 102900.0 1881450.0 ;
      RECT  99300.0 1880250.0 100500.0 1881450.0 ;
      RECT  94500.0 1871550.0 95700.0 1872750.0 ;
      RECT  96900.0 1871550.0 98100.0 1872750.0 ;
      RECT  96900.0 1871550.0 98100.0 1872750.0 ;
      RECT  94500.0 1871550.0 95700.0 1872750.0 ;
      RECT  96900.0 1871550.0 98100.0 1872750.0 ;
      RECT  99300.0 1871550.0 100500.0 1872750.0 ;
      RECT  99300.0 1871550.0 100500.0 1872750.0 ;
      RECT  96900.0 1871550.0 98100.0 1872750.0 ;
      RECT  99300.0 1871550.0 100500.0 1872750.0 ;
      RECT  101700.0 1871550.0 102900.0 1872750.0 ;
      RECT  101700.0 1871550.0 102900.0 1872750.0 ;
      RECT  99300.0 1871550.0 100500.0 1872750.0 ;
      RECT  104100.0 1880850.0 105300.0 1882050.0 ;
      RECT  104100.0 1870950.0 105300.0 1872150.0 ;
      RECT  101700.0 1873650.0 100500.0 1874850.0 ;
      RECT  99300.0 1875600.0 98100.0 1876800.0 ;
      RECT  96900.0 1877550.0 95700.0 1878750.0 ;
      RECT  96900.0 1880250.0 98100.0 1881450.0 ;
      RECT  101700.0 1880250.0 102900.0 1881450.0 ;
      RECT  101700.0 1871550.0 102900.0 1872750.0 ;
      RECT  101700.0 1877550.0 102900.0 1878750.0 ;
      RECT  95700.0 1877550.0 96900.0 1878750.0 ;
      RECT  98100.0 1875600.0 99300.0 1876800.0 ;
      RECT  100500.0 1873650.0 101700.0 1874850.0 ;
      RECT  101700.0 1877550.0 102900.0 1878750.0 ;
      RECT  92700.0 1882950.0 108300.0 1883850.0 ;
      RECT  92700.0 1869150.0 108300.0 1870050.0 ;
      RECT  94500.0 1895250.0 95700.0 1897650.0 ;
      RECT  94500.0 1886550.0 95700.0 1882950.0 ;
      RECT  99300.0 1886550.0 100500.0 1882950.0 ;
      RECT  104100.0 1885350.0 105300.0 1883400.0 ;
      RECT  104100.0 1897200.0 105300.0 1895250.0 ;
      RECT  94500.0 1886550.0 95700.0 1885350.0 ;
      RECT  96900.0 1886550.0 98100.0 1885350.0 ;
      RECT  96900.0 1886550.0 98100.0 1885350.0 ;
      RECT  94500.0 1886550.0 95700.0 1885350.0 ;
      RECT  96900.0 1886550.0 98100.0 1885350.0 ;
      RECT  99300.0 1886550.0 100500.0 1885350.0 ;
      RECT  99300.0 1886550.0 100500.0 1885350.0 ;
      RECT  96900.0 1886550.0 98100.0 1885350.0 ;
      RECT  99300.0 1886550.0 100500.0 1885350.0 ;
      RECT  101700.0 1886550.0 102900.0 1885350.0 ;
      RECT  101700.0 1886550.0 102900.0 1885350.0 ;
      RECT  99300.0 1886550.0 100500.0 1885350.0 ;
      RECT  94500.0 1895250.0 95700.0 1894050.0 ;
      RECT  96900.0 1895250.0 98100.0 1894050.0 ;
      RECT  96900.0 1895250.0 98100.0 1894050.0 ;
      RECT  94500.0 1895250.0 95700.0 1894050.0 ;
      RECT  96900.0 1895250.0 98100.0 1894050.0 ;
      RECT  99300.0 1895250.0 100500.0 1894050.0 ;
      RECT  99300.0 1895250.0 100500.0 1894050.0 ;
      RECT  96900.0 1895250.0 98100.0 1894050.0 ;
      RECT  99300.0 1895250.0 100500.0 1894050.0 ;
      RECT  101700.0 1895250.0 102900.0 1894050.0 ;
      RECT  101700.0 1895250.0 102900.0 1894050.0 ;
      RECT  99300.0 1895250.0 100500.0 1894050.0 ;
      RECT  104100.0 1885950.0 105300.0 1884750.0 ;
      RECT  104100.0 1895850.0 105300.0 1894650.0 ;
      RECT  101700.0 1893150.0 100500.0 1891950.0 ;
      RECT  99300.0 1891200.0 98100.0 1890000.0 ;
      RECT  96900.0 1889250.0 95700.0 1888050.0 ;
      RECT  96900.0 1886550.0 98100.0 1885350.0 ;
      RECT  101700.0 1886550.0 102900.0 1885350.0 ;
      RECT  101700.0 1895250.0 102900.0 1894050.0 ;
      RECT  101700.0 1889250.0 102900.0 1888050.0 ;
      RECT  95700.0 1889250.0 96900.0 1888050.0 ;
      RECT  98100.0 1891200.0 99300.0 1890000.0 ;
      RECT  100500.0 1893150.0 101700.0 1891950.0 ;
      RECT  101700.0 1889250.0 102900.0 1888050.0 ;
      RECT  92700.0 1883850.0 108300.0 1882950.0 ;
      RECT  92700.0 1897650.0 108300.0 1896750.0 ;
      RECT  94500.0 1899150.0 95700.0 1896750.0 ;
      RECT  94500.0 1907850.0 95700.0 1911450.0 ;
      RECT  99300.0 1907850.0 100500.0 1911450.0 ;
      RECT  104100.0 1909050.0 105300.0 1911000.0 ;
      RECT  104100.0 1897200.0 105300.0 1899150.0 ;
      RECT  94500.0 1907850.0 95700.0 1909050.0 ;
      RECT  96900.0 1907850.0 98100.0 1909050.0 ;
      RECT  96900.0 1907850.0 98100.0 1909050.0 ;
      RECT  94500.0 1907850.0 95700.0 1909050.0 ;
      RECT  96900.0 1907850.0 98100.0 1909050.0 ;
      RECT  99300.0 1907850.0 100500.0 1909050.0 ;
      RECT  99300.0 1907850.0 100500.0 1909050.0 ;
      RECT  96900.0 1907850.0 98100.0 1909050.0 ;
      RECT  99300.0 1907850.0 100500.0 1909050.0 ;
      RECT  101700.0 1907850.0 102900.0 1909050.0 ;
      RECT  101700.0 1907850.0 102900.0 1909050.0 ;
      RECT  99300.0 1907850.0 100500.0 1909050.0 ;
      RECT  94500.0 1899150.0 95700.0 1900350.0 ;
      RECT  96900.0 1899150.0 98100.0 1900350.0 ;
      RECT  96900.0 1899150.0 98100.0 1900350.0 ;
      RECT  94500.0 1899150.0 95700.0 1900350.0 ;
      RECT  96900.0 1899150.0 98100.0 1900350.0 ;
      RECT  99300.0 1899150.0 100500.0 1900350.0 ;
      RECT  99300.0 1899150.0 100500.0 1900350.0 ;
      RECT  96900.0 1899150.0 98100.0 1900350.0 ;
      RECT  99300.0 1899150.0 100500.0 1900350.0 ;
      RECT  101700.0 1899150.0 102900.0 1900350.0 ;
      RECT  101700.0 1899150.0 102900.0 1900350.0 ;
      RECT  99300.0 1899150.0 100500.0 1900350.0 ;
      RECT  104100.0 1908450.0 105300.0 1909650.0 ;
      RECT  104100.0 1898550.0 105300.0 1899750.0 ;
      RECT  101700.0 1901250.0 100500.0 1902450.0 ;
      RECT  99300.0 1903200.0 98100.0 1904400.0 ;
      RECT  96900.0 1905150.0 95700.0 1906350.0 ;
      RECT  96900.0 1907850.0 98100.0 1909050.0 ;
      RECT  101700.0 1907850.0 102900.0 1909050.0 ;
      RECT  101700.0 1899150.0 102900.0 1900350.0 ;
      RECT  101700.0 1905150.0 102900.0 1906350.0 ;
      RECT  95700.0 1905150.0 96900.0 1906350.0 ;
      RECT  98100.0 1903200.0 99300.0 1904400.0 ;
      RECT  100500.0 1901250.0 101700.0 1902450.0 ;
      RECT  101700.0 1905150.0 102900.0 1906350.0 ;
      RECT  92700.0 1910550.0 108300.0 1911450.0 ;
      RECT  92700.0 1896750.0 108300.0 1897650.0 ;
      RECT  94500.0 1922850.0 95700.0 1925250.0 ;
      RECT  94500.0 1914150.0 95700.0 1910550.0 ;
      RECT  99300.0 1914150.0 100500.0 1910550.0 ;
      RECT  104100.0 1912950.0 105300.0 1911000.0 ;
      RECT  104100.0 1924800.0 105300.0 1922850.0 ;
      RECT  94500.0 1914150.0 95700.0 1912950.0 ;
      RECT  96900.0 1914150.0 98100.0 1912950.0 ;
      RECT  96900.0 1914150.0 98100.0 1912950.0 ;
      RECT  94500.0 1914150.0 95700.0 1912950.0 ;
      RECT  96900.0 1914150.0 98100.0 1912950.0 ;
      RECT  99300.0 1914150.0 100500.0 1912950.0 ;
      RECT  99300.0 1914150.0 100500.0 1912950.0 ;
      RECT  96900.0 1914150.0 98100.0 1912950.0 ;
      RECT  99300.0 1914150.0 100500.0 1912950.0 ;
      RECT  101700.0 1914150.0 102900.0 1912950.0 ;
      RECT  101700.0 1914150.0 102900.0 1912950.0 ;
      RECT  99300.0 1914150.0 100500.0 1912950.0 ;
      RECT  94500.0 1922850.0 95700.0 1921650.0 ;
      RECT  96900.0 1922850.0 98100.0 1921650.0 ;
      RECT  96900.0 1922850.0 98100.0 1921650.0 ;
      RECT  94500.0 1922850.0 95700.0 1921650.0 ;
      RECT  96900.0 1922850.0 98100.0 1921650.0 ;
      RECT  99300.0 1922850.0 100500.0 1921650.0 ;
      RECT  99300.0 1922850.0 100500.0 1921650.0 ;
      RECT  96900.0 1922850.0 98100.0 1921650.0 ;
      RECT  99300.0 1922850.0 100500.0 1921650.0 ;
      RECT  101700.0 1922850.0 102900.0 1921650.0 ;
      RECT  101700.0 1922850.0 102900.0 1921650.0 ;
      RECT  99300.0 1922850.0 100500.0 1921650.0 ;
      RECT  104100.0 1913550.0 105300.0 1912350.0 ;
      RECT  104100.0 1923450.0 105300.0 1922250.0 ;
      RECT  101700.0 1920750.0 100500.0 1919550.0 ;
      RECT  99300.0 1918800.0 98100.0 1917600.0 ;
      RECT  96900.0 1916850.0 95700.0 1915650.0 ;
      RECT  96900.0 1914150.0 98100.0 1912950.0 ;
      RECT  101700.0 1914150.0 102900.0 1912950.0 ;
      RECT  101700.0 1922850.0 102900.0 1921650.0 ;
      RECT  101700.0 1916850.0 102900.0 1915650.0 ;
      RECT  95700.0 1916850.0 96900.0 1915650.0 ;
      RECT  98100.0 1918800.0 99300.0 1917600.0 ;
      RECT  100500.0 1920750.0 101700.0 1919550.0 ;
      RECT  101700.0 1916850.0 102900.0 1915650.0 ;
      RECT  92700.0 1911450.0 108300.0 1910550.0 ;
      RECT  92700.0 1925250.0 108300.0 1924350.0 ;
      RECT  94500.0 1926750.0 95700.0 1924350.0 ;
      RECT  94500.0 1935450.0 95700.0 1939050.0 ;
      RECT  99300.0 1935450.0 100500.0 1939050.0 ;
      RECT  104100.0 1936650.0 105300.0 1938600.0 ;
      RECT  104100.0 1924800.0 105300.0 1926750.0 ;
      RECT  94500.0 1935450.0 95700.0 1936650.0 ;
      RECT  96900.0 1935450.0 98100.0 1936650.0 ;
      RECT  96900.0 1935450.0 98100.0 1936650.0 ;
      RECT  94500.0 1935450.0 95700.0 1936650.0 ;
      RECT  96900.0 1935450.0 98100.0 1936650.0 ;
      RECT  99300.0 1935450.0 100500.0 1936650.0 ;
      RECT  99300.0 1935450.0 100500.0 1936650.0 ;
      RECT  96900.0 1935450.0 98100.0 1936650.0 ;
      RECT  99300.0 1935450.0 100500.0 1936650.0 ;
      RECT  101700.0 1935450.0 102900.0 1936650.0 ;
      RECT  101700.0 1935450.0 102900.0 1936650.0 ;
      RECT  99300.0 1935450.0 100500.0 1936650.0 ;
      RECT  94500.0 1926750.0 95700.0 1927950.0 ;
      RECT  96900.0 1926750.0 98100.0 1927950.0 ;
      RECT  96900.0 1926750.0 98100.0 1927950.0 ;
      RECT  94500.0 1926750.0 95700.0 1927950.0 ;
      RECT  96900.0 1926750.0 98100.0 1927950.0 ;
      RECT  99300.0 1926750.0 100500.0 1927950.0 ;
      RECT  99300.0 1926750.0 100500.0 1927950.0 ;
      RECT  96900.0 1926750.0 98100.0 1927950.0 ;
      RECT  99300.0 1926750.0 100500.0 1927950.0 ;
      RECT  101700.0 1926750.0 102900.0 1927950.0 ;
      RECT  101700.0 1926750.0 102900.0 1927950.0 ;
      RECT  99300.0 1926750.0 100500.0 1927950.0 ;
      RECT  104100.0 1936050.0 105300.0 1937250.0 ;
      RECT  104100.0 1926150.0 105300.0 1927350.0 ;
      RECT  101700.0 1928850.0 100500.0 1930050.0 ;
      RECT  99300.0 1930800.0 98100.0 1932000.0 ;
      RECT  96900.0 1932750.0 95700.0 1933950.0 ;
      RECT  96900.0 1935450.0 98100.0 1936650.0 ;
      RECT  101700.0 1935450.0 102900.0 1936650.0 ;
      RECT  101700.0 1926750.0 102900.0 1927950.0 ;
      RECT  101700.0 1932750.0 102900.0 1933950.0 ;
      RECT  95700.0 1932750.0 96900.0 1933950.0 ;
      RECT  98100.0 1930800.0 99300.0 1932000.0 ;
      RECT  100500.0 1928850.0 101700.0 1930050.0 ;
      RECT  101700.0 1932750.0 102900.0 1933950.0 ;
      RECT  92700.0 1938150.0 108300.0 1939050.0 ;
      RECT  92700.0 1924350.0 108300.0 1925250.0 ;
      RECT  94500.0 1950450.0 95700.0 1952850.0 ;
      RECT  94500.0 1941750.0 95700.0 1938150.0 ;
      RECT  99300.0 1941750.0 100500.0 1938150.0 ;
      RECT  104100.0 1940550.0 105300.0 1938600.0 ;
      RECT  104100.0 1952400.0 105300.0 1950450.0 ;
      RECT  94500.0 1941750.0 95700.0 1940550.0 ;
      RECT  96900.0 1941750.0 98100.0 1940550.0 ;
      RECT  96900.0 1941750.0 98100.0 1940550.0 ;
      RECT  94500.0 1941750.0 95700.0 1940550.0 ;
      RECT  96900.0 1941750.0 98100.0 1940550.0 ;
      RECT  99300.0 1941750.0 100500.0 1940550.0 ;
      RECT  99300.0 1941750.0 100500.0 1940550.0 ;
      RECT  96900.0 1941750.0 98100.0 1940550.0 ;
      RECT  99300.0 1941750.0 100500.0 1940550.0 ;
      RECT  101700.0 1941750.0 102900.0 1940550.0 ;
      RECT  101700.0 1941750.0 102900.0 1940550.0 ;
      RECT  99300.0 1941750.0 100500.0 1940550.0 ;
      RECT  94500.0 1950450.0 95700.0 1949250.0 ;
      RECT  96900.0 1950450.0 98100.0 1949250.0 ;
      RECT  96900.0 1950450.0 98100.0 1949250.0 ;
      RECT  94500.0 1950450.0 95700.0 1949250.0 ;
      RECT  96900.0 1950450.0 98100.0 1949250.0 ;
      RECT  99300.0 1950450.0 100500.0 1949250.0 ;
      RECT  99300.0 1950450.0 100500.0 1949250.0 ;
      RECT  96900.0 1950450.0 98100.0 1949250.0 ;
      RECT  99300.0 1950450.0 100500.0 1949250.0 ;
      RECT  101700.0 1950450.0 102900.0 1949250.0 ;
      RECT  101700.0 1950450.0 102900.0 1949250.0 ;
      RECT  99300.0 1950450.0 100500.0 1949250.0 ;
      RECT  104100.0 1941150.0 105300.0 1939950.0 ;
      RECT  104100.0 1951050.0 105300.0 1949850.0 ;
      RECT  101700.0 1948350.0 100500.0 1947150.0 ;
      RECT  99300.0 1946400.0 98100.0 1945200.0 ;
      RECT  96900.0 1944450.0 95700.0 1943250.0 ;
      RECT  96900.0 1941750.0 98100.0 1940550.0 ;
      RECT  101700.0 1941750.0 102900.0 1940550.0 ;
      RECT  101700.0 1950450.0 102900.0 1949250.0 ;
      RECT  101700.0 1944450.0 102900.0 1943250.0 ;
      RECT  95700.0 1944450.0 96900.0 1943250.0 ;
      RECT  98100.0 1946400.0 99300.0 1945200.0 ;
      RECT  100500.0 1948350.0 101700.0 1947150.0 ;
      RECT  101700.0 1944450.0 102900.0 1943250.0 ;
      RECT  92700.0 1939050.0 108300.0 1938150.0 ;
      RECT  92700.0 1952850.0 108300.0 1951950.0 ;
      RECT  94500.0 1954350.0 95700.0 1951950.0 ;
      RECT  94500.0 1963050.0 95700.0 1966650.0 ;
      RECT  99300.0 1963050.0 100500.0 1966650.0 ;
      RECT  104100.0 1964250.0 105300.0 1966200.0 ;
      RECT  104100.0 1952400.0 105300.0 1954350.0 ;
      RECT  94500.0 1963050.0 95700.0 1964250.0 ;
      RECT  96900.0 1963050.0 98100.0 1964250.0 ;
      RECT  96900.0 1963050.0 98100.0 1964250.0 ;
      RECT  94500.0 1963050.0 95700.0 1964250.0 ;
      RECT  96900.0 1963050.0 98100.0 1964250.0 ;
      RECT  99300.0 1963050.0 100500.0 1964250.0 ;
      RECT  99300.0 1963050.0 100500.0 1964250.0 ;
      RECT  96900.0 1963050.0 98100.0 1964250.0 ;
      RECT  99300.0 1963050.0 100500.0 1964250.0 ;
      RECT  101700.0 1963050.0 102900.0 1964250.0 ;
      RECT  101700.0 1963050.0 102900.0 1964250.0 ;
      RECT  99300.0 1963050.0 100500.0 1964250.0 ;
      RECT  94500.0 1954350.0 95700.0 1955550.0 ;
      RECT  96900.0 1954350.0 98100.0 1955550.0 ;
      RECT  96900.0 1954350.0 98100.0 1955550.0 ;
      RECT  94500.0 1954350.0 95700.0 1955550.0 ;
      RECT  96900.0 1954350.0 98100.0 1955550.0 ;
      RECT  99300.0 1954350.0 100500.0 1955550.0 ;
      RECT  99300.0 1954350.0 100500.0 1955550.0 ;
      RECT  96900.0 1954350.0 98100.0 1955550.0 ;
      RECT  99300.0 1954350.0 100500.0 1955550.0 ;
      RECT  101700.0 1954350.0 102900.0 1955550.0 ;
      RECT  101700.0 1954350.0 102900.0 1955550.0 ;
      RECT  99300.0 1954350.0 100500.0 1955550.0 ;
      RECT  104100.0 1963650.0 105300.0 1964850.0 ;
      RECT  104100.0 1953750.0 105300.0 1954950.0 ;
      RECT  101700.0 1956450.0 100500.0 1957650.0 ;
      RECT  99300.0 1958400.0 98100.0 1959600.0 ;
      RECT  96900.0 1960350.0 95700.0 1961550.0 ;
      RECT  96900.0 1963050.0 98100.0 1964250.0 ;
      RECT  101700.0 1963050.0 102900.0 1964250.0 ;
      RECT  101700.0 1954350.0 102900.0 1955550.0 ;
      RECT  101700.0 1960350.0 102900.0 1961550.0 ;
      RECT  95700.0 1960350.0 96900.0 1961550.0 ;
      RECT  98100.0 1958400.0 99300.0 1959600.0 ;
      RECT  100500.0 1956450.0 101700.0 1957650.0 ;
      RECT  101700.0 1960350.0 102900.0 1961550.0 ;
      RECT  92700.0 1965750.0 108300.0 1966650.0 ;
      RECT  92700.0 1951950.0 108300.0 1952850.0 ;
      RECT  94500.0 1978050.0 95700.0 1980450.0 ;
      RECT  94500.0 1969350.0 95700.0 1965750.0 ;
      RECT  99300.0 1969350.0 100500.0 1965750.0 ;
      RECT  104100.0 1968150.0 105300.0 1966200.0 ;
      RECT  104100.0 1980000.0 105300.0 1978050.0 ;
      RECT  94500.0 1969350.0 95700.0 1968150.0 ;
      RECT  96900.0 1969350.0 98100.0 1968150.0 ;
      RECT  96900.0 1969350.0 98100.0 1968150.0 ;
      RECT  94500.0 1969350.0 95700.0 1968150.0 ;
      RECT  96900.0 1969350.0 98100.0 1968150.0 ;
      RECT  99300.0 1969350.0 100500.0 1968150.0 ;
      RECT  99300.0 1969350.0 100500.0 1968150.0 ;
      RECT  96900.0 1969350.0 98100.0 1968150.0 ;
      RECT  99300.0 1969350.0 100500.0 1968150.0 ;
      RECT  101700.0 1969350.0 102900.0 1968150.0 ;
      RECT  101700.0 1969350.0 102900.0 1968150.0 ;
      RECT  99300.0 1969350.0 100500.0 1968150.0 ;
      RECT  94500.0 1978050.0 95700.0 1976850.0 ;
      RECT  96900.0 1978050.0 98100.0 1976850.0 ;
      RECT  96900.0 1978050.0 98100.0 1976850.0 ;
      RECT  94500.0 1978050.0 95700.0 1976850.0 ;
      RECT  96900.0 1978050.0 98100.0 1976850.0 ;
      RECT  99300.0 1978050.0 100500.0 1976850.0 ;
      RECT  99300.0 1978050.0 100500.0 1976850.0 ;
      RECT  96900.0 1978050.0 98100.0 1976850.0 ;
      RECT  99300.0 1978050.0 100500.0 1976850.0 ;
      RECT  101700.0 1978050.0 102900.0 1976850.0 ;
      RECT  101700.0 1978050.0 102900.0 1976850.0 ;
      RECT  99300.0 1978050.0 100500.0 1976850.0 ;
      RECT  104100.0 1968750.0 105300.0 1967550.0 ;
      RECT  104100.0 1978650.0 105300.0 1977450.0 ;
      RECT  101700.0 1975950.0 100500.0 1974750.0 ;
      RECT  99300.0 1974000.0 98100.0 1972800.0 ;
      RECT  96900.0 1972050.0 95700.0 1970850.0 ;
      RECT  96900.0 1969350.0 98100.0 1968150.0 ;
      RECT  101700.0 1969350.0 102900.0 1968150.0 ;
      RECT  101700.0 1978050.0 102900.0 1976850.0 ;
      RECT  101700.0 1972050.0 102900.0 1970850.0 ;
      RECT  95700.0 1972050.0 96900.0 1970850.0 ;
      RECT  98100.0 1974000.0 99300.0 1972800.0 ;
      RECT  100500.0 1975950.0 101700.0 1974750.0 ;
      RECT  101700.0 1972050.0 102900.0 1970850.0 ;
      RECT  92700.0 1966650.0 108300.0 1965750.0 ;
      RECT  92700.0 1980450.0 108300.0 1979550.0 ;
      RECT  94500.0 1981950.0 95700.0 1979550.0 ;
      RECT  94500.0 1990650.0 95700.0 1994250.0 ;
      RECT  99300.0 1990650.0 100500.0 1994250.0 ;
      RECT  104100.0 1991850.0 105300.0 1993800.0 ;
      RECT  104100.0 1980000.0 105300.0 1981950.0 ;
      RECT  94500.0 1990650.0 95700.0 1991850.0 ;
      RECT  96900.0 1990650.0 98100.0 1991850.0 ;
      RECT  96900.0 1990650.0 98100.0 1991850.0 ;
      RECT  94500.0 1990650.0 95700.0 1991850.0 ;
      RECT  96900.0 1990650.0 98100.0 1991850.0 ;
      RECT  99300.0 1990650.0 100500.0 1991850.0 ;
      RECT  99300.0 1990650.0 100500.0 1991850.0 ;
      RECT  96900.0 1990650.0 98100.0 1991850.0 ;
      RECT  99300.0 1990650.0 100500.0 1991850.0 ;
      RECT  101700.0 1990650.0 102900.0 1991850.0 ;
      RECT  101700.0 1990650.0 102900.0 1991850.0 ;
      RECT  99300.0 1990650.0 100500.0 1991850.0 ;
      RECT  94500.0 1981950.0 95700.0 1983150.0 ;
      RECT  96900.0 1981950.0 98100.0 1983150.0 ;
      RECT  96900.0 1981950.0 98100.0 1983150.0 ;
      RECT  94500.0 1981950.0 95700.0 1983150.0 ;
      RECT  96900.0 1981950.0 98100.0 1983150.0 ;
      RECT  99300.0 1981950.0 100500.0 1983150.0 ;
      RECT  99300.0 1981950.0 100500.0 1983150.0 ;
      RECT  96900.0 1981950.0 98100.0 1983150.0 ;
      RECT  99300.0 1981950.0 100500.0 1983150.0 ;
      RECT  101700.0 1981950.0 102900.0 1983150.0 ;
      RECT  101700.0 1981950.0 102900.0 1983150.0 ;
      RECT  99300.0 1981950.0 100500.0 1983150.0 ;
      RECT  104100.0 1991250.0 105300.0 1992450.0 ;
      RECT  104100.0 1981350.0 105300.0 1982550.0 ;
      RECT  101700.0 1984050.0 100500.0 1985250.0 ;
      RECT  99300.0 1986000.0 98100.0 1987200.0 ;
      RECT  96900.0 1987950.0 95700.0 1989150.0 ;
      RECT  96900.0 1990650.0 98100.0 1991850.0 ;
      RECT  101700.0 1990650.0 102900.0 1991850.0 ;
      RECT  101700.0 1981950.0 102900.0 1983150.0 ;
      RECT  101700.0 1987950.0 102900.0 1989150.0 ;
      RECT  95700.0 1987950.0 96900.0 1989150.0 ;
      RECT  98100.0 1986000.0 99300.0 1987200.0 ;
      RECT  100500.0 1984050.0 101700.0 1985250.0 ;
      RECT  101700.0 1987950.0 102900.0 1989150.0 ;
      RECT  92700.0 1993350.0 108300.0 1994250.0 ;
      RECT  92700.0 1979550.0 108300.0 1980450.0 ;
      RECT  94500.0 2005650.0 95700.0 2008050.0 ;
      RECT  94500.0 1996950.0 95700.0 1993350.0 ;
      RECT  99300.0 1996950.0 100500.0 1993350.0 ;
      RECT  104100.0 1995750.0 105300.0 1993800.0 ;
      RECT  104100.0 2007600.0 105300.0 2005650.0 ;
      RECT  94500.0 1996950.0 95700.0 1995750.0 ;
      RECT  96900.0 1996950.0 98100.0 1995750.0 ;
      RECT  96900.0 1996950.0 98100.0 1995750.0 ;
      RECT  94500.0 1996950.0 95700.0 1995750.0 ;
      RECT  96900.0 1996950.0 98100.0 1995750.0 ;
      RECT  99300.0 1996950.0 100500.0 1995750.0 ;
      RECT  99300.0 1996950.0 100500.0 1995750.0 ;
      RECT  96900.0 1996950.0 98100.0 1995750.0 ;
      RECT  99300.0 1996950.0 100500.0 1995750.0 ;
      RECT  101700.0 1996950.0 102900.0 1995750.0 ;
      RECT  101700.0 1996950.0 102900.0 1995750.0 ;
      RECT  99300.0 1996950.0 100500.0 1995750.0 ;
      RECT  94500.0 2005650.0 95700.0 2004450.0 ;
      RECT  96900.0 2005650.0 98100.0 2004450.0 ;
      RECT  96900.0 2005650.0 98100.0 2004450.0 ;
      RECT  94500.0 2005650.0 95700.0 2004450.0 ;
      RECT  96900.0 2005650.0 98100.0 2004450.0 ;
      RECT  99300.0 2005650.0 100500.0 2004450.0 ;
      RECT  99300.0 2005650.0 100500.0 2004450.0 ;
      RECT  96900.0 2005650.0 98100.0 2004450.0 ;
      RECT  99300.0 2005650.0 100500.0 2004450.0 ;
      RECT  101700.0 2005650.0 102900.0 2004450.0 ;
      RECT  101700.0 2005650.0 102900.0 2004450.0 ;
      RECT  99300.0 2005650.0 100500.0 2004450.0 ;
      RECT  104100.0 1996350.0 105300.0 1995150.0 ;
      RECT  104100.0 2006250.0 105300.0 2005050.0 ;
      RECT  101700.0 2003550.0 100500.0 2002350.0 ;
      RECT  99300.0 2001600.0 98100.0 2000400.0 ;
      RECT  96900.0 1999650.0 95700.0 1998450.0 ;
      RECT  96900.0 1996950.0 98100.0 1995750.0 ;
      RECT  101700.0 1996950.0 102900.0 1995750.0 ;
      RECT  101700.0 2005650.0 102900.0 2004450.0 ;
      RECT  101700.0 1999650.0 102900.0 1998450.0 ;
      RECT  95700.0 1999650.0 96900.0 1998450.0 ;
      RECT  98100.0 2001600.0 99300.0 2000400.0 ;
      RECT  100500.0 2003550.0 101700.0 2002350.0 ;
      RECT  101700.0 1999650.0 102900.0 1998450.0 ;
      RECT  92700.0 1994250.0 108300.0 1993350.0 ;
      RECT  92700.0 2008050.0 108300.0 2007150.0 ;
      RECT  94500.0 2009550.0 95700.0 2007150.0 ;
      RECT  94500.0 2018250.0 95700.0 2021850.0 ;
      RECT  99300.0 2018250.0 100500.0 2021850.0 ;
      RECT  104100.0 2019450.0 105300.0 2021400.0 ;
      RECT  104100.0 2007600.0 105300.0 2009550.0 ;
      RECT  94500.0 2018250.0 95700.0 2019450.0 ;
      RECT  96900.0 2018250.0 98100.0 2019450.0 ;
      RECT  96900.0 2018250.0 98100.0 2019450.0 ;
      RECT  94500.0 2018250.0 95700.0 2019450.0 ;
      RECT  96900.0 2018250.0 98100.0 2019450.0 ;
      RECT  99300.0 2018250.0 100500.0 2019450.0 ;
      RECT  99300.0 2018250.0 100500.0 2019450.0 ;
      RECT  96900.0 2018250.0 98100.0 2019450.0 ;
      RECT  99300.0 2018250.0 100500.0 2019450.0 ;
      RECT  101700.0 2018250.0 102900.0 2019450.0 ;
      RECT  101700.0 2018250.0 102900.0 2019450.0 ;
      RECT  99300.0 2018250.0 100500.0 2019450.0 ;
      RECT  94500.0 2009550.0 95700.0 2010750.0 ;
      RECT  96900.0 2009550.0 98100.0 2010750.0 ;
      RECT  96900.0 2009550.0 98100.0 2010750.0 ;
      RECT  94500.0 2009550.0 95700.0 2010750.0 ;
      RECT  96900.0 2009550.0 98100.0 2010750.0 ;
      RECT  99300.0 2009550.0 100500.0 2010750.0 ;
      RECT  99300.0 2009550.0 100500.0 2010750.0 ;
      RECT  96900.0 2009550.0 98100.0 2010750.0 ;
      RECT  99300.0 2009550.0 100500.0 2010750.0 ;
      RECT  101700.0 2009550.0 102900.0 2010750.0 ;
      RECT  101700.0 2009550.0 102900.0 2010750.0 ;
      RECT  99300.0 2009550.0 100500.0 2010750.0 ;
      RECT  104100.0 2018850.0 105300.0 2020050.0 ;
      RECT  104100.0 2008950.0 105300.0 2010150.0 ;
      RECT  101700.0 2011650.0 100500.0 2012850.0 ;
      RECT  99300.0 2013600.0 98100.0 2014800.0 ;
      RECT  96900.0 2015550.0 95700.0 2016750.0 ;
      RECT  96900.0 2018250.0 98100.0 2019450.0 ;
      RECT  101700.0 2018250.0 102900.0 2019450.0 ;
      RECT  101700.0 2009550.0 102900.0 2010750.0 ;
      RECT  101700.0 2015550.0 102900.0 2016750.0 ;
      RECT  95700.0 2015550.0 96900.0 2016750.0 ;
      RECT  98100.0 2013600.0 99300.0 2014800.0 ;
      RECT  100500.0 2011650.0 101700.0 2012850.0 ;
      RECT  101700.0 2015550.0 102900.0 2016750.0 ;
      RECT  92700.0 2020950.0 108300.0 2021850.0 ;
      RECT  92700.0 2007150.0 108300.0 2008050.0 ;
      RECT  94500.0 2033250.0 95700.0 2035650.0 ;
      RECT  94500.0 2024550.0 95700.0 2020950.0 ;
      RECT  99300.0 2024550.0 100500.0 2020950.0 ;
      RECT  104100.0 2023350.0 105300.0 2021400.0 ;
      RECT  104100.0 2035200.0 105300.0 2033250.0 ;
      RECT  94500.0 2024550.0 95700.0 2023350.0 ;
      RECT  96900.0 2024550.0 98100.0 2023350.0 ;
      RECT  96900.0 2024550.0 98100.0 2023350.0 ;
      RECT  94500.0 2024550.0 95700.0 2023350.0 ;
      RECT  96900.0 2024550.0 98100.0 2023350.0 ;
      RECT  99300.0 2024550.0 100500.0 2023350.0 ;
      RECT  99300.0 2024550.0 100500.0 2023350.0 ;
      RECT  96900.0 2024550.0 98100.0 2023350.0 ;
      RECT  99300.0 2024550.0 100500.0 2023350.0 ;
      RECT  101700.0 2024550.0 102900.0 2023350.0 ;
      RECT  101700.0 2024550.0 102900.0 2023350.0 ;
      RECT  99300.0 2024550.0 100500.0 2023350.0 ;
      RECT  94500.0 2033250.0 95700.0 2032050.0 ;
      RECT  96900.0 2033250.0 98100.0 2032050.0 ;
      RECT  96900.0 2033250.0 98100.0 2032050.0 ;
      RECT  94500.0 2033250.0 95700.0 2032050.0 ;
      RECT  96900.0 2033250.0 98100.0 2032050.0 ;
      RECT  99300.0 2033250.0 100500.0 2032050.0 ;
      RECT  99300.0 2033250.0 100500.0 2032050.0 ;
      RECT  96900.0 2033250.0 98100.0 2032050.0 ;
      RECT  99300.0 2033250.0 100500.0 2032050.0 ;
      RECT  101700.0 2033250.0 102900.0 2032050.0 ;
      RECT  101700.0 2033250.0 102900.0 2032050.0 ;
      RECT  99300.0 2033250.0 100500.0 2032050.0 ;
      RECT  104100.0 2023950.0 105300.0 2022750.0 ;
      RECT  104100.0 2033850.0 105300.0 2032650.0 ;
      RECT  101700.0 2031150.0 100500.0 2029950.0 ;
      RECT  99300.0 2029200.0 98100.0 2028000.0 ;
      RECT  96900.0 2027250.0 95700.0 2026050.0 ;
      RECT  96900.0 2024550.0 98100.0 2023350.0 ;
      RECT  101700.0 2024550.0 102900.0 2023350.0 ;
      RECT  101700.0 2033250.0 102900.0 2032050.0 ;
      RECT  101700.0 2027250.0 102900.0 2026050.0 ;
      RECT  95700.0 2027250.0 96900.0 2026050.0 ;
      RECT  98100.0 2029200.0 99300.0 2028000.0 ;
      RECT  100500.0 2031150.0 101700.0 2029950.0 ;
      RECT  101700.0 2027250.0 102900.0 2026050.0 ;
      RECT  92700.0 2021850.0 108300.0 2020950.0 ;
      RECT  92700.0 2035650.0 108300.0 2034750.0 ;
      RECT  94500.0 2037150.0 95700.0 2034750.0 ;
      RECT  94500.0 2045850.0 95700.0 2049450.0 ;
      RECT  99300.0 2045850.0 100500.0 2049450.0 ;
      RECT  104100.0 2047050.0 105300.0 2049000.0 ;
      RECT  104100.0 2035200.0 105300.0 2037150.0 ;
      RECT  94500.0 2045850.0 95700.0 2047050.0 ;
      RECT  96900.0 2045850.0 98100.0 2047050.0 ;
      RECT  96900.0 2045850.0 98100.0 2047050.0 ;
      RECT  94500.0 2045850.0 95700.0 2047050.0 ;
      RECT  96900.0 2045850.0 98100.0 2047050.0 ;
      RECT  99300.0 2045850.0 100500.0 2047050.0 ;
      RECT  99300.0 2045850.0 100500.0 2047050.0 ;
      RECT  96900.0 2045850.0 98100.0 2047050.0 ;
      RECT  99300.0 2045850.0 100500.0 2047050.0 ;
      RECT  101700.0 2045850.0 102900.0 2047050.0 ;
      RECT  101700.0 2045850.0 102900.0 2047050.0 ;
      RECT  99300.0 2045850.0 100500.0 2047050.0 ;
      RECT  94500.0 2037150.0 95700.0 2038350.0 ;
      RECT  96900.0 2037150.0 98100.0 2038350.0 ;
      RECT  96900.0 2037150.0 98100.0 2038350.0 ;
      RECT  94500.0 2037150.0 95700.0 2038350.0 ;
      RECT  96900.0 2037150.0 98100.0 2038350.0 ;
      RECT  99300.0 2037150.0 100500.0 2038350.0 ;
      RECT  99300.0 2037150.0 100500.0 2038350.0 ;
      RECT  96900.0 2037150.0 98100.0 2038350.0 ;
      RECT  99300.0 2037150.0 100500.0 2038350.0 ;
      RECT  101700.0 2037150.0 102900.0 2038350.0 ;
      RECT  101700.0 2037150.0 102900.0 2038350.0 ;
      RECT  99300.0 2037150.0 100500.0 2038350.0 ;
      RECT  104100.0 2046450.0 105300.0 2047650.0 ;
      RECT  104100.0 2036550.0 105300.0 2037750.0 ;
      RECT  101700.0 2039250.0 100500.0 2040450.0 ;
      RECT  99300.0 2041200.0 98100.0 2042400.0 ;
      RECT  96900.0 2043150.0 95700.0 2044350.0 ;
      RECT  96900.0 2045850.0 98100.0 2047050.0 ;
      RECT  101700.0 2045850.0 102900.0 2047050.0 ;
      RECT  101700.0 2037150.0 102900.0 2038350.0 ;
      RECT  101700.0 2043150.0 102900.0 2044350.0 ;
      RECT  95700.0 2043150.0 96900.0 2044350.0 ;
      RECT  98100.0 2041200.0 99300.0 2042400.0 ;
      RECT  100500.0 2039250.0 101700.0 2040450.0 ;
      RECT  101700.0 2043150.0 102900.0 2044350.0 ;
      RECT  92700.0 2048550.0 108300.0 2049450.0 ;
      RECT  92700.0 2034750.0 108300.0 2035650.0 ;
      RECT  94500.0 2060850.0 95700.0 2063250.0 ;
      RECT  94500.0 2052150.0 95700.0 2048550.0 ;
      RECT  99300.0 2052150.0 100500.0 2048550.0 ;
      RECT  104100.0 2050950.0 105300.0 2049000.0 ;
      RECT  104100.0 2062800.0 105300.0 2060850.0 ;
      RECT  94500.0 2052150.0 95700.0 2050950.0 ;
      RECT  96900.0 2052150.0 98100.0 2050950.0 ;
      RECT  96900.0 2052150.0 98100.0 2050950.0 ;
      RECT  94500.0 2052150.0 95700.0 2050950.0 ;
      RECT  96900.0 2052150.0 98100.0 2050950.0 ;
      RECT  99300.0 2052150.0 100500.0 2050950.0 ;
      RECT  99300.0 2052150.0 100500.0 2050950.0 ;
      RECT  96900.0 2052150.0 98100.0 2050950.0 ;
      RECT  99300.0 2052150.0 100500.0 2050950.0 ;
      RECT  101700.0 2052150.0 102900.0 2050950.0 ;
      RECT  101700.0 2052150.0 102900.0 2050950.0 ;
      RECT  99300.0 2052150.0 100500.0 2050950.0 ;
      RECT  94500.0 2060850.0 95700.0 2059650.0 ;
      RECT  96900.0 2060850.0 98100.0 2059650.0 ;
      RECT  96900.0 2060850.0 98100.0 2059650.0 ;
      RECT  94500.0 2060850.0 95700.0 2059650.0 ;
      RECT  96900.0 2060850.0 98100.0 2059650.0 ;
      RECT  99300.0 2060850.0 100500.0 2059650.0 ;
      RECT  99300.0 2060850.0 100500.0 2059650.0 ;
      RECT  96900.0 2060850.0 98100.0 2059650.0 ;
      RECT  99300.0 2060850.0 100500.0 2059650.0 ;
      RECT  101700.0 2060850.0 102900.0 2059650.0 ;
      RECT  101700.0 2060850.0 102900.0 2059650.0 ;
      RECT  99300.0 2060850.0 100500.0 2059650.0 ;
      RECT  104100.0 2051550.0 105300.0 2050350.0 ;
      RECT  104100.0 2061450.0 105300.0 2060250.0 ;
      RECT  101700.0 2058750.0 100500.0 2057550.0 ;
      RECT  99300.0 2056800.0 98100.0 2055600.0 ;
      RECT  96900.0 2054850.0 95700.0 2053650.0 ;
      RECT  96900.0 2052150.0 98100.0 2050950.0 ;
      RECT  101700.0 2052150.0 102900.0 2050950.0 ;
      RECT  101700.0 2060850.0 102900.0 2059650.0 ;
      RECT  101700.0 2054850.0 102900.0 2053650.0 ;
      RECT  95700.0 2054850.0 96900.0 2053650.0 ;
      RECT  98100.0 2056800.0 99300.0 2055600.0 ;
      RECT  100500.0 2058750.0 101700.0 2057550.0 ;
      RECT  101700.0 2054850.0 102900.0 2053650.0 ;
      RECT  92700.0 2049450.0 108300.0 2048550.0 ;
      RECT  92700.0 2063250.0 108300.0 2062350.0 ;
      RECT  94500.0 2064750.0 95700.0 2062350.0 ;
      RECT  94500.0 2073450.0 95700.0 2077050.0 ;
      RECT  99300.0 2073450.0 100500.0 2077050.0 ;
      RECT  104100.0 2074650.0 105300.0 2076600.0 ;
      RECT  104100.0 2062800.0 105300.0 2064750.0 ;
      RECT  94500.0 2073450.0 95700.0 2074650.0 ;
      RECT  96900.0 2073450.0 98100.0 2074650.0 ;
      RECT  96900.0 2073450.0 98100.0 2074650.0 ;
      RECT  94500.0 2073450.0 95700.0 2074650.0 ;
      RECT  96900.0 2073450.0 98100.0 2074650.0 ;
      RECT  99300.0 2073450.0 100500.0 2074650.0 ;
      RECT  99300.0 2073450.0 100500.0 2074650.0 ;
      RECT  96900.0 2073450.0 98100.0 2074650.0 ;
      RECT  99300.0 2073450.0 100500.0 2074650.0 ;
      RECT  101700.0 2073450.0 102900.0 2074650.0 ;
      RECT  101700.0 2073450.0 102900.0 2074650.0 ;
      RECT  99300.0 2073450.0 100500.0 2074650.0 ;
      RECT  94500.0 2064750.0 95700.0 2065950.0 ;
      RECT  96900.0 2064750.0 98100.0 2065950.0 ;
      RECT  96900.0 2064750.0 98100.0 2065950.0 ;
      RECT  94500.0 2064750.0 95700.0 2065950.0 ;
      RECT  96900.0 2064750.0 98100.0 2065950.0 ;
      RECT  99300.0 2064750.0 100500.0 2065950.0 ;
      RECT  99300.0 2064750.0 100500.0 2065950.0 ;
      RECT  96900.0 2064750.0 98100.0 2065950.0 ;
      RECT  99300.0 2064750.0 100500.0 2065950.0 ;
      RECT  101700.0 2064750.0 102900.0 2065950.0 ;
      RECT  101700.0 2064750.0 102900.0 2065950.0 ;
      RECT  99300.0 2064750.0 100500.0 2065950.0 ;
      RECT  104100.0 2074050.0 105300.0 2075250.0 ;
      RECT  104100.0 2064150.0 105300.0 2065350.0 ;
      RECT  101700.0 2066850.0 100500.0 2068050.0 ;
      RECT  99300.0 2068800.0 98100.0 2070000.0 ;
      RECT  96900.0 2070750.0 95700.0 2071950.0 ;
      RECT  96900.0 2073450.0 98100.0 2074650.0 ;
      RECT  101700.0 2073450.0 102900.0 2074650.0 ;
      RECT  101700.0 2064750.0 102900.0 2065950.0 ;
      RECT  101700.0 2070750.0 102900.0 2071950.0 ;
      RECT  95700.0 2070750.0 96900.0 2071950.0 ;
      RECT  98100.0 2068800.0 99300.0 2070000.0 ;
      RECT  100500.0 2066850.0 101700.0 2068050.0 ;
      RECT  101700.0 2070750.0 102900.0 2071950.0 ;
      RECT  92700.0 2076150.0 108300.0 2077050.0 ;
      RECT  92700.0 2062350.0 108300.0 2063250.0 ;
      RECT  94500.0 2088450.0 95700.0 2090850.0 ;
      RECT  94500.0 2079750.0 95700.0 2076150.0 ;
      RECT  99300.0 2079750.0 100500.0 2076150.0 ;
      RECT  104100.0 2078550.0 105300.0 2076600.0 ;
      RECT  104100.0 2090400.0 105300.0 2088450.0 ;
      RECT  94500.0 2079750.0 95700.0 2078550.0 ;
      RECT  96900.0 2079750.0 98100.0 2078550.0 ;
      RECT  96900.0 2079750.0 98100.0 2078550.0 ;
      RECT  94500.0 2079750.0 95700.0 2078550.0 ;
      RECT  96900.0 2079750.0 98100.0 2078550.0 ;
      RECT  99300.0 2079750.0 100500.0 2078550.0 ;
      RECT  99300.0 2079750.0 100500.0 2078550.0 ;
      RECT  96900.0 2079750.0 98100.0 2078550.0 ;
      RECT  99300.0 2079750.0 100500.0 2078550.0 ;
      RECT  101700.0 2079750.0 102900.0 2078550.0 ;
      RECT  101700.0 2079750.0 102900.0 2078550.0 ;
      RECT  99300.0 2079750.0 100500.0 2078550.0 ;
      RECT  94500.0 2088450.0 95700.0 2087250.0 ;
      RECT  96900.0 2088450.0 98100.0 2087250.0 ;
      RECT  96900.0 2088450.0 98100.0 2087250.0 ;
      RECT  94500.0 2088450.0 95700.0 2087250.0 ;
      RECT  96900.0 2088450.0 98100.0 2087250.0 ;
      RECT  99300.0 2088450.0 100500.0 2087250.0 ;
      RECT  99300.0 2088450.0 100500.0 2087250.0 ;
      RECT  96900.0 2088450.0 98100.0 2087250.0 ;
      RECT  99300.0 2088450.0 100500.0 2087250.0 ;
      RECT  101700.0 2088450.0 102900.0 2087250.0 ;
      RECT  101700.0 2088450.0 102900.0 2087250.0 ;
      RECT  99300.0 2088450.0 100500.0 2087250.0 ;
      RECT  104100.0 2079150.0 105300.0 2077950.0 ;
      RECT  104100.0 2089050.0 105300.0 2087850.0 ;
      RECT  101700.0 2086350.0 100500.0 2085150.0 ;
      RECT  99300.0 2084400.0 98100.0 2083200.0 ;
      RECT  96900.0 2082450.0 95700.0 2081250.0 ;
      RECT  96900.0 2079750.0 98100.0 2078550.0 ;
      RECT  101700.0 2079750.0 102900.0 2078550.0 ;
      RECT  101700.0 2088450.0 102900.0 2087250.0 ;
      RECT  101700.0 2082450.0 102900.0 2081250.0 ;
      RECT  95700.0 2082450.0 96900.0 2081250.0 ;
      RECT  98100.0 2084400.0 99300.0 2083200.0 ;
      RECT  100500.0 2086350.0 101700.0 2085150.0 ;
      RECT  101700.0 2082450.0 102900.0 2081250.0 ;
      RECT  92700.0 2077050.0 108300.0 2076150.0 ;
      RECT  92700.0 2090850.0 108300.0 2089950.0 ;
      RECT  94500.0 2092350.0 95700.0 2089950.0 ;
      RECT  94500.0 2101050.0 95700.0 2104650.0 ;
      RECT  99300.0 2101050.0 100500.0 2104650.0 ;
      RECT  104100.0 2102250.0 105300.0 2104200.0 ;
      RECT  104100.0 2090400.0 105300.0 2092350.0 ;
      RECT  94500.0 2101050.0 95700.0 2102250.0 ;
      RECT  96900.0 2101050.0 98100.0 2102250.0 ;
      RECT  96900.0 2101050.0 98100.0 2102250.0 ;
      RECT  94500.0 2101050.0 95700.0 2102250.0 ;
      RECT  96900.0 2101050.0 98100.0 2102250.0 ;
      RECT  99300.0 2101050.0 100500.0 2102250.0 ;
      RECT  99300.0 2101050.0 100500.0 2102250.0 ;
      RECT  96900.0 2101050.0 98100.0 2102250.0 ;
      RECT  99300.0 2101050.0 100500.0 2102250.0 ;
      RECT  101700.0 2101050.0 102900.0 2102250.0 ;
      RECT  101700.0 2101050.0 102900.0 2102250.0 ;
      RECT  99300.0 2101050.0 100500.0 2102250.0 ;
      RECT  94500.0 2092350.0 95700.0 2093550.0 ;
      RECT  96900.0 2092350.0 98100.0 2093550.0 ;
      RECT  96900.0 2092350.0 98100.0 2093550.0 ;
      RECT  94500.0 2092350.0 95700.0 2093550.0 ;
      RECT  96900.0 2092350.0 98100.0 2093550.0 ;
      RECT  99300.0 2092350.0 100500.0 2093550.0 ;
      RECT  99300.0 2092350.0 100500.0 2093550.0 ;
      RECT  96900.0 2092350.0 98100.0 2093550.0 ;
      RECT  99300.0 2092350.0 100500.0 2093550.0 ;
      RECT  101700.0 2092350.0 102900.0 2093550.0 ;
      RECT  101700.0 2092350.0 102900.0 2093550.0 ;
      RECT  99300.0 2092350.0 100500.0 2093550.0 ;
      RECT  104100.0 2101650.0 105300.0 2102850.0 ;
      RECT  104100.0 2091750.0 105300.0 2092950.0 ;
      RECT  101700.0 2094450.0 100500.0 2095650.0 ;
      RECT  99300.0 2096400.0 98100.0 2097600.0 ;
      RECT  96900.0 2098350.0 95700.0 2099550.0 ;
      RECT  96900.0 2101050.0 98100.0 2102250.0 ;
      RECT  101700.0 2101050.0 102900.0 2102250.0 ;
      RECT  101700.0 2092350.0 102900.0 2093550.0 ;
      RECT  101700.0 2098350.0 102900.0 2099550.0 ;
      RECT  95700.0 2098350.0 96900.0 2099550.0 ;
      RECT  98100.0 2096400.0 99300.0 2097600.0 ;
      RECT  100500.0 2094450.0 101700.0 2095650.0 ;
      RECT  101700.0 2098350.0 102900.0 2099550.0 ;
      RECT  92700.0 2103750.0 108300.0 2104650.0 ;
      RECT  92700.0 2089950.0 108300.0 2090850.0 ;
      RECT  94500.0 2116050.0 95700.0 2118450.0 ;
      RECT  94500.0 2107350.0 95700.0 2103750.0 ;
      RECT  99300.0 2107350.0 100500.0 2103750.0 ;
      RECT  104100.0 2106150.0 105300.0 2104200.0 ;
      RECT  104100.0 2118000.0 105300.0 2116050.0 ;
      RECT  94500.0 2107350.0 95700.0 2106150.0 ;
      RECT  96900.0 2107350.0 98100.0 2106150.0 ;
      RECT  96900.0 2107350.0 98100.0 2106150.0 ;
      RECT  94500.0 2107350.0 95700.0 2106150.0 ;
      RECT  96900.0 2107350.0 98100.0 2106150.0 ;
      RECT  99300.0 2107350.0 100500.0 2106150.0 ;
      RECT  99300.0 2107350.0 100500.0 2106150.0 ;
      RECT  96900.0 2107350.0 98100.0 2106150.0 ;
      RECT  99300.0 2107350.0 100500.0 2106150.0 ;
      RECT  101700.0 2107350.0 102900.0 2106150.0 ;
      RECT  101700.0 2107350.0 102900.0 2106150.0 ;
      RECT  99300.0 2107350.0 100500.0 2106150.0 ;
      RECT  94500.0 2116050.0 95700.0 2114850.0 ;
      RECT  96900.0 2116050.0 98100.0 2114850.0 ;
      RECT  96900.0 2116050.0 98100.0 2114850.0 ;
      RECT  94500.0 2116050.0 95700.0 2114850.0 ;
      RECT  96900.0 2116050.0 98100.0 2114850.0 ;
      RECT  99300.0 2116050.0 100500.0 2114850.0 ;
      RECT  99300.0 2116050.0 100500.0 2114850.0 ;
      RECT  96900.0 2116050.0 98100.0 2114850.0 ;
      RECT  99300.0 2116050.0 100500.0 2114850.0 ;
      RECT  101700.0 2116050.0 102900.0 2114850.0 ;
      RECT  101700.0 2116050.0 102900.0 2114850.0 ;
      RECT  99300.0 2116050.0 100500.0 2114850.0 ;
      RECT  104100.0 2106750.0 105300.0 2105550.0 ;
      RECT  104100.0 2116650.0 105300.0 2115450.0 ;
      RECT  101700.0 2113950.0 100500.0 2112750.0 ;
      RECT  99300.0 2112000.0 98100.0 2110800.0 ;
      RECT  96900.0 2110050.0 95700.0 2108850.0 ;
      RECT  96900.0 2107350.0 98100.0 2106150.0 ;
      RECT  101700.0 2107350.0 102900.0 2106150.0 ;
      RECT  101700.0 2116050.0 102900.0 2114850.0 ;
      RECT  101700.0 2110050.0 102900.0 2108850.0 ;
      RECT  95700.0 2110050.0 96900.0 2108850.0 ;
      RECT  98100.0 2112000.0 99300.0 2110800.0 ;
      RECT  100500.0 2113950.0 101700.0 2112750.0 ;
      RECT  101700.0 2110050.0 102900.0 2108850.0 ;
      RECT  92700.0 2104650.0 108300.0 2103750.0 ;
      RECT  92700.0 2118450.0 108300.0 2117550.0 ;
      RECT  94500.0 2119950.0 95700.0 2117550.0 ;
      RECT  94500.0 2128650.0 95700.0 2132250.0 ;
      RECT  99300.0 2128650.0 100500.0 2132250.0 ;
      RECT  104100.0 2129850.0 105300.0 2131800.0 ;
      RECT  104100.0 2118000.0 105300.0 2119950.0 ;
      RECT  94500.0 2128650.0 95700.0 2129850.0 ;
      RECT  96900.0 2128650.0 98100.0 2129850.0 ;
      RECT  96900.0 2128650.0 98100.0 2129850.0 ;
      RECT  94500.0 2128650.0 95700.0 2129850.0 ;
      RECT  96900.0 2128650.0 98100.0 2129850.0 ;
      RECT  99300.0 2128650.0 100500.0 2129850.0 ;
      RECT  99300.0 2128650.0 100500.0 2129850.0 ;
      RECT  96900.0 2128650.0 98100.0 2129850.0 ;
      RECT  99300.0 2128650.0 100500.0 2129850.0 ;
      RECT  101700.0 2128650.0 102900.0 2129850.0 ;
      RECT  101700.0 2128650.0 102900.0 2129850.0 ;
      RECT  99300.0 2128650.0 100500.0 2129850.0 ;
      RECT  94500.0 2119950.0 95700.0 2121150.0 ;
      RECT  96900.0 2119950.0 98100.0 2121150.0 ;
      RECT  96900.0 2119950.0 98100.0 2121150.0 ;
      RECT  94500.0 2119950.0 95700.0 2121150.0 ;
      RECT  96900.0 2119950.0 98100.0 2121150.0 ;
      RECT  99300.0 2119950.0 100500.0 2121150.0 ;
      RECT  99300.0 2119950.0 100500.0 2121150.0 ;
      RECT  96900.0 2119950.0 98100.0 2121150.0 ;
      RECT  99300.0 2119950.0 100500.0 2121150.0 ;
      RECT  101700.0 2119950.0 102900.0 2121150.0 ;
      RECT  101700.0 2119950.0 102900.0 2121150.0 ;
      RECT  99300.0 2119950.0 100500.0 2121150.0 ;
      RECT  104100.0 2129250.0 105300.0 2130450.0 ;
      RECT  104100.0 2119350.0 105300.0 2120550.0 ;
      RECT  101700.0 2122050.0 100500.0 2123250.0 ;
      RECT  99300.0 2124000.0 98100.0 2125200.0 ;
      RECT  96900.0 2125950.0 95700.0 2127150.0 ;
      RECT  96900.0 2128650.0 98100.0 2129850.0 ;
      RECT  101700.0 2128650.0 102900.0 2129850.0 ;
      RECT  101700.0 2119950.0 102900.0 2121150.0 ;
      RECT  101700.0 2125950.0 102900.0 2127150.0 ;
      RECT  95700.0 2125950.0 96900.0 2127150.0 ;
      RECT  98100.0 2124000.0 99300.0 2125200.0 ;
      RECT  100500.0 2122050.0 101700.0 2123250.0 ;
      RECT  101700.0 2125950.0 102900.0 2127150.0 ;
      RECT  92700.0 2131350.0 108300.0 2132250.0 ;
      RECT  92700.0 2117550.0 108300.0 2118450.0 ;
      RECT  94500.0 2143650.0 95700.0 2146050.0 ;
      RECT  94500.0 2134950.0 95700.0 2131350.0 ;
      RECT  99300.0 2134950.0 100500.0 2131350.0 ;
      RECT  104100.0 2133750.0 105300.0 2131800.0 ;
      RECT  104100.0 2145600.0 105300.0 2143650.0 ;
      RECT  94500.0 2134950.0 95700.0 2133750.0 ;
      RECT  96900.0 2134950.0 98100.0 2133750.0 ;
      RECT  96900.0 2134950.0 98100.0 2133750.0 ;
      RECT  94500.0 2134950.0 95700.0 2133750.0 ;
      RECT  96900.0 2134950.0 98100.0 2133750.0 ;
      RECT  99300.0 2134950.0 100500.0 2133750.0 ;
      RECT  99300.0 2134950.0 100500.0 2133750.0 ;
      RECT  96900.0 2134950.0 98100.0 2133750.0 ;
      RECT  99300.0 2134950.0 100500.0 2133750.0 ;
      RECT  101700.0 2134950.0 102900.0 2133750.0 ;
      RECT  101700.0 2134950.0 102900.0 2133750.0 ;
      RECT  99300.0 2134950.0 100500.0 2133750.0 ;
      RECT  94500.0 2143650.0 95700.0 2142450.0 ;
      RECT  96900.0 2143650.0 98100.0 2142450.0 ;
      RECT  96900.0 2143650.0 98100.0 2142450.0 ;
      RECT  94500.0 2143650.0 95700.0 2142450.0 ;
      RECT  96900.0 2143650.0 98100.0 2142450.0 ;
      RECT  99300.0 2143650.0 100500.0 2142450.0 ;
      RECT  99300.0 2143650.0 100500.0 2142450.0 ;
      RECT  96900.0 2143650.0 98100.0 2142450.0 ;
      RECT  99300.0 2143650.0 100500.0 2142450.0 ;
      RECT  101700.0 2143650.0 102900.0 2142450.0 ;
      RECT  101700.0 2143650.0 102900.0 2142450.0 ;
      RECT  99300.0 2143650.0 100500.0 2142450.0 ;
      RECT  104100.0 2134350.0 105300.0 2133150.0 ;
      RECT  104100.0 2144250.0 105300.0 2143050.0 ;
      RECT  101700.0 2141550.0 100500.0 2140350.0 ;
      RECT  99300.0 2139600.0 98100.0 2138400.0 ;
      RECT  96900.0 2137650.0 95700.0 2136450.0 ;
      RECT  96900.0 2134950.0 98100.0 2133750.0 ;
      RECT  101700.0 2134950.0 102900.0 2133750.0 ;
      RECT  101700.0 2143650.0 102900.0 2142450.0 ;
      RECT  101700.0 2137650.0 102900.0 2136450.0 ;
      RECT  95700.0 2137650.0 96900.0 2136450.0 ;
      RECT  98100.0 2139600.0 99300.0 2138400.0 ;
      RECT  100500.0 2141550.0 101700.0 2140350.0 ;
      RECT  101700.0 2137650.0 102900.0 2136450.0 ;
      RECT  92700.0 2132250.0 108300.0 2131350.0 ;
      RECT  92700.0 2146050.0 108300.0 2145150.0 ;
      RECT  114900.0 391050.0 116100.0 393000.0 ;
      RECT  114900.0 379200.0 116100.0 381150.0 ;
      RECT  110100.0 380550.0 111300.0 378750.0 ;
      RECT  110100.0 389850.0 111300.0 393450.0 ;
      RECT  112800.0 380550.0 113700.0 389850.0 ;
      RECT  110100.0 389850.0 111300.0 391050.0 ;
      RECT  112500.0 389850.0 113700.0 391050.0 ;
      RECT  112500.0 389850.0 113700.0 391050.0 ;
      RECT  110100.0 389850.0 111300.0 391050.0 ;
      RECT  110100.0 380550.0 111300.0 381750.0 ;
      RECT  112500.0 380550.0 113700.0 381750.0 ;
      RECT  112500.0 380550.0 113700.0 381750.0 ;
      RECT  110100.0 380550.0 111300.0 381750.0 ;
      RECT  114900.0 390450.0 116100.0 391650.0 ;
      RECT  114900.0 380550.0 116100.0 381750.0 ;
      RECT  110700.0 385200.0 111900.0 386400.0 ;
      RECT  110700.0 385200.0 111900.0 386400.0 ;
      RECT  113250.0 385350.0 114150.0 386250.0 ;
      RECT  108300.0 392550.0 117900.0 393450.0 ;
      RECT  108300.0 378750.0 117900.0 379650.0 ;
      RECT  114900.0 394950.0 116100.0 393000.0 ;
      RECT  114900.0 406800.0 116100.0 404850.0 ;
      RECT  110100.0 405450.0 111300.0 407250.0 ;
      RECT  110100.0 396150.0 111300.0 392550.0 ;
      RECT  112800.0 405450.0 113700.0 396150.0 ;
      RECT  110100.0 396150.0 111300.0 394950.0 ;
      RECT  112500.0 396150.0 113700.0 394950.0 ;
      RECT  112500.0 396150.0 113700.0 394950.0 ;
      RECT  110100.0 396150.0 111300.0 394950.0 ;
      RECT  110100.0 405450.0 111300.0 404250.0 ;
      RECT  112500.0 405450.0 113700.0 404250.0 ;
      RECT  112500.0 405450.0 113700.0 404250.0 ;
      RECT  110100.0 405450.0 111300.0 404250.0 ;
      RECT  114900.0 395550.0 116100.0 394350.0 ;
      RECT  114900.0 405450.0 116100.0 404250.0 ;
      RECT  110700.0 400800.0 111900.0 399600.0 ;
      RECT  110700.0 400800.0 111900.0 399600.0 ;
      RECT  113250.0 400650.0 114150.0 399750.0 ;
      RECT  108300.0 393450.0 117900.0 392550.0 ;
      RECT  108300.0 407250.0 117900.0 406350.0 ;
      RECT  114900.0 418650.0 116100.0 420600.0 ;
      RECT  114900.0 406800.0 116100.0 408750.0 ;
      RECT  110100.0 408150.0 111300.0 406350.0 ;
      RECT  110100.0 417450.0 111300.0 421050.0 ;
      RECT  112800.0 408150.0 113700.0 417450.0 ;
      RECT  110100.0 417450.0 111300.0 418650.0 ;
      RECT  112500.0 417450.0 113700.0 418650.0 ;
      RECT  112500.0 417450.0 113700.0 418650.0 ;
      RECT  110100.0 417450.0 111300.0 418650.0 ;
      RECT  110100.0 408150.0 111300.0 409350.0 ;
      RECT  112500.0 408150.0 113700.0 409350.0 ;
      RECT  112500.0 408150.0 113700.0 409350.0 ;
      RECT  110100.0 408150.0 111300.0 409350.0 ;
      RECT  114900.0 418050.0 116100.0 419250.0 ;
      RECT  114900.0 408150.0 116100.0 409350.0 ;
      RECT  110700.0 412800.0 111900.0 414000.0 ;
      RECT  110700.0 412800.0 111900.0 414000.0 ;
      RECT  113250.0 412950.0 114150.0 413850.0 ;
      RECT  108300.0 420150.0 117900.0 421050.0 ;
      RECT  108300.0 406350.0 117900.0 407250.0 ;
      RECT  114900.0 422550.0 116100.0 420600.0 ;
      RECT  114900.0 434400.0 116100.0 432450.0 ;
      RECT  110100.0 433050.0 111300.0 434850.0 ;
      RECT  110100.0 423750.0 111300.0 420150.0 ;
      RECT  112800.0 433050.0 113700.0 423750.0 ;
      RECT  110100.0 423750.0 111300.0 422550.0 ;
      RECT  112500.0 423750.0 113700.0 422550.0 ;
      RECT  112500.0 423750.0 113700.0 422550.0 ;
      RECT  110100.0 423750.0 111300.0 422550.0 ;
      RECT  110100.0 433050.0 111300.0 431850.0 ;
      RECT  112500.0 433050.0 113700.0 431850.0 ;
      RECT  112500.0 433050.0 113700.0 431850.0 ;
      RECT  110100.0 433050.0 111300.0 431850.0 ;
      RECT  114900.0 423150.0 116100.0 421950.0 ;
      RECT  114900.0 433050.0 116100.0 431850.0 ;
      RECT  110700.0 428400.0 111900.0 427200.0 ;
      RECT  110700.0 428400.0 111900.0 427200.0 ;
      RECT  113250.0 428250.0 114150.0 427350.0 ;
      RECT  108300.0 421050.0 117900.0 420150.0 ;
      RECT  108300.0 434850.0 117900.0 433950.0 ;
      RECT  114900.0 446250.0 116100.0 448200.0 ;
      RECT  114900.0 434400.0 116100.0 436350.0 ;
      RECT  110100.0 435750.0 111300.0 433950.0 ;
      RECT  110100.0 445050.0 111300.0 448650.0 ;
      RECT  112800.0 435750.0 113700.0 445050.0 ;
      RECT  110100.0 445050.0 111300.0 446250.0 ;
      RECT  112500.0 445050.0 113700.0 446250.0 ;
      RECT  112500.0 445050.0 113700.0 446250.0 ;
      RECT  110100.0 445050.0 111300.0 446250.0 ;
      RECT  110100.0 435750.0 111300.0 436950.0 ;
      RECT  112500.0 435750.0 113700.0 436950.0 ;
      RECT  112500.0 435750.0 113700.0 436950.0 ;
      RECT  110100.0 435750.0 111300.0 436950.0 ;
      RECT  114900.0 445650.0 116100.0 446850.0 ;
      RECT  114900.0 435750.0 116100.0 436950.0 ;
      RECT  110700.0 440400.0 111900.0 441600.0 ;
      RECT  110700.0 440400.0 111900.0 441600.0 ;
      RECT  113250.0 440550.0 114150.0 441450.0 ;
      RECT  108300.0 447750.0 117900.0 448650.0 ;
      RECT  108300.0 433950.0 117900.0 434850.0 ;
      RECT  114900.0 450150.0 116100.0 448200.0 ;
      RECT  114900.0 462000.0 116100.0 460050.0 ;
      RECT  110100.0 460650.0 111300.0 462450.0 ;
      RECT  110100.0 451350.0 111300.0 447750.0 ;
      RECT  112800.0 460650.0 113700.0 451350.0 ;
      RECT  110100.0 451350.0 111300.0 450150.0 ;
      RECT  112500.0 451350.0 113700.0 450150.0 ;
      RECT  112500.0 451350.0 113700.0 450150.0 ;
      RECT  110100.0 451350.0 111300.0 450150.0 ;
      RECT  110100.0 460650.0 111300.0 459450.0 ;
      RECT  112500.0 460650.0 113700.0 459450.0 ;
      RECT  112500.0 460650.0 113700.0 459450.0 ;
      RECT  110100.0 460650.0 111300.0 459450.0 ;
      RECT  114900.0 450750.0 116100.0 449550.0 ;
      RECT  114900.0 460650.0 116100.0 459450.0 ;
      RECT  110700.0 456000.0 111900.0 454800.0 ;
      RECT  110700.0 456000.0 111900.0 454800.0 ;
      RECT  113250.0 455850.0 114150.0 454950.0 ;
      RECT  108300.0 448650.0 117900.0 447750.0 ;
      RECT  108300.0 462450.0 117900.0 461550.0 ;
      RECT  114900.0 473850.0 116100.0 475800.0 ;
      RECT  114900.0 462000.0 116100.0 463950.0 ;
      RECT  110100.0 463350.0 111300.0 461550.0 ;
      RECT  110100.0 472650.0 111300.0 476250.0 ;
      RECT  112800.0 463350.0 113700.0 472650.0 ;
      RECT  110100.0 472650.0 111300.0 473850.0 ;
      RECT  112500.0 472650.0 113700.0 473850.0 ;
      RECT  112500.0 472650.0 113700.0 473850.0 ;
      RECT  110100.0 472650.0 111300.0 473850.0 ;
      RECT  110100.0 463350.0 111300.0 464550.0 ;
      RECT  112500.0 463350.0 113700.0 464550.0 ;
      RECT  112500.0 463350.0 113700.0 464550.0 ;
      RECT  110100.0 463350.0 111300.0 464550.0 ;
      RECT  114900.0 473250.0 116100.0 474450.0 ;
      RECT  114900.0 463350.0 116100.0 464550.0 ;
      RECT  110700.0 468000.0 111900.0 469200.0 ;
      RECT  110700.0 468000.0 111900.0 469200.0 ;
      RECT  113250.0 468150.0 114150.0 469050.0 ;
      RECT  108300.0 475350.0 117900.0 476250.0 ;
      RECT  108300.0 461550.0 117900.0 462450.0 ;
      RECT  114900.0 477750.0 116100.0 475800.0 ;
      RECT  114900.0 489600.0 116100.0 487650.0 ;
      RECT  110100.0 488250.0 111300.0 490050.0 ;
      RECT  110100.0 478950.0 111300.0 475350.0 ;
      RECT  112800.0 488250.0 113700.0 478950.0 ;
      RECT  110100.0 478950.0 111300.0 477750.0 ;
      RECT  112500.0 478950.0 113700.0 477750.0 ;
      RECT  112500.0 478950.0 113700.0 477750.0 ;
      RECT  110100.0 478950.0 111300.0 477750.0 ;
      RECT  110100.0 488250.0 111300.0 487050.0 ;
      RECT  112500.0 488250.0 113700.0 487050.0 ;
      RECT  112500.0 488250.0 113700.0 487050.0 ;
      RECT  110100.0 488250.0 111300.0 487050.0 ;
      RECT  114900.0 478350.0 116100.0 477150.0 ;
      RECT  114900.0 488250.0 116100.0 487050.0 ;
      RECT  110700.0 483600.0 111900.0 482400.0 ;
      RECT  110700.0 483600.0 111900.0 482400.0 ;
      RECT  113250.0 483450.0 114150.0 482550.0 ;
      RECT  108300.0 476250.0 117900.0 475350.0 ;
      RECT  108300.0 490050.0 117900.0 489150.0 ;
      RECT  114900.0 501450.0 116100.0 503400.0 ;
      RECT  114900.0 489600.0 116100.0 491550.0 ;
      RECT  110100.0 490950.0 111300.0 489150.0 ;
      RECT  110100.0 500250.0 111300.0 503850.0 ;
      RECT  112800.0 490950.0 113700.0 500250.0 ;
      RECT  110100.0 500250.0 111300.0 501450.0 ;
      RECT  112500.0 500250.0 113700.0 501450.0 ;
      RECT  112500.0 500250.0 113700.0 501450.0 ;
      RECT  110100.0 500250.0 111300.0 501450.0 ;
      RECT  110100.0 490950.0 111300.0 492150.0 ;
      RECT  112500.0 490950.0 113700.0 492150.0 ;
      RECT  112500.0 490950.0 113700.0 492150.0 ;
      RECT  110100.0 490950.0 111300.0 492150.0 ;
      RECT  114900.0 500850.0 116100.0 502050.0 ;
      RECT  114900.0 490950.0 116100.0 492150.0 ;
      RECT  110700.0 495600.0 111900.0 496800.0 ;
      RECT  110700.0 495600.0 111900.0 496800.0 ;
      RECT  113250.0 495750.0 114150.0 496650.0 ;
      RECT  108300.0 502950.0 117900.0 503850.0 ;
      RECT  108300.0 489150.0 117900.0 490050.0 ;
      RECT  114900.0 505350.0 116100.0 503400.0 ;
      RECT  114900.0 517200.0 116100.0 515250.0 ;
      RECT  110100.0 515850.0 111300.0 517650.0 ;
      RECT  110100.0 506550.0 111300.0 502950.0 ;
      RECT  112800.0 515850.0 113700.0 506550.0 ;
      RECT  110100.0 506550.0 111300.0 505350.0 ;
      RECT  112500.0 506550.0 113700.0 505350.0 ;
      RECT  112500.0 506550.0 113700.0 505350.0 ;
      RECT  110100.0 506550.0 111300.0 505350.0 ;
      RECT  110100.0 515850.0 111300.0 514650.0 ;
      RECT  112500.0 515850.0 113700.0 514650.0 ;
      RECT  112500.0 515850.0 113700.0 514650.0 ;
      RECT  110100.0 515850.0 111300.0 514650.0 ;
      RECT  114900.0 505950.0 116100.0 504750.0 ;
      RECT  114900.0 515850.0 116100.0 514650.0 ;
      RECT  110700.0 511200.0 111900.0 510000.0 ;
      RECT  110700.0 511200.0 111900.0 510000.0 ;
      RECT  113250.0 511050.0 114150.0 510150.0 ;
      RECT  108300.0 503850.0 117900.0 502950.0 ;
      RECT  108300.0 517650.0 117900.0 516750.0 ;
      RECT  114900.0 529050.0 116100.0 531000.0 ;
      RECT  114900.0 517200.0 116100.0 519150.0 ;
      RECT  110100.0 518550.0 111300.0 516750.0 ;
      RECT  110100.0 527850.0 111300.0 531450.0 ;
      RECT  112800.0 518550.0 113700.0 527850.0 ;
      RECT  110100.0 527850.0 111300.0 529050.0 ;
      RECT  112500.0 527850.0 113700.0 529050.0 ;
      RECT  112500.0 527850.0 113700.0 529050.0 ;
      RECT  110100.0 527850.0 111300.0 529050.0 ;
      RECT  110100.0 518550.0 111300.0 519750.0 ;
      RECT  112500.0 518550.0 113700.0 519750.0 ;
      RECT  112500.0 518550.0 113700.0 519750.0 ;
      RECT  110100.0 518550.0 111300.0 519750.0 ;
      RECT  114900.0 528450.0 116100.0 529650.0 ;
      RECT  114900.0 518550.0 116100.0 519750.0 ;
      RECT  110700.0 523200.0 111900.0 524400.0 ;
      RECT  110700.0 523200.0 111900.0 524400.0 ;
      RECT  113250.0 523350.0 114150.0 524250.0 ;
      RECT  108300.0 530550.0 117900.0 531450.0 ;
      RECT  108300.0 516750.0 117900.0 517650.0 ;
      RECT  114900.0 532950.0 116100.0 531000.0 ;
      RECT  114900.0 544800.0 116100.0 542850.0 ;
      RECT  110100.0 543450.0 111300.0 545250.0 ;
      RECT  110100.0 534150.0 111300.0 530550.0 ;
      RECT  112800.0 543450.0 113700.0 534150.0 ;
      RECT  110100.0 534150.0 111300.0 532950.0 ;
      RECT  112500.0 534150.0 113700.0 532950.0 ;
      RECT  112500.0 534150.0 113700.0 532950.0 ;
      RECT  110100.0 534150.0 111300.0 532950.0 ;
      RECT  110100.0 543450.0 111300.0 542250.0 ;
      RECT  112500.0 543450.0 113700.0 542250.0 ;
      RECT  112500.0 543450.0 113700.0 542250.0 ;
      RECT  110100.0 543450.0 111300.0 542250.0 ;
      RECT  114900.0 533550.0 116100.0 532350.0 ;
      RECT  114900.0 543450.0 116100.0 542250.0 ;
      RECT  110700.0 538800.0 111900.0 537600.0 ;
      RECT  110700.0 538800.0 111900.0 537600.0 ;
      RECT  113250.0 538650.0 114150.0 537750.0 ;
      RECT  108300.0 531450.0 117900.0 530550.0 ;
      RECT  108300.0 545250.0 117900.0 544350.0 ;
      RECT  114900.0 556650.0 116100.0 558600.0 ;
      RECT  114900.0 544800.0 116100.0 546750.0 ;
      RECT  110100.0 546150.0 111300.0 544350.0 ;
      RECT  110100.0 555450.0 111300.0 559050.0 ;
      RECT  112800.0 546150.0 113700.0 555450.0 ;
      RECT  110100.0 555450.0 111300.0 556650.0 ;
      RECT  112500.0 555450.0 113700.0 556650.0 ;
      RECT  112500.0 555450.0 113700.0 556650.0 ;
      RECT  110100.0 555450.0 111300.0 556650.0 ;
      RECT  110100.0 546150.0 111300.0 547350.0 ;
      RECT  112500.0 546150.0 113700.0 547350.0 ;
      RECT  112500.0 546150.0 113700.0 547350.0 ;
      RECT  110100.0 546150.0 111300.0 547350.0 ;
      RECT  114900.0 556050.0 116100.0 557250.0 ;
      RECT  114900.0 546150.0 116100.0 547350.0 ;
      RECT  110700.0 550800.0 111900.0 552000.0 ;
      RECT  110700.0 550800.0 111900.0 552000.0 ;
      RECT  113250.0 550950.0 114150.0 551850.0 ;
      RECT  108300.0 558150.0 117900.0 559050.0 ;
      RECT  108300.0 544350.0 117900.0 545250.0 ;
      RECT  114900.0 560550.0 116100.0 558600.0 ;
      RECT  114900.0 572400.0 116100.0 570450.0 ;
      RECT  110100.0 571050.0 111300.0 572850.0 ;
      RECT  110100.0 561750.0 111300.0 558150.0 ;
      RECT  112800.0 571050.0 113700.0 561750.0 ;
      RECT  110100.0 561750.0 111300.0 560550.0 ;
      RECT  112500.0 561750.0 113700.0 560550.0 ;
      RECT  112500.0 561750.0 113700.0 560550.0 ;
      RECT  110100.0 561750.0 111300.0 560550.0 ;
      RECT  110100.0 571050.0 111300.0 569850.0 ;
      RECT  112500.0 571050.0 113700.0 569850.0 ;
      RECT  112500.0 571050.0 113700.0 569850.0 ;
      RECT  110100.0 571050.0 111300.0 569850.0 ;
      RECT  114900.0 561150.0 116100.0 559950.0 ;
      RECT  114900.0 571050.0 116100.0 569850.0 ;
      RECT  110700.0 566400.0 111900.0 565200.0 ;
      RECT  110700.0 566400.0 111900.0 565200.0 ;
      RECT  113250.0 566250.0 114150.0 565350.0 ;
      RECT  108300.0 559050.0 117900.0 558150.0 ;
      RECT  108300.0 572850.0 117900.0 571950.0 ;
      RECT  114900.0 584250.0 116100.0 586200.0 ;
      RECT  114900.0 572400.0 116100.0 574350.0 ;
      RECT  110100.0 573750.0 111300.0 571950.0 ;
      RECT  110100.0 583050.0 111300.0 586650.0 ;
      RECT  112800.0 573750.0 113700.0 583050.0 ;
      RECT  110100.0 583050.0 111300.0 584250.0 ;
      RECT  112500.0 583050.0 113700.0 584250.0 ;
      RECT  112500.0 583050.0 113700.0 584250.0 ;
      RECT  110100.0 583050.0 111300.0 584250.0 ;
      RECT  110100.0 573750.0 111300.0 574950.0 ;
      RECT  112500.0 573750.0 113700.0 574950.0 ;
      RECT  112500.0 573750.0 113700.0 574950.0 ;
      RECT  110100.0 573750.0 111300.0 574950.0 ;
      RECT  114900.0 583650.0 116100.0 584850.0 ;
      RECT  114900.0 573750.0 116100.0 574950.0 ;
      RECT  110700.0 578400.0 111900.0 579600.0 ;
      RECT  110700.0 578400.0 111900.0 579600.0 ;
      RECT  113250.0 578550.0 114150.0 579450.0 ;
      RECT  108300.0 585750.0 117900.0 586650.0 ;
      RECT  108300.0 571950.0 117900.0 572850.0 ;
      RECT  114900.0 588150.0 116100.0 586200.0 ;
      RECT  114900.0 600000.0 116100.0 598050.0 ;
      RECT  110100.0 598650.0 111300.0 600450.0 ;
      RECT  110100.0 589350.0 111300.0 585750.0 ;
      RECT  112800.0 598650.0 113700.0 589350.0 ;
      RECT  110100.0 589350.0 111300.0 588150.0 ;
      RECT  112500.0 589350.0 113700.0 588150.0 ;
      RECT  112500.0 589350.0 113700.0 588150.0 ;
      RECT  110100.0 589350.0 111300.0 588150.0 ;
      RECT  110100.0 598650.0 111300.0 597450.0 ;
      RECT  112500.0 598650.0 113700.0 597450.0 ;
      RECT  112500.0 598650.0 113700.0 597450.0 ;
      RECT  110100.0 598650.0 111300.0 597450.0 ;
      RECT  114900.0 588750.0 116100.0 587550.0 ;
      RECT  114900.0 598650.0 116100.0 597450.0 ;
      RECT  110700.0 594000.0 111900.0 592800.0 ;
      RECT  110700.0 594000.0 111900.0 592800.0 ;
      RECT  113250.0 593850.0 114150.0 592950.0 ;
      RECT  108300.0 586650.0 117900.0 585750.0 ;
      RECT  108300.0 600450.0 117900.0 599550.0 ;
      RECT  114900.0 611850.0 116100.0 613800.0 ;
      RECT  114900.0 600000.0 116100.0 601950.0 ;
      RECT  110100.0 601350.0 111300.0 599550.0 ;
      RECT  110100.0 610650.0 111300.0 614250.0 ;
      RECT  112800.0 601350.0 113700.0 610650.0 ;
      RECT  110100.0 610650.0 111300.0 611850.0 ;
      RECT  112500.0 610650.0 113700.0 611850.0 ;
      RECT  112500.0 610650.0 113700.0 611850.0 ;
      RECT  110100.0 610650.0 111300.0 611850.0 ;
      RECT  110100.0 601350.0 111300.0 602550.0 ;
      RECT  112500.0 601350.0 113700.0 602550.0 ;
      RECT  112500.0 601350.0 113700.0 602550.0 ;
      RECT  110100.0 601350.0 111300.0 602550.0 ;
      RECT  114900.0 611250.0 116100.0 612450.0 ;
      RECT  114900.0 601350.0 116100.0 602550.0 ;
      RECT  110700.0 606000.0 111900.0 607200.0 ;
      RECT  110700.0 606000.0 111900.0 607200.0 ;
      RECT  113250.0 606150.0 114150.0 607050.0 ;
      RECT  108300.0 613350.0 117900.0 614250.0 ;
      RECT  108300.0 599550.0 117900.0 600450.0 ;
      RECT  114900.0 615750.0 116100.0 613800.0 ;
      RECT  114900.0 627600.0 116100.0 625650.0 ;
      RECT  110100.0 626250.0 111300.0 628050.0 ;
      RECT  110100.0 616950.0 111300.0 613350.0 ;
      RECT  112800.0 626250.0 113700.0 616950.0 ;
      RECT  110100.0 616950.0 111300.0 615750.0 ;
      RECT  112500.0 616950.0 113700.0 615750.0 ;
      RECT  112500.0 616950.0 113700.0 615750.0 ;
      RECT  110100.0 616950.0 111300.0 615750.0 ;
      RECT  110100.0 626250.0 111300.0 625050.0 ;
      RECT  112500.0 626250.0 113700.0 625050.0 ;
      RECT  112500.0 626250.0 113700.0 625050.0 ;
      RECT  110100.0 626250.0 111300.0 625050.0 ;
      RECT  114900.0 616350.0 116100.0 615150.0 ;
      RECT  114900.0 626250.0 116100.0 625050.0 ;
      RECT  110700.0 621600.0 111900.0 620400.0 ;
      RECT  110700.0 621600.0 111900.0 620400.0 ;
      RECT  113250.0 621450.0 114150.0 620550.0 ;
      RECT  108300.0 614250.0 117900.0 613350.0 ;
      RECT  108300.0 628050.0 117900.0 627150.0 ;
      RECT  114900.0 639450.0 116100.0 641400.0 ;
      RECT  114900.0 627600.0 116100.0 629550.0 ;
      RECT  110100.0 628950.0 111300.0 627150.0 ;
      RECT  110100.0 638250.0 111300.0 641850.0 ;
      RECT  112800.0 628950.0 113700.0 638250.0 ;
      RECT  110100.0 638250.0 111300.0 639450.0 ;
      RECT  112500.0 638250.0 113700.0 639450.0 ;
      RECT  112500.0 638250.0 113700.0 639450.0 ;
      RECT  110100.0 638250.0 111300.0 639450.0 ;
      RECT  110100.0 628950.0 111300.0 630150.0 ;
      RECT  112500.0 628950.0 113700.0 630150.0 ;
      RECT  112500.0 628950.0 113700.0 630150.0 ;
      RECT  110100.0 628950.0 111300.0 630150.0 ;
      RECT  114900.0 638850.0 116100.0 640050.0 ;
      RECT  114900.0 628950.0 116100.0 630150.0 ;
      RECT  110700.0 633600.0 111900.0 634800.0 ;
      RECT  110700.0 633600.0 111900.0 634800.0 ;
      RECT  113250.0 633750.0 114150.0 634650.0 ;
      RECT  108300.0 640950.0 117900.0 641850.0 ;
      RECT  108300.0 627150.0 117900.0 628050.0 ;
      RECT  114900.0 643350.0 116100.0 641400.0 ;
      RECT  114900.0 655200.0 116100.0 653250.0 ;
      RECT  110100.0 653850.0 111300.0 655650.0 ;
      RECT  110100.0 644550.0 111300.0 640950.0 ;
      RECT  112800.0 653850.0 113700.0 644550.0 ;
      RECT  110100.0 644550.0 111300.0 643350.0 ;
      RECT  112500.0 644550.0 113700.0 643350.0 ;
      RECT  112500.0 644550.0 113700.0 643350.0 ;
      RECT  110100.0 644550.0 111300.0 643350.0 ;
      RECT  110100.0 653850.0 111300.0 652650.0 ;
      RECT  112500.0 653850.0 113700.0 652650.0 ;
      RECT  112500.0 653850.0 113700.0 652650.0 ;
      RECT  110100.0 653850.0 111300.0 652650.0 ;
      RECT  114900.0 643950.0 116100.0 642750.0 ;
      RECT  114900.0 653850.0 116100.0 652650.0 ;
      RECT  110700.0 649200.0 111900.0 648000.0 ;
      RECT  110700.0 649200.0 111900.0 648000.0 ;
      RECT  113250.0 649050.0 114150.0 648150.0 ;
      RECT  108300.0 641850.0 117900.0 640950.0 ;
      RECT  108300.0 655650.0 117900.0 654750.0 ;
      RECT  114900.0 667050.0 116100.0 669000.0 ;
      RECT  114900.0 655200.0 116100.0 657150.0 ;
      RECT  110100.0 656550.0 111300.0 654750.0 ;
      RECT  110100.0 665850.0 111300.0 669450.0 ;
      RECT  112800.0 656550.0 113700.0 665850.0 ;
      RECT  110100.0 665850.0 111300.0 667050.0 ;
      RECT  112500.0 665850.0 113700.0 667050.0 ;
      RECT  112500.0 665850.0 113700.0 667050.0 ;
      RECT  110100.0 665850.0 111300.0 667050.0 ;
      RECT  110100.0 656550.0 111300.0 657750.0 ;
      RECT  112500.0 656550.0 113700.0 657750.0 ;
      RECT  112500.0 656550.0 113700.0 657750.0 ;
      RECT  110100.0 656550.0 111300.0 657750.0 ;
      RECT  114900.0 666450.0 116100.0 667650.0 ;
      RECT  114900.0 656550.0 116100.0 657750.0 ;
      RECT  110700.0 661200.0 111900.0 662400.0 ;
      RECT  110700.0 661200.0 111900.0 662400.0 ;
      RECT  113250.0 661350.0 114150.0 662250.0 ;
      RECT  108300.0 668550.0 117900.0 669450.0 ;
      RECT  108300.0 654750.0 117900.0 655650.0 ;
      RECT  114900.0 670950.0 116100.0 669000.0 ;
      RECT  114900.0 682800.0 116100.0 680850.0 ;
      RECT  110100.0 681450.0 111300.0 683250.0 ;
      RECT  110100.0 672150.0 111300.0 668550.0 ;
      RECT  112800.0 681450.0 113700.0 672150.0 ;
      RECT  110100.0 672150.0 111300.0 670950.0 ;
      RECT  112500.0 672150.0 113700.0 670950.0 ;
      RECT  112500.0 672150.0 113700.0 670950.0 ;
      RECT  110100.0 672150.0 111300.0 670950.0 ;
      RECT  110100.0 681450.0 111300.0 680250.0 ;
      RECT  112500.0 681450.0 113700.0 680250.0 ;
      RECT  112500.0 681450.0 113700.0 680250.0 ;
      RECT  110100.0 681450.0 111300.0 680250.0 ;
      RECT  114900.0 671550.0 116100.0 670350.0 ;
      RECT  114900.0 681450.0 116100.0 680250.0 ;
      RECT  110700.0 676800.0 111900.0 675600.0 ;
      RECT  110700.0 676800.0 111900.0 675600.0 ;
      RECT  113250.0 676650.0 114150.0 675750.0 ;
      RECT  108300.0 669450.0 117900.0 668550.0 ;
      RECT  108300.0 683250.0 117900.0 682350.0 ;
      RECT  114900.0 694650.0 116100.0 696600.0 ;
      RECT  114900.0 682800.0 116100.0 684750.0 ;
      RECT  110100.0 684150.0 111300.0 682350.0 ;
      RECT  110100.0 693450.0 111300.0 697050.0 ;
      RECT  112800.0 684150.0 113700.0 693450.0 ;
      RECT  110100.0 693450.0 111300.0 694650.0 ;
      RECT  112500.0 693450.0 113700.0 694650.0 ;
      RECT  112500.0 693450.0 113700.0 694650.0 ;
      RECT  110100.0 693450.0 111300.0 694650.0 ;
      RECT  110100.0 684150.0 111300.0 685350.0 ;
      RECT  112500.0 684150.0 113700.0 685350.0 ;
      RECT  112500.0 684150.0 113700.0 685350.0 ;
      RECT  110100.0 684150.0 111300.0 685350.0 ;
      RECT  114900.0 694050.0 116100.0 695250.0 ;
      RECT  114900.0 684150.0 116100.0 685350.0 ;
      RECT  110700.0 688800.0 111900.0 690000.0 ;
      RECT  110700.0 688800.0 111900.0 690000.0 ;
      RECT  113250.0 688950.0 114150.0 689850.0 ;
      RECT  108300.0 696150.0 117900.0 697050.0 ;
      RECT  108300.0 682350.0 117900.0 683250.0 ;
      RECT  114900.0 698550.0 116100.0 696600.0 ;
      RECT  114900.0 710400.0 116100.0 708450.0 ;
      RECT  110100.0 709050.0 111300.0 710850.0 ;
      RECT  110100.0 699750.0 111300.0 696150.0 ;
      RECT  112800.0 709050.0 113700.0 699750.0 ;
      RECT  110100.0 699750.0 111300.0 698550.0 ;
      RECT  112500.0 699750.0 113700.0 698550.0 ;
      RECT  112500.0 699750.0 113700.0 698550.0 ;
      RECT  110100.0 699750.0 111300.0 698550.0 ;
      RECT  110100.0 709050.0 111300.0 707850.0 ;
      RECT  112500.0 709050.0 113700.0 707850.0 ;
      RECT  112500.0 709050.0 113700.0 707850.0 ;
      RECT  110100.0 709050.0 111300.0 707850.0 ;
      RECT  114900.0 699150.0 116100.0 697950.0 ;
      RECT  114900.0 709050.0 116100.0 707850.0 ;
      RECT  110700.0 704400.0 111900.0 703200.0 ;
      RECT  110700.0 704400.0 111900.0 703200.0 ;
      RECT  113250.0 704250.0 114150.0 703350.0 ;
      RECT  108300.0 697050.0 117900.0 696150.0 ;
      RECT  108300.0 710850.0 117900.0 709950.0 ;
      RECT  114900.0 722250.0 116100.0 724200.0 ;
      RECT  114900.0 710400.0 116100.0 712350.0 ;
      RECT  110100.0 711750.0 111300.0 709950.0 ;
      RECT  110100.0 721050.0 111300.0 724650.0 ;
      RECT  112800.0 711750.0 113700.0 721050.0 ;
      RECT  110100.0 721050.0 111300.0 722250.0 ;
      RECT  112500.0 721050.0 113700.0 722250.0 ;
      RECT  112500.0 721050.0 113700.0 722250.0 ;
      RECT  110100.0 721050.0 111300.0 722250.0 ;
      RECT  110100.0 711750.0 111300.0 712950.0 ;
      RECT  112500.0 711750.0 113700.0 712950.0 ;
      RECT  112500.0 711750.0 113700.0 712950.0 ;
      RECT  110100.0 711750.0 111300.0 712950.0 ;
      RECT  114900.0 721650.0 116100.0 722850.0 ;
      RECT  114900.0 711750.0 116100.0 712950.0 ;
      RECT  110700.0 716400.0 111900.0 717600.0 ;
      RECT  110700.0 716400.0 111900.0 717600.0 ;
      RECT  113250.0 716550.0 114150.0 717450.0 ;
      RECT  108300.0 723750.0 117900.0 724650.0 ;
      RECT  108300.0 709950.0 117900.0 710850.0 ;
      RECT  114900.0 726150.0 116100.0 724200.0 ;
      RECT  114900.0 738000.0 116100.0 736050.0 ;
      RECT  110100.0 736650.0 111300.0 738450.0 ;
      RECT  110100.0 727350.0 111300.0 723750.0 ;
      RECT  112800.0 736650.0 113700.0 727350.0 ;
      RECT  110100.0 727350.0 111300.0 726150.0 ;
      RECT  112500.0 727350.0 113700.0 726150.0 ;
      RECT  112500.0 727350.0 113700.0 726150.0 ;
      RECT  110100.0 727350.0 111300.0 726150.0 ;
      RECT  110100.0 736650.0 111300.0 735450.0 ;
      RECT  112500.0 736650.0 113700.0 735450.0 ;
      RECT  112500.0 736650.0 113700.0 735450.0 ;
      RECT  110100.0 736650.0 111300.0 735450.0 ;
      RECT  114900.0 726750.0 116100.0 725550.0 ;
      RECT  114900.0 736650.0 116100.0 735450.0 ;
      RECT  110700.0 732000.0 111900.0 730800.0 ;
      RECT  110700.0 732000.0 111900.0 730800.0 ;
      RECT  113250.0 731850.0 114150.0 730950.0 ;
      RECT  108300.0 724650.0 117900.0 723750.0 ;
      RECT  108300.0 738450.0 117900.0 737550.0 ;
      RECT  114900.0 749850.0 116100.0 751800.0 ;
      RECT  114900.0 738000.0 116100.0 739950.0 ;
      RECT  110100.0 739350.0 111300.0 737550.0 ;
      RECT  110100.0 748650.0 111300.0 752250.0 ;
      RECT  112800.0 739350.0 113700.0 748650.0 ;
      RECT  110100.0 748650.0 111300.0 749850.0 ;
      RECT  112500.0 748650.0 113700.0 749850.0 ;
      RECT  112500.0 748650.0 113700.0 749850.0 ;
      RECT  110100.0 748650.0 111300.0 749850.0 ;
      RECT  110100.0 739350.0 111300.0 740550.0 ;
      RECT  112500.0 739350.0 113700.0 740550.0 ;
      RECT  112500.0 739350.0 113700.0 740550.0 ;
      RECT  110100.0 739350.0 111300.0 740550.0 ;
      RECT  114900.0 749250.0 116100.0 750450.0 ;
      RECT  114900.0 739350.0 116100.0 740550.0 ;
      RECT  110700.0 744000.0 111900.0 745200.0 ;
      RECT  110700.0 744000.0 111900.0 745200.0 ;
      RECT  113250.0 744150.0 114150.0 745050.0 ;
      RECT  108300.0 751350.0 117900.0 752250.0 ;
      RECT  108300.0 737550.0 117900.0 738450.0 ;
      RECT  114900.0 753750.0 116100.0 751800.0 ;
      RECT  114900.0 765600.0 116100.0 763650.0 ;
      RECT  110100.0 764250.0 111300.0 766050.0 ;
      RECT  110100.0 754950.0 111300.0 751350.0 ;
      RECT  112800.0 764250.0 113700.0 754950.0 ;
      RECT  110100.0 754950.0 111300.0 753750.0 ;
      RECT  112500.0 754950.0 113700.0 753750.0 ;
      RECT  112500.0 754950.0 113700.0 753750.0 ;
      RECT  110100.0 754950.0 111300.0 753750.0 ;
      RECT  110100.0 764250.0 111300.0 763050.0 ;
      RECT  112500.0 764250.0 113700.0 763050.0 ;
      RECT  112500.0 764250.0 113700.0 763050.0 ;
      RECT  110100.0 764250.0 111300.0 763050.0 ;
      RECT  114900.0 754350.0 116100.0 753150.0 ;
      RECT  114900.0 764250.0 116100.0 763050.0 ;
      RECT  110700.0 759600.0 111900.0 758400.0 ;
      RECT  110700.0 759600.0 111900.0 758400.0 ;
      RECT  113250.0 759450.0 114150.0 758550.0 ;
      RECT  108300.0 752250.0 117900.0 751350.0 ;
      RECT  108300.0 766050.0 117900.0 765150.0 ;
      RECT  114900.0 777450.0 116100.0 779400.0 ;
      RECT  114900.0 765600.0 116100.0 767550.0 ;
      RECT  110100.0 766950.0 111300.0 765150.0 ;
      RECT  110100.0 776250.0 111300.0 779850.0 ;
      RECT  112800.0 766950.0 113700.0 776250.0 ;
      RECT  110100.0 776250.0 111300.0 777450.0 ;
      RECT  112500.0 776250.0 113700.0 777450.0 ;
      RECT  112500.0 776250.0 113700.0 777450.0 ;
      RECT  110100.0 776250.0 111300.0 777450.0 ;
      RECT  110100.0 766950.0 111300.0 768150.0 ;
      RECT  112500.0 766950.0 113700.0 768150.0 ;
      RECT  112500.0 766950.0 113700.0 768150.0 ;
      RECT  110100.0 766950.0 111300.0 768150.0 ;
      RECT  114900.0 776850.0 116100.0 778050.0 ;
      RECT  114900.0 766950.0 116100.0 768150.0 ;
      RECT  110700.0 771600.0 111900.0 772800.0 ;
      RECT  110700.0 771600.0 111900.0 772800.0 ;
      RECT  113250.0 771750.0 114150.0 772650.0 ;
      RECT  108300.0 778950.0 117900.0 779850.0 ;
      RECT  108300.0 765150.0 117900.0 766050.0 ;
      RECT  114900.0 781350.0 116100.0 779400.0 ;
      RECT  114900.0 793200.0 116100.0 791250.0 ;
      RECT  110100.0 791850.0 111300.0 793650.0 ;
      RECT  110100.0 782550.0 111300.0 778950.0 ;
      RECT  112800.0 791850.0 113700.0 782550.0 ;
      RECT  110100.0 782550.0 111300.0 781350.0 ;
      RECT  112500.0 782550.0 113700.0 781350.0 ;
      RECT  112500.0 782550.0 113700.0 781350.0 ;
      RECT  110100.0 782550.0 111300.0 781350.0 ;
      RECT  110100.0 791850.0 111300.0 790650.0 ;
      RECT  112500.0 791850.0 113700.0 790650.0 ;
      RECT  112500.0 791850.0 113700.0 790650.0 ;
      RECT  110100.0 791850.0 111300.0 790650.0 ;
      RECT  114900.0 781950.0 116100.0 780750.0 ;
      RECT  114900.0 791850.0 116100.0 790650.0 ;
      RECT  110700.0 787200.0 111900.0 786000.0 ;
      RECT  110700.0 787200.0 111900.0 786000.0 ;
      RECT  113250.0 787050.0 114150.0 786150.0 ;
      RECT  108300.0 779850.0 117900.0 778950.0 ;
      RECT  108300.0 793650.0 117900.0 792750.0 ;
      RECT  114900.0 805050.0 116100.0 807000.0 ;
      RECT  114900.0 793200.0 116100.0 795150.0 ;
      RECT  110100.0 794550.0 111300.0 792750.0 ;
      RECT  110100.0 803850.0 111300.0 807450.0 ;
      RECT  112800.0 794550.0 113700.0 803850.0 ;
      RECT  110100.0 803850.0 111300.0 805050.0 ;
      RECT  112500.0 803850.0 113700.0 805050.0 ;
      RECT  112500.0 803850.0 113700.0 805050.0 ;
      RECT  110100.0 803850.0 111300.0 805050.0 ;
      RECT  110100.0 794550.0 111300.0 795750.0 ;
      RECT  112500.0 794550.0 113700.0 795750.0 ;
      RECT  112500.0 794550.0 113700.0 795750.0 ;
      RECT  110100.0 794550.0 111300.0 795750.0 ;
      RECT  114900.0 804450.0 116100.0 805650.0 ;
      RECT  114900.0 794550.0 116100.0 795750.0 ;
      RECT  110700.0 799200.0 111900.0 800400.0 ;
      RECT  110700.0 799200.0 111900.0 800400.0 ;
      RECT  113250.0 799350.0 114150.0 800250.0 ;
      RECT  108300.0 806550.0 117900.0 807450.0 ;
      RECT  108300.0 792750.0 117900.0 793650.0 ;
      RECT  114900.0 808950.0 116100.0 807000.0 ;
      RECT  114900.0 820800.0 116100.0 818850.0 ;
      RECT  110100.0 819450.0 111300.0 821250.0 ;
      RECT  110100.0 810150.0 111300.0 806550.0 ;
      RECT  112800.0 819450.0 113700.0 810150.0 ;
      RECT  110100.0 810150.0 111300.0 808950.0 ;
      RECT  112500.0 810150.0 113700.0 808950.0 ;
      RECT  112500.0 810150.0 113700.0 808950.0 ;
      RECT  110100.0 810150.0 111300.0 808950.0 ;
      RECT  110100.0 819450.0 111300.0 818250.0 ;
      RECT  112500.0 819450.0 113700.0 818250.0 ;
      RECT  112500.0 819450.0 113700.0 818250.0 ;
      RECT  110100.0 819450.0 111300.0 818250.0 ;
      RECT  114900.0 809550.0 116100.0 808350.0 ;
      RECT  114900.0 819450.0 116100.0 818250.0 ;
      RECT  110700.0 814800.0 111900.0 813600.0 ;
      RECT  110700.0 814800.0 111900.0 813600.0 ;
      RECT  113250.0 814650.0 114150.0 813750.0 ;
      RECT  108300.0 807450.0 117900.0 806550.0 ;
      RECT  108300.0 821250.0 117900.0 820350.0 ;
      RECT  114900.0 832650.0 116100.0 834600.0 ;
      RECT  114900.0 820800.0 116100.0 822750.0 ;
      RECT  110100.0 822150.0 111300.0 820350.0 ;
      RECT  110100.0 831450.0 111300.0 835050.0 ;
      RECT  112800.0 822150.0 113700.0 831450.0 ;
      RECT  110100.0 831450.0 111300.0 832650.0 ;
      RECT  112500.0 831450.0 113700.0 832650.0 ;
      RECT  112500.0 831450.0 113700.0 832650.0 ;
      RECT  110100.0 831450.0 111300.0 832650.0 ;
      RECT  110100.0 822150.0 111300.0 823350.0 ;
      RECT  112500.0 822150.0 113700.0 823350.0 ;
      RECT  112500.0 822150.0 113700.0 823350.0 ;
      RECT  110100.0 822150.0 111300.0 823350.0 ;
      RECT  114900.0 832050.0 116100.0 833250.0 ;
      RECT  114900.0 822150.0 116100.0 823350.0 ;
      RECT  110700.0 826800.0 111900.0 828000.0 ;
      RECT  110700.0 826800.0 111900.0 828000.0 ;
      RECT  113250.0 826950.0 114150.0 827850.0 ;
      RECT  108300.0 834150.0 117900.0 835050.0 ;
      RECT  108300.0 820350.0 117900.0 821250.0 ;
      RECT  114900.0 836550.0 116100.0 834600.0 ;
      RECT  114900.0 848400.0 116100.0 846450.0 ;
      RECT  110100.0 847050.0 111300.0 848850.0 ;
      RECT  110100.0 837750.0 111300.0 834150.0 ;
      RECT  112800.0 847050.0 113700.0 837750.0 ;
      RECT  110100.0 837750.0 111300.0 836550.0 ;
      RECT  112500.0 837750.0 113700.0 836550.0 ;
      RECT  112500.0 837750.0 113700.0 836550.0 ;
      RECT  110100.0 837750.0 111300.0 836550.0 ;
      RECT  110100.0 847050.0 111300.0 845850.0 ;
      RECT  112500.0 847050.0 113700.0 845850.0 ;
      RECT  112500.0 847050.0 113700.0 845850.0 ;
      RECT  110100.0 847050.0 111300.0 845850.0 ;
      RECT  114900.0 837150.0 116100.0 835950.0 ;
      RECT  114900.0 847050.0 116100.0 845850.0 ;
      RECT  110700.0 842400.0 111900.0 841200.0 ;
      RECT  110700.0 842400.0 111900.0 841200.0 ;
      RECT  113250.0 842250.0 114150.0 841350.0 ;
      RECT  108300.0 835050.0 117900.0 834150.0 ;
      RECT  108300.0 848850.0 117900.0 847950.0 ;
      RECT  114900.0 860250.0 116100.0 862200.0 ;
      RECT  114900.0 848400.0 116100.0 850350.0 ;
      RECT  110100.0 849750.0 111300.0 847950.0 ;
      RECT  110100.0 859050.0 111300.0 862650.0 ;
      RECT  112800.0 849750.0 113700.0 859050.0 ;
      RECT  110100.0 859050.0 111300.0 860250.0 ;
      RECT  112500.0 859050.0 113700.0 860250.0 ;
      RECT  112500.0 859050.0 113700.0 860250.0 ;
      RECT  110100.0 859050.0 111300.0 860250.0 ;
      RECT  110100.0 849750.0 111300.0 850950.0 ;
      RECT  112500.0 849750.0 113700.0 850950.0 ;
      RECT  112500.0 849750.0 113700.0 850950.0 ;
      RECT  110100.0 849750.0 111300.0 850950.0 ;
      RECT  114900.0 859650.0 116100.0 860850.0 ;
      RECT  114900.0 849750.0 116100.0 850950.0 ;
      RECT  110700.0 854400.0 111900.0 855600.0 ;
      RECT  110700.0 854400.0 111900.0 855600.0 ;
      RECT  113250.0 854550.0 114150.0 855450.0 ;
      RECT  108300.0 861750.0 117900.0 862650.0 ;
      RECT  108300.0 847950.0 117900.0 848850.0 ;
      RECT  114900.0 864150.0 116100.0 862200.0 ;
      RECT  114900.0 876000.0 116100.0 874050.0 ;
      RECT  110100.0 874650.0 111300.0 876450.0 ;
      RECT  110100.0 865350.0 111300.0 861750.0 ;
      RECT  112800.0 874650.0 113700.0 865350.0 ;
      RECT  110100.0 865350.0 111300.0 864150.0 ;
      RECT  112500.0 865350.0 113700.0 864150.0 ;
      RECT  112500.0 865350.0 113700.0 864150.0 ;
      RECT  110100.0 865350.0 111300.0 864150.0 ;
      RECT  110100.0 874650.0 111300.0 873450.0 ;
      RECT  112500.0 874650.0 113700.0 873450.0 ;
      RECT  112500.0 874650.0 113700.0 873450.0 ;
      RECT  110100.0 874650.0 111300.0 873450.0 ;
      RECT  114900.0 864750.0 116100.0 863550.0 ;
      RECT  114900.0 874650.0 116100.0 873450.0 ;
      RECT  110700.0 870000.0 111900.0 868800.0 ;
      RECT  110700.0 870000.0 111900.0 868800.0 ;
      RECT  113250.0 869850.0 114150.0 868950.0 ;
      RECT  108300.0 862650.0 117900.0 861750.0 ;
      RECT  108300.0 876450.0 117900.0 875550.0 ;
      RECT  114900.0 887850.0 116100.0 889800.0 ;
      RECT  114900.0 876000.0 116100.0 877950.0 ;
      RECT  110100.0 877350.0 111300.0 875550.0 ;
      RECT  110100.0 886650.0 111300.0 890250.0 ;
      RECT  112800.0 877350.0 113700.0 886650.0 ;
      RECT  110100.0 886650.0 111300.0 887850.0 ;
      RECT  112500.0 886650.0 113700.0 887850.0 ;
      RECT  112500.0 886650.0 113700.0 887850.0 ;
      RECT  110100.0 886650.0 111300.0 887850.0 ;
      RECT  110100.0 877350.0 111300.0 878550.0 ;
      RECT  112500.0 877350.0 113700.0 878550.0 ;
      RECT  112500.0 877350.0 113700.0 878550.0 ;
      RECT  110100.0 877350.0 111300.0 878550.0 ;
      RECT  114900.0 887250.0 116100.0 888450.0 ;
      RECT  114900.0 877350.0 116100.0 878550.0 ;
      RECT  110700.0 882000.0 111900.0 883200.0 ;
      RECT  110700.0 882000.0 111900.0 883200.0 ;
      RECT  113250.0 882150.0 114150.0 883050.0 ;
      RECT  108300.0 889350.0 117900.0 890250.0 ;
      RECT  108300.0 875550.0 117900.0 876450.0 ;
      RECT  114900.0 891750.0 116100.0 889800.0 ;
      RECT  114900.0 903600.0 116100.0 901650.0 ;
      RECT  110100.0 902250.0 111300.0 904050.0 ;
      RECT  110100.0 892950.0 111300.0 889350.0 ;
      RECT  112800.0 902250.0 113700.0 892950.0 ;
      RECT  110100.0 892950.0 111300.0 891750.0 ;
      RECT  112500.0 892950.0 113700.0 891750.0 ;
      RECT  112500.0 892950.0 113700.0 891750.0 ;
      RECT  110100.0 892950.0 111300.0 891750.0 ;
      RECT  110100.0 902250.0 111300.0 901050.0 ;
      RECT  112500.0 902250.0 113700.0 901050.0 ;
      RECT  112500.0 902250.0 113700.0 901050.0 ;
      RECT  110100.0 902250.0 111300.0 901050.0 ;
      RECT  114900.0 892350.0 116100.0 891150.0 ;
      RECT  114900.0 902250.0 116100.0 901050.0 ;
      RECT  110700.0 897600.0 111900.0 896400.0 ;
      RECT  110700.0 897600.0 111900.0 896400.0 ;
      RECT  113250.0 897450.0 114150.0 896550.0 ;
      RECT  108300.0 890250.0 117900.0 889350.0 ;
      RECT  108300.0 904050.0 117900.0 903150.0 ;
      RECT  114900.0 915450.0 116100.0 917400.0 ;
      RECT  114900.0 903600.0 116100.0 905550.0 ;
      RECT  110100.0 904950.0 111300.0 903150.0 ;
      RECT  110100.0 914250.0 111300.0 917850.0 ;
      RECT  112800.0 904950.0 113700.0 914250.0 ;
      RECT  110100.0 914250.0 111300.0 915450.0 ;
      RECT  112500.0 914250.0 113700.0 915450.0 ;
      RECT  112500.0 914250.0 113700.0 915450.0 ;
      RECT  110100.0 914250.0 111300.0 915450.0 ;
      RECT  110100.0 904950.0 111300.0 906150.0 ;
      RECT  112500.0 904950.0 113700.0 906150.0 ;
      RECT  112500.0 904950.0 113700.0 906150.0 ;
      RECT  110100.0 904950.0 111300.0 906150.0 ;
      RECT  114900.0 914850.0 116100.0 916050.0 ;
      RECT  114900.0 904950.0 116100.0 906150.0 ;
      RECT  110700.0 909600.0 111900.0 910800.0 ;
      RECT  110700.0 909600.0 111900.0 910800.0 ;
      RECT  113250.0 909750.0 114150.0 910650.0 ;
      RECT  108300.0 916950.0 117900.0 917850.0 ;
      RECT  108300.0 903150.0 117900.0 904050.0 ;
      RECT  114900.0 919350.0 116100.0 917400.0 ;
      RECT  114900.0 931200.0 116100.0 929250.0 ;
      RECT  110100.0 929850.0 111300.0 931650.0 ;
      RECT  110100.0 920550.0 111300.0 916950.0 ;
      RECT  112800.0 929850.0 113700.0 920550.0 ;
      RECT  110100.0 920550.0 111300.0 919350.0 ;
      RECT  112500.0 920550.0 113700.0 919350.0 ;
      RECT  112500.0 920550.0 113700.0 919350.0 ;
      RECT  110100.0 920550.0 111300.0 919350.0 ;
      RECT  110100.0 929850.0 111300.0 928650.0 ;
      RECT  112500.0 929850.0 113700.0 928650.0 ;
      RECT  112500.0 929850.0 113700.0 928650.0 ;
      RECT  110100.0 929850.0 111300.0 928650.0 ;
      RECT  114900.0 919950.0 116100.0 918750.0 ;
      RECT  114900.0 929850.0 116100.0 928650.0 ;
      RECT  110700.0 925200.0 111900.0 924000.0 ;
      RECT  110700.0 925200.0 111900.0 924000.0 ;
      RECT  113250.0 925050.0 114150.0 924150.0 ;
      RECT  108300.0 917850.0 117900.0 916950.0 ;
      RECT  108300.0 931650.0 117900.0 930750.0 ;
      RECT  114900.0 943050.0 116100.0 945000.0 ;
      RECT  114900.0 931200.0 116100.0 933150.0 ;
      RECT  110100.0 932550.0 111300.0 930750.0 ;
      RECT  110100.0 941850.0 111300.0 945450.0 ;
      RECT  112800.0 932550.0 113700.0 941850.0 ;
      RECT  110100.0 941850.0 111300.0 943050.0 ;
      RECT  112500.0 941850.0 113700.0 943050.0 ;
      RECT  112500.0 941850.0 113700.0 943050.0 ;
      RECT  110100.0 941850.0 111300.0 943050.0 ;
      RECT  110100.0 932550.0 111300.0 933750.0 ;
      RECT  112500.0 932550.0 113700.0 933750.0 ;
      RECT  112500.0 932550.0 113700.0 933750.0 ;
      RECT  110100.0 932550.0 111300.0 933750.0 ;
      RECT  114900.0 942450.0 116100.0 943650.0 ;
      RECT  114900.0 932550.0 116100.0 933750.0 ;
      RECT  110700.0 937200.0 111900.0 938400.0 ;
      RECT  110700.0 937200.0 111900.0 938400.0 ;
      RECT  113250.0 937350.0 114150.0 938250.0 ;
      RECT  108300.0 944550.0 117900.0 945450.0 ;
      RECT  108300.0 930750.0 117900.0 931650.0 ;
      RECT  114900.0 946950.0 116100.0 945000.0 ;
      RECT  114900.0 958800.0 116100.0 956850.0 ;
      RECT  110100.0 957450.0 111300.0 959250.0 ;
      RECT  110100.0 948150.0 111300.0 944550.0 ;
      RECT  112800.0 957450.0 113700.0 948150.0 ;
      RECT  110100.0 948150.0 111300.0 946950.0 ;
      RECT  112500.0 948150.0 113700.0 946950.0 ;
      RECT  112500.0 948150.0 113700.0 946950.0 ;
      RECT  110100.0 948150.0 111300.0 946950.0 ;
      RECT  110100.0 957450.0 111300.0 956250.0 ;
      RECT  112500.0 957450.0 113700.0 956250.0 ;
      RECT  112500.0 957450.0 113700.0 956250.0 ;
      RECT  110100.0 957450.0 111300.0 956250.0 ;
      RECT  114900.0 947550.0 116100.0 946350.0 ;
      RECT  114900.0 957450.0 116100.0 956250.0 ;
      RECT  110700.0 952800.0 111900.0 951600.0 ;
      RECT  110700.0 952800.0 111900.0 951600.0 ;
      RECT  113250.0 952650.0 114150.0 951750.0 ;
      RECT  108300.0 945450.0 117900.0 944550.0 ;
      RECT  108300.0 959250.0 117900.0 958350.0 ;
      RECT  114900.0 970650.0 116100.0 972600.0 ;
      RECT  114900.0 958800.0 116100.0 960750.0 ;
      RECT  110100.0 960150.0 111300.0 958350.0 ;
      RECT  110100.0 969450.0 111300.0 973050.0 ;
      RECT  112800.0 960150.0 113700.0 969450.0 ;
      RECT  110100.0 969450.0 111300.0 970650.0 ;
      RECT  112500.0 969450.0 113700.0 970650.0 ;
      RECT  112500.0 969450.0 113700.0 970650.0 ;
      RECT  110100.0 969450.0 111300.0 970650.0 ;
      RECT  110100.0 960150.0 111300.0 961350.0 ;
      RECT  112500.0 960150.0 113700.0 961350.0 ;
      RECT  112500.0 960150.0 113700.0 961350.0 ;
      RECT  110100.0 960150.0 111300.0 961350.0 ;
      RECT  114900.0 970050.0 116100.0 971250.0 ;
      RECT  114900.0 960150.0 116100.0 961350.0 ;
      RECT  110700.0 964800.0 111900.0 966000.0 ;
      RECT  110700.0 964800.0 111900.0 966000.0 ;
      RECT  113250.0 964950.0 114150.0 965850.0 ;
      RECT  108300.0 972150.0 117900.0 973050.0 ;
      RECT  108300.0 958350.0 117900.0 959250.0 ;
      RECT  114900.0 974550.0 116100.0 972600.0 ;
      RECT  114900.0 986400.0 116100.0 984450.0 ;
      RECT  110100.0 985050.0 111300.0 986850.0 ;
      RECT  110100.0 975750.0 111300.0 972150.0 ;
      RECT  112800.0 985050.0 113700.0 975750.0 ;
      RECT  110100.0 975750.0 111300.0 974550.0 ;
      RECT  112500.0 975750.0 113700.0 974550.0 ;
      RECT  112500.0 975750.0 113700.0 974550.0 ;
      RECT  110100.0 975750.0 111300.0 974550.0 ;
      RECT  110100.0 985050.0 111300.0 983850.0 ;
      RECT  112500.0 985050.0 113700.0 983850.0 ;
      RECT  112500.0 985050.0 113700.0 983850.0 ;
      RECT  110100.0 985050.0 111300.0 983850.0 ;
      RECT  114900.0 975150.0 116100.0 973950.0 ;
      RECT  114900.0 985050.0 116100.0 983850.0 ;
      RECT  110700.0 980400.0 111900.0 979200.0 ;
      RECT  110700.0 980400.0 111900.0 979200.0 ;
      RECT  113250.0 980250.0 114150.0 979350.0 ;
      RECT  108300.0 973050.0 117900.0 972150.0 ;
      RECT  108300.0 986850.0 117900.0 985950.0 ;
      RECT  114900.0 998250.0 116100.0 1000200.0 ;
      RECT  114900.0 986400.0 116100.0 988350.0 ;
      RECT  110100.0 987750.0 111300.0 985950.0 ;
      RECT  110100.0 997050.0 111300.0 1000650.0 ;
      RECT  112800.0 987750.0 113700.0 997050.0 ;
      RECT  110100.0 997050.0 111300.0 998250.0 ;
      RECT  112500.0 997050.0 113700.0 998250.0 ;
      RECT  112500.0 997050.0 113700.0 998250.0 ;
      RECT  110100.0 997050.0 111300.0 998250.0 ;
      RECT  110100.0 987750.0 111300.0 988950.0 ;
      RECT  112500.0 987750.0 113700.0 988950.0 ;
      RECT  112500.0 987750.0 113700.0 988950.0 ;
      RECT  110100.0 987750.0 111300.0 988950.0 ;
      RECT  114900.0 997650.0 116100.0 998850.0 ;
      RECT  114900.0 987750.0 116100.0 988950.0 ;
      RECT  110700.0 992400.0 111900.0 993600.0 ;
      RECT  110700.0 992400.0 111900.0 993600.0 ;
      RECT  113250.0 992550.0 114150.0 993450.0 ;
      RECT  108300.0 999750.0 117900.0 1000650.0 ;
      RECT  108300.0 985950.0 117900.0 986850.0 ;
      RECT  114900.0 1002150.0 116100.0 1000200.0 ;
      RECT  114900.0 1014000.0 116100.0 1012050.0 ;
      RECT  110100.0 1012650.0 111300.0 1014450.0 ;
      RECT  110100.0 1003350.0 111300.0 999750.0 ;
      RECT  112800.0 1012650.0 113700.0 1003350.0 ;
      RECT  110100.0 1003350.0 111300.0 1002150.0 ;
      RECT  112500.0 1003350.0 113700.0 1002150.0 ;
      RECT  112500.0 1003350.0 113700.0 1002150.0 ;
      RECT  110100.0 1003350.0 111300.0 1002150.0 ;
      RECT  110100.0 1012650.0 111300.0 1011450.0 ;
      RECT  112500.0 1012650.0 113700.0 1011450.0 ;
      RECT  112500.0 1012650.0 113700.0 1011450.0 ;
      RECT  110100.0 1012650.0 111300.0 1011450.0 ;
      RECT  114900.0 1002750.0 116100.0 1001550.0 ;
      RECT  114900.0 1012650.0 116100.0 1011450.0 ;
      RECT  110700.0 1008000.0 111900.0 1006800.0 ;
      RECT  110700.0 1008000.0 111900.0 1006800.0 ;
      RECT  113250.0 1007850.0 114150.0 1006950.0 ;
      RECT  108300.0 1000650.0 117900.0 999750.0 ;
      RECT  108300.0 1014450.0 117900.0 1013550.0 ;
      RECT  114900.0 1025850.0 116100.0 1027800.0 ;
      RECT  114900.0 1014000.0 116100.0 1015950.0 ;
      RECT  110100.0 1015350.0 111300.0 1013550.0 ;
      RECT  110100.0 1024650.0 111300.0 1028250.0 ;
      RECT  112800.0 1015350.0 113700.0 1024650.0 ;
      RECT  110100.0 1024650.0 111300.0 1025850.0 ;
      RECT  112500.0 1024650.0 113700.0 1025850.0 ;
      RECT  112500.0 1024650.0 113700.0 1025850.0 ;
      RECT  110100.0 1024650.0 111300.0 1025850.0 ;
      RECT  110100.0 1015350.0 111300.0 1016550.0 ;
      RECT  112500.0 1015350.0 113700.0 1016550.0 ;
      RECT  112500.0 1015350.0 113700.0 1016550.0 ;
      RECT  110100.0 1015350.0 111300.0 1016550.0 ;
      RECT  114900.0 1025250.0 116100.0 1026450.0 ;
      RECT  114900.0 1015350.0 116100.0 1016550.0 ;
      RECT  110700.0 1020000.0 111900.0 1021200.0 ;
      RECT  110700.0 1020000.0 111900.0 1021200.0 ;
      RECT  113250.0 1020150.0 114150.0 1021050.0 ;
      RECT  108300.0 1027350.0 117900.0 1028250.0 ;
      RECT  108300.0 1013550.0 117900.0 1014450.0 ;
      RECT  114900.0 1029750.0 116100.0 1027800.0 ;
      RECT  114900.0 1041600.0 116100.0 1039650.0 ;
      RECT  110100.0 1040250.0 111300.0 1042050.0 ;
      RECT  110100.0 1030950.0 111300.0 1027350.0 ;
      RECT  112800.0 1040250.0 113700.0 1030950.0 ;
      RECT  110100.0 1030950.0 111300.0 1029750.0 ;
      RECT  112500.0 1030950.0 113700.0 1029750.0 ;
      RECT  112500.0 1030950.0 113700.0 1029750.0 ;
      RECT  110100.0 1030950.0 111300.0 1029750.0 ;
      RECT  110100.0 1040250.0 111300.0 1039050.0 ;
      RECT  112500.0 1040250.0 113700.0 1039050.0 ;
      RECT  112500.0 1040250.0 113700.0 1039050.0 ;
      RECT  110100.0 1040250.0 111300.0 1039050.0 ;
      RECT  114900.0 1030350.0 116100.0 1029150.0 ;
      RECT  114900.0 1040250.0 116100.0 1039050.0 ;
      RECT  110700.0 1035600.0 111900.0 1034400.0 ;
      RECT  110700.0 1035600.0 111900.0 1034400.0 ;
      RECT  113250.0 1035450.0 114150.0 1034550.0 ;
      RECT  108300.0 1028250.0 117900.0 1027350.0 ;
      RECT  108300.0 1042050.0 117900.0 1041150.0 ;
      RECT  114900.0 1053450.0 116100.0 1055400.0 ;
      RECT  114900.0 1041600.0 116100.0 1043550.0 ;
      RECT  110100.0 1042950.0 111300.0 1041150.0 ;
      RECT  110100.0 1052250.0 111300.0 1055850.0 ;
      RECT  112800.0 1042950.0 113700.0 1052250.0 ;
      RECT  110100.0 1052250.0 111300.0 1053450.0 ;
      RECT  112500.0 1052250.0 113700.0 1053450.0 ;
      RECT  112500.0 1052250.0 113700.0 1053450.0 ;
      RECT  110100.0 1052250.0 111300.0 1053450.0 ;
      RECT  110100.0 1042950.0 111300.0 1044150.0 ;
      RECT  112500.0 1042950.0 113700.0 1044150.0 ;
      RECT  112500.0 1042950.0 113700.0 1044150.0 ;
      RECT  110100.0 1042950.0 111300.0 1044150.0 ;
      RECT  114900.0 1052850.0 116100.0 1054050.0 ;
      RECT  114900.0 1042950.0 116100.0 1044150.0 ;
      RECT  110700.0 1047600.0 111900.0 1048800.0 ;
      RECT  110700.0 1047600.0 111900.0 1048800.0 ;
      RECT  113250.0 1047750.0 114150.0 1048650.0 ;
      RECT  108300.0 1054950.0 117900.0 1055850.0 ;
      RECT  108300.0 1041150.0 117900.0 1042050.0 ;
      RECT  114900.0 1057350.0 116100.0 1055400.0 ;
      RECT  114900.0 1069200.0 116100.0 1067250.0 ;
      RECT  110100.0 1067850.0 111300.0 1069650.0 ;
      RECT  110100.0 1058550.0 111300.0 1054950.0 ;
      RECT  112800.0 1067850.0 113700.0 1058550.0 ;
      RECT  110100.0 1058550.0 111300.0 1057350.0 ;
      RECT  112500.0 1058550.0 113700.0 1057350.0 ;
      RECT  112500.0 1058550.0 113700.0 1057350.0 ;
      RECT  110100.0 1058550.0 111300.0 1057350.0 ;
      RECT  110100.0 1067850.0 111300.0 1066650.0 ;
      RECT  112500.0 1067850.0 113700.0 1066650.0 ;
      RECT  112500.0 1067850.0 113700.0 1066650.0 ;
      RECT  110100.0 1067850.0 111300.0 1066650.0 ;
      RECT  114900.0 1057950.0 116100.0 1056750.0 ;
      RECT  114900.0 1067850.0 116100.0 1066650.0 ;
      RECT  110700.0 1063200.0 111900.0 1062000.0 ;
      RECT  110700.0 1063200.0 111900.0 1062000.0 ;
      RECT  113250.0 1063050.0 114150.0 1062150.0 ;
      RECT  108300.0 1055850.0 117900.0 1054950.0 ;
      RECT  108300.0 1069650.0 117900.0 1068750.0 ;
      RECT  114900.0 1081050.0 116100.0 1083000.0 ;
      RECT  114900.0 1069200.0 116100.0 1071150.0 ;
      RECT  110100.0 1070550.0 111300.0 1068750.0 ;
      RECT  110100.0 1079850.0 111300.0 1083450.0 ;
      RECT  112800.0 1070550.0 113700.0 1079850.0 ;
      RECT  110100.0 1079850.0 111300.0 1081050.0 ;
      RECT  112500.0 1079850.0 113700.0 1081050.0 ;
      RECT  112500.0 1079850.0 113700.0 1081050.0 ;
      RECT  110100.0 1079850.0 111300.0 1081050.0 ;
      RECT  110100.0 1070550.0 111300.0 1071750.0 ;
      RECT  112500.0 1070550.0 113700.0 1071750.0 ;
      RECT  112500.0 1070550.0 113700.0 1071750.0 ;
      RECT  110100.0 1070550.0 111300.0 1071750.0 ;
      RECT  114900.0 1080450.0 116100.0 1081650.0 ;
      RECT  114900.0 1070550.0 116100.0 1071750.0 ;
      RECT  110700.0 1075200.0 111900.0 1076400.0 ;
      RECT  110700.0 1075200.0 111900.0 1076400.0 ;
      RECT  113250.0 1075350.0 114150.0 1076250.0 ;
      RECT  108300.0 1082550.0 117900.0 1083450.0 ;
      RECT  108300.0 1068750.0 117900.0 1069650.0 ;
      RECT  114900.0 1084950.0 116100.0 1083000.0 ;
      RECT  114900.0 1096800.0 116100.0 1094850.0 ;
      RECT  110100.0 1095450.0 111300.0 1097250.0 ;
      RECT  110100.0 1086150.0 111300.0 1082550.0 ;
      RECT  112800.0 1095450.0 113700.0 1086150.0 ;
      RECT  110100.0 1086150.0 111300.0 1084950.0 ;
      RECT  112500.0 1086150.0 113700.0 1084950.0 ;
      RECT  112500.0 1086150.0 113700.0 1084950.0 ;
      RECT  110100.0 1086150.0 111300.0 1084950.0 ;
      RECT  110100.0 1095450.0 111300.0 1094250.0 ;
      RECT  112500.0 1095450.0 113700.0 1094250.0 ;
      RECT  112500.0 1095450.0 113700.0 1094250.0 ;
      RECT  110100.0 1095450.0 111300.0 1094250.0 ;
      RECT  114900.0 1085550.0 116100.0 1084350.0 ;
      RECT  114900.0 1095450.0 116100.0 1094250.0 ;
      RECT  110700.0 1090800.0 111900.0 1089600.0 ;
      RECT  110700.0 1090800.0 111900.0 1089600.0 ;
      RECT  113250.0 1090650.0 114150.0 1089750.0 ;
      RECT  108300.0 1083450.0 117900.0 1082550.0 ;
      RECT  108300.0 1097250.0 117900.0 1096350.0 ;
      RECT  114900.0 1108650.0 116100.0 1110600.0 ;
      RECT  114900.0 1096800.0 116100.0 1098750.0 ;
      RECT  110100.0 1098150.0 111300.0 1096350.0 ;
      RECT  110100.0 1107450.0 111300.0 1111050.0 ;
      RECT  112800.0 1098150.0 113700.0 1107450.0 ;
      RECT  110100.0 1107450.0 111300.0 1108650.0 ;
      RECT  112500.0 1107450.0 113700.0 1108650.0 ;
      RECT  112500.0 1107450.0 113700.0 1108650.0 ;
      RECT  110100.0 1107450.0 111300.0 1108650.0 ;
      RECT  110100.0 1098150.0 111300.0 1099350.0 ;
      RECT  112500.0 1098150.0 113700.0 1099350.0 ;
      RECT  112500.0 1098150.0 113700.0 1099350.0 ;
      RECT  110100.0 1098150.0 111300.0 1099350.0 ;
      RECT  114900.0 1108050.0 116100.0 1109250.0 ;
      RECT  114900.0 1098150.0 116100.0 1099350.0 ;
      RECT  110700.0 1102800.0 111900.0 1104000.0 ;
      RECT  110700.0 1102800.0 111900.0 1104000.0 ;
      RECT  113250.0 1102950.0 114150.0 1103850.0 ;
      RECT  108300.0 1110150.0 117900.0 1111050.0 ;
      RECT  108300.0 1096350.0 117900.0 1097250.0 ;
      RECT  114900.0 1112550.0 116100.0 1110600.0 ;
      RECT  114900.0 1124400.0 116100.0 1122450.0 ;
      RECT  110100.0 1123050.0 111300.0 1124850.0 ;
      RECT  110100.0 1113750.0 111300.0 1110150.0 ;
      RECT  112800.0 1123050.0 113700.0 1113750.0 ;
      RECT  110100.0 1113750.0 111300.0 1112550.0 ;
      RECT  112500.0 1113750.0 113700.0 1112550.0 ;
      RECT  112500.0 1113750.0 113700.0 1112550.0 ;
      RECT  110100.0 1113750.0 111300.0 1112550.0 ;
      RECT  110100.0 1123050.0 111300.0 1121850.0 ;
      RECT  112500.0 1123050.0 113700.0 1121850.0 ;
      RECT  112500.0 1123050.0 113700.0 1121850.0 ;
      RECT  110100.0 1123050.0 111300.0 1121850.0 ;
      RECT  114900.0 1113150.0 116100.0 1111950.0 ;
      RECT  114900.0 1123050.0 116100.0 1121850.0 ;
      RECT  110700.0 1118400.0 111900.0 1117200.0 ;
      RECT  110700.0 1118400.0 111900.0 1117200.0 ;
      RECT  113250.0 1118250.0 114150.0 1117350.0 ;
      RECT  108300.0 1111050.0 117900.0 1110150.0 ;
      RECT  108300.0 1124850.0 117900.0 1123950.0 ;
      RECT  114900.0 1136250.0 116100.0 1138200.0 ;
      RECT  114900.0 1124400.0 116100.0 1126350.0 ;
      RECT  110100.0 1125750.0 111300.0 1123950.0 ;
      RECT  110100.0 1135050.0 111300.0 1138650.0 ;
      RECT  112800.0 1125750.0 113700.0 1135050.0 ;
      RECT  110100.0 1135050.0 111300.0 1136250.0 ;
      RECT  112500.0 1135050.0 113700.0 1136250.0 ;
      RECT  112500.0 1135050.0 113700.0 1136250.0 ;
      RECT  110100.0 1135050.0 111300.0 1136250.0 ;
      RECT  110100.0 1125750.0 111300.0 1126950.0 ;
      RECT  112500.0 1125750.0 113700.0 1126950.0 ;
      RECT  112500.0 1125750.0 113700.0 1126950.0 ;
      RECT  110100.0 1125750.0 111300.0 1126950.0 ;
      RECT  114900.0 1135650.0 116100.0 1136850.0 ;
      RECT  114900.0 1125750.0 116100.0 1126950.0 ;
      RECT  110700.0 1130400.0 111900.0 1131600.0 ;
      RECT  110700.0 1130400.0 111900.0 1131600.0 ;
      RECT  113250.0 1130550.0 114150.0 1131450.0 ;
      RECT  108300.0 1137750.0 117900.0 1138650.0 ;
      RECT  108300.0 1123950.0 117900.0 1124850.0 ;
      RECT  114900.0 1140150.0 116100.0 1138200.0 ;
      RECT  114900.0 1152000.0 116100.0 1150050.0 ;
      RECT  110100.0 1150650.0 111300.0 1152450.0 ;
      RECT  110100.0 1141350.0 111300.0 1137750.0 ;
      RECT  112800.0 1150650.0 113700.0 1141350.0 ;
      RECT  110100.0 1141350.0 111300.0 1140150.0 ;
      RECT  112500.0 1141350.0 113700.0 1140150.0 ;
      RECT  112500.0 1141350.0 113700.0 1140150.0 ;
      RECT  110100.0 1141350.0 111300.0 1140150.0 ;
      RECT  110100.0 1150650.0 111300.0 1149450.0 ;
      RECT  112500.0 1150650.0 113700.0 1149450.0 ;
      RECT  112500.0 1150650.0 113700.0 1149450.0 ;
      RECT  110100.0 1150650.0 111300.0 1149450.0 ;
      RECT  114900.0 1140750.0 116100.0 1139550.0 ;
      RECT  114900.0 1150650.0 116100.0 1149450.0 ;
      RECT  110700.0 1146000.0 111900.0 1144800.0 ;
      RECT  110700.0 1146000.0 111900.0 1144800.0 ;
      RECT  113250.0 1145850.0 114150.0 1144950.0 ;
      RECT  108300.0 1138650.0 117900.0 1137750.0 ;
      RECT  108300.0 1152450.0 117900.0 1151550.0 ;
      RECT  114900.0 1163850.0 116100.0 1165800.0 ;
      RECT  114900.0 1152000.0 116100.0 1153950.0 ;
      RECT  110100.0 1153350.0 111300.0 1151550.0 ;
      RECT  110100.0 1162650.0 111300.0 1166250.0 ;
      RECT  112800.0 1153350.0 113700.0 1162650.0 ;
      RECT  110100.0 1162650.0 111300.0 1163850.0 ;
      RECT  112500.0 1162650.0 113700.0 1163850.0 ;
      RECT  112500.0 1162650.0 113700.0 1163850.0 ;
      RECT  110100.0 1162650.0 111300.0 1163850.0 ;
      RECT  110100.0 1153350.0 111300.0 1154550.0 ;
      RECT  112500.0 1153350.0 113700.0 1154550.0 ;
      RECT  112500.0 1153350.0 113700.0 1154550.0 ;
      RECT  110100.0 1153350.0 111300.0 1154550.0 ;
      RECT  114900.0 1163250.0 116100.0 1164450.0 ;
      RECT  114900.0 1153350.0 116100.0 1154550.0 ;
      RECT  110700.0 1158000.0 111900.0 1159200.0 ;
      RECT  110700.0 1158000.0 111900.0 1159200.0 ;
      RECT  113250.0 1158150.0 114150.0 1159050.0 ;
      RECT  108300.0 1165350.0 117900.0 1166250.0 ;
      RECT  108300.0 1151550.0 117900.0 1152450.0 ;
      RECT  114900.0 1167750.0 116100.0 1165800.0 ;
      RECT  114900.0 1179600.0 116100.0 1177650.0 ;
      RECT  110100.0 1178250.0 111300.0 1180050.0 ;
      RECT  110100.0 1168950.0 111300.0 1165350.0 ;
      RECT  112800.0 1178250.0 113700.0 1168950.0 ;
      RECT  110100.0 1168950.0 111300.0 1167750.0 ;
      RECT  112500.0 1168950.0 113700.0 1167750.0 ;
      RECT  112500.0 1168950.0 113700.0 1167750.0 ;
      RECT  110100.0 1168950.0 111300.0 1167750.0 ;
      RECT  110100.0 1178250.0 111300.0 1177050.0 ;
      RECT  112500.0 1178250.0 113700.0 1177050.0 ;
      RECT  112500.0 1178250.0 113700.0 1177050.0 ;
      RECT  110100.0 1178250.0 111300.0 1177050.0 ;
      RECT  114900.0 1168350.0 116100.0 1167150.0 ;
      RECT  114900.0 1178250.0 116100.0 1177050.0 ;
      RECT  110700.0 1173600.0 111900.0 1172400.0 ;
      RECT  110700.0 1173600.0 111900.0 1172400.0 ;
      RECT  113250.0 1173450.0 114150.0 1172550.0 ;
      RECT  108300.0 1166250.0 117900.0 1165350.0 ;
      RECT  108300.0 1180050.0 117900.0 1179150.0 ;
      RECT  114900.0 1191450.0 116100.0 1193400.0 ;
      RECT  114900.0 1179600.0 116100.0 1181550.0 ;
      RECT  110100.0 1180950.0 111300.0 1179150.0 ;
      RECT  110100.0 1190250.0 111300.0 1193850.0 ;
      RECT  112800.0 1180950.0 113700.0 1190250.0 ;
      RECT  110100.0 1190250.0 111300.0 1191450.0 ;
      RECT  112500.0 1190250.0 113700.0 1191450.0 ;
      RECT  112500.0 1190250.0 113700.0 1191450.0 ;
      RECT  110100.0 1190250.0 111300.0 1191450.0 ;
      RECT  110100.0 1180950.0 111300.0 1182150.0 ;
      RECT  112500.0 1180950.0 113700.0 1182150.0 ;
      RECT  112500.0 1180950.0 113700.0 1182150.0 ;
      RECT  110100.0 1180950.0 111300.0 1182150.0 ;
      RECT  114900.0 1190850.0 116100.0 1192050.0 ;
      RECT  114900.0 1180950.0 116100.0 1182150.0 ;
      RECT  110700.0 1185600.0 111900.0 1186800.0 ;
      RECT  110700.0 1185600.0 111900.0 1186800.0 ;
      RECT  113250.0 1185750.0 114150.0 1186650.0 ;
      RECT  108300.0 1192950.0 117900.0 1193850.0 ;
      RECT  108300.0 1179150.0 117900.0 1180050.0 ;
      RECT  114900.0 1195350.0 116100.0 1193400.0 ;
      RECT  114900.0 1207200.0 116100.0 1205250.0 ;
      RECT  110100.0 1205850.0 111300.0 1207650.0 ;
      RECT  110100.0 1196550.0 111300.0 1192950.0 ;
      RECT  112800.0 1205850.0 113700.0 1196550.0 ;
      RECT  110100.0 1196550.0 111300.0 1195350.0 ;
      RECT  112500.0 1196550.0 113700.0 1195350.0 ;
      RECT  112500.0 1196550.0 113700.0 1195350.0 ;
      RECT  110100.0 1196550.0 111300.0 1195350.0 ;
      RECT  110100.0 1205850.0 111300.0 1204650.0 ;
      RECT  112500.0 1205850.0 113700.0 1204650.0 ;
      RECT  112500.0 1205850.0 113700.0 1204650.0 ;
      RECT  110100.0 1205850.0 111300.0 1204650.0 ;
      RECT  114900.0 1195950.0 116100.0 1194750.0 ;
      RECT  114900.0 1205850.0 116100.0 1204650.0 ;
      RECT  110700.0 1201200.0 111900.0 1200000.0 ;
      RECT  110700.0 1201200.0 111900.0 1200000.0 ;
      RECT  113250.0 1201050.0 114150.0 1200150.0 ;
      RECT  108300.0 1193850.0 117900.0 1192950.0 ;
      RECT  108300.0 1207650.0 117900.0 1206750.0 ;
      RECT  114900.0 1219050.0 116100.0 1221000.0 ;
      RECT  114900.0 1207200.0 116100.0 1209150.0 ;
      RECT  110100.0 1208550.0 111300.0 1206750.0 ;
      RECT  110100.0 1217850.0 111300.0 1221450.0 ;
      RECT  112800.0 1208550.0 113700.0 1217850.0 ;
      RECT  110100.0 1217850.0 111300.0 1219050.0 ;
      RECT  112500.0 1217850.0 113700.0 1219050.0 ;
      RECT  112500.0 1217850.0 113700.0 1219050.0 ;
      RECT  110100.0 1217850.0 111300.0 1219050.0 ;
      RECT  110100.0 1208550.0 111300.0 1209750.0 ;
      RECT  112500.0 1208550.0 113700.0 1209750.0 ;
      RECT  112500.0 1208550.0 113700.0 1209750.0 ;
      RECT  110100.0 1208550.0 111300.0 1209750.0 ;
      RECT  114900.0 1218450.0 116100.0 1219650.0 ;
      RECT  114900.0 1208550.0 116100.0 1209750.0 ;
      RECT  110700.0 1213200.0 111900.0 1214400.0 ;
      RECT  110700.0 1213200.0 111900.0 1214400.0 ;
      RECT  113250.0 1213350.0 114150.0 1214250.0 ;
      RECT  108300.0 1220550.0 117900.0 1221450.0 ;
      RECT  108300.0 1206750.0 117900.0 1207650.0 ;
      RECT  114900.0 1222950.0 116100.0 1221000.0 ;
      RECT  114900.0 1234800.0 116100.0 1232850.0 ;
      RECT  110100.0 1233450.0 111300.0 1235250.0 ;
      RECT  110100.0 1224150.0 111300.0 1220550.0 ;
      RECT  112800.0 1233450.0 113700.0 1224150.0 ;
      RECT  110100.0 1224150.0 111300.0 1222950.0 ;
      RECT  112500.0 1224150.0 113700.0 1222950.0 ;
      RECT  112500.0 1224150.0 113700.0 1222950.0 ;
      RECT  110100.0 1224150.0 111300.0 1222950.0 ;
      RECT  110100.0 1233450.0 111300.0 1232250.0 ;
      RECT  112500.0 1233450.0 113700.0 1232250.0 ;
      RECT  112500.0 1233450.0 113700.0 1232250.0 ;
      RECT  110100.0 1233450.0 111300.0 1232250.0 ;
      RECT  114900.0 1223550.0 116100.0 1222350.0 ;
      RECT  114900.0 1233450.0 116100.0 1232250.0 ;
      RECT  110700.0 1228800.0 111900.0 1227600.0 ;
      RECT  110700.0 1228800.0 111900.0 1227600.0 ;
      RECT  113250.0 1228650.0 114150.0 1227750.0 ;
      RECT  108300.0 1221450.0 117900.0 1220550.0 ;
      RECT  108300.0 1235250.0 117900.0 1234350.0 ;
      RECT  114900.0 1246650.0 116100.0 1248600.0 ;
      RECT  114900.0 1234800.0 116100.0 1236750.0 ;
      RECT  110100.0 1236150.0 111300.0 1234350.0 ;
      RECT  110100.0 1245450.0 111300.0 1249050.0 ;
      RECT  112800.0 1236150.0 113700.0 1245450.0 ;
      RECT  110100.0 1245450.0 111300.0 1246650.0 ;
      RECT  112500.0 1245450.0 113700.0 1246650.0 ;
      RECT  112500.0 1245450.0 113700.0 1246650.0 ;
      RECT  110100.0 1245450.0 111300.0 1246650.0 ;
      RECT  110100.0 1236150.0 111300.0 1237350.0 ;
      RECT  112500.0 1236150.0 113700.0 1237350.0 ;
      RECT  112500.0 1236150.0 113700.0 1237350.0 ;
      RECT  110100.0 1236150.0 111300.0 1237350.0 ;
      RECT  114900.0 1246050.0 116100.0 1247250.0 ;
      RECT  114900.0 1236150.0 116100.0 1237350.0 ;
      RECT  110700.0 1240800.0 111900.0 1242000.0 ;
      RECT  110700.0 1240800.0 111900.0 1242000.0 ;
      RECT  113250.0 1240950.0 114150.0 1241850.0 ;
      RECT  108300.0 1248150.0 117900.0 1249050.0 ;
      RECT  108300.0 1234350.0 117900.0 1235250.0 ;
      RECT  114900.0 1250550.0 116100.0 1248600.0 ;
      RECT  114900.0 1262400.0 116100.0 1260450.0 ;
      RECT  110100.0 1261050.0 111300.0 1262850.0 ;
      RECT  110100.0 1251750.0 111300.0 1248150.0 ;
      RECT  112800.0 1261050.0 113700.0 1251750.0 ;
      RECT  110100.0 1251750.0 111300.0 1250550.0 ;
      RECT  112500.0 1251750.0 113700.0 1250550.0 ;
      RECT  112500.0 1251750.0 113700.0 1250550.0 ;
      RECT  110100.0 1251750.0 111300.0 1250550.0 ;
      RECT  110100.0 1261050.0 111300.0 1259850.0 ;
      RECT  112500.0 1261050.0 113700.0 1259850.0 ;
      RECT  112500.0 1261050.0 113700.0 1259850.0 ;
      RECT  110100.0 1261050.0 111300.0 1259850.0 ;
      RECT  114900.0 1251150.0 116100.0 1249950.0 ;
      RECT  114900.0 1261050.0 116100.0 1259850.0 ;
      RECT  110700.0 1256400.0 111900.0 1255200.0 ;
      RECT  110700.0 1256400.0 111900.0 1255200.0 ;
      RECT  113250.0 1256250.0 114150.0 1255350.0 ;
      RECT  108300.0 1249050.0 117900.0 1248150.0 ;
      RECT  108300.0 1262850.0 117900.0 1261950.0 ;
      RECT  114900.0 1274250.0 116100.0 1276200.0 ;
      RECT  114900.0 1262400.0 116100.0 1264350.0 ;
      RECT  110100.0 1263750.0 111300.0 1261950.0 ;
      RECT  110100.0 1273050.0 111300.0 1276650.0 ;
      RECT  112800.0 1263750.0 113700.0 1273050.0 ;
      RECT  110100.0 1273050.0 111300.0 1274250.0 ;
      RECT  112500.0 1273050.0 113700.0 1274250.0 ;
      RECT  112500.0 1273050.0 113700.0 1274250.0 ;
      RECT  110100.0 1273050.0 111300.0 1274250.0 ;
      RECT  110100.0 1263750.0 111300.0 1264950.0 ;
      RECT  112500.0 1263750.0 113700.0 1264950.0 ;
      RECT  112500.0 1263750.0 113700.0 1264950.0 ;
      RECT  110100.0 1263750.0 111300.0 1264950.0 ;
      RECT  114900.0 1273650.0 116100.0 1274850.0 ;
      RECT  114900.0 1263750.0 116100.0 1264950.0 ;
      RECT  110700.0 1268400.0 111900.0 1269600.0 ;
      RECT  110700.0 1268400.0 111900.0 1269600.0 ;
      RECT  113250.0 1268550.0 114150.0 1269450.0 ;
      RECT  108300.0 1275750.0 117900.0 1276650.0 ;
      RECT  108300.0 1261950.0 117900.0 1262850.0 ;
      RECT  114900.0 1278150.0 116100.0 1276200.0 ;
      RECT  114900.0 1290000.0 116100.0 1288050.0 ;
      RECT  110100.0 1288650.0 111300.0 1290450.0 ;
      RECT  110100.0 1279350.0 111300.0 1275750.0 ;
      RECT  112800.0 1288650.0 113700.0 1279350.0 ;
      RECT  110100.0 1279350.0 111300.0 1278150.0 ;
      RECT  112500.0 1279350.0 113700.0 1278150.0 ;
      RECT  112500.0 1279350.0 113700.0 1278150.0 ;
      RECT  110100.0 1279350.0 111300.0 1278150.0 ;
      RECT  110100.0 1288650.0 111300.0 1287450.0 ;
      RECT  112500.0 1288650.0 113700.0 1287450.0 ;
      RECT  112500.0 1288650.0 113700.0 1287450.0 ;
      RECT  110100.0 1288650.0 111300.0 1287450.0 ;
      RECT  114900.0 1278750.0 116100.0 1277550.0 ;
      RECT  114900.0 1288650.0 116100.0 1287450.0 ;
      RECT  110700.0 1284000.0 111900.0 1282800.0 ;
      RECT  110700.0 1284000.0 111900.0 1282800.0 ;
      RECT  113250.0 1283850.0 114150.0 1282950.0 ;
      RECT  108300.0 1276650.0 117900.0 1275750.0 ;
      RECT  108300.0 1290450.0 117900.0 1289550.0 ;
      RECT  114900.0 1301850.0 116100.0 1303800.0 ;
      RECT  114900.0 1290000.0 116100.0 1291950.0 ;
      RECT  110100.0 1291350.0 111300.0 1289550.0 ;
      RECT  110100.0 1300650.0 111300.0 1304250.0 ;
      RECT  112800.0 1291350.0 113700.0 1300650.0 ;
      RECT  110100.0 1300650.0 111300.0 1301850.0 ;
      RECT  112500.0 1300650.0 113700.0 1301850.0 ;
      RECT  112500.0 1300650.0 113700.0 1301850.0 ;
      RECT  110100.0 1300650.0 111300.0 1301850.0 ;
      RECT  110100.0 1291350.0 111300.0 1292550.0 ;
      RECT  112500.0 1291350.0 113700.0 1292550.0 ;
      RECT  112500.0 1291350.0 113700.0 1292550.0 ;
      RECT  110100.0 1291350.0 111300.0 1292550.0 ;
      RECT  114900.0 1301250.0 116100.0 1302450.0 ;
      RECT  114900.0 1291350.0 116100.0 1292550.0 ;
      RECT  110700.0 1296000.0 111900.0 1297200.0 ;
      RECT  110700.0 1296000.0 111900.0 1297200.0 ;
      RECT  113250.0 1296150.0 114150.0 1297050.0 ;
      RECT  108300.0 1303350.0 117900.0 1304250.0 ;
      RECT  108300.0 1289550.0 117900.0 1290450.0 ;
      RECT  114900.0 1305750.0 116100.0 1303800.0 ;
      RECT  114900.0 1317600.0 116100.0 1315650.0 ;
      RECT  110100.0 1316250.0 111300.0 1318050.0 ;
      RECT  110100.0 1306950.0 111300.0 1303350.0 ;
      RECT  112800.0 1316250.0 113700.0 1306950.0 ;
      RECT  110100.0 1306950.0 111300.0 1305750.0 ;
      RECT  112500.0 1306950.0 113700.0 1305750.0 ;
      RECT  112500.0 1306950.0 113700.0 1305750.0 ;
      RECT  110100.0 1306950.0 111300.0 1305750.0 ;
      RECT  110100.0 1316250.0 111300.0 1315050.0 ;
      RECT  112500.0 1316250.0 113700.0 1315050.0 ;
      RECT  112500.0 1316250.0 113700.0 1315050.0 ;
      RECT  110100.0 1316250.0 111300.0 1315050.0 ;
      RECT  114900.0 1306350.0 116100.0 1305150.0 ;
      RECT  114900.0 1316250.0 116100.0 1315050.0 ;
      RECT  110700.0 1311600.0 111900.0 1310400.0 ;
      RECT  110700.0 1311600.0 111900.0 1310400.0 ;
      RECT  113250.0 1311450.0 114150.0 1310550.0 ;
      RECT  108300.0 1304250.0 117900.0 1303350.0 ;
      RECT  108300.0 1318050.0 117900.0 1317150.0 ;
      RECT  114900.0 1329450.0 116100.0 1331400.0 ;
      RECT  114900.0 1317600.0 116100.0 1319550.0 ;
      RECT  110100.0 1318950.0 111300.0 1317150.0 ;
      RECT  110100.0 1328250.0 111300.0 1331850.0 ;
      RECT  112800.0 1318950.0 113700.0 1328250.0 ;
      RECT  110100.0 1328250.0 111300.0 1329450.0 ;
      RECT  112500.0 1328250.0 113700.0 1329450.0 ;
      RECT  112500.0 1328250.0 113700.0 1329450.0 ;
      RECT  110100.0 1328250.0 111300.0 1329450.0 ;
      RECT  110100.0 1318950.0 111300.0 1320150.0 ;
      RECT  112500.0 1318950.0 113700.0 1320150.0 ;
      RECT  112500.0 1318950.0 113700.0 1320150.0 ;
      RECT  110100.0 1318950.0 111300.0 1320150.0 ;
      RECT  114900.0 1328850.0 116100.0 1330050.0 ;
      RECT  114900.0 1318950.0 116100.0 1320150.0 ;
      RECT  110700.0 1323600.0 111900.0 1324800.0 ;
      RECT  110700.0 1323600.0 111900.0 1324800.0 ;
      RECT  113250.0 1323750.0 114150.0 1324650.0 ;
      RECT  108300.0 1330950.0 117900.0 1331850.0 ;
      RECT  108300.0 1317150.0 117900.0 1318050.0 ;
      RECT  114900.0 1333350.0 116100.0 1331400.0 ;
      RECT  114900.0 1345200.0 116100.0 1343250.0 ;
      RECT  110100.0 1343850.0 111300.0 1345650.0 ;
      RECT  110100.0 1334550.0 111300.0 1330950.0 ;
      RECT  112800.0 1343850.0 113700.0 1334550.0 ;
      RECT  110100.0 1334550.0 111300.0 1333350.0 ;
      RECT  112500.0 1334550.0 113700.0 1333350.0 ;
      RECT  112500.0 1334550.0 113700.0 1333350.0 ;
      RECT  110100.0 1334550.0 111300.0 1333350.0 ;
      RECT  110100.0 1343850.0 111300.0 1342650.0 ;
      RECT  112500.0 1343850.0 113700.0 1342650.0 ;
      RECT  112500.0 1343850.0 113700.0 1342650.0 ;
      RECT  110100.0 1343850.0 111300.0 1342650.0 ;
      RECT  114900.0 1333950.0 116100.0 1332750.0 ;
      RECT  114900.0 1343850.0 116100.0 1342650.0 ;
      RECT  110700.0 1339200.0 111900.0 1338000.0 ;
      RECT  110700.0 1339200.0 111900.0 1338000.0 ;
      RECT  113250.0 1339050.0 114150.0 1338150.0 ;
      RECT  108300.0 1331850.0 117900.0 1330950.0 ;
      RECT  108300.0 1345650.0 117900.0 1344750.0 ;
      RECT  114900.0 1357050.0 116100.0 1359000.0 ;
      RECT  114900.0 1345200.0 116100.0 1347150.0 ;
      RECT  110100.0 1346550.0 111300.0 1344750.0 ;
      RECT  110100.0 1355850.0 111300.0 1359450.0 ;
      RECT  112800.0 1346550.0 113700.0 1355850.0 ;
      RECT  110100.0 1355850.0 111300.0 1357050.0 ;
      RECT  112500.0 1355850.0 113700.0 1357050.0 ;
      RECT  112500.0 1355850.0 113700.0 1357050.0 ;
      RECT  110100.0 1355850.0 111300.0 1357050.0 ;
      RECT  110100.0 1346550.0 111300.0 1347750.0 ;
      RECT  112500.0 1346550.0 113700.0 1347750.0 ;
      RECT  112500.0 1346550.0 113700.0 1347750.0 ;
      RECT  110100.0 1346550.0 111300.0 1347750.0 ;
      RECT  114900.0 1356450.0 116100.0 1357650.0 ;
      RECT  114900.0 1346550.0 116100.0 1347750.0 ;
      RECT  110700.0 1351200.0 111900.0 1352400.0 ;
      RECT  110700.0 1351200.0 111900.0 1352400.0 ;
      RECT  113250.0 1351350.0 114150.0 1352250.0 ;
      RECT  108300.0 1358550.0 117900.0 1359450.0 ;
      RECT  108300.0 1344750.0 117900.0 1345650.0 ;
      RECT  114900.0 1360950.0 116100.0 1359000.0 ;
      RECT  114900.0 1372800.0 116100.0 1370850.0 ;
      RECT  110100.0 1371450.0 111300.0 1373250.0 ;
      RECT  110100.0 1362150.0 111300.0 1358550.0 ;
      RECT  112800.0 1371450.0 113700.0 1362150.0 ;
      RECT  110100.0 1362150.0 111300.0 1360950.0 ;
      RECT  112500.0 1362150.0 113700.0 1360950.0 ;
      RECT  112500.0 1362150.0 113700.0 1360950.0 ;
      RECT  110100.0 1362150.0 111300.0 1360950.0 ;
      RECT  110100.0 1371450.0 111300.0 1370250.0 ;
      RECT  112500.0 1371450.0 113700.0 1370250.0 ;
      RECT  112500.0 1371450.0 113700.0 1370250.0 ;
      RECT  110100.0 1371450.0 111300.0 1370250.0 ;
      RECT  114900.0 1361550.0 116100.0 1360350.0 ;
      RECT  114900.0 1371450.0 116100.0 1370250.0 ;
      RECT  110700.0 1366800.0 111900.0 1365600.0 ;
      RECT  110700.0 1366800.0 111900.0 1365600.0 ;
      RECT  113250.0 1366650.0 114150.0 1365750.0 ;
      RECT  108300.0 1359450.0 117900.0 1358550.0 ;
      RECT  108300.0 1373250.0 117900.0 1372350.0 ;
      RECT  114900.0 1384650.0 116100.0 1386600.0 ;
      RECT  114900.0 1372800.0 116100.0 1374750.0 ;
      RECT  110100.0 1374150.0 111300.0 1372350.0 ;
      RECT  110100.0 1383450.0 111300.0 1387050.0 ;
      RECT  112800.0 1374150.0 113700.0 1383450.0 ;
      RECT  110100.0 1383450.0 111300.0 1384650.0 ;
      RECT  112500.0 1383450.0 113700.0 1384650.0 ;
      RECT  112500.0 1383450.0 113700.0 1384650.0 ;
      RECT  110100.0 1383450.0 111300.0 1384650.0 ;
      RECT  110100.0 1374150.0 111300.0 1375350.0 ;
      RECT  112500.0 1374150.0 113700.0 1375350.0 ;
      RECT  112500.0 1374150.0 113700.0 1375350.0 ;
      RECT  110100.0 1374150.0 111300.0 1375350.0 ;
      RECT  114900.0 1384050.0 116100.0 1385250.0 ;
      RECT  114900.0 1374150.0 116100.0 1375350.0 ;
      RECT  110700.0 1378800.0 111900.0 1380000.0 ;
      RECT  110700.0 1378800.0 111900.0 1380000.0 ;
      RECT  113250.0 1378950.0 114150.0 1379850.0 ;
      RECT  108300.0 1386150.0 117900.0 1387050.0 ;
      RECT  108300.0 1372350.0 117900.0 1373250.0 ;
      RECT  114900.0 1388550.0 116100.0 1386600.0 ;
      RECT  114900.0 1400400.0 116100.0 1398450.0 ;
      RECT  110100.0 1399050.0 111300.0 1400850.0 ;
      RECT  110100.0 1389750.0 111300.0 1386150.0 ;
      RECT  112800.0 1399050.0 113700.0 1389750.0 ;
      RECT  110100.0 1389750.0 111300.0 1388550.0 ;
      RECT  112500.0 1389750.0 113700.0 1388550.0 ;
      RECT  112500.0 1389750.0 113700.0 1388550.0 ;
      RECT  110100.0 1389750.0 111300.0 1388550.0 ;
      RECT  110100.0 1399050.0 111300.0 1397850.0 ;
      RECT  112500.0 1399050.0 113700.0 1397850.0 ;
      RECT  112500.0 1399050.0 113700.0 1397850.0 ;
      RECT  110100.0 1399050.0 111300.0 1397850.0 ;
      RECT  114900.0 1389150.0 116100.0 1387950.0 ;
      RECT  114900.0 1399050.0 116100.0 1397850.0 ;
      RECT  110700.0 1394400.0 111900.0 1393200.0 ;
      RECT  110700.0 1394400.0 111900.0 1393200.0 ;
      RECT  113250.0 1394250.0 114150.0 1393350.0 ;
      RECT  108300.0 1387050.0 117900.0 1386150.0 ;
      RECT  108300.0 1400850.0 117900.0 1399950.0 ;
      RECT  114900.0 1412250.0 116100.0 1414200.0 ;
      RECT  114900.0 1400400.0 116100.0 1402350.0 ;
      RECT  110100.0 1401750.0 111300.0 1399950.0 ;
      RECT  110100.0 1411050.0 111300.0 1414650.0 ;
      RECT  112800.0 1401750.0 113700.0 1411050.0 ;
      RECT  110100.0 1411050.0 111300.0 1412250.0 ;
      RECT  112500.0 1411050.0 113700.0 1412250.0 ;
      RECT  112500.0 1411050.0 113700.0 1412250.0 ;
      RECT  110100.0 1411050.0 111300.0 1412250.0 ;
      RECT  110100.0 1401750.0 111300.0 1402950.0 ;
      RECT  112500.0 1401750.0 113700.0 1402950.0 ;
      RECT  112500.0 1401750.0 113700.0 1402950.0 ;
      RECT  110100.0 1401750.0 111300.0 1402950.0 ;
      RECT  114900.0 1411650.0 116100.0 1412850.0 ;
      RECT  114900.0 1401750.0 116100.0 1402950.0 ;
      RECT  110700.0 1406400.0 111900.0 1407600.0 ;
      RECT  110700.0 1406400.0 111900.0 1407600.0 ;
      RECT  113250.0 1406550.0 114150.0 1407450.0 ;
      RECT  108300.0 1413750.0 117900.0 1414650.0 ;
      RECT  108300.0 1399950.0 117900.0 1400850.0 ;
      RECT  114900.0 1416150.0 116100.0 1414200.0 ;
      RECT  114900.0 1428000.0 116100.0 1426050.0 ;
      RECT  110100.0 1426650.0 111300.0 1428450.0 ;
      RECT  110100.0 1417350.0 111300.0 1413750.0 ;
      RECT  112800.0 1426650.0 113700.0 1417350.0 ;
      RECT  110100.0 1417350.0 111300.0 1416150.0 ;
      RECT  112500.0 1417350.0 113700.0 1416150.0 ;
      RECT  112500.0 1417350.0 113700.0 1416150.0 ;
      RECT  110100.0 1417350.0 111300.0 1416150.0 ;
      RECT  110100.0 1426650.0 111300.0 1425450.0 ;
      RECT  112500.0 1426650.0 113700.0 1425450.0 ;
      RECT  112500.0 1426650.0 113700.0 1425450.0 ;
      RECT  110100.0 1426650.0 111300.0 1425450.0 ;
      RECT  114900.0 1416750.0 116100.0 1415550.0 ;
      RECT  114900.0 1426650.0 116100.0 1425450.0 ;
      RECT  110700.0 1422000.0 111900.0 1420800.0 ;
      RECT  110700.0 1422000.0 111900.0 1420800.0 ;
      RECT  113250.0 1421850.0 114150.0 1420950.0 ;
      RECT  108300.0 1414650.0 117900.0 1413750.0 ;
      RECT  108300.0 1428450.0 117900.0 1427550.0 ;
      RECT  114900.0 1439850.0 116100.0 1441800.0 ;
      RECT  114900.0 1428000.0 116100.0 1429950.0 ;
      RECT  110100.0 1429350.0 111300.0 1427550.0 ;
      RECT  110100.0 1438650.0 111300.0 1442250.0 ;
      RECT  112800.0 1429350.0 113700.0 1438650.0 ;
      RECT  110100.0 1438650.0 111300.0 1439850.0 ;
      RECT  112500.0 1438650.0 113700.0 1439850.0 ;
      RECT  112500.0 1438650.0 113700.0 1439850.0 ;
      RECT  110100.0 1438650.0 111300.0 1439850.0 ;
      RECT  110100.0 1429350.0 111300.0 1430550.0 ;
      RECT  112500.0 1429350.0 113700.0 1430550.0 ;
      RECT  112500.0 1429350.0 113700.0 1430550.0 ;
      RECT  110100.0 1429350.0 111300.0 1430550.0 ;
      RECT  114900.0 1439250.0 116100.0 1440450.0 ;
      RECT  114900.0 1429350.0 116100.0 1430550.0 ;
      RECT  110700.0 1434000.0 111900.0 1435200.0 ;
      RECT  110700.0 1434000.0 111900.0 1435200.0 ;
      RECT  113250.0 1434150.0 114150.0 1435050.0 ;
      RECT  108300.0 1441350.0 117900.0 1442250.0 ;
      RECT  108300.0 1427550.0 117900.0 1428450.0 ;
      RECT  114900.0 1443750.0 116100.0 1441800.0 ;
      RECT  114900.0 1455600.0 116100.0 1453650.0 ;
      RECT  110100.0 1454250.0 111300.0 1456050.0 ;
      RECT  110100.0 1444950.0 111300.0 1441350.0 ;
      RECT  112800.0 1454250.0 113700.0 1444950.0 ;
      RECT  110100.0 1444950.0 111300.0 1443750.0 ;
      RECT  112500.0 1444950.0 113700.0 1443750.0 ;
      RECT  112500.0 1444950.0 113700.0 1443750.0 ;
      RECT  110100.0 1444950.0 111300.0 1443750.0 ;
      RECT  110100.0 1454250.0 111300.0 1453050.0 ;
      RECT  112500.0 1454250.0 113700.0 1453050.0 ;
      RECT  112500.0 1454250.0 113700.0 1453050.0 ;
      RECT  110100.0 1454250.0 111300.0 1453050.0 ;
      RECT  114900.0 1444350.0 116100.0 1443150.0 ;
      RECT  114900.0 1454250.0 116100.0 1453050.0 ;
      RECT  110700.0 1449600.0 111900.0 1448400.0 ;
      RECT  110700.0 1449600.0 111900.0 1448400.0 ;
      RECT  113250.0 1449450.0 114150.0 1448550.0 ;
      RECT  108300.0 1442250.0 117900.0 1441350.0 ;
      RECT  108300.0 1456050.0 117900.0 1455150.0 ;
      RECT  114900.0 1467450.0 116100.0 1469400.0 ;
      RECT  114900.0 1455600.0 116100.0 1457550.0 ;
      RECT  110100.0 1456950.0 111300.0 1455150.0 ;
      RECT  110100.0 1466250.0 111300.0 1469850.0 ;
      RECT  112800.0 1456950.0 113700.0 1466250.0 ;
      RECT  110100.0 1466250.0 111300.0 1467450.0 ;
      RECT  112500.0 1466250.0 113700.0 1467450.0 ;
      RECT  112500.0 1466250.0 113700.0 1467450.0 ;
      RECT  110100.0 1466250.0 111300.0 1467450.0 ;
      RECT  110100.0 1456950.0 111300.0 1458150.0 ;
      RECT  112500.0 1456950.0 113700.0 1458150.0 ;
      RECT  112500.0 1456950.0 113700.0 1458150.0 ;
      RECT  110100.0 1456950.0 111300.0 1458150.0 ;
      RECT  114900.0 1466850.0 116100.0 1468050.0 ;
      RECT  114900.0 1456950.0 116100.0 1458150.0 ;
      RECT  110700.0 1461600.0 111900.0 1462800.0 ;
      RECT  110700.0 1461600.0 111900.0 1462800.0 ;
      RECT  113250.0 1461750.0 114150.0 1462650.0 ;
      RECT  108300.0 1468950.0 117900.0 1469850.0 ;
      RECT  108300.0 1455150.0 117900.0 1456050.0 ;
      RECT  114900.0 1471350.0 116100.0 1469400.0 ;
      RECT  114900.0 1483200.0 116100.0 1481250.0 ;
      RECT  110100.0 1481850.0 111300.0 1483650.0 ;
      RECT  110100.0 1472550.0 111300.0 1468950.0 ;
      RECT  112800.0 1481850.0 113700.0 1472550.0 ;
      RECT  110100.0 1472550.0 111300.0 1471350.0 ;
      RECT  112500.0 1472550.0 113700.0 1471350.0 ;
      RECT  112500.0 1472550.0 113700.0 1471350.0 ;
      RECT  110100.0 1472550.0 111300.0 1471350.0 ;
      RECT  110100.0 1481850.0 111300.0 1480650.0 ;
      RECT  112500.0 1481850.0 113700.0 1480650.0 ;
      RECT  112500.0 1481850.0 113700.0 1480650.0 ;
      RECT  110100.0 1481850.0 111300.0 1480650.0 ;
      RECT  114900.0 1471950.0 116100.0 1470750.0 ;
      RECT  114900.0 1481850.0 116100.0 1480650.0 ;
      RECT  110700.0 1477200.0 111900.0 1476000.0 ;
      RECT  110700.0 1477200.0 111900.0 1476000.0 ;
      RECT  113250.0 1477050.0 114150.0 1476150.0 ;
      RECT  108300.0 1469850.0 117900.0 1468950.0 ;
      RECT  108300.0 1483650.0 117900.0 1482750.0 ;
      RECT  114900.0 1495050.0 116100.0 1497000.0 ;
      RECT  114900.0 1483200.0 116100.0 1485150.0 ;
      RECT  110100.0 1484550.0 111300.0 1482750.0 ;
      RECT  110100.0 1493850.0 111300.0 1497450.0 ;
      RECT  112800.0 1484550.0 113700.0 1493850.0 ;
      RECT  110100.0 1493850.0 111300.0 1495050.0 ;
      RECT  112500.0 1493850.0 113700.0 1495050.0 ;
      RECT  112500.0 1493850.0 113700.0 1495050.0 ;
      RECT  110100.0 1493850.0 111300.0 1495050.0 ;
      RECT  110100.0 1484550.0 111300.0 1485750.0 ;
      RECT  112500.0 1484550.0 113700.0 1485750.0 ;
      RECT  112500.0 1484550.0 113700.0 1485750.0 ;
      RECT  110100.0 1484550.0 111300.0 1485750.0 ;
      RECT  114900.0 1494450.0 116100.0 1495650.0 ;
      RECT  114900.0 1484550.0 116100.0 1485750.0 ;
      RECT  110700.0 1489200.0 111900.0 1490400.0 ;
      RECT  110700.0 1489200.0 111900.0 1490400.0 ;
      RECT  113250.0 1489350.0 114150.0 1490250.0 ;
      RECT  108300.0 1496550.0 117900.0 1497450.0 ;
      RECT  108300.0 1482750.0 117900.0 1483650.0 ;
      RECT  114900.0 1498950.0 116100.0 1497000.0 ;
      RECT  114900.0 1510800.0 116100.0 1508850.0 ;
      RECT  110100.0 1509450.0 111300.0 1511250.0 ;
      RECT  110100.0 1500150.0 111300.0 1496550.0 ;
      RECT  112800.0 1509450.0 113700.0 1500150.0 ;
      RECT  110100.0 1500150.0 111300.0 1498950.0 ;
      RECT  112500.0 1500150.0 113700.0 1498950.0 ;
      RECT  112500.0 1500150.0 113700.0 1498950.0 ;
      RECT  110100.0 1500150.0 111300.0 1498950.0 ;
      RECT  110100.0 1509450.0 111300.0 1508250.0 ;
      RECT  112500.0 1509450.0 113700.0 1508250.0 ;
      RECT  112500.0 1509450.0 113700.0 1508250.0 ;
      RECT  110100.0 1509450.0 111300.0 1508250.0 ;
      RECT  114900.0 1499550.0 116100.0 1498350.0 ;
      RECT  114900.0 1509450.0 116100.0 1508250.0 ;
      RECT  110700.0 1504800.0 111900.0 1503600.0 ;
      RECT  110700.0 1504800.0 111900.0 1503600.0 ;
      RECT  113250.0 1504650.0 114150.0 1503750.0 ;
      RECT  108300.0 1497450.0 117900.0 1496550.0 ;
      RECT  108300.0 1511250.0 117900.0 1510350.0 ;
      RECT  114900.0 1522650.0 116100.0 1524600.0 ;
      RECT  114900.0 1510800.0 116100.0 1512750.0 ;
      RECT  110100.0 1512150.0 111300.0 1510350.0 ;
      RECT  110100.0 1521450.0 111300.0 1525050.0 ;
      RECT  112800.0 1512150.0 113700.0 1521450.0 ;
      RECT  110100.0 1521450.0 111300.0 1522650.0 ;
      RECT  112500.0 1521450.0 113700.0 1522650.0 ;
      RECT  112500.0 1521450.0 113700.0 1522650.0 ;
      RECT  110100.0 1521450.0 111300.0 1522650.0 ;
      RECT  110100.0 1512150.0 111300.0 1513350.0 ;
      RECT  112500.0 1512150.0 113700.0 1513350.0 ;
      RECT  112500.0 1512150.0 113700.0 1513350.0 ;
      RECT  110100.0 1512150.0 111300.0 1513350.0 ;
      RECT  114900.0 1522050.0 116100.0 1523250.0 ;
      RECT  114900.0 1512150.0 116100.0 1513350.0 ;
      RECT  110700.0 1516800.0 111900.0 1518000.0 ;
      RECT  110700.0 1516800.0 111900.0 1518000.0 ;
      RECT  113250.0 1516950.0 114150.0 1517850.0 ;
      RECT  108300.0 1524150.0 117900.0 1525050.0 ;
      RECT  108300.0 1510350.0 117900.0 1511250.0 ;
      RECT  114900.0 1526550.0 116100.0 1524600.0 ;
      RECT  114900.0 1538400.0 116100.0 1536450.0 ;
      RECT  110100.0 1537050.0 111300.0 1538850.0 ;
      RECT  110100.0 1527750.0 111300.0 1524150.0 ;
      RECT  112800.0 1537050.0 113700.0 1527750.0 ;
      RECT  110100.0 1527750.0 111300.0 1526550.0 ;
      RECT  112500.0 1527750.0 113700.0 1526550.0 ;
      RECT  112500.0 1527750.0 113700.0 1526550.0 ;
      RECT  110100.0 1527750.0 111300.0 1526550.0 ;
      RECT  110100.0 1537050.0 111300.0 1535850.0 ;
      RECT  112500.0 1537050.0 113700.0 1535850.0 ;
      RECT  112500.0 1537050.0 113700.0 1535850.0 ;
      RECT  110100.0 1537050.0 111300.0 1535850.0 ;
      RECT  114900.0 1527150.0 116100.0 1525950.0 ;
      RECT  114900.0 1537050.0 116100.0 1535850.0 ;
      RECT  110700.0 1532400.0 111900.0 1531200.0 ;
      RECT  110700.0 1532400.0 111900.0 1531200.0 ;
      RECT  113250.0 1532250.0 114150.0 1531350.0 ;
      RECT  108300.0 1525050.0 117900.0 1524150.0 ;
      RECT  108300.0 1538850.0 117900.0 1537950.0 ;
      RECT  114900.0 1550250.0 116100.0 1552200.0 ;
      RECT  114900.0 1538400.0 116100.0 1540350.0 ;
      RECT  110100.0 1539750.0 111300.0 1537950.0 ;
      RECT  110100.0 1549050.0 111300.0 1552650.0 ;
      RECT  112800.0 1539750.0 113700.0 1549050.0 ;
      RECT  110100.0 1549050.0 111300.0 1550250.0 ;
      RECT  112500.0 1549050.0 113700.0 1550250.0 ;
      RECT  112500.0 1549050.0 113700.0 1550250.0 ;
      RECT  110100.0 1549050.0 111300.0 1550250.0 ;
      RECT  110100.0 1539750.0 111300.0 1540950.0 ;
      RECT  112500.0 1539750.0 113700.0 1540950.0 ;
      RECT  112500.0 1539750.0 113700.0 1540950.0 ;
      RECT  110100.0 1539750.0 111300.0 1540950.0 ;
      RECT  114900.0 1549650.0 116100.0 1550850.0 ;
      RECT  114900.0 1539750.0 116100.0 1540950.0 ;
      RECT  110700.0 1544400.0 111900.0 1545600.0 ;
      RECT  110700.0 1544400.0 111900.0 1545600.0 ;
      RECT  113250.0 1544550.0 114150.0 1545450.0 ;
      RECT  108300.0 1551750.0 117900.0 1552650.0 ;
      RECT  108300.0 1537950.0 117900.0 1538850.0 ;
      RECT  114900.0 1554150.0 116100.0 1552200.0 ;
      RECT  114900.0 1566000.0 116100.0 1564050.0 ;
      RECT  110100.0 1564650.0 111300.0 1566450.0 ;
      RECT  110100.0 1555350.0 111300.0 1551750.0 ;
      RECT  112800.0 1564650.0 113700.0 1555350.0 ;
      RECT  110100.0 1555350.0 111300.0 1554150.0 ;
      RECT  112500.0 1555350.0 113700.0 1554150.0 ;
      RECT  112500.0 1555350.0 113700.0 1554150.0 ;
      RECT  110100.0 1555350.0 111300.0 1554150.0 ;
      RECT  110100.0 1564650.0 111300.0 1563450.0 ;
      RECT  112500.0 1564650.0 113700.0 1563450.0 ;
      RECT  112500.0 1564650.0 113700.0 1563450.0 ;
      RECT  110100.0 1564650.0 111300.0 1563450.0 ;
      RECT  114900.0 1554750.0 116100.0 1553550.0 ;
      RECT  114900.0 1564650.0 116100.0 1563450.0 ;
      RECT  110700.0 1560000.0 111900.0 1558800.0 ;
      RECT  110700.0 1560000.0 111900.0 1558800.0 ;
      RECT  113250.0 1559850.0 114150.0 1558950.0 ;
      RECT  108300.0 1552650.0 117900.0 1551750.0 ;
      RECT  108300.0 1566450.0 117900.0 1565550.0 ;
      RECT  114900.0 1577850.0 116100.0 1579800.0 ;
      RECT  114900.0 1566000.0 116100.0 1567950.0 ;
      RECT  110100.0 1567350.0 111300.0 1565550.0 ;
      RECT  110100.0 1576650.0 111300.0 1580250.0 ;
      RECT  112800.0 1567350.0 113700.0 1576650.0 ;
      RECT  110100.0 1576650.0 111300.0 1577850.0 ;
      RECT  112500.0 1576650.0 113700.0 1577850.0 ;
      RECT  112500.0 1576650.0 113700.0 1577850.0 ;
      RECT  110100.0 1576650.0 111300.0 1577850.0 ;
      RECT  110100.0 1567350.0 111300.0 1568550.0 ;
      RECT  112500.0 1567350.0 113700.0 1568550.0 ;
      RECT  112500.0 1567350.0 113700.0 1568550.0 ;
      RECT  110100.0 1567350.0 111300.0 1568550.0 ;
      RECT  114900.0 1577250.0 116100.0 1578450.0 ;
      RECT  114900.0 1567350.0 116100.0 1568550.0 ;
      RECT  110700.0 1572000.0 111900.0 1573200.0 ;
      RECT  110700.0 1572000.0 111900.0 1573200.0 ;
      RECT  113250.0 1572150.0 114150.0 1573050.0 ;
      RECT  108300.0 1579350.0 117900.0 1580250.0 ;
      RECT  108300.0 1565550.0 117900.0 1566450.0 ;
      RECT  114900.0 1581750.0 116100.0 1579800.0 ;
      RECT  114900.0 1593600.0 116100.0 1591650.0 ;
      RECT  110100.0 1592250.0 111300.0 1594050.0 ;
      RECT  110100.0 1582950.0 111300.0 1579350.0 ;
      RECT  112800.0 1592250.0 113700.0 1582950.0 ;
      RECT  110100.0 1582950.0 111300.0 1581750.0 ;
      RECT  112500.0 1582950.0 113700.0 1581750.0 ;
      RECT  112500.0 1582950.0 113700.0 1581750.0 ;
      RECT  110100.0 1582950.0 111300.0 1581750.0 ;
      RECT  110100.0 1592250.0 111300.0 1591050.0 ;
      RECT  112500.0 1592250.0 113700.0 1591050.0 ;
      RECT  112500.0 1592250.0 113700.0 1591050.0 ;
      RECT  110100.0 1592250.0 111300.0 1591050.0 ;
      RECT  114900.0 1582350.0 116100.0 1581150.0 ;
      RECT  114900.0 1592250.0 116100.0 1591050.0 ;
      RECT  110700.0 1587600.0 111900.0 1586400.0 ;
      RECT  110700.0 1587600.0 111900.0 1586400.0 ;
      RECT  113250.0 1587450.0 114150.0 1586550.0 ;
      RECT  108300.0 1580250.0 117900.0 1579350.0 ;
      RECT  108300.0 1594050.0 117900.0 1593150.0 ;
      RECT  114900.0 1605450.0 116100.0 1607400.0 ;
      RECT  114900.0 1593600.0 116100.0 1595550.0 ;
      RECT  110100.0 1594950.0 111300.0 1593150.0 ;
      RECT  110100.0 1604250.0 111300.0 1607850.0 ;
      RECT  112800.0 1594950.0 113700.0 1604250.0 ;
      RECT  110100.0 1604250.0 111300.0 1605450.0 ;
      RECT  112500.0 1604250.0 113700.0 1605450.0 ;
      RECT  112500.0 1604250.0 113700.0 1605450.0 ;
      RECT  110100.0 1604250.0 111300.0 1605450.0 ;
      RECT  110100.0 1594950.0 111300.0 1596150.0 ;
      RECT  112500.0 1594950.0 113700.0 1596150.0 ;
      RECT  112500.0 1594950.0 113700.0 1596150.0 ;
      RECT  110100.0 1594950.0 111300.0 1596150.0 ;
      RECT  114900.0 1604850.0 116100.0 1606050.0 ;
      RECT  114900.0 1594950.0 116100.0 1596150.0 ;
      RECT  110700.0 1599600.0 111900.0 1600800.0 ;
      RECT  110700.0 1599600.0 111900.0 1600800.0 ;
      RECT  113250.0 1599750.0 114150.0 1600650.0 ;
      RECT  108300.0 1606950.0 117900.0 1607850.0 ;
      RECT  108300.0 1593150.0 117900.0 1594050.0 ;
      RECT  114900.0 1609350.0 116100.0 1607400.0 ;
      RECT  114900.0 1621200.0 116100.0 1619250.0 ;
      RECT  110100.0 1619850.0 111300.0 1621650.0 ;
      RECT  110100.0 1610550.0 111300.0 1606950.0 ;
      RECT  112800.0 1619850.0 113700.0 1610550.0 ;
      RECT  110100.0 1610550.0 111300.0 1609350.0 ;
      RECT  112500.0 1610550.0 113700.0 1609350.0 ;
      RECT  112500.0 1610550.0 113700.0 1609350.0 ;
      RECT  110100.0 1610550.0 111300.0 1609350.0 ;
      RECT  110100.0 1619850.0 111300.0 1618650.0 ;
      RECT  112500.0 1619850.0 113700.0 1618650.0 ;
      RECT  112500.0 1619850.0 113700.0 1618650.0 ;
      RECT  110100.0 1619850.0 111300.0 1618650.0 ;
      RECT  114900.0 1609950.0 116100.0 1608750.0 ;
      RECT  114900.0 1619850.0 116100.0 1618650.0 ;
      RECT  110700.0 1615200.0 111900.0 1614000.0 ;
      RECT  110700.0 1615200.0 111900.0 1614000.0 ;
      RECT  113250.0 1615050.0 114150.0 1614150.0 ;
      RECT  108300.0 1607850.0 117900.0 1606950.0 ;
      RECT  108300.0 1621650.0 117900.0 1620750.0 ;
      RECT  114900.0 1633050.0 116100.0 1635000.0 ;
      RECT  114900.0 1621200.0 116100.0 1623150.0 ;
      RECT  110100.0 1622550.0 111300.0 1620750.0 ;
      RECT  110100.0 1631850.0 111300.0 1635450.0 ;
      RECT  112800.0 1622550.0 113700.0 1631850.0 ;
      RECT  110100.0 1631850.0 111300.0 1633050.0 ;
      RECT  112500.0 1631850.0 113700.0 1633050.0 ;
      RECT  112500.0 1631850.0 113700.0 1633050.0 ;
      RECT  110100.0 1631850.0 111300.0 1633050.0 ;
      RECT  110100.0 1622550.0 111300.0 1623750.0 ;
      RECT  112500.0 1622550.0 113700.0 1623750.0 ;
      RECT  112500.0 1622550.0 113700.0 1623750.0 ;
      RECT  110100.0 1622550.0 111300.0 1623750.0 ;
      RECT  114900.0 1632450.0 116100.0 1633650.0 ;
      RECT  114900.0 1622550.0 116100.0 1623750.0 ;
      RECT  110700.0 1627200.0 111900.0 1628400.0 ;
      RECT  110700.0 1627200.0 111900.0 1628400.0 ;
      RECT  113250.0 1627350.0 114150.0 1628250.0 ;
      RECT  108300.0 1634550.0 117900.0 1635450.0 ;
      RECT  108300.0 1620750.0 117900.0 1621650.0 ;
      RECT  114900.0 1636950.0 116100.0 1635000.0 ;
      RECT  114900.0 1648800.0 116100.0 1646850.0 ;
      RECT  110100.0 1647450.0 111300.0 1649250.0 ;
      RECT  110100.0 1638150.0 111300.0 1634550.0 ;
      RECT  112800.0 1647450.0 113700.0 1638150.0 ;
      RECT  110100.0 1638150.0 111300.0 1636950.0 ;
      RECT  112500.0 1638150.0 113700.0 1636950.0 ;
      RECT  112500.0 1638150.0 113700.0 1636950.0 ;
      RECT  110100.0 1638150.0 111300.0 1636950.0 ;
      RECT  110100.0 1647450.0 111300.0 1646250.0 ;
      RECT  112500.0 1647450.0 113700.0 1646250.0 ;
      RECT  112500.0 1647450.0 113700.0 1646250.0 ;
      RECT  110100.0 1647450.0 111300.0 1646250.0 ;
      RECT  114900.0 1637550.0 116100.0 1636350.0 ;
      RECT  114900.0 1647450.0 116100.0 1646250.0 ;
      RECT  110700.0 1642800.0 111900.0 1641600.0 ;
      RECT  110700.0 1642800.0 111900.0 1641600.0 ;
      RECT  113250.0 1642650.0 114150.0 1641750.0 ;
      RECT  108300.0 1635450.0 117900.0 1634550.0 ;
      RECT  108300.0 1649250.0 117900.0 1648350.0 ;
      RECT  114900.0 1660650.0 116100.0 1662600.0 ;
      RECT  114900.0 1648800.0 116100.0 1650750.0 ;
      RECT  110100.0 1650150.0 111300.0 1648350.0 ;
      RECT  110100.0 1659450.0 111300.0 1663050.0 ;
      RECT  112800.0 1650150.0 113700.0 1659450.0 ;
      RECT  110100.0 1659450.0 111300.0 1660650.0 ;
      RECT  112500.0 1659450.0 113700.0 1660650.0 ;
      RECT  112500.0 1659450.0 113700.0 1660650.0 ;
      RECT  110100.0 1659450.0 111300.0 1660650.0 ;
      RECT  110100.0 1650150.0 111300.0 1651350.0 ;
      RECT  112500.0 1650150.0 113700.0 1651350.0 ;
      RECT  112500.0 1650150.0 113700.0 1651350.0 ;
      RECT  110100.0 1650150.0 111300.0 1651350.0 ;
      RECT  114900.0 1660050.0 116100.0 1661250.0 ;
      RECT  114900.0 1650150.0 116100.0 1651350.0 ;
      RECT  110700.0 1654800.0 111900.0 1656000.0 ;
      RECT  110700.0 1654800.0 111900.0 1656000.0 ;
      RECT  113250.0 1654950.0 114150.0 1655850.0 ;
      RECT  108300.0 1662150.0 117900.0 1663050.0 ;
      RECT  108300.0 1648350.0 117900.0 1649250.0 ;
      RECT  114900.0 1664550.0 116100.0 1662600.0 ;
      RECT  114900.0 1676400.0 116100.0 1674450.0 ;
      RECT  110100.0 1675050.0 111300.0 1676850.0 ;
      RECT  110100.0 1665750.0 111300.0 1662150.0 ;
      RECT  112800.0 1675050.0 113700.0 1665750.0 ;
      RECT  110100.0 1665750.0 111300.0 1664550.0 ;
      RECT  112500.0 1665750.0 113700.0 1664550.0 ;
      RECT  112500.0 1665750.0 113700.0 1664550.0 ;
      RECT  110100.0 1665750.0 111300.0 1664550.0 ;
      RECT  110100.0 1675050.0 111300.0 1673850.0 ;
      RECT  112500.0 1675050.0 113700.0 1673850.0 ;
      RECT  112500.0 1675050.0 113700.0 1673850.0 ;
      RECT  110100.0 1675050.0 111300.0 1673850.0 ;
      RECT  114900.0 1665150.0 116100.0 1663950.0 ;
      RECT  114900.0 1675050.0 116100.0 1673850.0 ;
      RECT  110700.0 1670400.0 111900.0 1669200.0 ;
      RECT  110700.0 1670400.0 111900.0 1669200.0 ;
      RECT  113250.0 1670250.0 114150.0 1669350.0 ;
      RECT  108300.0 1663050.0 117900.0 1662150.0 ;
      RECT  108300.0 1676850.0 117900.0 1675950.0 ;
      RECT  114900.0 1688250.0 116100.0 1690200.0 ;
      RECT  114900.0 1676400.0 116100.0 1678350.0 ;
      RECT  110100.0 1677750.0 111300.0 1675950.0 ;
      RECT  110100.0 1687050.0 111300.0 1690650.0 ;
      RECT  112800.0 1677750.0 113700.0 1687050.0 ;
      RECT  110100.0 1687050.0 111300.0 1688250.0 ;
      RECT  112500.0 1687050.0 113700.0 1688250.0 ;
      RECT  112500.0 1687050.0 113700.0 1688250.0 ;
      RECT  110100.0 1687050.0 111300.0 1688250.0 ;
      RECT  110100.0 1677750.0 111300.0 1678950.0 ;
      RECT  112500.0 1677750.0 113700.0 1678950.0 ;
      RECT  112500.0 1677750.0 113700.0 1678950.0 ;
      RECT  110100.0 1677750.0 111300.0 1678950.0 ;
      RECT  114900.0 1687650.0 116100.0 1688850.0 ;
      RECT  114900.0 1677750.0 116100.0 1678950.0 ;
      RECT  110700.0 1682400.0 111900.0 1683600.0 ;
      RECT  110700.0 1682400.0 111900.0 1683600.0 ;
      RECT  113250.0 1682550.0 114150.0 1683450.0 ;
      RECT  108300.0 1689750.0 117900.0 1690650.0 ;
      RECT  108300.0 1675950.0 117900.0 1676850.0 ;
      RECT  114900.0 1692150.0 116100.0 1690200.0 ;
      RECT  114900.0 1704000.0 116100.0 1702050.0 ;
      RECT  110100.0 1702650.0 111300.0 1704450.0 ;
      RECT  110100.0 1693350.0 111300.0 1689750.0 ;
      RECT  112800.0 1702650.0 113700.0 1693350.0 ;
      RECT  110100.0 1693350.0 111300.0 1692150.0 ;
      RECT  112500.0 1693350.0 113700.0 1692150.0 ;
      RECT  112500.0 1693350.0 113700.0 1692150.0 ;
      RECT  110100.0 1693350.0 111300.0 1692150.0 ;
      RECT  110100.0 1702650.0 111300.0 1701450.0 ;
      RECT  112500.0 1702650.0 113700.0 1701450.0 ;
      RECT  112500.0 1702650.0 113700.0 1701450.0 ;
      RECT  110100.0 1702650.0 111300.0 1701450.0 ;
      RECT  114900.0 1692750.0 116100.0 1691550.0 ;
      RECT  114900.0 1702650.0 116100.0 1701450.0 ;
      RECT  110700.0 1698000.0 111900.0 1696800.0 ;
      RECT  110700.0 1698000.0 111900.0 1696800.0 ;
      RECT  113250.0 1697850.0 114150.0 1696950.0 ;
      RECT  108300.0 1690650.0 117900.0 1689750.0 ;
      RECT  108300.0 1704450.0 117900.0 1703550.0 ;
      RECT  114900.0 1715850.0 116100.0 1717800.0 ;
      RECT  114900.0 1704000.0 116100.0 1705950.0 ;
      RECT  110100.0 1705350.0 111300.0 1703550.0 ;
      RECT  110100.0 1714650.0 111300.0 1718250.0 ;
      RECT  112800.0 1705350.0 113700.0 1714650.0 ;
      RECT  110100.0 1714650.0 111300.0 1715850.0 ;
      RECT  112500.0 1714650.0 113700.0 1715850.0 ;
      RECT  112500.0 1714650.0 113700.0 1715850.0 ;
      RECT  110100.0 1714650.0 111300.0 1715850.0 ;
      RECT  110100.0 1705350.0 111300.0 1706550.0 ;
      RECT  112500.0 1705350.0 113700.0 1706550.0 ;
      RECT  112500.0 1705350.0 113700.0 1706550.0 ;
      RECT  110100.0 1705350.0 111300.0 1706550.0 ;
      RECT  114900.0 1715250.0 116100.0 1716450.0 ;
      RECT  114900.0 1705350.0 116100.0 1706550.0 ;
      RECT  110700.0 1710000.0 111900.0 1711200.0 ;
      RECT  110700.0 1710000.0 111900.0 1711200.0 ;
      RECT  113250.0 1710150.0 114150.0 1711050.0 ;
      RECT  108300.0 1717350.0 117900.0 1718250.0 ;
      RECT  108300.0 1703550.0 117900.0 1704450.0 ;
      RECT  114900.0 1719750.0 116100.0 1717800.0 ;
      RECT  114900.0 1731600.0 116100.0 1729650.0 ;
      RECT  110100.0 1730250.0 111300.0 1732050.0 ;
      RECT  110100.0 1720950.0 111300.0 1717350.0 ;
      RECT  112800.0 1730250.0 113700.0 1720950.0 ;
      RECT  110100.0 1720950.0 111300.0 1719750.0 ;
      RECT  112500.0 1720950.0 113700.0 1719750.0 ;
      RECT  112500.0 1720950.0 113700.0 1719750.0 ;
      RECT  110100.0 1720950.0 111300.0 1719750.0 ;
      RECT  110100.0 1730250.0 111300.0 1729050.0 ;
      RECT  112500.0 1730250.0 113700.0 1729050.0 ;
      RECT  112500.0 1730250.0 113700.0 1729050.0 ;
      RECT  110100.0 1730250.0 111300.0 1729050.0 ;
      RECT  114900.0 1720350.0 116100.0 1719150.0 ;
      RECT  114900.0 1730250.0 116100.0 1729050.0 ;
      RECT  110700.0 1725600.0 111900.0 1724400.0 ;
      RECT  110700.0 1725600.0 111900.0 1724400.0 ;
      RECT  113250.0 1725450.0 114150.0 1724550.0 ;
      RECT  108300.0 1718250.0 117900.0 1717350.0 ;
      RECT  108300.0 1732050.0 117900.0 1731150.0 ;
      RECT  114900.0 1743450.0 116100.0 1745400.0 ;
      RECT  114900.0 1731600.0 116100.0 1733550.0 ;
      RECT  110100.0 1732950.0 111300.0 1731150.0 ;
      RECT  110100.0 1742250.0 111300.0 1745850.0 ;
      RECT  112800.0 1732950.0 113700.0 1742250.0 ;
      RECT  110100.0 1742250.0 111300.0 1743450.0 ;
      RECT  112500.0 1742250.0 113700.0 1743450.0 ;
      RECT  112500.0 1742250.0 113700.0 1743450.0 ;
      RECT  110100.0 1742250.0 111300.0 1743450.0 ;
      RECT  110100.0 1732950.0 111300.0 1734150.0 ;
      RECT  112500.0 1732950.0 113700.0 1734150.0 ;
      RECT  112500.0 1732950.0 113700.0 1734150.0 ;
      RECT  110100.0 1732950.0 111300.0 1734150.0 ;
      RECT  114900.0 1742850.0 116100.0 1744050.0 ;
      RECT  114900.0 1732950.0 116100.0 1734150.0 ;
      RECT  110700.0 1737600.0 111900.0 1738800.0 ;
      RECT  110700.0 1737600.0 111900.0 1738800.0 ;
      RECT  113250.0 1737750.0 114150.0 1738650.0 ;
      RECT  108300.0 1744950.0 117900.0 1745850.0 ;
      RECT  108300.0 1731150.0 117900.0 1732050.0 ;
      RECT  114900.0 1747350.0 116100.0 1745400.0 ;
      RECT  114900.0 1759200.0 116100.0 1757250.0 ;
      RECT  110100.0 1757850.0 111300.0 1759650.0 ;
      RECT  110100.0 1748550.0 111300.0 1744950.0 ;
      RECT  112800.0 1757850.0 113700.0 1748550.0 ;
      RECT  110100.0 1748550.0 111300.0 1747350.0 ;
      RECT  112500.0 1748550.0 113700.0 1747350.0 ;
      RECT  112500.0 1748550.0 113700.0 1747350.0 ;
      RECT  110100.0 1748550.0 111300.0 1747350.0 ;
      RECT  110100.0 1757850.0 111300.0 1756650.0 ;
      RECT  112500.0 1757850.0 113700.0 1756650.0 ;
      RECT  112500.0 1757850.0 113700.0 1756650.0 ;
      RECT  110100.0 1757850.0 111300.0 1756650.0 ;
      RECT  114900.0 1747950.0 116100.0 1746750.0 ;
      RECT  114900.0 1757850.0 116100.0 1756650.0 ;
      RECT  110700.0 1753200.0 111900.0 1752000.0 ;
      RECT  110700.0 1753200.0 111900.0 1752000.0 ;
      RECT  113250.0 1753050.0 114150.0 1752150.0 ;
      RECT  108300.0 1745850.0 117900.0 1744950.0 ;
      RECT  108300.0 1759650.0 117900.0 1758750.0 ;
      RECT  114900.0 1771050.0 116100.0 1773000.0 ;
      RECT  114900.0 1759200.0 116100.0 1761150.0 ;
      RECT  110100.0 1760550.0 111300.0 1758750.0 ;
      RECT  110100.0 1769850.0 111300.0 1773450.0 ;
      RECT  112800.0 1760550.0 113700.0 1769850.0 ;
      RECT  110100.0 1769850.0 111300.0 1771050.0 ;
      RECT  112500.0 1769850.0 113700.0 1771050.0 ;
      RECT  112500.0 1769850.0 113700.0 1771050.0 ;
      RECT  110100.0 1769850.0 111300.0 1771050.0 ;
      RECT  110100.0 1760550.0 111300.0 1761750.0 ;
      RECT  112500.0 1760550.0 113700.0 1761750.0 ;
      RECT  112500.0 1760550.0 113700.0 1761750.0 ;
      RECT  110100.0 1760550.0 111300.0 1761750.0 ;
      RECT  114900.0 1770450.0 116100.0 1771650.0 ;
      RECT  114900.0 1760550.0 116100.0 1761750.0 ;
      RECT  110700.0 1765200.0 111900.0 1766400.0 ;
      RECT  110700.0 1765200.0 111900.0 1766400.0 ;
      RECT  113250.0 1765350.0 114150.0 1766250.0 ;
      RECT  108300.0 1772550.0 117900.0 1773450.0 ;
      RECT  108300.0 1758750.0 117900.0 1759650.0 ;
      RECT  114900.0 1774950.0 116100.0 1773000.0 ;
      RECT  114900.0 1786800.0 116100.0 1784850.0 ;
      RECT  110100.0 1785450.0 111300.0 1787250.0 ;
      RECT  110100.0 1776150.0 111300.0 1772550.0 ;
      RECT  112800.0 1785450.0 113700.0 1776150.0 ;
      RECT  110100.0 1776150.0 111300.0 1774950.0 ;
      RECT  112500.0 1776150.0 113700.0 1774950.0 ;
      RECT  112500.0 1776150.0 113700.0 1774950.0 ;
      RECT  110100.0 1776150.0 111300.0 1774950.0 ;
      RECT  110100.0 1785450.0 111300.0 1784250.0 ;
      RECT  112500.0 1785450.0 113700.0 1784250.0 ;
      RECT  112500.0 1785450.0 113700.0 1784250.0 ;
      RECT  110100.0 1785450.0 111300.0 1784250.0 ;
      RECT  114900.0 1775550.0 116100.0 1774350.0 ;
      RECT  114900.0 1785450.0 116100.0 1784250.0 ;
      RECT  110700.0 1780800.0 111900.0 1779600.0 ;
      RECT  110700.0 1780800.0 111900.0 1779600.0 ;
      RECT  113250.0 1780650.0 114150.0 1779750.0 ;
      RECT  108300.0 1773450.0 117900.0 1772550.0 ;
      RECT  108300.0 1787250.0 117900.0 1786350.0 ;
      RECT  114900.0 1798650.0 116100.0 1800600.0 ;
      RECT  114900.0 1786800.0 116100.0 1788750.0 ;
      RECT  110100.0 1788150.0 111300.0 1786350.0 ;
      RECT  110100.0 1797450.0 111300.0 1801050.0 ;
      RECT  112800.0 1788150.0 113700.0 1797450.0 ;
      RECT  110100.0 1797450.0 111300.0 1798650.0 ;
      RECT  112500.0 1797450.0 113700.0 1798650.0 ;
      RECT  112500.0 1797450.0 113700.0 1798650.0 ;
      RECT  110100.0 1797450.0 111300.0 1798650.0 ;
      RECT  110100.0 1788150.0 111300.0 1789350.0 ;
      RECT  112500.0 1788150.0 113700.0 1789350.0 ;
      RECT  112500.0 1788150.0 113700.0 1789350.0 ;
      RECT  110100.0 1788150.0 111300.0 1789350.0 ;
      RECT  114900.0 1798050.0 116100.0 1799250.0 ;
      RECT  114900.0 1788150.0 116100.0 1789350.0 ;
      RECT  110700.0 1792800.0 111900.0 1794000.0 ;
      RECT  110700.0 1792800.0 111900.0 1794000.0 ;
      RECT  113250.0 1792950.0 114150.0 1793850.0 ;
      RECT  108300.0 1800150.0 117900.0 1801050.0 ;
      RECT  108300.0 1786350.0 117900.0 1787250.0 ;
      RECT  114900.0 1802550.0 116100.0 1800600.0 ;
      RECT  114900.0 1814400.0 116100.0 1812450.0 ;
      RECT  110100.0 1813050.0 111300.0 1814850.0 ;
      RECT  110100.0 1803750.0 111300.0 1800150.0 ;
      RECT  112800.0 1813050.0 113700.0 1803750.0 ;
      RECT  110100.0 1803750.0 111300.0 1802550.0 ;
      RECT  112500.0 1803750.0 113700.0 1802550.0 ;
      RECT  112500.0 1803750.0 113700.0 1802550.0 ;
      RECT  110100.0 1803750.0 111300.0 1802550.0 ;
      RECT  110100.0 1813050.0 111300.0 1811850.0 ;
      RECT  112500.0 1813050.0 113700.0 1811850.0 ;
      RECT  112500.0 1813050.0 113700.0 1811850.0 ;
      RECT  110100.0 1813050.0 111300.0 1811850.0 ;
      RECT  114900.0 1803150.0 116100.0 1801950.0 ;
      RECT  114900.0 1813050.0 116100.0 1811850.0 ;
      RECT  110700.0 1808400.0 111900.0 1807200.0 ;
      RECT  110700.0 1808400.0 111900.0 1807200.0 ;
      RECT  113250.0 1808250.0 114150.0 1807350.0 ;
      RECT  108300.0 1801050.0 117900.0 1800150.0 ;
      RECT  108300.0 1814850.0 117900.0 1813950.0 ;
      RECT  114900.0 1826250.0 116100.0 1828200.0 ;
      RECT  114900.0 1814400.0 116100.0 1816350.0 ;
      RECT  110100.0 1815750.0 111300.0 1813950.0 ;
      RECT  110100.0 1825050.0 111300.0 1828650.0 ;
      RECT  112800.0 1815750.0 113700.0 1825050.0 ;
      RECT  110100.0 1825050.0 111300.0 1826250.0 ;
      RECT  112500.0 1825050.0 113700.0 1826250.0 ;
      RECT  112500.0 1825050.0 113700.0 1826250.0 ;
      RECT  110100.0 1825050.0 111300.0 1826250.0 ;
      RECT  110100.0 1815750.0 111300.0 1816950.0 ;
      RECT  112500.0 1815750.0 113700.0 1816950.0 ;
      RECT  112500.0 1815750.0 113700.0 1816950.0 ;
      RECT  110100.0 1815750.0 111300.0 1816950.0 ;
      RECT  114900.0 1825650.0 116100.0 1826850.0 ;
      RECT  114900.0 1815750.0 116100.0 1816950.0 ;
      RECT  110700.0 1820400.0 111900.0 1821600.0 ;
      RECT  110700.0 1820400.0 111900.0 1821600.0 ;
      RECT  113250.0 1820550.0 114150.0 1821450.0 ;
      RECT  108300.0 1827750.0 117900.0 1828650.0 ;
      RECT  108300.0 1813950.0 117900.0 1814850.0 ;
      RECT  114900.0 1830150.0 116100.0 1828200.0 ;
      RECT  114900.0 1842000.0 116100.0 1840050.0 ;
      RECT  110100.0 1840650.0 111300.0 1842450.0 ;
      RECT  110100.0 1831350.0 111300.0 1827750.0 ;
      RECT  112800.0 1840650.0 113700.0 1831350.0 ;
      RECT  110100.0 1831350.0 111300.0 1830150.0 ;
      RECT  112500.0 1831350.0 113700.0 1830150.0 ;
      RECT  112500.0 1831350.0 113700.0 1830150.0 ;
      RECT  110100.0 1831350.0 111300.0 1830150.0 ;
      RECT  110100.0 1840650.0 111300.0 1839450.0 ;
      RECT  112500.0 1840650.0 113700.0 1839450.0 ;
      RECT  112500.0 1840650.0 113700.0 1839450.0 ;
      RECT  110100.0 1840650.0 111300.0 1839450.0 ;
      RECT  114900.0 1830750.0 116100.0 1829550.0 ;
      RECT  114900.0 1840650.0 116100.0 1839450.0 ;
      RECT  110700.0 1836000.0 111900.0 1834800.0 ;
      RECT  110700.0 1836000.0 111900.0 1834800.0 ;
      RECT  113250.0 1835850.0 114150.0 1834950.0 ;
      RECT  108300.0 1828650.0 117900.0 1827750.0 ;
      RECT  108300.0 1842450.0 117900.0 1841550.0 ;
      RECT  114900.0 1853850.0 116100.0 1855800.0 ;
      RECT  114900.0 1842000.0 116100.0 1843950.0 ;
      RECT  110100.0 1843350.0 111300.0 1841550.0 ;
      RECT  110100.0 1852650.0 111300.0 1856250.0 ;
      RECT  112800.0 1843350.0 113700.0 1852650.0 ;
      RECT  110100.0 1852650.0 111300.0 1853850.0 ;
      RECT  112500.0 1852650.0 113700.0 1853850.0 ;
      RECT  112500.0 1852650.0 113700.0 1853850.0 ;
      RECT  110100.0 1852650.0 111300.0 1853850.0 ;
      RECT  110100.0 1843350.0 111300.0 1844550.0 ;
      RECT  112500.0 1843350.0 113700.0 1844550.0 ;
      RECT  112500.0 1843350.0 113700.0 1844550.0 ;
      RECT  110100.0 1843350.0 111300.0 1844550.0 ;
      RECT  114900.0 1853250.0 116100.0 1854450.0 ;
      RECT  114900.0 1843350.0 116100.0 1844550.0 ;
      RECT  110700.0 1848000.0 111900.0 1849200.0 ;
      RECT  110700.0 1848000.0 111900.0 1849200.0 ;
      RECT  113250.0 1848150.0 114150.0 1849050.0 ;
      RECT  108300.0 1855350.0 117900.0 1856250.0 ;
      RECT  108300.0 1841550.0 117900.0 1842450.0 ;
      RECT  114900.0 1857750.0 116100.0 1855800.0 ;
      RECT  114900.0 1869600.0 116100.0 1867650.0 ;
      RECT  110100.0 1868250.0 111300.0 1870050.0 ;
      RECT  110100.0 1858950.0 111300.0 1855350.0 ;
      RECT  112800.0 1868250.0 113700.0 1858950.0 ;
      RECT  110100.0 1858950.0 111300.0 1857750.0 ;
      RECT  112500.0 1858950.0 113700.0 1857750.0 ;
      RECT  112500.0 1858950.0 113700.0 1857750.0 ;
      RECT  110100.0 1858950.0 111300.0 1857750.0 ;
      RECT  110100.0 1868250.0 111300.0 1867050.0 ;
      RECT  112500.0 1868250.0 113700.0 1867050.0 ;
      RECT  112500.0 1868250.0 113700.0 1867050.0 ;
      RECT  110100.0 1868250.0 111300.0 1867050.0 ;
      RECT  114900.0 1858350.0 116100.0 1857150.0 ;
      RECT  114900.0 1868250.0 116100.0 1867050.0 ;
      RECT  110700.0 1863600.0 111900.0 1862400.0 ;
      RECT  110700.0 1863600.0 111900.0 1862400.0 ;
      RECT  113250.0 1863450.0 114150.0 1862550.0 ;
      RECT  108300.0 1856250.0 117900.0 1855350.0 ;
      RECT  108300.0 1870050.0 117900.0 1869150.0 ;
      RECT  114900.0 1881450.0 116100.0 1883400.0 ;
      RECT  114900.0 1869600.0 116100.0 1871550.0 ;
      RECT  110100.0 1870950.0 111300.0 1869150.0 ;
      RECT  110100.0 1880250.0 111300.0 1883850.0 ;
      RECT  112800.0 1870950.0 113700.0 1880250.0 ;
      RECT  110100.0 1880250.0 111300.0 1881450.0 ;
      RECT  112500.0 1880250.0 113700.0 1881450.0 ;
      RECT  112500.0 1880250.0 113700.0 1881450.0 ;
      RECT  110100.0 1880250.0 111300.0 1881450.0 ;
      RECT  110100.0 1870950.0 111300.0 1872150.0 ;
      RECT  112500.0 1870950.0 113700.0 1872150.0 ;
      RECT  112500.0 1870950.0 113700.0 1872150.0 ;
      RECT  110100.0 1870950.0 111300.0 1872150.0 ;
      RECT  114900.0 1880850.0 116100.0 1882050.0 ;
      RECT  114900.0 1870950.0 116100.0 1872150.0 ;
      RECT  110700.0 1875600.0 111900.0 1876800.0 ;
      RECT  110700.0 1875600.0 111900.0 1876800.0 ;
      RECT  113250.0 1875750.0 114150.0 1876650.0 ;
      RECT  108300.0 1882950.0 117900.0 1883850.0 ;
      RECT  108300.0 1869150.0 117900.0 1870050.0 ;
      RECT  114900.0 1885350.0 116100.0 1883400.0 ;
      RECT  114900.0 1897200.0 116100.0 1895250.0 ;
      RECT  110100.0 1895850.0 111300.0 1897650.0 ;
      RECT  110100.0 1886550.0 111300.0 1882950.0 ;
      RECT  112800.0 1895850.0 113700.0 1886550.0 ;
      RECT  110100.0 1886550.0 111300.0 1885350.0 ;
      RECT  112500.0 1886550.0 113700.0 1885350.0 ;
      RECT  112500.0 1886550.0 113700.0 1885350.0 ;
      RECT  110100.0 1886550.0 111300.0 1885350.0 ;
      RECT  110100.0 1895850.0 111300.0 1894650.0 ;
      RECT  112500.0 1895850.0 113700.0 1894650.0 ;
      RECT  112500.0 1895850.0 113700.0 1894650.0 ;
      RECT  110100.0 1895850.0 111300.0 1894650.0 ;
      RECT  114900.0 1885950.0 116100.0 1884750.0 ;
      RECT  114900.0 1895850.0 116100.0 1894650.0 ;
      RECT  110700.0 1891200.0 111900.0 1890000.0 ;
      RECT  110700.0 1891200.0 111900.0 1890000.0 ;
      RECT  113250.0 1891050.0 114150.0 1890150.0 ;
      RECT  108300.0 1883850.0 117900.0 1882950.0 ;
      RECT  108300.0 1897650.0 117900.0 1896750.0 ;
      RECT  114900.0 1909050.0 116100.0 1911000.0 ;
      RECT  114900.0 1897200.0 116100.0 1899150.0 ;
      RECT  110100.0 1898550.0 111300.0 1896750.0 ;
      RECT  110100.0 1907850.0 111300.0 1911450.0 ;
      RECT  112800.0 1898550.0 113700.0 1907850.0 ;
      RECT  110100.0 1907850.0 111300.0 1909050.0 ;
      RECT  112500.0 1907850.0 113700.0 1909050.0 ;
      RECT  112500.0 1907850.0 113700.0 1909050.0 ;
      RECT  110100.0 1907850.0 111300.0 1909050.0 ;
      RECT  110100.0 1898550.0 111300.0 1899750.0 ;
      RECT  112500.0 1898550.0 113700.0 1899750.0 ;
      RECT  112500.0 1898550.0 113700.0 1899750.0 ;
      RECT  110100.0 1898550.0 111300.0 1899750.0 ;
      RECT  114900.0 1908450.0 116100.0 1909650.0 ;
      RECT  114900.0 1898550.0 116100.0 1899750.0 ;
      RECT  110700.0 1903200.0 111900.0 1904400.0 ;
      RECT  110700.0 1903200.0 111900.0 1904400.0 ;
      RECT  113250.0 1903350.0 114150.0 1904250.0 ;
      RECT  108300.0 1910550.0 117900.0 1911450.0 ;
      RECT  108300.0 1896750.0 117900.0 1897650.0 ;
      RECT  114900.0 1912950.0 116100.0 1911000.0 ;
      RECT  114900.0 1924800.0 116100.0 1922850.0 ;
      RECT  110100.0 1923450.0 111300.0 1925250.0 ;
      RECT  110100.0 1914150.0 111300.0 1910550.0 ;
      RECT  112800.0 1923450.0 113700.0 1914150.0 ;
      RECT  110100.0 1914150.0 111300.0 1912950.0 ;
      RECT  112500.0 1914150.0 113700.0 1912950.0 ;
      RECT  112500.0 1914150.0 113700.0 1912950.0 ;
      RECT  110100.0 1914150.0 111300.0 1912950.0 ;
      RECT  110100.0 1923450.0 111300.0 1922250.0 ;
      RECT  112500.0 1923450.0 113700.0 1922250.0 ;
      RECT  112500.0 1923450.0 113700.0 1922250.0 ;
      RECT  110100.0 1923450.0 111300.0 1922250.0 ;
      RECT  114900.0 1913550.0 116100.0 1912350.0 ;
      RECT  114900.0 1923450.0 116100.0 1922250.0 ;
      RECT  110700.0 1918800.0 111900.0 1917600.0 ;
      RECT  110700.0 1918800.0 111900.0 1917600.0 ;
      RECT  113250.0 1918650.0 114150.0 1917750.0 ;
      RECT  108300.0 1911450.0 117900.0 1910550.0 ;
      RECT  108300.0 1925250.0 117900.0 1924350.0 ;
      RECT  114900.0 1936650.0 116100.0 1938600.0 ;
      RECT  114900.0 1924800.0 116100.0 1926750.0 ;
      RECT  110100.0 1926150.0 111300.0 1924350.0 ;
      RECT  110100.0 1935450.0 111300.0 1939050.0 ;
      RECT  112800.0 1926150.0 113700.0 1935450.0 ;
      RECT  110100.0 1935450.0 111300.0 1936650.0 ;
      RECT  112500.0 1935450.0 113700.0 1936650.0 ;
      RECT  112500.0 1935450.0 113700.0 1936650.0 ;
      RECT  110100.0 1935450.0 111300.0 1936650.0 ;
      RECT  110100.0 1926150.0 111300.0 1927350.0 ;
      RECT  112500.0 1926150.0 113700.0 1927350.0 ;
      RECT  112500.0 1926150.0 113700.0 1927350.0 ;
      RECT  110100.0 1926150.0 111300.0 1927350.0 ;
      RECT  114900.0 1936050.0 116100.0 1937250.0 ;
      RECT  114900.0 1926150.0 116100.0 1927350.0 ;
      RECT  110700.0 1930800.0 111900.0 1932000.0 ;
      RECT  110700.0 1930800.0 111900.0 1932000.0 ;
      RECT  113250.0 1930950.0 114150.0 1931850.0 ;
      RECT  108300.0 1938150.0 117900.0 1939050.0 ;
      RECT  108300.0 1924350.0 117900.0 1925250.0 ;
      RECT  114900.0 1940550.0 116100.0 1938600.0 ;
      RECT  114900.0 1952400.0 116100.0 1950450.0 ;
      RECT  110100.0 1951050.0 111300.0 1952850.0 ;
      RECT  110100.0 1941750.0 111300.0 1938150.0 ;
      RECT  112800.0 1951050.0 113700.0 1941750.0 ;
      RECT  110100.0 1941750.0 111300.0 1940550.0 ;
      RECT  112500.0 1941750.0 113700.0 1940550.0 ;
      RECT  112500.0 1941750.0 113700.0 1940550.0 ;
      RECT  110100.0 1941750.0 111300.0 1940550.0 ;
      RECT  110100.0 1951050.0 111300.0 1949850.0 ;
      RECT  112500.0 1951050.0 113700.0 1949850.0 ;
      RECT  112500.0 1951050.0 113700.0 1949850.0 ;
      RECT  110100.0 1951050.0 111300.0 1949850.0 ;
      RECT  114900.0 1941150.0 116100.0 1939950.0 ;
      RECT  114900.0 1951050.0 116100.0 1949850.0 ;
      RECT  110700.0 1946400.0 111900.0 1945200.0 ;
      RECT  110700.0 1946400.0 111900.0 1945200.0 ;
      RECT  113250.0 1946250.0 114150.0 1945350.0 ;
      RECT  108300.0 1939050.0 117900.0 1938150.0 ;
      RECT  108300.0 1952850.0 117900.0 1951950.0 ;
      RECT  114900.0 1964250.0 116100.0 1966200.0 ;
      RECT  114900.0 1952400.0 116100.0 1954350.0 ;
      RECT  110100.0 1953750.0 111300.0 1951950.0 ;
      RECT  110100.0 1963050.0 111300.0 1966650.0 ;
      RECT  112800.0 1953750.0 113700.0 1963050.0 ;
      RECT  110100.0 1963050.0 111300.0 1964250.0 ;
      RECT  112500.0 1963050.0 113700.0 1964250.0 ;
      RECT  112500.0 1963050.0 113700.0 1964250.0 ;
      RECT  110100.0 1963050.0 111300.0 1964250.0 ;
      RECT  110100.0 1953750.0 111300.0 1954950.0 ;
      RECT  112500.0 1953750.0 113700.0 1954950.0 ;
      RECT  112500.0 1953750.0 113700.0 1954950.0 ;
      RECT  110100.0 1953750.0 111300.0 1954950.0 ;
      RECT  114900.0 1963650.0 116100.0 1964850.0 ;
      RECT  114900.0 1953750.0 116100.0 1954950.0 ;
      RECT  110700.0 1958400.0 111900.0 1959600.0 ;
      RECT  110700.0 1958400.0 111900.0 1959600.0 ;
      RECT  113250.0 1958550.0 114150.0 1959450.0 ;
      RECT  108300.0 1965750.0 117900.0 1966650.0 ;
      RECT  108300.0 1951950.0 117900.0 1952850.0 ;
      RECT  114900.0 1968150.0 116100.0 1966200.0 ;
      RECT  114900.0 1980000.0 116100.0 1978050.0 ;
      RECT  110100.0 1978650.0 111300.0 1980450.0 ;
      RECT  110100.0 1969350.0 111300.0 1965750.0 ;
      RECT  112800.0 1978650.0 113700.0 1969350.0 ;
      RECT  110100.0 1969350.0 111300.0 1968150.0 ;
      RECT  112500.0 1969350.0 113700.0 1968150.0 ;
      RECT  112500.0 1969350.0 113700.0 1968150.0 ;
      RECT  110100.0 1969350.0 111300.0 1968150.0 ;
      RECT  110100.0 1978650.0 111300.0 1977450.0 ;
      RECT  112500.0 1978650.0 113700.0 1977450.0 ;
      RECT  112500.0 1978650.0 113700.0 1977450.0 ;
      RECT  110100.0 1978650.0 111300.0 1977450.0 ;
      RECT  114900.0 1968750.0 116100.0 1967550.0 ;
      RECT  114900.0 1978650.0 116100.0 1977450.0 ;
      RECT  110700.0 1974000.0 111900.0 1972800.0 ;
      RECT  110700.0 1974000.0 111900.0 1972800.0 ;
      RECT  113250.0 1973850.0 114150.0 1972950.0 ;
      RECT  108300.0 1966650.0 117900.0 1965750.0 ;
      RECT  108300.0 1980450.0 117900.0 1979550.0 ;
      RECT  114900.0 1991850.0 116100.0 1993800.0 ;
      RECT  114900.0 1980000.0 116100.0 1981950.0 ;
      RECT  110100.0 1981350.0 111300.0 1979550.0 ;
      RECT  110100.0 1990650.0 111300.0 1994250.0 ;
      RECT  112800.0 1981350.0 113700.0 1990650.0 ;
      RECT  110100.0 1990650.0 111300.0 1991850.0 ;
      RECT  112500.0 1990650.0 113700.0 1991850.0 ;
      RECT  112500.0 1990650.0 113700.0 1991850.0 ;
      RECT  110100.0 1990650.0 111300.0 1991850.0 ;
      RECT  110100.0 1981350.0 111300.0 1982550.0 ;
      RECT  112500.0 1981350.0 113700.0 1982550.0 ;
      RECT  112500.0 1981350.0 113700.0 1982550.0 ;
      RECT  110100.0 1981350.0 111300.0 1982550.0 ;
      RECT  114900.0 1991250.0 116100.0 1992450.0 ;
      RECT  114900.0 1981350.0 116100.0 1982550.0 ;
      RECT  110700.0 1986000.0 111900.0 1987200.0 ;
      RECT  110700.0 1986000.0 111900.0 1987200.0 ;
      RECT  113250.0 1986150.0 114150.0 1987050.0 ;
      RECT  108300.0 1993350.0 117900.0 1994250.0 ;
      RECT  108300.0 1979550.0 117900.0 1980450.0 ;
      RECT  114900.0 1995750.0 116100.0 1993800.0 ;
      RECT  114900.0 2007600.0 116100.0 2005650.0 ;
      RECT  110100.0 2006250.0 111300.0 2008050.0 ;
      RECT  110100.0 1996950.0 111300.0 1993350.0 ;
      RECT  112800.0 2006250.0 113700.0 1996950.0 ;
      RECT  110100.0 1996950.0 111300.0 1995750.0 ;
      RECT  112500.0 1996950.0 113700.0 1995750.0 ;
      RECT  112500.0 1996950.0 113700.0 1995750.0 ;
      RECT  110100.0 1996950.0 111300.0 1995750.0 ;
      RECT  110100.0 2006250.0 111300.0 2005050.0 ;
      RECT  112500.0 2006250.0 113700.0 2005050.0 ;
      RECT  112500.0 2006250.0 113700.0 2005050.0 ;
      RECT  110100.0 2006250.0 111300.0 2005050.0 ;
      RECT  114900.0 1996350.0 116100.0 1995150.0 ;
      RECT  114900.0 2006250.0 116100.0 2005050.0 ;
      RECT  110700.0 2001600.0 111900.0 2000400.0 ;
      RECT  110700.0 2001600.0 111900.0 2000400.0 ;
      RECT  113250.0 2001450.0 114150.0 2000550.0 ;
      RECT  108300.0 1994250.0 117900.0 1993350.0 ;
      RECT  108300.0 2008050.0 117900.0 2007150.0 ;
      RECT  114900.0 2019450.0 116100.0 2021400.0 ;
      RECT  114900.0 2007600.0 116100.0 2009550.0 ;
      RECT  110100.0 2008950.0 111300.0 2007150.0 ;
      RECT  110100.0 2018250.0 111300.0 2021850.0 ;
      RECT  112800.0 2008950.0 113700.0 2018250.0 ;
      RECT  110100.0 2018250.0 111300.0 2019450.0 ;
      RECT  112500.0 2018250.0 113700.0 2019450.0 ;
      RECT  112500.0 2018250.0 113700.0 2019450.0 ;
      RECT  110100.0 2018250.0 111300.0 2019450.0 ;
      RECT  110100.0 2008950.0 111300.0 2010150.0 ;
      RECT  112500.0 2008950.0 113700.0 2010150.0 ;
      RECT  112500.0 2008950.0 113700.0 2010150.0 ;
      RECT  110100.0 2008950.0 111300.0 2010150.0 ;
      RECT  114900.0 2018850.0 116100.0 2020050.0 ;
      RECT  114900.0 2008950.0 116100.0 2010150.0 ;
      RECT  110700.0 2013600.0 111900.0 2014800.0 ;
      RECT  110700.0 2013600.0 111900.0 2014800.0 ;
      RECT  113250.0 2013750.0 114150.0 2014650.0 ;
      RECT  108300.0 2020950.0 117900.0 2021850.0 ;
      RECT  108300.0 2007150.0 117900.0 2008050.0 ;
      RECT  114900.0 2023350.0 116100.0 2021400.0 ;
      RECT  114900.0 2035200.0 116100.0 2033250.0 ;
      RECT  110100.0 2033850.0 111300.0 2035650.0 ;
      RECT  110100.0 2024550.0 111300.0 2020950.0 ;
      RECT  112800.0 2033850.0 113700.0 2024550.0 ;
      RECT  110100.0 2024550.0 111300.0 2023350.0 ;
      RECT  112500.0 2024550.0 113700.0 2023350.0 ;
      RECT  112500.0 2024550.0 113700.0 2023350.0 ;
      RECT  110100.0 2024550.0 111300.0 2023350.0 ;
      RECT  110100.0 2033850.0 111300.0 2032650.0 ;
      RECT  112500.0 2033850.0 113700.0 2032650.0 ;
      RECT  112500.0 2033850.0 113700.0 2032650.0 ;
      RECT  110100.0 2033850.0 111300.0 2032650.0 ;
      RECT  114900.0 2023950.0 116100.0 2022750.0 ;
      RECT  114900.0 2033850.0 116100.0 2032650.0 ;
      RECT  110700.0 2029200.0 111900.0 2028000.0 ;
      RECT  110700.0 2029200.0 111900.0 2028000.0 ;
      RECT  113250.0 2029050.0 114150.0 2028150.0 ;
      RECT  108300.0 2021850.0 117900.0 2020950.0 ;
      RECT  108300.0 2035650.0 117900.0 2034750.0 ;
      RECT  114900.0 2047050.0 116100.0 2049000.0 ;
      RECT  114900.0 2035200.0 116100.0 2037150.0 ;
      RECT  110100.0 2036550.0 111300.0 2034750.0 ;
      RECT  110100.0 2045850.0 111300.0 2049450.0 ;
      RECT  112800.0 2036550.0 113700.0 2045850.0 ;
      RECT  110100.0 2045850.0 111300.0 2047050.0 ;
      RECT  112500.0 2045850.0 113700.0 2047050.0 ;
      RECT  112500.0 2045850.0 113700.0 2047050.0 ;
      RECT  110100.0 2045850.0 111300.0 2047050.0 ;
      RECT  110100.0 2036550.0 111300.0 2037750.0 ;
      RECT  112500.0 2036550.0 113700.0 2037750.0 ;
      RECT  112500.0 2036550.0 113700.0 2037750.0 ;
      RECT  110100.0 2036550.0 111300.0 2037750.0 ;
      RECT  114900.0 2046450.0 116100.0 2047650.0 ;
      RECT  114900.0 2036550.0 116100.0 2037750.0 ;
      RECT  110700.0 2041200.0 111900.0 2042400.0 ;
      RECT  110700.0 2041200.0 111900.0 2042400.0 ;
      RECT  113250.0 2041350.0 114150.0 2042250.0 ;
      RECT  108300.0 2048550.0 117900.0 2049450.0 ;
      RECT  108300.0 2034750.0 117900.0 2035650.0 ;
      RECT  114900.0 2050950.0 116100.0 2049000.0 ;
      RECT  114900.0 2062800.0 116100.0 2060850.0 ;
      RECT  110100.0 2061450.0 111300.0 2063250.0 ;
      RECT  110100.0 2052150.0 111300.0 2048550.0 ;
      RECT  112800.0 2061450.0 113700.0 2052150.0 ;
      RECT  110100.0 2052150.0 111300.0 2050950.0 ;
      RECT  112500.0 2052150.0 113700.0 2050950.0 ;
      RECT  112500.0 2052150.0 113700.0 2050950.0 ;
      RECT  110100.0 2052150.0 111300.0 2050950.0 ;
      RECT  110100.0 2061450.0 111300.0 2060250.0 ;
      RECT  112500.0 2061450.0 113700.0 2060250.0 ;
      RECT  112500.0 2061450.0 113700.0 2060250.0 ;
      RECT  110100.0 2061450.0 111300.0 2060250.0 ;
      RECT  114900.0 2051550.0 116100.0 2050350.0 ;
      RECT  114900.0 2061450.0 116100.0 2060250.0 ;
      RECT  110700.0 2056800.0 111900.0 2055600.0 ;
      RECT  110700.0 2056800.0 111900.0 2055600.0 ;
      RECT  113250.0 2056650.0 114150.0 2055750.0 ;
      RECT  108300.0 2049450.0 117900.0 2048550.0 ;
      RECT  108300.0 2063250.0 117900.0 2062350.0 ;
      RECT  114900.0 2074650.0 116100.0 2076600.0 ;
      RECT  114900.0 2062800.0 116100.0 2064750.0 ;
      RECT  110100.0 2064150.0 111300.0 2062350.0 ;
      RECT  110100.0 2073450.0 111300.0 2077050.0 ;
      RECT  112800.0 2064150.0 113700.0 2073450.0 ;
      RECT  110100.0 2073450.0 111300.0 2074650.0 ;
      RECT  112500.0 2073450.0 113700.0 2074650.0 ;
      RECT  112500.0 2073450.0 113700.0 2074650.0 ;
      RECT  110100.0 2073450.0 111300.0 2074650.0 ;
      RECT  110100.0 2064150.0 111300.0 2065350.0 ;
      RECT  112500.0 2064150.0 113700.0 2065350.0 ;
      RECT  112500.0 2064150.0 113700.0 2065350.0 ;
      RECT  110100.0 2064150.0 111300.0 2065350.0 ;
      RECT  114900.0 2074050.0 116100.0 2075250.0 ;
      RECT  114900.0 2064150.0 116100.0 2065350.0 ;
      RECT  110700.0 2068800.0 111900.0 2070000.0 ;
      RECT  110700.0 2068800.0 111900.0 2070000.0 ;
      RECT  113250.0 2068950.0 114150.0 2069850.0 ;
      RECT  108300.0 2076150.0 117900.0 2077050.0 ;
      RECT  108300.0 2062350.0 117900.0 2063250.0 ;
      RECT  114900.0 2078550.0 116100.0 2076600.0 ;
      RECT  114900.0 2090400.0 116100.0 2088450.0 ;
      RECT  110100.0 2089050.0 111300.0 2090850.0 ;
      RECT  110100.0 2079750.0 111300.0 2076150.0 ;
      RECT  112800.0 2089050.0 113700.0 2079750.0 ;
      RECT  110100.0 2079750.0 111300.0 2078550.0 ;
      RECT  112500.0 2079750.0 113700.0 2078550.0 ;
      RECT  112500.0 2079750.0 113700.0 2078550.0 ;
      RECT  110100.0 2079750.0 111300.0 2078550.0 ;
      RECT  110100.0 2089050.0 111300.0 2087850.0 ;
      RECT  112500.0 2089050.0 113700.0 2087850.0 ;
      RECT  112500.0 2089050.0 113700.0 2087850.0 ;
      RECT  110100.0 2089050.0 111300.0 2087850.0 ;
      RECT  114900.0 2079150.0 116100.0 2077950.0 ;
      RECT  114900.0 2089050.0 116100.0 2087850.0 ;
      RECT  110700.0 2084400.0 111900.0 2083200.0 ;
      RECT  110700.0 2084400.0 111900.0 2083200.0 ;
      RECT  113250.0 2084250.0 114150.0 2083350.0 ;
      RECT  108300.0 2077050.0 117900.0 2076150.0 ;
      RECT  108300.0 2090850.0 117900.0 2089950.0 ;
      RECT  114900.0 2102250.0 116100.0 2104200.0 ;
      RECT  114900.0 2090400.0 116100.0 2092350.0 ;
      RECT  110100.0 2091750.0 111300.0 2089950.0 ;
      RECT  110100.0 2101050.0 111300.0 2104650.0 ;
      RECT  112800.0 2091750.0 113700.0 2101050.0 ;
      RECT  110100.0 2101050.0 111300.0 2102250.0 ;
      RECT  112500.0 2101050.0 113700.0 2102250.0 ;
      RECT  112500.0 2101050.0 113700.0 2102250.0 ;
      RECT  110100.0 2101050.0 111300.0 2102250.0 ;
      RECT  110100.0 2091750.0 111300.0 2092950.0 ;
      RECT  112500.0 2091750.0 113700.0 2092950.0 ;
      RECT  112500.0 2091750.0 113700.0 2092950.0 ;
      RECT  110100.0 2091750.0 111300.0 2092950.0 ;
      RECT  114900.0 2101650.0 116100.0 2102850.0 ;
      RECT  114900.0 2091750.0 116100.0 2092950.0 ;
      RECT  110700.0 2096400.0 111900.0 2097600.0 ;
      RECT  110700.0 2096400.0 111900.0 2097600.0 ;
      RECT  113250.0 2096550.0 114150.0 2097450.0 ;
      RECT  108300.0 2103750.0 117900.0 2104650.0 ;
      RECT  108300.0 2089950.0 117900.0 2090850.0 ;
      RECT  114900.0 2106150.0 116100.0 2104200.0 ;
      RECT  114900.0 2118000.0 116100.0 2116050.0 ;
      RECT  110100.0 2116650.0 111300.0 2118450.0 ;
      RECT  110100.0 2107350.0 111300.0 2103750.0 ;
      RECT  112800.0 2116650.0 113700.0 2107350.0 ;
      RECT  110100.0 2107350.0 111300.0 2106150.0 ;
      RECT  112500.0 2107350.0 113700.0 2106150.0 ;
      RECT  112500.0 2107350.0 113700.0 2106150.0 ;
      RECT  110100.0 2107350.0 111300.0 2106150.0 ;
      RECT  110100.0 2116650.0 111300.0 2115450.0 ;
      RECT  112500.0 2116650.0 113700.0 2115450.0 ;
      RECT  112500.0 2116650.0 113700.0 2115450.0 ;
      RECT  110100.0 2116650.0 111300.0 2115450.0 ;
      RECT  114900.0 2106750.0 116100.0 2105550.0 ;
      RECT  114900.0 2116650.0 116100.0 2115450.0 ;
      RECT  110700.0 2112000.0 111900.0 2110800.0 ;
      RECT  110700.0 2112000.0 111900.0 2110800.0 ;
      RECT  113250.0 2111850.0 114150.0 2110950.0 ;
      RECT  108300.0 2104650.0 117900.0 2103750.0 ;
      RECT  108300.0 2118450.0 117900.0 2117550.0 ;
      RECT  114900.0 2129850.0 116100.0 2131800.0 ;
      RECT  114900.0 2118000.0 116100.0 2119950.0 ;
      RECT  110100.0 2119350.0 111300.0 2117550.0 ;
      RECT  110100.0 2128650.0 111300.0 2132250.0 ;
      RECT  112800.0 2119350.0 113700.0 2128650.0 ;
      RECT  110100.0 2128650.0 111300.0 2129850.0 ;
      RECT  112500.0 2128650.0 113700.0 2129850.0 ;
      RECT  112500.0 2128650.0 113700.0 2129850.0 ;
      RECT  110100.0 2128650.0 111300.0 2129850.0 ;
      RECT  110100.0 2119350.0 111300.0 2120550.0 ;
      RECT  112500.0 2119350.0 113700.0 2120550.0 ;
      RECT  112500.0 2119350.0 113700.0 2120550.0 ;
      RECT  110100.0 2119350.0 111300.0 2120550.0 ;
      RECT  114900.0 2129250.0 116100.0 2130450.0 ;
      RECT  114900.0 2119350.0 116100.0 2120550.0 ;
      RECT  110700.0 2124000.0 111900.0 2125200.0 ;
      RECT  110700.0 2124000.0 111900.0 2125200.0 ;
      RECT  113250.0 2124150.0 114150.0 2125050.0 ;
      RECT  108300.0 2131350.0 117900.0 2132250.0 ;
      RECT  108300.0 2117550.0 117900.0 2118450.0 ;
      RECT  114900.0 2133750.0 116100.0 2131800.0 ;
      RECT  114900.0 2145600.0 116100.0 2143650.0 ;
      RECT  110100.0 2144250.0 111300.0 2146050.0 ;
      RECT  110100.0 2134950.0 111300.0 2131350.0 ;
      RECT  112800.0 2144250.0 113700.0 2134950.0 ;
      RECT  110100.0 2134950.0 111300.0 2133750.0 ;
      RECT  112500.0 2134950.0 113700.0 2133750.0 ;
      RECT  112500.0 2134950.0 113700.0 2133750.0 ;
      RECT  110100.0 2134950.0 111300.0 2133750.0 ;
      RECT  110100.0 2144250.0 111300.0 2143050.0 ;
      RECT  112500.0 2144250.0 113700.0 2143050.0 ;
      RECT  112500.0 2144250.0 113700.0 2143050.0 ;
      RECT  110100.0 2144250.0 111300.0 2143050.0 ;
      RECT  114900.0 2134350.0 116100.0 2133150.0 ;
      RECT  114900.0 2144250.0 116100.0 2143050.0 ;
      RECT  110700.0 2139600.0 111900.0 2138400.0 ;
      RECT  110700.0 2139600.0 111900.0 2138400.0 ;
      RECT  113250.0 2139450.0 114150.0 2138550.0 ;
      RECT  108300.0 2132250.0 117900.0 2131350.0 ;
      RECT  108300.0 2146050.0 117900.0 2145150.0 ;
      RECT  60150.0 164400.0 58950.0 165600.0 ;
      RECT  62250.0 178800.0 61050.0 180000.0 ;
      RECT  64350.0 192000.0 63150.0 193200.0 ;
      RECT  66450.0 206400.0 65250.0 207600.0 ;
      RECT  68550.0 219600.0 67350.0 220800.0 ;
      RECT  70650.0 234000.0 69450.0 235200.0 ;
      RECT  72750.0 247200.0 71550.0 248400.0 ;
      RECT  74850.0 261600.0 73650.0 262800.0 ;
      RECT  76950.0 274800.0 75750.0 276000.0 ;
      RECT  79050.0 289200.0 77850.0 290400.0 ;
      RECT  81150.0 302400.0 79950.0 303600.0 ;
      RECT  83250.0 316800.0 82050.0 318000.0 ;
      RECT  85350.0 330000.0 84150.0 331200.0 ;
      RECT  87450.0 344400.0 86250.0 345600.0 ;
      RECT  89550.0 357600.0 88350.0 358800.0 ;
      RECT  91650.0 372000.0 90450.0 373200.0 ;
      RECT  60150.0 387150.0 58950.0 388350.0 ;
      RECT  68550.0 385200.0 67350.0 386400.0 ;
      RECT  76950.0 383250.0 75750.0 384450.0 ;
      RECT  60150.0 397650.0 58950.0 398850.0 ;
      RECT  68550.0 399600.0 67350.0 400800.0 ;
      RECT  79050.0 401550.0 77850.0 402750.0 ;
      RECT  60150.0 414750.0 58950.0 415950.0 ;
      RECT  68550.0 412800.0 67350.0 414000.0 ;
      RECT  81150.0 410850.0 79950.0 412050.0 ;
      RECT  60150.0 425250.0 58950.0 426450.0 ;
      RECT  68550.0 427200.0 67350.0 428400.0 ;
      RECT  83250.0 429150.0 82050.0 430350.0 ;
      RECT  60150.0 442350.0 58950.0 443550.0 ;
      RECT  68550.0 440400.0 67350.0 441600.0 ;
      RECT  85350.0 438450.0 84150.0 439650.0 ;
      RECT  60150.0 452850.0 58950.0 454050.0 ;
      RECT  68550.0 454800.0 67350.0 456000.0 ;
      RECT  87450.0 456750.0 86250.0 457950.0 ;
      RECT  60150.0 469950.0 58950.0 471150.0 ;
      RECT  68550.0 468000.0 67350.0 469200.0 ;
      RECT  89550.0 466050.0 88350.0 467250.0 ;
      RECT  60150.0 480450.0 58950.0 481650.0 ;
      RECT  68550.0 482400.0 67350.0 483600.0 ;
      RECT  91650.0 484350.0 90450.0 485550.0 ;
      RECT  60150.0 497550.0 58950.0 498750.0 ;
      RECT  70650.0 495600.0 69450.0 496800.0 ;
      RECT  76950.0 493650.0 75750.0 494850.0 ;
      RECT  60150.0 508050.0 58950.0 509250.0 ;
      RECT  70650.0 510000.0 69450.0 511200.0 ;
      RECT  79050.0 511950.0 77850.0 513150.0 ;
      RECT  60150.0 525150.0 58950.0 526350.0 ;
      RECT  70650.0 523200.0 69450.0 524400.0 ;
      RECT  81150.0 521250.0 79950.0 522450.0 ;
      RECT  60150.0 535650.0 58950.0 536850.0 ;
      RECT  70650.0 537600.0 69450.0 538800.0 ;
      RECT  83250.0 539550.0 82050.0 540750.0 ;
      RECT  60150.0 552750.0 58950.0 553950.0 ;
      RECT  70650.0 550800.0 69450.0 552000.0 ;
      RECT  85350.0 548850.0 84150.0 550050.0 ;
      RECT  60150.0 563250.0 58950.0 564450.0 ;
      RECT  70650.0 565200.0 69450.0 566400.0 ;
      RECT  87450.0 567150.0 86250.0 568350.0 ;
      RECT  60150.0 580350.0 58950.0 581550.0 ;
      RECT  70650.0 578400.0 69450.0 579600.0 ;
      RECT  89550.0 576450.0 88350.0 577650.0 ;
      RECT  60150.0 590850.0 58950.0 592050.0 ;
      RECT  70650.0 592800.0 69450.0 594000.0 ;
      RECT  91650.0 594750.0 90450.0 595950.0 ;
      RECT  60150.0 607950.0 58950.0 609150.0 ;
      RECT  72750.0 606000.0 71550.0 607200.0 ;
      RECT  76950.0 604050.0 75750.0 605250.0 ;
      RECT  60150.0 618450.0 58950.0 619650.0 ;
      RECT  72750.0 620400.0 71550.0 621600.0 ;
      RECT  79050.0 622350.0 77850.0 623550.0 ;
      RECT  60150.0 635550.0 58950.0 636750.0 ;
      RECT  72750.0 633600.0 71550.0 634800.0 ;
      RECT  81150.0 631650.0 79950.0 632850.0 ;
      RECT  60150.0 646050.0 58950.0 647250.0 ;
      RECT  72750.0 648000.0 71550.0 649200.0 ;
      RECT  83250.0 649950.0 82050.0 651150.0 ;
      RECT  60150.0 663150.0 58950.0 664350.0 ;
      RECT  72750.0 661200.0 71550.0 662400.0 ;
      RECT  85350.0 659250.0 84150.0 660450.0 ;
      RECT  60150.0 673650.0 58950.0 674850.0 ;
      RECT  72750.0 675600.0 71550.0 676800.0 ;
      RECT  87450.0 677550.0 86250.0 678750.0 ;
      RECT  60150.0 690750.0 58950.0 691950.0 ;
      RECT  72750.0 688800.0 71550.0 690000.0 ;
      RECT  89550.0 686850.0 88350.0 688050.0 ;
      RECT  60150.0 701250.0 58950.0 702450.0 ;
      RECT  72750.0 703200.0 71550.0 704400.0 ;
      RECT  91650.0 705150.0 90450.0 706350.0 ;
      RECT  60150.0 718350.0 58950.0 719550.0 ;
      RECT  74850.0 716400.0 73650.0 717600.0 ;
      RECT  76950.0 714450.0 75750.0 715650.0 ;
      RECT  60150.0 728850.0 58950.0 730050.0 ;
      RECT  74850.0 730800.0 73650.0 732000.0 ;
      RECT  79050.0 732750.0 77850.0 733950.0 ;
      RECT  60150.0 745950.0 58950.0 747150.0 ;
      RECT  74850.0 744000.0 73650.0 745200.0 ;
      RECT  81150.0 742050.0 79950.0 743250.0 ;
      RECT  60150.0 756450.0 58950.0 757650.0 ;
      RECT  74850.0 758400.0 73650.0 759600.0 ;
      RECT  83250.0 760350.0 82050.0 761550.0 ;
      RECT  60150.0 773550.0 58950.0 774750.0 ;
      RECT  74850.0 771600.0 73650.0 772800.0 ;
      RECT  85350.0 769650.0 84150.0 770850.0 ;
      RECT  60150.0 784050.0 58950.0 785250.0 ;
      RECT  74850.0 786000.0 73650.0 787200.0 ;
      RECT  87450.0 787950.0 86250.0 789150.0 ;
      RECT  60150.0 801150.0 58950.0 802350.0 ;
      RECT  74850.0 799200.0 73650.0 800400.0 ;
      RECT  89550.0 797250.0 88350.0 798450.0 ;
      RECT  60150.0 811650.0 58950.0 812850.0 ;
      RECT  74850.0 813600.0 73650.0 814800.0 ;
      RECT  91650.0 815550.0 90450.0 816750.0 ;
      RECT  62250.0 828750.0 61050.0 829950.0 ;
      RECT  68550.0 826800.0 67350.0 828000.0 ;
      RECT  76950.0 824850.0 75750.0 826050.0 ;
      RECT  62250.0 839250.0 61050.0 840450.0 ;
      RECT  68550.0 841200.0 67350.0 842400.0 ;
      RECT  79050.0 843150.0 77850.0 844350.0 ;
      RECT  62250.0 856350.0 61050.0 857550.0 ;
      RECT  68550.0 854400.0 67350.0 855600.0 ;
      RECT  81150.0 852450.0 79950.0 853650.0 ;
      RECT  62250.0 866850.0 61050.0 868050.0 ;
      RECT  68550.0 868800.0 67350.0 870000.0 ;
      RECT  83250.0 870750.0 82050.0 871950.0 ;
      RECT  62250.0 883950.0 61050.0 885150.0 ;
      RECT  68550.0 882000.0 67350.0 883200.0 ;
      RECT  85350.0 880050.0 84150.0 881250.0 ;
      RECT  62250.0 894450.0 61050.0 895650.0 ;
      RECT  68550.0 896400.0 67350.0 897600.0 ;
      RECT  87450.0 898350.0 86250.0 899550.0 ;
      RECT  62250.0 911550.0 61050.0 912750.0 ;
      RECT  68550.0 909600.0 67350.0 910800.0 ;
      RECT  89550.0 907650.0 88350.0 908850.0 ;
      RECT  62250.0 922050.0 61050.0 923250.0 ;
      RECT  68550.0 924000.0 67350.0 925200.0 ;
      RECT  91650.0 925950.0 90450.0 927150.0 ;
      RECT  62250.0 939150.0 61050.0 940350.0 ;
      RECT  70650.0 937200.0 69450.0 938400.0 ;
      RECT  76950.0 935250.0 75750.0 936450.0 ;
      RECT  62250.0 949650.0 61050.0 950850.0 ;
      RECT  70650.0 951600.0 69450.0 952800.0 ;
      RECT  79050.0 953550.0 77850.0 954750.0 ;
      RECT  62250.0 966750.0 61050.0 967950.0 ;
      RECT  70650.0 964800.0 69450.0 966000.0 ;
      RECT  81150.0 962850.0 79950.0 964050.0 ;
      RECT  62250.0 977250.0 61050.0 978450.0 ;
      RECT  70650.0 979200.0 69450.0 980400.0 ;
      RECT  83250.0 981150.0 82050.0 982350.0 ;
      RECT  62250.0 994350.0 61050.0 995550.0 ;
      RECT  70650.0 992400.0 69450.0 993600.0 ;
      RECT  85350.0 990450.0 84150.0 991650.0 ;
      RECT  62250.0 1004850.0 61050.0 1006050.0 ;
      RECT  70650.0 1006800.0 69450.0 1008000.0 ;
      RECT  87450.0 1008750.0 86250.0 1009950.0 ;
      RECT  62250.0 1021950.0 61050.0 1023150.0 ;
      RECT  70650.0 1020000.0 69450.0 1021200.0 ;
      RECT  89550.0 1018050.0 88350.0 1019250.0 ;
      RECT  62250.0 1032450.0 61050.0 1033650.0 ;
      RECT  70650.0 1034400.0 69450.0 1035600.0 ;
      RECT  91650.0 1036350.0 90450.0 1037550.0 ;
      RECT  62250.0 1049550.0 61050.0 1050750.0 ;
      RECT  72750.0 1047600.0 71550.0 1048800.0 ;
      RECT  76950.0 1045650.0 75750.0 1046850.0 ;
      RECT  62250.0 1060050.0 61050.0 1061250.0 ;
      RECT  72750.0 1062000.0 71550.0 1063200.0 ;
      RECT  79050.0 1063950.0 77850.0 1065150.0 ;
      RECT  62250.0 1077150.0 61050.0 1078350.0 ;
      RECT  72750.0 1075200.0 71550.0 1076400.0 ;
      RECT  81150.0 1073250.0 79950.0 1074450.0 ;
      RECT  62250.0 1087650.0 61050.0 1088850.0 ;
      RECT  72750.0 1089600.0 71550.0 1090800.0 ;
      RECT  83250.0 1091550.0 82050.0 1092750.0 ;
      RECT  62250.0 1104750.0 61050.0 1105950.0 ;
      RECT  72750.0 1102800.0 71550.0 1104000.0 ;
      RECT  85350.0 1100850.0 84150.0 1102050.0 ;
      RECT  62250.0 1115250.0 61050.0 1116450.0 ;
      RECT  72750.0 1117200.0 71550.0 1118400.0 ;
      RECT  87450.0 1119150.0 86250.0 1120350.0 ;
      RECT  62250.0 1132350.0 61050.0 1133550.0 ;
      RECT  72750.0 1130400.0 71550.0 1131600.0 ;
      RECT  89550.0 1128450.0 88350.0 1129650.0 ;
      RECT  62250.0 1142850.0 61050.0 1144050.0 ;
      RECT  72750.0 1144800.0 71550.0 1146000.0 ;
      RECT  91650.0 1146750.0 90450.0 1147950.0 ;
      RECT  62250.0 1159950.0 61050.0 1161150.0 ;
      RECT  74850.0 1158000.0 73650.0 1159200.0 ;
      RECT  76950.0 1156050.0 75750.0 1157250.0 ;
      RECT  62250.0 1170450.0 61050.0 1171650.0 ;
      RECT  74850.0 1172400.0 73650.0 1173600.0 ;
      RECT  79050.0 1174350.0 77850.0 1175550.0 ;
      RECT  62250.0 1187550.0 61050.0 1188750.0 ;
      RECT  74850.0 1185600.0 73650.0 1186800.0 ;
      RECT  81150.0 1183650.0 79950.0 1184850.0 ;
      RECT  62250.0 1198050.0 61050.0 1199250.0 ;
      RECT  74850.0 1200000.0 73650.0 1201200.0 ;
      RECT  83250.0 1201950.0 82050.0 1203150.0 ;
      RECT  62250.0 1215150.0 61050.0 1216350.0 ;
      RECT  74850.0 1213200.0 73650.0 1214400.0 ;
      RECT  85350.0 1211250.0 84150.0 1212450.0 ;
      RECT  62250.0 1225650.0 61050.0 1226850.0 ;
      RECT  74850.0 1227600.0 73650.0 1228800.0 ;
      RECT  87450.0 1229550.0 86250.0 1230750.0 ;
      RECT  62250.0 1242750.0 61050.0 1243950.0 ;
      RECT  74850.0 1240800.0 73650.0 1242000.0 ;
      RECT  89550.0 1238850.0 88350.0 1240050.0 ;
      RECT  62250.0 1253250.0 61050.0 1254450.0 ;
      RECT  74850.0 1255200.0 73650.0 1256400.0 ;
      RECT  91650.0 1257150.0 90450.0 1258350.0 ;
      RECT  64350.0 1270350.0 63150.0 1271550.0 ;
      RECT  68550.0 1268400.0 67350.0 1269600.0 ;
      RECT  76950.0 1266450.0 75750.0 1267650.0 ;
      RECT  64350.0 1280850.0 63150.0 1282050.0 ;
      RECT  68550.0 1282800.0 67350.0 1284000.0 ;
      RECT  79050.0 1284750.0 77850.0 1285950.0 ;
      RECT  64350.0 1297950.0 63150.0 1299150.0 ;
      RECT  68550.0 1296000.0 67350.0 1297200.0 ;
      RECT  81150.0 1294050.0 79950.0 1295250.0 ;
      RECT  64350.0 1308450.0 63150.0 1309650.0 ;
      RECT  68550.0 1310400.0 67350.0 1311600.0 ;
      RECT  83250.0 1312350.0 82050.0 1313550.0 ;
      RECT  64350.0 1325550.0 63150.0 1326750.0 ;
      RECT  68550.0 1323600.0 67350.0 1324800.0 ;
      RECT  85350.0 1321650.0 84150.0 1322850.0 ;
      RECT  64350.0 1336050.0 63150.0 1337250.0 ;
      RECT  68550.0 1338000.0 67350.0 1339200.0 ;
      RECT  87450.0 1339950.0 86250.0 1341150.0 ;
      RECT  64350.0 1353150.0 63150.0 1354350.0 ;
      RECT  68550.0 1351200.0 67350.0 1352400.0 ;
      RECT  89550.0 1349250.0 88350.0 1350450.0 ;
      RECT  64350.0 1363650.0 63150.0 1364850.0 ;
      RECT  68550.0 1365600.0 67350.0 1366800.0 ;
      RECT  91650.0 1367550.0 90450.0 1368750.0 ;
      RECT  64350.0 1380750.0 63150.0 1381950.0 ;
      RECT  70650.0 1378800.0 69450.0 1380000.0 ;
      RECT  76950.0 1376850.0 75750.0 1378050.0 ;
      RECT  64350.0 1391250.0 63150.0 1392450.0 ;
      RECT  70650.0 1393200.0 69450.0 1394400.0 ;
      RECT  79050.0 1395150.0 77850.0 1396350.0 ;
      RECT  64350.0 1408350.0 63150.0 1409550.0 ;
      RECT  70650.0 1406400.0 69450.0 1407600.0 ;
      RECT  81150.0 1404450.0 79950.0 1405650.0 ;
      RECT  64350.0 1418850.0 63150.0 1420050.0 ;
      RECT  70650.0 1420800.0 69450.0 1422000.0 ;
      RECT  83250.0 1422750.0 82050.0 1423950.0 ;
      RECT  64350.0 1435950.0 63150.0 1437150.0 ;
      RECT  70650.0 1434000.0 69450.0 1435200.0 ;
      RECT  85350.0 1432050.0 84150.0 1433250.0 ;
      RECT  64350.0 1446450.0 63150.0 1447650.0 ;
      RECT  70650.0 1448400.0 69450.0 1449600.0 ;
      RECT  87450.0 1450350.0 86250.0 1451550.0 ;
      RECT  64350.0 1463550.0 63150.0 1464750.0 ;
      RECT  70650.0 1461600.0 69450.0 1462800.0 ;
      RECT  89550.0 1459650.0 88350.0 1460850.0 ;
      RECT  64350.0 1474050.0 63150.0 1475250.0 ;
      RECT  70650.0 1476000.0 69450.0 1477200.0 ;
      RECT  91650.0 1477950.0 90450.0 1479150.0 ;
      RECT  64350.0 1491150.0 63150.0 1492350.0 ;
      RECT  72750.0 1489200.0 71550.0 1490400.0 ;
      RECT  76950.0 1487250.0 75750.0 1488450.0 ;
      RECT  64350.0 1501650.0 63150.0 1502850.0 ;
      RECT  72750.0 1503600.0 71550.0 1504800.0 ;
      RECT  79050.0 1505550.0 77850.0 1506750.0 ;
      RECT  64350.0 1518750.0 63150.0 1519950.0 ;
      RECT  72750.0 1516800.0 71550.0 1518000.0 ;
      RECT  81150.0 1514850.0 79950.0 1516050.0 ;
      RECT  64350.0 1529250.0 63150.0 1530450.0 ;
      RECT  72750.0 1531200.0 71550.0 1532400.0 ;
      RECT  83250.0 1533150.0 82050.0 1534350.0 ;
      RECT  64350.0 1546350.0 63150.0 1547550.0 ;
      RECT  72750.0 1544400.0 71550.0 1545600.0 ;
      RECT  85350.0 1542450.0 84150.0 1543650.0 ;
      RECT  64350.0 1556850.0 63150.0 1558050.0 ;
      RECT  72750.0 1558800.0 71550.0 1560000.0 ;
      RECT  87450.0 1560750.0 86250.0 1561950.0 ;
      RECT  64350.0 1573950.0 63150.0 1575150.0 ;
      RECT  72750.0 1572000.0 71550.0 1573200.0 ;
      RECT  89550.0 1570050.0 88350.0 1571250.0 ;
      RECT  64350.0 1584450.0 63150.0 1585650.0 ;
      RECT  72750.0 1586400.0 71550.0 1587600.0 ;
      RECT  91650.0 1588350.0 90450.0 1589550.0 ;
      RECT  64350.0 1601550.0 63150.0 1602750.0 ;
      RECT  74850.0 1599600.0 73650.0 1600800.0 ;
      RECT  76950.0 1597650.0 75750.0 1598850.0 ;
      RECT  64350.0 1612050.0 63150.0 1613250.0 ;
      RECT  74850.0 1614000.0 73650.0 1615200.0 ;
      RECT  79050.0 1615950.0 77850.0 1617150.0 ;
      RECT  64350.0 1629150.0 63150.0 1630350.0 ;
      RECT  74850.0 1627200.0 73650.0 1628400.0 ;
      RECT  81150.0 1625250.0 79950.0 1626450.0 ;
      RECT  64350.0 1639650.0 63150.0 1640850.0 ;
      RECT  74850.0 1641600.0 73650.0 1642800.0 ;
      RECT  83250.0 1643550.0 82050.0 1644750.0 ;
      RECT  64350.0 1656750.0 63150.0 1657950.0 ;
      RECT  74850.0 1654800.0 73650.0 1656000.0 ;
      RECT  85350.0 1652850.0 84150.0 1654050.0 ;
      RECT  64350.0 1667250.0 63150.0 1668450.0 ;
      RECT  74850.0 1669200.0 73650.0 1670400.0 ;
      RECT  87450.0 1671150.0 86250.0 1672350.0 ;
      RECT  64350.0 1684350.0 63150.0 1685550.0 ;
      RECT  74850.0 1682400.0 73650.0 1683600.0 ;
      RECT  89550.0 1680450.0 88350.0 1681650.0 ;
      RECT  64350.0 1694850.0 63150.0 1696050.0 ;
      RECT  74850.0 1696800.0 73650.0 1698000.0 ;
      RECT  91650.0 1698750.0 90450.0 1699950.0 ;
      RECT  66450.0 1711950.0 65250.0 1713150.0 ;
      RECT  68550.0 1710000.0 67350.0 1711200.0 ;
      RECT  76950.0 1708050.0 75750.0 1709250.0 ;
      RECT  66450.0 1722450.0 65250.0 1723650.0 ;
      RECT  68550.0 1724400.0 67350.0 1725600.0 ;
      RECT  79050.0 1726350.0 77850.0 1727550.0 ;
      RECT  66450.0 1739550.0 65250.0 1740750.0 ;
      RECT  68550.0 1737600.0 67350.0 1738800.0 ;
      RECT  81150.0 1735650.0 79950.0 1736850.0 ;
      RECT  66450.0 1750050.0 65250.0 1751250.0 ;
      RECT  68550.0 1752000.0 67350.0 1753200.0 ;
      RECT  83250.0 1753950.0 82050.0 1755150.0 ;
      RECT  66450.0 1767150.0 65250.0 1768350.0 ;
      RECT  68550.0 1765200.0 67350.0 1766400.0 ;
      RECT  85350.0 1763250.0 84150.0 1764450.0 ;
      RECT  66450.0 1777650.0 65250.0 1778850.0 ;
      RECT  68550.0 1779600.0 67350.0 1780800.0 ;
      RECT  87450.0 1781550.0 86250.0 1782750.0 ;
      RECT  66450.0 1794750.0 65250.0 1795950.0 ;
      RECT  68550.0 1792800.0 67350.0 1794000.0 ;
      RECT  89550.0 1790850.0 88350.0 1792050.0 ;
      RECT  66450.0 1805250.0 65250.0 1806450.0 ;
      RECT  68550.0 1807200.0 67350.0 1808400.0 ;
      RECT  91650.0 1809150.0 90450.0 1810350.0 ;
      RECT  66450.0 1822350.0 65250.0 1823550.0 ;
      RECT  70650.0 1820400.0 69450.0 1821600.0 ;
      RECT  76950.0 1818450.0 75750.0 1819650.0 ;
      RECT  66450.0 1832850.0 65250.0 1834050.0 ;
      RECT  70650.0 1834800.0 69450.0 1836000.0 ;
      RECT  79050.0 1836750.0 77850.0 1837950.0 ;
      RECT  66450.0 1849950.0 65250.0 1851150.0 ;
      RECT  70650.0 1848000.0 69450.0 1849200.0 ;
      RECT  81150.0 1846050.0 79950.0 1847250.0 ;
      RECT  66450.0 1860450.0 65250.0 1861650.0 ;
      RECT  70650.0 1862400.0 69450.0 1863600.0 ;
      RECT  83250.0 1864350.0 82050.0 1865550.0 ;
      RECT  66450.0 1877550.0 65250.0 1878750.0 ;
      RECT  70650.0 1875600.0 69450.0 1876800.0 ;
      RECT  85350.0 1873650.0 84150.0 1874850.0 ;
      RECT  66450.0 1888050.0 65250.0 1889250.0 ;
      RECT  70650.0 1890000.0 69450.0 1891200.0 ;
      RECT  87450.0 1891950.0 86250.0 1893150.0 ;
      RECT  66450.0 1905150.0 65250.0 1906350.0 ;
      RECT  70650.0 1903200.0 69450.0 1904400.0 ;
      RECT  89550.0 1901250.0 88350.0 1902450.0 ;
      RECT  66450.0 1915650.0 65250.0 1916850.0 ;
      RECT  70650.0 1917600.0 69450.0 1918800.0 ;
      RECT  91650.0 1919550.0 90450.0 1920750.0 ;
      RECT  66450.0 1932750.0 65250.0 1933950.0 ;
      RECT  72750.0 1930800.0 71550.0 1932000.0 ;
      RECT  76950.0 1928850.0 75750.0 1930050.0 ;
      RECT  66450.0 1943250.0 65250.0 1944450.0 ;
      RECT  72750.0 1945200.0 71550.0 1946400.0 ;
      RECT  79050.0 1947150.0 77850.0 1948350.0 ;
      RECT  66450.0 1960350.0 65250.0 1961550.0 ;
      RECT  72750.0 1958400.0 71550.0 1959600.0 ;
      RECT  81150.0 1956450.0 79950.0 1957650.0 ;
      RECT  66450.0 1970850.0 65250.0 1972050.0 ;
      RECT  72750.0 1972800.0 71550.0 1974000.0 ;
      RECT  83250.0 1974750.0 82050.0 1975950.0 ;
      RECT  66450.0 1987950.0 65250.0 1989150.0 ;
      RECT  72750.0 1986000.0 71550.0 1987200.0 ;
      RECT  85350.0 1984050.0 84150.0 1985250.0 ;
      RECT  66450.0 1998450.0 65250.0 1999650.0 ;
      RECT  72750.0 2000400.0 71550.0 2001600.0 ;
      RECT  87450.0 2002350.0 86250.0 2003550.0 ;
      RECT  66450.0 2015550.0 65250.0 2016750.0 ;
      RECT  72750.0 2013600.0 71550.0 2014800.0 ;
      RECT  89550.0 2011650.0 88350.0 2012850.0 ;
      RECT  66450.0 2026050.0 65250.0 2027250.0 ;
      RECT  72750.0 2028000.0 71550.0 2029200.0 ;
      RECT  91650.0 2029950.0 90450.0 2031150.0 ;
      RECT  66450.0 2043150.0 65250.0 2044350.0 ;
      RECT  74850.0 2041200.0 73650.0 2042400.0 ;
      RECT  76950.0 2039250.0 75750.0 2040450.0 ;
      RECT  66450.0 2053650.0 65250.0 2054850.0 ;
      RECT  74850.0 2055600.0 73650.0 2056800.0 ;
      RECT  79050.0 2057550.0 77850.0 2058750.0 ;
      RECT  66450.0 2070750.0 65250.0 2071950.0 ;
      RECT  74850.0 2068800.0 73650.0 2070000.0 ;
      RECT  81150.0 2066850.0 79950.0 2068050.0 ;
      RECT  66450.0 2081250.0 65250.0 2082450.0 ;
      RECT  74850.0 2083200.0 73650.0 2084400.0 ;
      RECT  83250.0 2085150.0 82050.0 2086350.0 ;
      RECT  66450.0 2098350.0 65250.0 2099550.0 ;
      RECT  74850.0 2096400.0 73650.0 2097600.0 ;
      RECT  85350.0 2094450.0 84150.0 2095650.0 ;
      RECT  66450.0 2108850.0 65250.0 2110050.0 ;
      RECT  74850.0 2110800.0 73650.0 2112000.0 ;
      RECT  87450.0 2112750.0 86250.0 2113950.0 ;
      RECT  66450.0 2125950.0 65250.0 2127150.0 ;
      RECT  74850.0 2124000.0 73650.0 2125200.0 ;
      RECT  89550.0 2122050.0 88350.0 2123250.0 ;
      RECT  66450.0 2136450.0 65250.0 2137650.0 ;
      RECT  74850.0 2138400.0 73650.0 2139600.0 ;
      RECT  91650.0 2140350.0 90450.0 2141550.0 ;
      RECT  113250.0 385350.0 114150.0 386250.0 ;
      RECT  113250.0 399750.0 114150.0 400650.0 ;
      RECT  113250.0 412950.0 114150.0 413850.0 ;
      RECT  113250.0 427350.0 114150.0 428250.0 ;
      RECT  113250.0 440550.0 114150.0 441450.0 ;
      RECT  113250.0 454950.0 114150.0 455850.0 ;
      RECT  113250.0 468150.0 114150.0 469050.0 ;
      RECT  113250.0 482550.0 114150.0 483450.0 ;
      RECT  113250.0 495750.0 114150.0 496650.0 ;
      RECT  113250.0 510150.0 114150.0 511050.0 ;
      RECT  113250.0 523350.0 114150.0 524250.0 ;
      RECT  113250.0 537750.0 114150.0 538650.0 ;
      RECT  113250.0 550950.0 114150.0 551850.0 ;
      RECT  113250.0 565350.0 114150.0 566250.0 ;
      RECT  113250.0 578550.0 114150.0 579450.0 ;
      RECT  113250.0 592950.0 114150.0 593850.0 ;
      RECT  113250.0 606150.0 114150.0 607050.0 ;
      RECT  113250.0 620550.0 114150.0 621450.0 ;
      RECT  113250.0 633750.0 114150.0 634650.0 ;
      RECT  113250.0 648150.0 114150.0 649050.0 ;
      RECT  113250.0 661350.0 114150.0 662250.0 ;
      RECT  113250.0 675750.0 114150.0 676650.0 ;
      RECT  113250.0 688950.0 114150.0 689850.0 ;
      RECT  113250.0 703350.0 114150.0 704250.0 ;
      RECT  113250.0 716550.0 114150.0 717450.0 ;
      RECT  113250.0 730950.0 114150.0 731850.0 ;
      RECT  113250.0 744150.0 114150.0 745050.0 ;
      RECT  113250.0 758550.0 114150.0 759450.0 ;
      RECT  113250.0 771750.0 114150.0 772650.0 ;
      RECT  113250.0 786150.0 114150.0 787050.0 ;
      RECT  113250.0 799350.0 114150.0 800250.0 ;
      RECT  113250.0 813750.0 114150.0 814650.0 ;
      RECT  113250.0 826950.0 114150.0 827850.0 ;
      RECT  113250.0 841350.0 114150.0 842250.0 ;
      RECT  113250.0 854550.0 114150.0 855450.0 ;
      RECT  113250.0 868950.0 114150.0 869850.0 ;
      RECT  113250.0 882150.0 114150.0 883050.0 ;
      RECT  113250.0 896550.0 114150.0 897450.0 ;
      RECT  113250.0 909750.0 114150.0 910650.0 ;
      RECT  113250.0 924150.0 114150.0 925050.0 ;
      RECT  113250.0 937350.0 114150.0 938250.0 ;
      RECT  113250.0 951750.0 114150.0 952650.0 ;
      RECT  113250.0 964950.0 114150.0 965850.0 ;
      RECT  113250.0 979350.0 114150.0 980250.0 ;
      RECT  113250.0 992550.0 114150.0 993450.0 ;
      RECT  113250.0 1006950.0 114150.0 1007850.0 ;
      RECT  113250.0 1020150.0 114150.0 1021050.0 ;
      RECT  113250.0 1034550.0 114150.0 1035450.0 ;
      RECT  113250.0 1047750.0 114150.0 1048650.0 ;
      RECT  113250.0 1062150.0 114150.0 1063050.0 ;
      RECT  113250.0 1075350.0 114150.0 1076250.0 ;
      RECT  113250.0 1089750.0 114150.0 1090650.0 ;
      RECT  113250.0 1102950.0 114150.0 1103850.0 ;
      RECT  113250.0 1117350.0 114150.0 1118250.0 ;
      RECT  113250.0 1130550.0 114150.0 1131450.0 ;
      RECT  113250.0 1144950.0 114150.0 1145850.0 ;
      RECT  113250.0 1158150.0 114150.0 1159050.0 ;
      RECT  113250.0 1172550.0 114150.0 1173450.0 ;
      RECT  113250.0 1185750.0 114150.0 1186650.0 ;
      RECT  113250.0 1200150.0 114150.0 1201050.0 ;
      RECT  113250.0 1213350.0 114150.0 1214250.0 ;
      RECT  113250.0 1227750.0 114150.0 1228650.0 ;
      RECT  113250.0 1240950.0 114150.0 1241850.0 ;
      RECT  113250.0 1255350.0 114150.0 1256250.0 ;
      RECT  113250.0 1268550.0 114150.0 1269450.0 ;
      RECT  113250.0 1282950.0 114150.0 1283850.0 ;
      RECT  113250.0 1296150.0 114150.0 1297050.0 ;
      RECT  113250.0 1310550.0 114150.0 1311450.0 ;
      RECT  113250.0 1323750.0 114150.0 1324650.0 ;
      RECT  113250.0 1338150.0 114150.0 1339050.0 ;
      RECT  113250.0 1351350.0 114150.0 1352250.0 ;
      RECT  113250.0 1365750.0 114150.0 1366650.0 ;
      RECT  113250.0 1378950.0 114150.0 1379850.0 ;
      RECT  113250.0 1393350.0 114150.0 1394250.0 ;
      RECT  113250.0 1406550.0 114150.0 1407450.0 ;
      RECT  113250.0 1420950.0 114150.0 1421850.0 ;
      RECT  113250.0 1434150.0 114150.0 1435050.0 ;
      RECT  113250.0 1448550.0 114150.0 1449450.0 ;
      RECT  113250.0 1461750.0 114150.0 1462650.0 ;
      RECT  113250.0 1476150.0 114150.0 1477050.0 ;
      RECT  113250.0 1489350.0 114150.0 1490250.0 ;
      RECT  113250.0 1503750.0 114150.0 1504650.0 ;
      RECT  113250.0 1516950.0 114150.0 1517850.0 ;
      RECT  113250.0 1531350.0 114150.0 1532250.0 ;
      RECT  113250.0 1544550.0 114150.0 1545450.0 ;
      RECT  113250.0 1558950.0 114150.0 1559850.0 ;
      RECT  113250.0 1572150.0 114150.0 1573050.0 ;
      RECT  113250.0 1586550.0 114150.0 1587450.0 ;
      RECT  113250.0 1599750.0 114150.0 1600650.0 ;
      RECT  113250.0 1614150.0 114150.0 1615050.0 ;
      RECT  113250.0 1627350.0 114150.0 1628250.0 ;
      RECT  113250.0 1641750.0 114150.0 1642650.0 ;
      RECT  113250.0 1654950.0 114150.0 1655850.0 ;
      RECT  113250.0 1669350.0 114150.0 1670250.0 ;
      RECT  113250.0 1682550.0 114150.0 1683450.0 ;
      RECT  113250.0 1696950.0 114150.0 1697850.0 ;
      RECT  113250.0 1710150.0 114150.0 1711050.0 ;
      RECT  113250.0 1724550.0 114150.0 1725450.0 ;
      RECT  113250.0 1737750.0 114150.0 1738650.0 ;
      RECT  113250.0 1752150.0 114150.0 1753050.0 ;
      RECT  113250.0 1765350.0 114150.0 1766250.0 ;
      RECT  113250.0 1779750.0 114150.0 1780650.0 ;
      RECT  113250.0 1792950.0 114150.0 1793850.0 ;
      RECT  113250.0 1807350.0 114150.0 1808250.0 ;
      RECT  113250.0 1820550.0 114150.0 1821450.0 ;
      RECT  113250.0 1834950.0 114150.0 1835850.0 ;
      RECT  113250.0 1848150.0 114150.0 1849050.0 ;
      RECT  113250.0 1862550.0 114150.0 1863450.0 ;
      RECT  113250.0 1875750.0 114150.0 1876650.0 ;
      RECT  113250.0 1890150.0 114150.0 1891050.0 ;
      RECT  113250.0 1903350.0 114150.0 1904250.0 ;
      RECT  113250.0 1917750.0 114150.0 1918650.0 ;
      RECT  113250.0 1930950.0 114150.0 1931850.0 ;
      RECT  113250.0 1945350.0 114150.0 1946250.0 ;
      RECT  113250.0 1958550.0 114150.0 1959450.0 ;
      RECT  113250.0 1972950.0 114150.0 1973850.0 ;
      RECT  113250.0 1986150.0 114150.0 1987050.0 ;
      RECT  113250.0 2000550.0 114150.0 2001450.0 ;
      RECT  113250.0 2013750.0 114150.0 2014650.0 ;
      RECT  113250.0 2028150.0 114150.0 2029050.0 ;
      RECT  113250.0 2041350.0 114150.0 2042250.0 ;
      RECT  113250.0 2055750.0 114150.0 2056650.0 ;
      RECT  113250.0 2068950.0 114150.0 2069850.0 ;
      RECT  113250.0 2083350.0 114150.0 2084250.0 ;
      RECT  113250.0 2096550.0 114150.0 2097450.0 ;
      RECT  113250.0 2110950.0 114150.0 2111850.0 ;
      RECT  113250.0 2124150.0 114150.0 2125050.0 ;
      RECT  113250.0 2138550.0 114150.0 2139450.0 ;
      RECT  59100.0 171750.0 157500.0 172650.0 ;
      RECT  59100.0 199350.0 157500.0 200250.0 ;
      RECT  59100.0 226950.0 157500.0 227850.0 ;
      RECT  59100.0 254550.0 157500.0 255450.0 ;
      RECT  59100.0 282150.0 157500.0 283050.0 ;
      RECT  59100.0 309750.0 157500.0 310650.0 ;
      RECT  59100.0 337350.0 157500.0 338250.0 ;
      RECT  59100.0 364950.0 157500.0 365850.0 ;
      RECT  59100.0 392550.0 157500.0 393450.0 ;
      RECT  59100.0 420150.0 157500.0 421050.0 ;
      RECT  59100.0 447750.0 157500.0 448650.0 ;
      RECT  59100.0 475350.0 157500.0 476250.0 ;
      RECT  59100.0 502950.0 157500.0 503850.0 ;
      RECT  59100.0 530550.0 157500.0 531450.0 ;
      RECT  59100.0 558150.0 157500.0 559050.0 ;
      RECT  59100.0 585750.0 157500.0 586650.0 ;
      RECT  59100.0 613350.0 157500.0 614250.0 ;
      RECT  59100.0 640950.0 157500.0 641850.0 ;
      RECT  59100.0 668550.0 157500.0 669450.0 ;
      RECT  59100.0 696150.0 157500.0 697050.0 ;
      RECT  59100.0 723750.0 157500.0 724650.0 ;
      RECT  59100.0 751350.0 157500.0 752250.0 ;
      RECT  59100.0 778950.0 157500.0 779850.0 ;
      RECT  59100.0 806550.0 157500.0 807450.0 ;
      RECT  59100.0 834150.0 157500.0 835050.0 ;
      RECT  59100.0 861750.0 157500.0 862650.0 ;
      RECT  59100.0 889350.0 157500.0 890250.0 ;
      RECT  59100.0 916950.0 157500.0 917850.0 ;
      RECT  59100.0 944550.0 157500.0 945450.0 ;
      RECT  59100.0 972150.0 157500.0 973050.0 ;
      RECT  59100.0 999750.0 157500.0 1000650.0 ;
      RECT  59100.0 1027350.0 157500.0 1028250.0 ;
      RECT  59100.0 1054950.0 157500.0 1055850.0 ;
      RECT  59100.0 1082550.0 157500.0 1083450.0 ;
      RECT  59100.0 1110150.0 157500.0 1111050.0 ;
      RECT  59100.0 1137750.0 157500.0 1138650.0 ;
      RECT  59100.0 1165350.0 157500.0 1166250.0 ;
      RECT  59100.0 1192950.0 157500.0 1193850.0 ;
      RECT  59100.0 1220550.0 157500.0 1221450.0 ;
      RECT  59100.0 1248150.0 157500.0 1249050.0 ;
      RECT  59100.0 1275750.0 157500.0 1276650.0 ;
      RECT  59100.0 1303350.0 157500.0 1304250.0 ;
      RECT  59100.0 1330950.0 157500.0 1331850.0 ;
      RECT  59100.0 1358550.0 157500.0 1359450.0 ;
      RECT  59100.0 1386150.0 157500.0 1387050.0 ;
      RECT  59100.0 1413750.0 157500.0 1414650.0 ;
      RECT  59100.0 1441350.0 157500.0 1442250.0 ;
      RECT  59100.0 1468950.0 157500.0 1469850.0 ;
      RECT  59100.0 1496550.0 157500.0 1497450.0 ;
      RECT  59100.0 1524150.0 157500.0 1525050.0 ;
      RECT  59100.0 1551750.0 157500.0 1552650.0 ;
      RECT  59100.0 1579350.0 157500.0 1580250.0 ;
      RECT  59100.0 1606950.0 157500.0 1607850.0 ;
      RECT  59100.0 1634550.0 157500.0 1635450.0 ;
      RECT  59100.0 1662150.0 157500.0 1663050.0 ;
      RECT  59100.0 1689750.0 157500.0 1690650.0 ;
      RECT  59100.0 1717350.0 157500.0 1718250.0 ;
      RECT  59100.0 1744950.0 157500.0 1745850.0 ;
      RECT  59100.0 1772550.0 157500.0 1773450.0 ;
      RECT  59100.0 1800150.0 157500.0 1801050.0 ;
      RECT  59100.0 1827750.0 157500.0 1828650.0 ;
      RECT  59100.0 1855350.0 157500.0 1856250.0 ;
      RECT  59100.0 1882950.0 157500.0 1883850.0 ;
      RECT  59100.0 1910550.0 157500.0 1911450.0 ;
      RECT  59100.0 1938150.0 157500.0 1939050.0 ;
      RECT  59100.0 1965750.0 157500.0 1966650.0 ;
      RECT  59100.0 1993350.0 157500.0 1994250.0 ;
      RECT  59100.0 2020950.0 157500.0 2021850.0 ;
      RECT  59100.0 2048550.0 157500.0 2049450.0 ;
      RECT  59100.0 2076150.0 157500.0 2077050.0 ;
      RECT  59100.0 2103750.0 157500.0 2104650.0 ;
      RECT  59100.0 2131350.0 157500.0 2132250.0 ;
      RECT  59100.0 157950.0 157500.0 158850.0 ;
      RECT  59100.0 185550.0 157500.0 186450.0 ;
      RECT  59100.0 213150.0 157500.0 214050.0 ;
      RECT  59100.0 240750.0 157500.0 241650.0 ;
      RECT  59100.0 268350.0 157500.0 269250.0 ;
      RECT  59100.0 295950.0 157500.0 296850.0 ;
      RECT  59100.0 323550.0 157500.0 324450.0 ;
      RECT  59100.0 351150.0 157500.0 352050.0 ;
      RECT  59100.0 378750.0 157500.0 379650.0 ;
      RECT  59100.0 406350.0 157500.0 407250.0 ;
      RECT  59100.0 433950.0 157500.0 434850.0 ;
      RECT  59100.0 461550.0 157500.0 462450.0 ;
      RECT  59100.0 489150.0 157500.0 490050.0 ;
      RECT  59100.0 516750.0 157500.0 517650.0 ;
      RECT  59100.0 544350.0 157500.0 545250.0 ;
      RECT  59100.0 571950.0 157500.0 572850.0 ;
      RECT  59100.0 599550.0 157500.0 600450.0 ;
      RECT  59100.0 627150.0 157500.0 628050.0 ;
      RECT  59100.0 654750.0 157500.0 655650.0 ;
      RECT  59100.0 682350.0 157500.0 683250.0 ;
      RECT  59100.0 709950.0 157500.0 710850.0 ;
      RECT  59100.0 737550.0 157500.0 738450.0 ;
      RECT  59100.0 765150.0 157500.0 766050.0 ;
      RECT  59100.0 792750.0 157500.0 793650.0 ;
      RECT  59100.0 820350.0 157500.0 821250.0 ;
      RECT  59100.0 847950.0 157500.0 848850.0 ;
      RECT  59100.0 875550.0 157500.0 876450.0 ;
      RECT  59100.0 903150.0 157500.0 904050.0 ;
      RECT  59100.0 930750.0 157500.0 931650.0 ;
      RECT  59100.0 958350.0 157500.0 959250.0 ;
      RECT  59100.0 985950.0 157500.0 986850.0 ;
      RECT  59100.0 1013550.0 157500.0 1014450.0 ;
      RECT  59100.0 1041150.0 157500.0 1042050.0 ;
      RECT  59100.0 1068750.0 157500.0 1069650.0 ;
      RECT  59100.0 1096350.0 157500.0 1097250.0 ;
      RECT  59100.0 1123950.0 157500.0 1124850.0 ;
      RECT  59100.0 1151550.0 157500.0 1152450.0 ;
      RECT  59100.0 1179150.0 157500.0 1180050.0 ;
      RECT  59100.0 1206750.0 157500.0 1207650.0 ;
      RECT  59100.0 1234350.0 157500.0 1235250.0 ;
      RECT  59100.0 1261950.0 157500.0 1262850.0 ;
      RECT  59100.0 1289550.0 157500.0 1290450.0 ;
      RECT  59100.0 1317150.0 157500.0 1318050.0 ;
      RECT  59100.0 1344750.0 157500.0 1345650.0 ;
      RECT  59100.0 1372350.0 157500.0 1373250.0 ;
      RECT  59100.0 1399950.0 157500.0 1400850.0 ;
      RECT  59100.0 1427550.0 157500.0 1428450.0 ;
      RECT  59100.0 1455150.0 157500.0 1456050.0 ;
      RECT  59100.0 1482750.0 157500.0 1483650.0 ;
      RECT  59100.0 1510350.0 157500.0 1511250.0 ;
      RECT  59100.0 1537950.0 157500.0 1538850.0 ;
      RECT  59100.0 1565550.0 157500.0 1566450.0 ;
      RECT  59100.0 1593150.0 157500.0 1594050.0 ;
      RECT  59100.0 1620750.0 157500.0 1621650.0 ;
      RECT  59100.0 1648350.0 157500.0 1649250.0 ;
      RECT  59100.0 1675950.0 157500.0 1676850.0 ;
      RECT  59100.0 1703550.0 157500.0 1704450.0 ;
      RECT  59100.0 1731150.0 157500.0 1732050.0 ;
      RECT  59100.0 1758750.0 157500.0 1759650.0 ;
      RECT  59100.0 1786350.0 157500.0 1787250.0 ;
      RECT  59100.0 1813950.0 157500.0 1814850.0 ;
      RECT  59100.0 1841550.0 157500.0 1842450.0 ;
      RECT  59100.0 1869150.0 157500.0 1870050.0 ;
      RECT  59100.0 1896750.0 157500.0 1897650.0 ;
      RECT  59100.0 1924350.0 157500.0 1925250.0 ;
      RECT  59100.0 1951950.0 157500.0 1952850.0 ;
      RECT  59100.0 1979550.0 157500.0 1980450.0 ;
      RECT  59100.0 2007150.0 157500.0 2008050.0 ;
      RECT  59100.0 2034750.0 157500.0 2035650.0 ;
      RECT  59100.0 2062350.0 157500.0 2063250.0 ;
      RECT  59100.0 2089950.0 157500.0 2090850.0 ;
      RECT  59100.0 2117550.0 157500.0 2118450.0 ;
      RECT  59100.0 2145150.0 157500.0 2146050.0 ;
      RECT  121050.0 385350.0 126600.0 386250.0 ;
      RECT  129150.0 386550.0 130050.0 387450.0 ;
      RECT  129150.0 385350.0 130050.0 386250.0 ;
      RECT  129150.0 386250.0 130050.0 387000.0 ;
      RECT  129600.0 386550.0 136200.0 387450.0 ;
      RECT  136200.0 386550.0 137400.0 387450.0 ;
      RECT  145650.0 386550.0 146550.0 387450.0 ;
      RECT  145650.0 385350.0 146550.0 386250.0 ;
      RECT  141600.0 386550.0 146100.0 387450.0 ;
      RECT  145650.0 385800.0 146550.0 387000.0 ;
      RECT  146100.0 385350.0 150600.0 386250.0 ;
      RECT  121050.0 399750.0 126600.0 400650.0 ;
      RECT  129150.0 398550.0 130050.0 399450.0 ;
      RECT  129150.0 399750.0 130050.0 400650.0 ;
      RECT  129150.0 399000.0 130050.0 400650.0 ;
      RECT  129600.0 398550.0 136200.0 399450.0 ;
      RECT  136200.0 398550.0 137400.0 399450.0 ;
      RECT  145650.0 398550.0 146550.0 399450.0 ;
      RECT  145650.0 399750.0 146550.0 400650.0 ;
      RECT  141600.0 398550.0 146100.0 399450.0 ;
      RECT  145650.0 399000.0 146550.0 400200.0 ;
      RECT  146100.0 399750.0 150600.0 400650.0 ;
      RECT  121050.0 412950.0 126600.0 413850.0 ;
      RECT  129150.0 414150.0 130050.0 415050.0 ;
      RECT  129150.0 412950.0 130050.0 413850.0 ;
      RECT  129150.0 413850.0 130050.0 414600.0 ;
      RECT  129600.0 414150.0 136200.0 415050.0 ;
      RECT  136200.0 414150.0 137400.0 415050.0 ;
      RECT  145650.0 414150.0 146550.0 415050.0 ;
      RECT  145650.0 412950.0 146550.0 413850.0 ;
      RECT  141600.0 414150.0 146100.0 415050.0 ;
      RECT  145650.0 413400.0 146550.0 414600.0 ;
      RECT  146100.0 412950.0 150600.0 413850.0 ;
      RECT  121050.0 427350.0 126600.0 428250.0 ;
      RECT  129150.0 426150.0 130050.0 427050.0 ;
      RECT  129150.0 427350.0 130050.0 428250.0 ;
      RECT  129150.0 426600.0 130050.0 428250.0 ;
      RECT  129600.0 426150.0 136200.0 427050.0 ;
      RECT  136200.0 426150.0 137400.0 427050.0 ;
      RECT  145650.0 426150.0 146550.0 427050.0 ;
      RECT  145650.0 427350.0 146550.0 428250.0 ;
      RECT  141600.0 426150.0 146100.0 427050.0 ;
      RECT  145650.0 426600.0 146550.0 427800.0 ;
      RECT  146100.0 427350.0 150600.0 428250.0 ;
      RECT  121050.0 440550.0 126600.0 441450.0 ;
      RECT  129150.0 441750.0 130050.0 442650.0 ;
      RECT  129150.0 440550.0 130050.0 441450.0 ;
      RECT  129150.0 441450.0 130050.0 442200.0 ;
      RECT  129600.0 441750.0 136200.0 442650.0 ;
      RECT  136200.0 441750.0 137400.0 442650.0 ;
      RECT  145650.0 441750.0 146550.0 442650.0 ;
      RECT  145650.0 440550.0 146550.0 441450.0 ;
      RECT  141600.0 441750.0 146100.0 442650.0 ;
      RECT  145650.0 441000.0 146550.0 442200.0 ;
      RECT  146100.0 440550.0 150600.0 441450.0 ;
      RECT  121050.0 454950.0 126600.0 455850.0 ;
      RECT  129150.0 453750.0 130050.0 454650.0 ;
      RECT  129150.0 454950.0 130050.0 455850.0 ;
      RECT  129150.0 454200.0 130050.0 455850.0 ;
      RECT  129600.0 453750.0 136200.0 454650.0 ;
      RECT  136200.0 453750.0 137400.0 454650.0 ;
      RECT  145650.0 453750.0 146550.0 454650.0 ;
      RECT  145650.0 454950.0 146550.0 455850.0 ;
      RECT  141600.0 453750.0 146100.0 454650.0 ;
      RECT  145650.0 454200.0 146550.0 455400.0 ;
      RECT  146100.0 454950.0 150600.0 455850.0 ;
      RECT  121050.0 468150.0 126600.0 469050.0 ;
      RECT  129150.0 469350.0 130050.0 470250.0 ;
      RECT  129150.0 468150.0 130050.0 469050.0 ;
      RECT  129150.0 469050.0 130050.0 469800.0 ;
      RECT  129600.0 469350.0 136200.0 470250.0 ;
      RECT  136200.0 469350.0 137400.0 470250.0 ;
      RECT  145650.0 469350.0 146550.0 470250.0 ;
      RECT  145650.0 468150.0 146550.0 469050.0 ;
      RECT  141600.0 469350.0 146100.0 470250.0 ;
      RECT  145650.0 468600.0 146550.0 469800.0 ;
      RECT  146100.0 468150.0 150600.0 469050.0 ;
      RECT  121050.0 482550.0 126600.0 483450.0 ;
      RECT  129150.0 481350.0 130050.0 482250.0 ;
      RECT  129150.0 482550.0 130050.0 483450.0 ;
      RECT  129150.0 481800.0 130050.0 483450.0 ;
      RECT  129600.0 481350.0 136200.0 482250.0 ;
      RECT  136200.0 481350.0 137400.0 482250.0 ;
      RECT  145650.0 481350.0 146550.0 482250.0 ;
      RECT  145650.0 482550.0 146550.0 483450.0 ;
      RECT  141600.0 481350.0 146100.0 482250.0 ;
      RECT  145650.0 481800.0 146550.0 483000.0 ;
      RECT  146100.0 482550.0 150600.0 483450.0 ;
      RECT  121050.0 495750.0 126600.0 496650.0 ;
      RECT  129150.0 496950.0 130050.0 497850.0 ;
      RECT  129150.0 495750.0 130050.0 496650.0 ;
      RECT  129150.0 496650.0 130050.0 497400.0 ;
      RECT  129600.0 496950.0 136200.0 497850.0 ;
      RECT  136200.0 496950.0 137400.0 497850.0 ;
      RECT  145650.0 496950.0 146550.0 497850.0 ;
      RECT  145650.0 495750.0 146550.0 496650.0 ;
      RECT  141600.0 496950.0 146100.0 497850.0 ;
      RECT  145650.0 496200.0 146550.0 497400.0 ;
      RECT  146100.0 495750.0 150600.0 496650.0 ;
      RECT  121050.0 510150.0 126600.0 511050.0 ;
      RECT  129150.0 508950.0 130050.0 509850.0 ;
      RECT  129150.0 510150.0 130050.0 511050.0 ;
      RECT  129150.0 509400.0 130050.0 511050.0 ;
      RECT  129600.0 508950.0 136200.0 509850.0 ;
      RECT  136200.0 508950.0 137400.0 509850.0 ;
      RECT  145650.0 508950.0 146550.0 509850.0 ;
      RECT  145650.0 510150.0 146550.0 511050.0 ;
      RECT  141600.0 508950.0 146100.0 509850.0 ;
      RECT  145650.0 509400.0 146550.0 510600.0 ;
      RECT  146100.0 510150.0 150600.0 511050.0 ;
      RECT  121050.0 523350.0 126600.0 524250.0 ;
      RECT  129150.0 524550.0 130050.0 525450.0 ;
      RECT  129150.0 523350.0 130050.0 524250.0 ;
      RECT  129150.0 524250.0 130050.0 525000.0 ;
      RECT  129600.0 524550.0 136200.0 525450.0 ;
      RECT  136200.0 524550.0 137400.0 525450.0 ;
      RECT  145650.0 524550.0 146550.0 525450.0 ;
      RECT  145650.0 523350.0 146550.0 524250.0 ;
      RECT  141600.0 524550.0 146100.0 525450.0 ;
      RECT  145650.0 523800.0 146550.0 525000.0 ;
      RECT  146100.0 523350.0 150600.0 524250.0 ;
      RECT  121050.0 537750.0 126600.0 538650.0 ;
      RECT  129150.0 536550.0 130050.0 537450.0 ;
      RECT  129150.0 537750.0 130050.0 538650.0 ;
      RECT  129150.0 537000.0 130050.0 538650.0 ;
      RECT  129600.0 536550.0 136200.0 537450.0 ;
      RECT  136200.0 536550.0 137400.0 537450.0 ;
      RECT  145650.0 536550.0 146550.0 537450.0 ;
      RECT  145650.0 537750.0 146550.0 538650.0 ;
      RECT  141600.0 536550.0 146100.0 537450.0 ;
      RECT  145650.0 537000.0 146550.0 538200.0 ;
      RECT  146100.0 537750.0 150600.0 538650.0 ;
      RECT  121050.0 550950.0 126600.0 551850.0 ;
      RECT  129150.0 552150.0 130050.0 553050.0 ;
      RECT  129150.0 550950.0 130050.0 551850.0 ;
      RECT  129150.0 551850.0 130050.0 552600.0 ;
      RECT  129600.0 552150.0 136200.0 553050.0 ;
      RECT  136200.0 552150.0 137400.0 553050.0 ;
      RECT  145650.0 552150.0 146550.0 553050.0 ;
      RECT  145650.0 550950.0 146550.0 551850.0 ;
      RECT  141600.0 552150.0 146100.0 553050.0 ;
      RECT  145650.0 551400.0 146550.0 552600.0 ;
      RECT  146100.0 550950.0 150600.0 551850.0 ;
      RECT  121050.0 565350.0 126600.0 566250.0 ;
      RECT  129150.0 564150.0 130050.0 565050.0 ;
      RECT  129150.0 565350.0 130050.0 566250.0 ;
      RECT  129150.0 564600.0 130050.0 566250.0 ;
      RECT  129600.0 564150.0 136200.0 565050.0 ;
      RECT  136200.0 564150.0 137400.0 565050.0 ;
      RECT  145650.0 564150.0 146550.0 565050.0 ;
      RECT  145650.0 565350.0 146550.0 566250.0 ;
      RECT  141600.0 564150.0 146100.0 565050.0 ;
      RECT  145650.0 564600.0 146550.0 565800.0 ;
      RECT  146100.0 565350.0 150600.0 566250.0 ;
      RECT  121050.0 578550.0 126600.0 579450.0 ;
      RECT  129150.0 579750.0 130050.0 580650.0 ;
      RECT  129150.0 578550.0 130050.0 579450.0 ;
      RECT  129150.0 579450.0 130050.0 580200.0 ;
      RECT  129600.0 579750.0 136200.0 580650.0 ;
      RECT  136200.0 579750.0 137400.0 580650.0 ;
      RECT  145650.0 579750.0 146550.0 580650.0 ;
      RECT  145650.0 578550.0 146550.0 579450.0 ;
      RECT  141600.0 579750.0 146100.0 580650.0 ;
      RECT  145650.0 579000.0 146550.0 580200.0 ;
      RECT  146100.0 578550.0 150600.0 579450.0 ;
      RECT  121050.0 592950.0 126600.0 593850.0 ;
      RECT  129150.0 591750.0 130050.0 592650.0 ;
      RECT  129150.0 592950.0 130050.0 593850.0 ;
      RECT  129150.0 592200.0 130050.0 593850.0 ;
      RECT  129600.0 591750.0 136200.0 592650.0 ;
      RECT  136200.0 591750.0 137400.0 592650.0 ;
      RECT  145650.0 591750.0 146550.0 592650.0 ;
      RECT  145650.0 592950.0 146550.0 593850.0 ;
      RECT  141600.0 591750.0 146100.0 592650.0 ;
      RECT  145650.0 592200.0 146550.0 593400.0 ;
      RECT  146100.0 592950.0 150600.0 593850.0 ;
      RECT  121050.0 606150.0 126600.0 607050.0 ;
      RECT  129150.0 607350.0 130050.0 608250.0 ;
      RECT  129150.0 606150.0 130050.0 607050.0 ;
      RECT  129150.0 607050.0 130050.0 607800.0 ;
      RECT  129600.0 607350.0 136200.0 608250.0 ;
      RECT  136200.0 607350.0 137400.0 608250.0 ;
      RECT  145650.0 607350.0 146550.0 608250.0 ;
      RECT  145650.0 606150.0 146550.0 607050.0 ;
      RECT  141600.0 607350.0 146100.0 608250.0 ;
      RECT  145650.0 606600.0 146550.0 607800.0 ;
      RECT  146100.0 606150.0 150600.0 607050.0 ;
      RECT  121050.0 620550.0 126600.0 621450.0 ;
      RECT  129150.0 619350.0 130050.0 620250.0 ;
      RECT  129150.0 620550.0 130050.0 621450.0 ;
      RECT  129150.0 619800.0 130050.0 621450.0 ;
      RECT  129600.0 619350.0 136200.0 620250.0 ;
      RECT  136200.0 619350.0 137400.0 620250.0 ;
      RECT  145650.0 619350.0 146550.0 620250.0 ;
      RECT  145650.0 620550.0 146550.0 621450.0 ;
      RECT  141600.0 619350.0 146100.0 620250.0 ;
      RECT  145650.0 619800.0 146550.0 621000.0 ;
      RECT  146100.0 620550.0 150600.0 621450.0 ;
      RECT  121050.0 633750.0 126600.0 634650.0 ;
      RECT  129150.0 634950.0 130050.0 635850.0 ;
      RECT  129150.0 633750.0 130050.0 634650.0 ;
      RECT  129150.0 634650.0 130050.0 635400.0 ;
      RECT  129600.0 634950.0 136200.0 635850.0 ;
      RECT  136200.0 634950.0 137400.0 635850.0 ;
      RECT  145650.0 634950.0 146550.0 635850.0 ;
      RECT  145650.0 633750.0 146550.0 634650.0 ;
      RECT  141600.0 634950.0 146100.0 635850.0 ;
      RECT  145650.0 634200.0 146550.0 635400.0 ;
      RECT  146100.0 633750.0 150600.0 634650.0 ;
      RECT  121050.0 648150.0 126600.0 649050.0 ;
      RECT  129150.0 646950.0 130050.0 647850.0 ;
      RECT  129150.0 648150.0 130050.0 649050.0 ;
      RECT  129150.0 647400.0 130050.0 649050.0 ;
      RECT  129600.0 646950.0 136200.0 647850.0 ;
      RECT  136200.0 646950.0 137400.0 647850.0 ;
      RECT  145650.0 646950.0 146550.0 647850.0 ;
      RECT  145650.0 648150.0 146550.0 649050.0 ;
      RECT  141600.0 646950.0 146100.0 647850.0 ;
      RECT  145650.0 647400.0 146550.0 648600.0 ;
      RECT  146100.0 648150.0 150600.0 649050.0 ;
      RECT  121050.0 661350.0 126600.0 662250.0 ;
      RECT  129150.0 662550.0 130050.0 663450.0 ;
      RECT  129150.0 661350.0 130050.0 662250.0 ;
      RECT  129150.0 662250.0 130050.0 663000.0 ;
      RECT  129600.0 662550.0 136200.0 663450.0 ;
      RECT  136200.0 662550.0 137400.0 663450.0 ;
      RECT  145650.0 662550.0 146550.0 663450.0 ;
      RECT  145650.0 661350.0 146550.0 662250.0 ;
      RECT  141600.0 662550.0 146100.0 663450.0 ;
      RECT  145650.0 661800.0 146550.0 663000.0 ;
      RECT  146100.0 661350.0 150600.0 662250.0 ;
      RECT  121050.0 675750.0 126600.0 676650.0 ;
      RECT  129150.0 674550.0 130050.0 675450.0 ;
      RECT  129150.0 675750.0 130050.0 676650.0 ;
      RECT  129150.0 675000.0 130050.0 676650.0 ;
      RECT  129600.0 674550.0 136200.0 675450.0 ;
      RECT  136200.0 674550.0 137400.0 675450.0 ;
      RECT  145650.0 674550.0 146550.0 675450.0 ;
      RECT  145650.0 675750.0 146550.0 676650.0 ;
      RECT  141600.0 674550.0 146100.0 675450.0 ;
      RECT  145650.0 675000.0 146550.0 676200.0 ;
      RECT  146100.0 675750.0 150600.0 676650.0 ;
      RECT  121050.0 688950.0 126600.0 689850.0 ;
      RECT  129150.0 690150.0 130050.0 691050.0 ;
      RECT  129150.0 688950.0 130050.0 689850.0 ;
      RECT  129150.0 689850.0 130050.0 690600.0 ;
      RECT  129600.0 690150.0 136200.0 691050.0 ;
      RECT  136200.0 690150.0 137400.0 691050.0 ;
      RECT  145650.0 690150.0 146550.0 691050.0 ;
      RECT  145650.0 688950.0 146550.0 689850.0 ;
      RECT  141600.0 690150.0 146100.0 691050.0 ;
      RECT  145650.0 689400.0 146550.0 690600.0 ;
      RECT  146100.0 688950.0 150600.0 689850.0 ;
      RECT  121050.0 703350.0 126600.0 704250.0 ;
      RECT  129150.0 702150.0 130050.0 703050.0 ;
      RECT  129150.0 703350.0 130050.0 704250.0 ;
      RECT  129150.0 702600.0 130050.0 704250.0 ;
      RECT  129600.0 702150.0 136200.0 703050.0 ;
      RECT  136200.0 702150.0 137400.0 703050.0 ;
      RECT  145650.0 702150.0 146550.0 703050.0 ;
      RECT  145650.0 703350.0 146550.0 704250.0 ;
      RECT  141600.0 702150.0 146100.0 703050.0 ;
      RECT  145650.0 702600.0 146550.0 703800.0 ;
      RECT  146100.0 703350.0 150600.0 704250.0 ;
      RECT  121050.0 716550.0 126600.0 717450.0 ;
      RECT  129150.0 717750.0 130050.0 718650.0 ;
      RECT  129150.0 716550.0 130050.0 717450.0 ;
      RECT  129150.0 717450.0 130050.0 718200.0 ;
      RECT  129600.0 717750.0 136200.0 718650.0 ;
      RECT  136200.0 717750.0 137400.0 718650.0 ;
      RECT  145650.0 717750.0 146550.0 718650.0 ;
      RECT  145650.0 716550.0 146550.0 717450.0 ;
      RECT  141600.0 717750.0 146100.0 718650.0 ;
      RECT  145650.0 717000.0 146550.0 718200.0 ;
      RECT  146100.0 716550.0 150600.0 717450.0 ;
      RECT  121050.0 730950.0 126600.0 731850.0 ;
      RECT  129150.0 729750.0 130050.0 730650.0 ;
      RECT  129150.0 730950.0 130050.0 731850.0 ;
      RECT  129150.0 730200.0 130050.0 731850.0 ;
      RECT  129600.0 729750.0 136200.0 730650.0 ;
      RECT  136200.0 729750.0 137400.0 730650.0 ;
      RECT  145650.0 729750.0 146550.0 730650.0 ;
      RECT  145650.0 730950.0 146550.0 731850.0 ;
      RECT  141600.0 729750.0 146100.0 730650.0 ;
      RECT  145650.0 730200.0 146550.0 731400.0 ;
      RECT  146100.0 730950.0 150600.0 731850.0 ;
      RECT  121050.0 744150.0 126600.0 745050.0 ;
      RECT  129150.0 745350.0 130050.0 746250.0 ;
      RECT  129150.0 744150.0 130050.0 745050.0 ;
      RECT  129150.0 745050.0 130050.0 745800.0 ;
      RECT  129600.0 745350.0 136200.0 746250.0 ;
      RECT  136200.0 745350.0 137400.0 746250.0 ;
      RECT  145650.0 745350.0 146550.0 746250.0 ;
      RECT  145650.0 744150.0 146550.0 745050.0 ;
      RECT  141600.0 745350.0 146100.0 746250.0 ;
      RECT  145650.0 744600.0 146550.0 745800.0 ;
      RECT  146100.0 744150.0 150600.0 745050.0 ;
      RECT  121050.0 758550.0 126600.0 759450.0 ;
      RECT  129150.0 757350.0 130050.0 758250.0 ;
      RECT  129150.0 758550.0 130050.0 759450.0 ;
      RECT  129150.0 757800.0 130050.0 759450.0 ;
      RECT  129600.0 757350.0 136200.0 758250.0 ;
      RECT  136200.0 757350.0 137400.0 758250.0 ;
      RECT  145650.0 757350.0 146550.0 758250.0 ;
      RECT  145650.0 758550.0 146550.0 759450.0 ;
      RECT  141600.0 757350.0 146100.0 758250.0 ;
      RECT  145650.0 757800.0 146550.0 759000.0 ;
      RECT  146100.0 758550.0 150600.0 759450.0 ;
      RECT  121050.0 771750.0 126600.0 772650.0 ;
      RECT  129150.0 772950.0 130050.0 773850.0 ;
      RECT  129150.0 771750.0 130050.0 772650.0 ;
      RECT  129150.0 772650.0 130050.0 773400.0 ;
      RECT  129600.0 772950.0 136200.0 773850.0 ;
      RECT  136200.0 772950.0 137400.0 773850.0 ;
      RECT  145650.0 772950.0 146550.0 773850.0 ;
      RECT  145650.0 771750.0 146550.0 772650.0 ;
      RECT  141600.0 772950.0 146100.0 773850.0 ;
      RECT  145650.0 772200.0 146550.0 773400.0 ;
      RECT  146100.0 771750.0 150600.0 772650.0 ;
      RECT  121050.0 786150.0 126600.0 787050.0 ;
      RECT  129150.0 784950.0 130050.0 785850.0 ;
      RECT  129150.0 786150.0 130050.0 787050.0 ;
      RECT  129150.0 785400.0 130050.0 787050.0 ;
      RECT  129600.0 784950.0 136200.0 785850.0 ;
      RECT  136200.0 784950.0 137400.0 785850.0 ;
      RECT  145650.0 784950.0 146550.0 785850.0 ;
      RECT  145650.0 786150.0 146550.0 787050.0 ;
      RECT  141600.0 784950.0 146100.0 785850.0 ;
      RECT  145650.0 785400.0 146550.0 786600.0 ;
      RECT  146100.0 786150.0 150600.0 787050.0 ;
      RECT  121050.0 799350.0 126600.0 800250.0 ;
      RECT  129150.0 800550.0 130050.0 801450.0 ;
      RECT  129150.0 799350.0 130050.0 800250.0 ;
      RECT  129150.0 800250.0 130050.0 801000.0 ;
      RECT  129600.0 800550.0 136200.0 801450.0 ;
      RECT  136200.0 800550.0 137400.0 801450.0 ;
      RECT  145650.0 800550.0 146550.0 801450.0 ;
      RECT  145650.0 799350.0 146550.0 800250.0 ;
      RECT  141600.0 800550.0 146100.0 801450.0 ;
      RECT  145650.0 799800.0 146550.0 801000.0 ;
      RECT  146100.0 799350.0 150600.0 800250.0 ;
      RECT  121050.0 813750.0 126600.0 814650.0 ;
      RECT  129150.0 812550.0 130050.0 813450.0 ;
      RECT  129150.0 813750.0 130050.0 814650.0 ;
      RECT  129150.0 813000.0 130050.0 814650.0 ;
      RECT  129600.0 812550.0 136200.0 813450.0 ;
      RECT  136200.0 812550.0 137400.0 813450.0 ;
      RECT  145650.0 812550.0 146550.0 813450.0 ;
      RECT  145650.0 813750.0 146550.0 814650.0 ;
      RECT  141600.0 812550.0 146100.0 813450.0 ;
      RECT  145650.0 813000.0 146550.0 814200.0 ;
      RECT  146100.0 813750.0 150600.0 814650.0 ;
      RECT  121050.0 826950.0 126600.0 827850.0 ;
      RECT  129150.0 828150.0 130050.0 829050.0 ;
      RECT  129150.0 826950.0 130050.0 827850.0 ;
      RECT  129150.0 827850.0 130050.0 828600.0 ;
      RECT  129600.0 828150.0 136200.0 829050.0 ;
      RECT  136200.0 828150.0 137400.0 829050.0 ;
      RECT  145650.0 828150.0 146550.0 829050.0 ;
      RECT  145650.0 826950.0 146550.0 827850.0 ;
      RECT  141600.0 828150.0 146100.0 829050.0 ;
      RECT  145650.0 827400.0 146550.0 828600.0 ;
      RECT  146100.0 826950.0 150600.0 827850.0 ;
      RECT  121050.0 841350.0 126600.0 842250.0 ;
      RECT  129150.0 840150.0 130050.0 841050.0 ;
      RECT  129150.0 841350.0 130050.0 842250.0 ;
      RECT  129150.0 840600.0 130050.0 842250.0 ;
      RECT  129600.0 840150.0 136200.0 841050.0 ;
      RECT  136200.0 840150.0 137400.0 841050.0 ;
      RECT  145650.0 840150.0 146550.0 841050.0 ;
      RECT  145650.0 841350.0 146550.0 842250.0 ;
      RECT  141600.0 840150.0 146100.0 841050.0 ;
      RECT  145650.0 840600.0 146550.0 841800.0 ;
      RECT  146100.0 841350.0 150600.0 842250.0 ;
      RECT  121050.0 854550.0 126600.0 855450.0 ;
      RECT  129150.0 855750.0 130050.0 856650.0 ;
      RECT  129150.0 854550.0 130050.0 855450.0 ;
      RECT  129150.0 855450.0 130050.0 856200.0 ;
      RECT  129600.0 855750.0 136200.0 856650.0 ;
      RECT  136200.0 855750.0 137400.0 856650.0 ;
      RECT  145650.0 855750.0 146550.0 856650.0 ;
      RECT  145650.0 854550.0 146550.0 855450.0 ;
      RECT  141600.0 855750.0 146100.0 856650.0 ;
      RECT  145650.0 855000.0 146550.0 856200.0 ;
      RECT  146100.0 854550.0 150600.0 855450.0 ;
      RECT  121050.0 868950.0 126600.0 869850.0 ;
      RECT  129150.0 867750.0 130050.0 868650.0 ;
      RECT  129150.0 868950.0 130050.0 869850.0 ;
      RECT  129150.0 868200.0 130050.0 869850.0 ;
      RECT  129600.0 867750.0 136200.0 868650.0 ;
      RECT  136200.0 867750.0 137400.0 868650.0 ;
      RECT  145650.0 867750.0 146550.0 868650.0 ;
      RECT  145650.0 868950.0 146550.0 869850.0 ;
      RECT  141600.0 867750.0 146100.0 868650.0 ;
      RECT  145650.0 868200.0 146550.0 869400.0 ;
      RECT  146100.0 868950.0 150600.0 869850.0 ;
      RECT  121050.0 882150.0 126600.0 883050.0 ;
      RECT  129150.0 883350.0 130050.0 884250.0 ;
      RECT  129150.0 882150.0 130050.0 883050.0 ;
      RECT  129150.0 883050.0 130050.0 883800.0 ;
      RECT  129600.0 883350.0 136200.0 884250.0 ;
      RECT  136200.0 883350.0 137400.0 884250.0 ;
      RECT  145650.0 883350.0 146550.0 884250.0 ;
      RECT  145650.0 882150.0 146550.0 883050.0 ;
      RECT  141600.0 883350.0 146100.0 884250.0 ;
      RECT  145650.0 882600.0 146550.0 883800.0 ;
      RECT  146100.0 882150.0 150600.0 883050.0 ;
      RECT  121050.0 896550.0 126600.0 897450.0 ;
      RECT  129150.0 895350.0 130050.0 896250.0 ;
      RECT  129150.0 896550.0 130050.0 897450.0 ;
      RECT  129150.0 895800.0 130050.0 897450.0 ;
      RECT  129600.0 895350.0 136200.0 896250.0 ;
      RECT  136200.0 895350.0 137400.0 896250.0 ;
      RECT  145650.0 895350.0 146550.0 896250.0 ;
      RECT  145650.0 896550.0 146550.0 897450.0 ;
      RECT  141600.0 895350.0 146100.0 896250.0 ;
      RECT  145650.0 895800.0 146550.0 897000.0 ;
      RECT  146100.0 896550.0 150600.0 897450.0 ;
      RECT  121050.0 909750.0 126600.0 910650.0 ;
      RECT  129150.0 910950.0 130050.0 911850.0 ;
      RECT  129150.0 909750.0 130050.0 910650.0 ;
      RECT  129150.0 910650.0 130050.0 911400.0 ;
      RECT  129600.0 910950.0 136200.0 911850.0 ;
      RECT  136200.0 910950.0 137400.0 911850.0 ;
      RECT  145650.0 910950.0 146550.0 911850.0 ;
      RECT  145650.0 909750.0 146550.0 910650.0 ;
      RECT  141600.0 910950.0 146100.0 911850.0 ;
      RECT  145650.0 910200.0 146550.0 911400.0 ;
      RECT  146100.0 909750.0 150600.0 910650.0 ;
      RECT  121050.0 924150.0 126600.0 925050.0 ;
      RECT  129150.0 922950.0 130050.0 923850.0 ;
      RECT  129150.0 924150.0 130050.0 925050.0 ;
      RECT  129150.0 923400.0 130050.0 925050.0 ;
      RECT  129600.0 922950.0 136200.0 923850.0 ;
      RECT  136200.0 922950.0 137400.0 923850.0 ;
      RECT  145650.0 922950.0 146550.0 923850.0 ;
      RECT  145650.0 924150.0 146550.0 925050.0 ;
      RECT  141600.0 922950.0 146100.0 923850.0 ;
      RECT  145650.0 923400.0 146550.0 924600.0 ;
      RECT  146100.0 924150.0 150600.0 925050.0 ;
      RECT  121050.0 937350.0 126600.0 938250.0 ;
      RECT  129150.0 938550.0 130050.0 939450.0 ;
      RECT  129150.0 937350.0 130050.0 938250.0 ;
      RECT  129150.0 938250.0 130050.0 939000.0 ;
      RECT  129600.0 938550.0 136200.0 939450.0 ;
      RECT  136200.0 938550.0 137400.0 939450.0 ;
      RECT  145650.0 938550.0 146550.0 939450.0 ;
      RECT  145650.0 937350.0 146550.0 938250.0 ;
      RECT  141600.0 938550.0 146100.0 939450.0 ;
      RECT  145650.0 937800.0 146550.0 939000.0 ;
      RECT  146100.0 937350.0 150600.0 938250.0 ;
      RECT  121050.0 951750.0 126600.0 952650.0 ;
      RECT  129150.0 950550.0 130050.0 951450.0 ;
      RECT  129150.0 951750.0 130050.0 952650.0 ;
      RECT  129150.0 951000.0 130050.0 952650.0 ;
      RECT  129600.0 950550.0 136200.0 951450.0 ;
      RECT  136200.0 950550.0 137400.0 951450.0 ;
      RECT  145650.0 950550.0 146550.0 951450.0 ;
      RECT  145650.0 951750.0 146550.0 952650.0 ;
      RECT  141600.0 950550.0 146100.0 951450.0 ;
      RECT  145650.0 951000.0 146550.0 952200.0 ;
      RECT  146100.0 951750.0 150600.0 952650.0 ;
      RECT  121050.0 964950.0 126600.0 965850.0 ;
      RECT  129150.0 966150.0 130050.0 967050.0 ;
      RECT  129150.0 964950.0 130050.0 965850.0 ;
      RECT  129150.0 965850.0 130050.0 966600.0 ;
      RECT  129600.0 966150.0 136200.0 967050.0 ;
      RECT  136200.0 966150.0 137400.0 967050.0 ;
      RECT  145650.0 966150.0 146550.0 967050.0 ;
      RECT  145650.0 964950.0 146550.0 965850.0 ;
      RECT  141600.0 966150.0 146100.0 967050.0 ;
      RECT  145650.0 965400.0 146550.0 966600.0 ;
      RECT  146100.0 964950.0 150600.0 965850.0 ;
      RECT  121050.0 979350.0 126600.0 980250.0 ;
      RECT  129150.0 978150.0 130050.0 979050.0 ;
      RECT  129150.0 979350.0 130050.0 980250.0 ;
      RECT  129150.0 978600.0 130050.0 980250.0 ;
      RECT  129600.0 978150.0 136200.0 979050.0 ;
      RECT  136200.0 978150.0 137400.0 979050.0 ;
      RECT  145650.0 978150.0 146550.0 979050.0 ;
      RECT  145650.0 979350.0 146550.0 980250.0 ;
      RECT  141600.0 978150.0 146100.0 979050.0 ;
      RECT  145650.0 978600.0 146550.0 979800.0 ;
      RECT  146100.0 979350.0 150600.0 980250.0 ;
      RECT  121050.0 992550.0 126600.0 993450.0 ;
      RECT  129150.0 993750.0 130050.0 994650.0 ;
      RECT  129150.0 992550.0 130050.0 993450.0 ;
      RECT  129150.0 993450.0 130050.0 994200.0 ;
      RECT  129600.0 993750.0 136200.0 994650.0 ;
      RECT  136200.0 993750.0 137400.0 994650.0 ;
      RECT  145650.0 993750.0 146550.0 994650.0 ;
      RECT  145650.0 992550.0 146550.0 993450.0 ;
      RECT  141600.0 993750.0 146100.0 994650.0 ;
      RECT  145650.0 993000.0 146550.0 994200.0 ;
      RECT  146100.0 992550.0 150600.0 993450.0 ;
      RECT  121050.0 1006950.0 126600.0 1007850.0 ;
      RECT  129150.0 1005750.0 130050.0 1006650.0 ;
      RECT  129150.0 1006950.0 130050.0 1007850.0 ;
      RECT  129150.0 1006200.0 130050.0 1007850.0 ;
      RECT  129600.0 1005750.0 136200.0 1006650.0 ;
      RECT  136200.0 1005750.0 137400.0 1006650.0 ;
      RECT  145650.0 1005750.0 146550.0 1006650.0 ;
      RECT  145650.0 1006950.0 146550.0 1007850.0 ;
      RECT  141600.0 1005750.0 146100.0 1006650.0 ;
      RECT  145650.0 1006200.0 146550.0 1007400.0 ;
      RECT  146100.0 1006950.0 150600.0 1007850.0 ;
      RECT  121050.0 1020150.0 126600.0 1021050.0 ;
      RECT  129150.0 1021350.0 130050.0 1022250.0 ;
      RECT  129150.0 1020150.0 130050.0 1021050.0 ;
      RECT  129150.0 1021050.0 130050.0 1021800.0 ;
      RECT  129600.0 1021350.0 136200.0 1022250.0 ;
      RECT  136200.0 1021350.0 137400.0 1022250.0 ;
      RECT  145650.0 1021350.0 146550.0 1022250.0 ;
      RECT  145650.0 1020150.0 146550.0 1021050.0 ;
      RECT  141600.0 1021350.0 146100.0 1022250.0 ;
      RECT  145650.0 1020600.0 146550.0 1021800.0 ;
      RECT  146100.0 1020150.0 150600.0 1021050.0 ;
      RECT  121050.0 1034550.0 126600.0 1035450.0 ;
      RECT  129150.0 1033350.0 130050.0 1034250.0 ;
      RECT  129150.0 1034550.0 130050.0 1035450.0 ;
      RECT  129150.0 1033800.0 130050.0 1035450.0 ;
      RECT  129600.0 1033350.0 136200.0 1034250.0 ;
      RECT  136200.0 1033350.0 137400.0 1034250.0 ;
      RECT  145650.0 1033350.0 146550.0 1034250.0 ;
      RECT  145650.0 1034550.0 146550.0 1035450.0 ;
      RECT  141600.0 1033350.0 146100.0 1034250.0 ;
      RECT  145650.0 1033800.0 146550.0 1035000.0 ;
      RECT  146100.0 1034550.0 150600.0 1035450.0 ;
      RECT  121050.0 1047750.0 126600.0 1048650.0 ;
      RECT  129150.0 1048950.0 130050.0 1049850.0 ;
      RECT  129150.0 1047750.0 130050.0 1048650.0 ;
      RECT  129150.0 1048650.0 130050.0 1049400.0 ;
      RECT  129600.0 1048950.0 136200.0 1049850.0 ;
      RECT  136200.0 1048950.0 137400.0 1049850.0 ;
      RECT  145650.0 1048950.0 146550.0 1049850.0 ;
      RECT  145650.0 1047750.0 146550.0 1048650.0 ;
      RECT  141600.0 1048950.0 146100.0 1049850.0 ;
      RECT  145650.0 1048200.0 146550.0 1049400.0 ;
      RECT  146100.0 1047750.0 150600.0 1048650.0 ;
      RECT  121050.0 1062150.0 126600.0 1063050.0 ;
      RECT  129150.0 1060950.0 130050.0 1061850.0 ;
      RECT  129150.0 1062150.0 130050.0 1063050.0 ;
      RECT  129150.0 1061400.0 130050.0 1063050.0 ;
      RECT  129600.0 1060950.0 136200.0 1061850.0 ;
      RECT  136200.0 1060950.0 137400.0 1061850.0 ;
      RECT  145650.0 1060950.0 146550.0 1061850.0 ;
      RECT  145650.0 1062150.0 146550.0 1063050.0 ;
      RECT  141600.0 1060950.0 146100.0 1061850.0 ;
      RECT  145650.0 1061400.0 146550.0 1062600.0 ;
      RECT  146100.0 1062150.0 150600.0 1063050.0 ;
      RECT  121050.0 1075350.0 126600.0 1076250.0 ;
      RECT  129150.0 1076550.0 130050.0 1077450.0 ;
      RECT  129150.0 1075350.0 130050.0 1076250.0 ;
      RECT  129150.0 1076250.0 130050.0 1077000.0 ;
      RECT  129600.0 1076550.0 136200.0 1077450.0 ;
      RECT  136200.0 1076550.0 137400.0 1077450.0 ;
      RECT  145650.0 1076550.0 146550.0 1077450.0 ;
      RECT  145650.0 1075350.0 146550.0 1076250.0 ;
      RECT  141600.0 1076550.0 146100.0 1077450.0 ;
      RECT  145650.0 1075800.0 146550.0 1077000.0 ;
      RECT  146100.0 1075350.0 150600.0 1076250.0 ;
      RECT  121050.0 1089750.0 126600.0 1090650.0 ;
      RECT  129150.0 1088550.0 130050.0 1089450.0 ;
      RECT  129150.0 1089750.0 130050.0 1090650.0 ;
      RECT  129150.0 1089000.0 130050.0 1090650.0 ;
      RECT  129600.0 1088550.0 136200.0 1089450.0 ;
      RECT  136200.0 1088550.0 137400.0 1089450.0 ;
      RECT  145650.0 1088550.0 146550.0 1089450.0 ;
      RECT  145650.0 1089750.0 146550.0 1090650.0 ;
      RECT  141600.0 1088550.0 146100.0 1089450.0 ;
      RECT  145650.0 1089000.0 146550.0 1090200.0 ;
      RECT  146100.0 1089750.0 150600.0 1090650.0 ;
      RECT  121050.0 1102950.0 126600.0 1103850.0 ;
      RECT  129150.0 1104150.0 130050.0 1105050.0 ;
      RECT  129150.0 1102950.0 130050.0 1103850.0 ;
      RECT  129150.0 1103850.0 130050.0 1104600.0 ;
      RECT  129600.0 1104150.0 136200.0 1105050.0 ;
      RECT  136200.0 1104150.0 137400.0 1105050.0 ;
      RECT  145650.0 1104150.0 146550.0 1105050.0 ;
      RECT  145650.0 1102950.0 146550.0 1103850.0 ;
      RECT  141600.0 1104150.0 146100.0 1105050.0 ;
      RECT  145650.0 1103400.0 146550.0 1104600.0 ;
      RECT  146100.0 1102950.0 150600.0 1103850.0 ;
      RECT  121050.0 1117350.0 126600.0 1118250.0 ;
      RECT  129150.0 1116150.0 130050.0 1117050.0 ;
      RECT  129150.0 1117350.0 130050.0 1118250.0 ;
      RECT  129150.0 1116600.0 130050.0 1118250.0 ;
      RECT  129600.0 1116150.0 136200.0 1117050.0 ;
      RECT  136200.0 1116150.0 137400.0 1117050.0 ;
      RECT  145650.0 1116150.0 146550.0 1117050.0 ;
      RECT  145650.0 1117350.0 146550.0 1118250.0 ;
      RECT  141600.0 1116150.0 146100.0 1117050.0 ;
      RECT  145650.0 1116600.0 146550.0 1117800.0 ;
      RECT  146100.0 1117350.0 150600.0 1118250.0 ;
      RECT  121050.0 1130550.0 126600.0 1131450.0 ;
      RECT  129150.0 1131750.0 130050.0 1132650.0 ;
      RECT  129150.0 1130550.0 130050.0 1131450.0 ;
      RECT  129150.0 1131450.0 130050.0 1132200.0 ;
      RECT  129600.0 1131750.0 136200.0 1132650.0 ;
      RECT  136200.0 1131750.0 137400.0 1132650.0 ;
      RECT  145650.0 1131750.0 146550.0 1132650.0 ;
      RECT  145650.0 1130550.0 146550.0 1131450.0 ;
      RECT  141600.0 1131750.0 146100.0 1132650.0 ;
      RECT  145650.0 1131000.0 146550.0 1132200.0 ;
      RECT  146100.0 1130550.0 150600.0 1131450.0 ;
      RECT  121050.0 1144950.0 126600.0 1145850.0 ;
      RECT  129150.0 1143750.0 130050.0 1144650.0 ;
      RECT  129150.0 1144950.0 130050.0 1145850.0 ;
      RECT  129150.0 1144200.0 130050.0 1145850.0 ;
      RECT  129600.0 1143750.0 136200.0 1144650.0 ;
      RECT  136200.0 1143750.0 137400.0 1144650.0 ;
      RECT  145650.0 1143750.0 146550.0 1144650.0 ;
      RECT  145650.0 1144950.0 146550.0 1145850.0 ;
      RECT  141600.0 1143750.0 146100.0 1144650.0 ;
      RECT  145650.0 1144200.0 146550.0 1145400.0 ;
      RECT  146100.0 1144950.0 150600.0 1145850.0 ;
      RECT  121050.0 1158150.0 126600.0 1159050.0 ;
      RECT  129150.0 1159350.0 130050.0 1160250.0 ;
      RECT  129150.0 1158150.0 130050.0 1159050.0 ;
      RECT  129150.0 1159050.0 130050.0 1159800.0 ;
      RECT  129600.0 1159350.0 136200.0 1160250.0 ;
      RECT  136200.0 1159350.0 137400.0 1160250.0 ;
      RECT  145650.0 1159350.0 146550.0 1160250.0 ;
      RECT  145650.0 1158150.0 146550.0 1159050.0 ;
      RECT  141600.0 1159350.0 146100.0 1160250.0 ;
      RECT  145650.0 1158600.0 146550.0 1159800.0 ;
      RECT  146100.0 1158150.0 150600.0 1159050.0 ;
      RECT  121050.0 1172550.0 126600.0 1173450.0 ;
      RECT  129150.0 1171350.0 130050.0 1172250.0 ;
      RECT  129150.0 1172550.0 130050.0 1173450.0 ;
      RECT  129150.0 1171800.0 130050.0 1173450.0 ;
      RECT  129600.0 1171350.0 136200.0 1172250.0 ;
      RECT  136200.0 1171350.0 137400.0 1172250.0 ;
      RECT  145650.0 1171350.0 146550.0 1172250.0 ;
      RECT  145650.0 1172550.0 146550.0 1173450.0 ;
      RECT  141600.0 1171350.0 146100.0 1172250.0 ;
      RECT  145650.0 1171800.0 146550.0 1173000.0 ;
      RECT  146100.0 1172550.0 150600.0 1173450.0 ;
      RECT  121050.0 1185750.0 126600.0 1186650.0 ;
      RECT  129150.0 1186950.0 130050.0 1187850.0 ;
      RECT  129150.0 1185750.0 130050.0 1186650.0 ;
      RECT  129150.0 1186650.0 130050.0 1187400.0 ;
      RECT  129600.0 1186950.0 136200.0 1187850.0 ;
      RECT  136200.0 1186950.0 137400.0 1187850.0 ;
      RECT  145650.0 1186950.0 146550.0 1187850.0 ;
      RECT  145650.0 1185750.0 146550.0 1186650.0 ;
      RECT  141600.0 1186950.0 146100.0 1187850.0 ;
      RECT  145650.0 1186200.0 146550.0 1187400.0 ;
      RECT  146100.0 1185750.0 150600.0 1186650.0 ;
      RECT  121050.0 1200150.0 126600.0 1201050.0 ;
      RECT  129150.0 1198950.0 130050.0 1199850.0 ;
      RECT  129150.0 1200150.0 130050.0 1201050.0 ;
      RECT  129150.0 1199400.0 130050.0 1201050.0 ;
      RECT  129600.0 1198950.0 136200.0 1199850.0 ;
      RECT  136200.0 1198950.0 137400.0 1199850.0 ;
      RECT  145650.0 1198950.0 146550.0 1199850.0 ;
      RECT  145650.0 1200150.0 146550.0 1201050.0 ;
      RECT  141600.0 1198950.0 146100.0 1199850.0 ;
      RECT  145650.0 1199400.0 146550.0 1200600.0 ;
      RECT  146100.0 1200150.0 150600.0 1201050.0 ;
      RECT  121050.0 1213350.0 126600.0 1214250.0 ;
      RECT  129150.0 1214550.0 130050.0 1215450.0 ;
      RECT  129150.0 1213350.0 130050.0 1214250.0 ;
      RECT  129150.0 1214250.0 130050.0 1215000.0 ;
      RECT  129600.0 1214550.0 136200.0 1215450.0 ;
      RECT  136200.0 1214550.0 137400.0 1215450.0 ;
      RECT  145650.0 1214550.0 146550.0 1215450.0 ;
      RECT  145650.0 1213350.0 146550.0 1214250.0 ;
      RECT  141600.0 1214550.0 146100.0 1215450.0 ;
      RECT  145650.0 1213800.0 146550.0 1215000.0 ;
      RECT  146100.0 1213350.0 150600.0 1214250.0 ;
      RECT  121050.0 1227750.0 126600.0 1228650.0 ;
      RECT  129150.0 1226550.0 130050.0 1227450.0 ;
      RECT  129150.0 1227750.0 130050.0 1228650.0 ;
      RECT  129150.0 1227000.0 130050.0 1228650.0 ;
      RECT  129600.0 1226550.0 136200.0 1227450.0 ;
      RECT  136200.0 1226550.0 137400.0 1227450.0 ;
      RECT  145650.0 1226550.0 146550.0 1227450.0 ;
      RECT  145650.0 1227750.0 146550.0 1228650.0 ;
      RECT  141600.0 1226550.0 146100.0 1227450.0 ;
      RECT  145650.0 1227000.0 146550.0 1228200.0 ;
      RECT  146100.0 1227750.0 150600.0 1228650.0 ;
      RECT  121050.0 1240950.0 126600.0 1241850.0 ;
      RECT  129150.0 1242150.0 130050.0 1243050.0 ;
      RECT  129150.0 1240950.0 130050.0 1241850.0 ;
      RECT  129150.0 1241850.0 130050.0 1242600.0 ;
      RECT  129600.0 1242150.0 136200.0 1243050.0 ;
      RECT  136200.0 1242150.0 137400.0 1243050.0 ;
      RECT  145650.0 1242150.0 146550.0 1243050.0 ;
      RECT  145650.0 1240950.0 146550.0 1241850.0 ;
      RECT  141600.0 1242150.0 146100.0 1243050.0 ;
      RECT  145650.0 1241400.0 146550.0 1242600.0 ;
      RECT  146100.0 1240950.0 150600.0 1241850.0 ;
      RECT  121050.0 1255350.0 126600.0 1256250.0 ;
      RECT  129150.0 1254150.0 130050.0 1255050.0 ;
      RECT  129150.0 1255350.0 130050.0 1256250.0 ;
      RECT  129150.0 1254600.0 130050.0 1256250.0 ;
      RECT  129600.0 1254150.0 136200.0 1255050.0 ;
      RECT  136200.0 1254150.0 137400.0 1255050.0 ;
      RECT  145650.0 1254150.0 146550.0 1255050.0 ;
      RECT  145650.0 1255350.0 146550.0 1256250.0 ;
      RECT  141600.0 1254150.0 146100.0 1255050.0 ;
      RECT  145650.0 1254600.0 146550.0 1255800.0 ;
      RECT  146100.0 1255350.0 150600.0 1256250.0 ;
      RECT  121050.0 1268550.0 126600.0 1269450.0 ;
      RECT  129150.0 1269750.0 130050.0 1270650.0 ;
      RECT  129150.0 1268550.0 130050.0 1269450.0 ;
      RECT  129150.0 1269450.0 130050.0 1270200.0 ;
      RECT  129600.0 1269750.0 136200.0 1270650.0 ;
      RECT  136200.0 1269750.0 137400.0 1270650.0 ;
      RECT  145650.0 1269750.0 146550.0 1270650.0 ;
      RECT  145650.0 1268550.0 146550.0 1269450.0 ;
      RECT  141600.0 1269750.0 146100.0 1270650.0 ;
      RECT  145650.0 1269000.0 146550.0 1270200.0 ;
      RECT  146100.0 1268550.0 150600.0 1269450.0 ;
      RECT  121050.0 1282950.0 126600.0 1283850.0 ;
      RECT  129150.0 1281750.0 130050.0 1282650.0 ;
      RECT  129150.0 1282950.0 130050.0 1283850.0 ;
      RECT  129150.0 1282200.0 130050.0 1283850.0 ;
      RECT  129600.0 1281750.0 136200.0 1282650.0 ;
      RECT  136200.0 1281750.0 137400.0 1282650.0 ;
      RECT  145650.0 1281750.0 146550.0 1282650.0 ;
      RECT  145650.0 1282950.0 146550.0 1283850.0 ;
      RECT  141600.0 1281750.0 146100.0 1282650.0 ;
      RECT  145650.0 1282200.0 146550.0 1283400.0 ;
      RECT  146100.0 1282950.0 150600.0 1283850.0 ;
      RECT  121050.0 1296150.0 126600.0 1297050.0 ;
      RECT  129150.0 1297350.0 130050.0 1298250.0 ;
      RECT  129150.0 1296150.0 130050.0 1297050.0 ;
      RECT  129150.0 1297050.0 130050.0 1297800.0 ;
      RECT  129600.0 1297350.0 136200.0 1298250.0 ;
      RECT  136200.0 1297350.0 137400.0 1298250.0 ;
      RECT  145650.0 1297350.0 146550.0 1298250.0 ;
      RECT  145650.0 1296150.0 146550.0 1297050.0 ;
      RECT  141600.0 1297350.0 146100.0 1298250.0 ;
      RECT  145650.0 1296600.0 146550.0 1297800.0 ;
      RECT  146100.0 1296150.0 150600.0 1297050.0 ;
      RECT  121050.0 1310550.0 126600.0 1311450.0 ;
      RECT  129150.0 1309350.0 130050.0 1310250.0 ;
      RECT  129150.0 1310550.0 130050.0 1311450.0 ;
      RECT  129150.0 1309800.0 130050.0 1311450.0 ;
      RECT  129600.0 1309350.0 136200.0 1310250.0 ;
      RECT  136200.0 1309350.0 137400.0 1310250.0 ;
      RECT  145650.0 1309350.0 146550.0 1310250.0 ;
      RECT  145650.0 1310550.0 146550.0 1311450.0 ;
      RECT  141600.0 1309350.0 146100.0 1310250.0 ;
      RECT  145650.0 1309800.0 146550.0 1311000.0 ;
      RECT  146100.0 1310550.0 150600.0 1311450.0 ;
      RECT  121050.0 1323750.0 126600.0 1324650.0 ;
      RECT  129150.0 1324950.0 130050.0 1325850.0 ;
      RECT  129150.0 1323750.0 130050.0 1324650.0 ;
      RECT  129150.0 1324650.0 130050.0 1325400.0 ;
      RECT  129600.0 1324950.0 136200.0 1325850.0 ;
      RECT  136200.0 1324950.0 137400.0 1325850.0 ;
      RECT  145650.0 1324950.0 146550.0 1325850.0 ;
      RECT  145650.0 1323750.0 146550.0 1324650.0 ;
      RECT  141600.0 1324950.0 146100.0 1325850.0 ;
      RECT  145650.0 1324200.0 146550.0 1325400.0 ;
      RECT  146100.0 1323750.0 150600.0 1324650.0 ;
      RECT  121050.0 1338150.0 126600.0 1339050.0 ;
      RECT  129150.0 1336950.0 130050.0 1337850.0 ;
      RECT  129150.0 1338150.0 130050.0 1339050.0 ;
      RECT  129150.0 1337400.0 130050.0 1339050.0 ;
      RECT  129600.0 1336950.0 136200.0 1337850.0 ;
      RECT  136200.0 1336950.0 137400.0 1337850.0 ;
      RECT  145650.0 1336950.0 146550.0 1337850.0 ;
      RECT  145650.0 1338150.0 146550.0 1339050.0 ;
      RECT  141600.0 1336950.0 146100.0 1337850.0 ;
      RECT  145650.0 1337400.0 146550.0 1338600.0 ;
      RECT  146100.0 1338150.0 150600.0 1339050.0 ;
      RECT  121050.0 1351350.0 126600.0 1352250.0 ;
      RECT  129150.0 1352550.0 130050.0 1353450.0 ;
      RECT  129150.0 1351350.0 130050.0 1352250.0 ;
      RECT  129150.0 1352250.0 130050.0 1353000.0 ;
      RECT  129600.0 1352550.0 136200.0 1353450.0 ;
      RECT  136200.0 1352550.0 137400.0 1353450.0 ;
      RECT  145650.0 1352550.0 146550.0 1353450.0 ;
      RECT  145650.0 1351350.0 146550.0 1352250.0 ;
      RECT  141600.0 1352550.0 146100.0 1353450.0 ;
      RECT  145650.0 1351800.0 146550.0 1353000.0 ;
      RECT  146100.0 1351350.0 150600.0 1352250.0 ;
      RECT  121050.0 1365750.0 126600.0 1366650.0 ;
      RECT  129150.0 1364550.0 130050.0 1365450.0 ;
      RECT  129150.0 1365750.0 130050.0 1366650.0 ;
      RECT  129150.0 1365000.0 130050.0 1366650.0 ;
      RECT  129600.0 1364550.0 136200.0 1365450.0 ;
      RECT  136200.0 1364550.0 137400.0 1365450.0 ;
      RECT  145650.0 1364550.0 146550.0 1365450.0 ;
      RECT  145650.0 1365750.0 146550.0 1366650.0 ;
      RECT  141600.0 1364550.0 146100.0 1365450.0 ;
      RECT  145650.0 1365000.0 146550.0 1366200.0 ;
      RECT  146100.0 1365750.0 150600.0 1366650.0 ;
      RECT  121050.0 1378950.0 126600.0 1379850.0 ;
      RECT  129150.0 1380150.0 130050.0 1381050.0 ;
      RECT  129150.0 1378950.0 130050.0 1379850.0 ;
      RECT  129150.0 1379850.0 130050.0 1380600.0 ;
      RECT  129600.0 1380150.0 136200.0 1381050.0 ;
      RECT  136200.0 1380150.0 137400.0 1381050.0 ;
      RECT  145650.0 1380150.0 146550.0 1381050.0 ;
      RECT  145650.0 1378950.0 146550.0 1379850.0 ;
      RECT  141600.0 1380150.0 146100.0 1381050.0 ;
      RECT  145650.0 1379400.0 146550.0 1380600.0 ;
      RECT  146100.0 1378950.0 150600.0 1379850.0 ;
      RECT  121050.0 1393350.0 126600.0 1394250.0 ;
      RECT  129150.0 1392150.0 130050.0 1393050.0 ;
      RECT  129150.0 1393350.0 130050.0 1394250.0 ;
      RECT  129150.0 1392600.0 130050.0 1394250.0 ;
      RECT  129600.0 1392150.0 136200.0 1393050.0 ;
      RECT  136200.0 1392150.0 137400.0 1393050.0 ;
      RECT  145650.0 1392150.0 146550.0 1393050.0 ;
      RECT  145650.0 1393350.0 146550.0 1394250.0 ;
      RECT  141600.0 1392150.0 146100.0 1393050.0 ;
      RECT  145650.0 1392600.0 146550.0 1393800.0 ;
      RECT  146100.0 1393350.0 150600.0 1394250.0 ;
      RECT  121050.0 1406550.0 126600.0 1407450.0 ;
      RECT  129150.0 1407750.0 130050.0 1408650.0 ;
      RECT  129150.0 1406550.0 130050.0 1407450.0 ;
      RECT  129150.0 1407450.0 130050.0 1408200.0 ;
      RECT  129600.0 1407750.0 136200.0 1408650.0 ;
      RECT  136200.0 1407750.0 137400.0 1408650.0 ;
      RECT  145650.0 1407750.0 146550.0 1408650.0 ;
      RECT  145650.0 1406550.0 146550.0 1407450.0 ;
      RECT  141600.0 1407750.0 146100.0 1408650.0 ;
      RECT  145650.0 1407000.0 146550.0 1408200.0 ;
      RECT  146100.0 1406550.0 150600.0 1407450.0 ;
      RECT  121050.0 1420950.0 126600.0 1421850.0 ;
      RECT  129150.0 1419750.0 130050.0 1420650.0 ;
      RECT  129150.0 1420950.0 130050.0 1421850.0 ;
      RECT  129150.0 1420200.0 130050.0 1421850.0 ;
      RECT  129600.0 1419750.0 136200.0 1420650.0 ;
      RECT  136200.0 1419750.0 137400.0 1420650.0 ;
      RECT  145650.0 1419750.0 146550.0 1420650.0 ;
      RECT  145650.0 1420950.0 146550.0 1421850.0 ;
      RECT  141600.0 1419750.0 146100.0 1420650.0 ;
      RECT  145650.0 1420200.0 146550.0 1421400.0 ;
      RECT  146100.0 1420950.0 150600.0 1421850.0 ;
      RECT  121050.0 1434150.0 126600.0 1435050.0 ;
      RECT  129150.0 1435350.0 130050.0 1436250.0 ;
      RECT  129150.0 1434150.0 130050.0 1435050.0 ;
      RECT  129150.0 1435050.0 130050.0 1435800.0 ;
      RECT  129600.0 1435350.0 136200.0 1436250.0 ;
      RECT  136200.0 1435350.0 137400.0 1436250.0 ;
      RECT  145650.0 1435350.0 146550.0 1436250.0 ;
      RECT  145650.0 1434150.0 146550.0 1435050.0 ;
      RECT  141600.0 1435350.0 146100.0 1436250.0 ;
      RECT  145650.0 1434600.0 146550.0 1435800.0 ;
      RECT  146100.0 1434150.0 150600.0 1435050.0 ;
      RECT  121050.0 1448550.0 126600.0 1449450.0 ;
      RECT  129150.0 1447350.0 130050.0 1448250.0 ;
      RECT  129150.0 1448550.0 130050.0 1449450.0 ;
      RECT  129150.0 1447800.0 130050.0 1449450.0 ;
      RECT  129600.0 1447350.0 136200.0 1448250.0 ;
      RECT  136200.0 1447350.0 137400.0 1448250.0 ;
      RECT  145650.0 1447350.0 146550.0 1448250.0 ;
      RECT  145650.0 1448550.0 146550.0 1449450.0 ;
      RECT  141600.0 1447350.0 146100.0 1448250.0 ;
      RECT  145650.0 1447800.0 146550.0 1449000.0 ;
      RECT  146100.0 1448550.0 150600.0 1449450.0 ;
      RECT  121050.0 1461750.0 126600.0 1462650.0 ;
      RECT  129150.0 1462950.0 130050.0 1463850.0 ;
      RECT  129150.0 1461750.0 130050.0 1462650.0 ;
      RECT  129150.0 1462650.0 130050.0 1463400.0 ;
      RECT  129600.0 1462950.0 136200.0 1463850.0 ;
      RECT  136200.0 1462950.0 137400.0 1463850.0 ;
      RECT  145650.0 1462950.0 146550.0 1463850.0 ;
      RECT  145650.0 1461750.0 146550.0 1462650.0 ;
      RECT  141600.0 1462950.0 146100.0 1463850.0 ;
      RECT  145650.0 1462200.0 146550.0 1463400.0 ;
      RECT  146100.0 1461750.0 150600.0 1462650.0 ;
      RECT  121050.0 1476150.0 126600.0 1477050.0 ;
      RECT  129150.0 1474950.0 130050.0 1475850.0 ;
      RECT  129150.0 1476150.0 130050.0 1477050.0 ;
      RECT  129150.0 1475400.0 130050.0 1477050.0 ;
      RECT  129600.0 1474950.0 136200.0 1475850.0 ;
      RECT  136200.0 1474950.0 137400.0 1475850.0 ;
      RECT  145650.0 1474950.0 146550.0 1475850.0 ;
      RECT  145650.0 1476150.0 146550.0 1477050.0 ;
      RECT  141600.0 1474950.0 146100.0 1475850.0 ;
      RECT  145650.0 1475400.0 146550.0 1476600.0 ;
      RECT  146100.0 1476150.0 150600.0 1477050.0 ;
      RECT  121050.0 1489350.0 126600.0 1490250.0 ;
      RECT  129150.0 1490550.0 130050.0 1491450.0 ;
      RECT  129150.0 1489350.0 130050.0 1490250.0 ;
      RECT  129150.0 1490250.0 130050.0 1491000.0 ;
      RECT  129600.0 1490550.0 136200.0 1491450.0 ;
      RECT  136200.0 1490550.0 137400.0 1491450.0 ;
      RECT  145650.0 1490550.0 146550.0 1491450.0 ;
      RECT  145650.0 1489350.0 146550.0 1490250.0 ;
      RECT  141600.0 1490550.0 146100.0 1491450.0 ;
      RECT  145650.0 1489800.0 146550.0 1491000.0 ;
      RECT  146100.0 1489350.0 150600.0 1490250.0 ;
      RECT  121050.0 1503750.0 126600.0 1504650.0 ;
      RECT  129150.0 1502550.0 130050.0 1503450.0 ;
      RECT  129150.0 1503750.0 130050.0 1504650.0 ;
      RECT  129150.0 1503000.0 130050.0 1504650.0 ;
      RECT  129600.0 1502550.0 136200.0 1503450.0 ;
      RECT  136200.0 1502550.0 137400.0 1503450.0 ;
      RECT  145650.0 1502550.0 146550.0 1503450.0 ;
      RECT  145650.0 1503750.0 146550.0 1504650.0 ;
      RECT  141600.0 1502550.0 146100.0 1503450.0 ;
      RECT  145650.0 1503000.0 146550.0 1504200.0 ;
      RECT  146100.0 1503750.0 150600.0 1504650.0 ;
      RECT  121050.0 1516950.0 126600.0 1517850.0 ;
      RECT  129150.0 1518150.0 130050.0 1519050.0 ;
      RECT  129150.0 1516950.0 130050.0 1517850.0 ;
      RECT  129150.0 1517850.0 130050.0 1518600.0 ;
      RECT  129600.0 1518150.0 136200.0 1519050.0 ;
      RECT  136200.0 1518150.0 137400.0 1519050.0 ;
      RECT  145650.0 1518150.0 146550.0 1519050.0 ;
      RECT  145650.0 1516950.0 146550.0 1517850.0 ;
      RECT  141600.0 1518150.0 146100.0 1519050.0 ;
      RECT  145650.0 1517400.0 146550.0 1518600.0 ;
      RECT  146100.0 1516950.0 150600.0 1517850.0 ;
      RECT  121050.0 1531350.0 126600.0 1532250.0 ;
      RECT  129150.0 1530150.0 130050.0 1531050.0 ;
      RECT  129150.0 1531350.0 130050.0 1532250.0 ;
      RECT  129150.0 1530600.0 130050.0 1532250.0 ;
      RECT  129600.0 1530150.0 136200.0 1531050.0 ;
      RECT  136200.0 1530150.0 137400.0 1531050.0 ;
      RECT  145650.0 1530150.0 146550.0 1531050.0 ;
      RECT  145650.0 1531350.0 146550.0 1532250.0 ;
      RECT  141600.0 1530150.0 146100.0 1531050.0 ;
      RECT  145650.0 1530600.0 146550.0 1531800.0 ;
      RECT  146100.0 1531350.0 150600.0 1532250.0 ;
      RECT  121050.0 1544550.0 126600.0 1545450.0 ;
      RECT  129150.0 1545750.0 130050.0 1546650.0 ;
      RECT  129150.0 1544550.0 130050.0 1545450.0 ;
      RECT  129150.0 1545450.0 130050.0 1546200.0 ;
      RECT  129600.0 1545750.0 136200.0 1546650.0 ;
      RECT  136200.0 1545750.0 137400.0 1546650.0 ;
      RECT  145650.0 1545750.0 146550.0 1546650.0 ;
      RECT  145650.0 1544550.0 146550.0 1545450.0 ;
      RECT  141600.0 1545750.0 146100.0 1546650.0 ;
      RECT  145650.0 1545000.0 146550.0 1546200.0 ;
      RECT  146100.0 1544550.0 150600.0 1545450.0 ;
      RECT  121050.0 1558950.0 126600.0 1559850.0 ;
      RECT  129150.0 1557750.0 130050.0 1558650.0 ;
      RECT  129150.0 1558950.0 130050.0 1559850.0 ;
      RECT  129150.0 1558200.0 130050.0 1559850.0 ;
      RECT  129600.0 1557750.0 136200.0 1558650.0 ;
      RECT  136200.0 1557750.0 137400.0 1558650.0 ;
      RECT  145650.0 1557750.0 146550.0 1558650.0 ;
      RECT  145650.0 1558950.0 146550.0 1559850.0 ;
      RECT  141600.0 1557750.0 146100.0 1558650.0 ;
      RECT  145650.0 1558200.0 146550.0 1559400.0 ;
      RECT  146100.0 1558950.0 150600.0 1559850.0 ;
      RECT  121050.0 1572150.0 126600.0 1573050.0 ;
      RECT  129150.0 1573350.0 130050.0 1574250.0 ;
      RECT  129150.0 1572150.0 130050.0 1573050.0 ;
      RECT  129150.0 1573050.0 130050.0 1573800.0 ;
      RECT  129600.0 1573350.0 136200.0 1574250.0 ;
      RECT  136200.0 1573350.0 137400.0 1574250.0 ;
      RECT  145650.0 1573350.0 146550.0 1574250.0 ;
      RECT  145650.0 1572150.0 146550.0 1573050.0 ;
      RECT  141600.0 1573350.0 146100.0 1574250.0 ;
      RECT  145650.0 1572600.0 146550.0 1573800.0 ;
      RECT  146100.0 1572150.0 150600.0 1573050.0 ;
      RECT  121050.0 1586550.0 126600.0 1587450.0 ;
      RECT  129150.0 1585350.0 130050.0 1586250.0 ;
      RECT  129150.0 1586550.0 130050.0 1587450.0 ;
      RECT  129150.0 1585800.0 130050.0 1587450.0 ;
      RECT  129600.0 1585350.0 136200.0 1586250.0 ;
      RECT  136200.0 1585350.0 137400.0 1586250.0 ;
      RECT  145650.0 1585350.0 146550.0 1586250.0 ;
      RECT  145650.0 1586550.0 146550.0 1587450.0 ;
      RECT  141600.0 1585350.0 146100.0 1586250.0 ;
      RECT  145650.0 1585800.0 146550.0 1587000.0 ;
      RECT  146100.0 1586550.0 150600.0 1587450.0 ;
      RECT  121050.0 1599750.0 126600.0 1600650.0 ;
      RECT  129150.0 1600950.0 130050.0 1601850.0 ;
      RECT  129150.0 1599750.0 130050.0 1600650.0 ;
      RECT  129150.0 1600650.0 130050.0 1601400.0 ;
      RECT  129600.0 1600950.0 136200.0 1601850.0 ;
      RECT  136200.0 1600950.0 137400.0 1601850.0 ;
      RECT  145650.0 1600950.0 146550.0 1601850.0 ;
      RECT  145650.0 1599750.0 146550.0 1600650.0 ;
      RECT  141600.0 1600950.0 146100.0 1601850.0 ;
      RECT  145650.0 1600200.0 146550.0 1601400.0 ;
      RECT  146100.0 1599750.0 150600.0 1600650.0 ;
      RECT  121050.0 1614150.0 126600.0 1615050.0 ;
      RECT  129150.0 1612950.0 130050.0 1613850.0 ;
      RECT  129150.0 1614150.0 130050.0 1615050.0 ;
      RECT  129150.0 1613400.0 130050.0 1615050.0 ;
      RECT  129600.0 1612950.0 136200.0 1613850.0 ;
      RECT  136200.0 1612950.0 137400.0 1613850.0 ;
      RECT  145650.0 1612950.0 146550.0 1613850.0 ;
      RECT  145650.0 1614150.0 146550.0 1615050.0 ;
      RECT  141600.0 1612950.0 146100.0 1613850.0 ;
      RECT  145650.0 1613400.0 146550.0 1614600.0 ;
      RECT  146100.0 1614150.0 150600.0 1615050.0 ;
      RECT  121050.0 1627350.0 126600.0 1628250.0 ;
      RECT  129150.0 1628550.0 130050.0 1629450.0 ;
      RECT  129150.0 1627350.0 130050.0 1628250.0 ;
      RECT  129150.0 1628250.0 130050.0 1629000.0 ;
      RECT  129600.0 1628550.0 136200.0 1629450.0 ;
      RECT  136200.0 1628550.0 137400.0 1629450.0 ;
      RECT  145650.0 1628550.0 146550.0 1629450.0 ;
      RECT  145650.0 1627350.0 146550.0 1628250.0 ;
      RECT  141600.0 1628550.0 146100.0 1629450.0 ;
      RECT  145650.0 1627800.0 146550.0 1629000.0 ;
      RECT  146100.0 1627350.0 150600.0 1628250.0 ;
      RECT  121050.0 1641750.0 126600.0 1642650.0 ;
      RECT  129150.0 1640550.0 130050.0 1641450.0 ;
      RECT  129150.0 1641750.0 130050.0 1642650.0 ;
      RECT  129150.0 1641000.0 130050.0 1642650.0 ;
      RECT  129600.0 1640550.0 136200.0 1641450.0 ;
      RECT  136200.0 1640550.0 137400.0 1641450.0 ;
      RECT  145650.0 1640550.0 146550.0 1641450.0 ;
      RECT  145650.0 1641750.0 146550.0 1642650.0 ;
      RECT  141600.0 1640550.0 146100.0 1641450.0 ;
      RECT  145650.0 1641000.0 146550.0 1642200.0 ;
      RECT  146100.0 1641750.0 150600.0 1642650.0 ;
      RECT  121050.0 1654950.0 126600.0 1655850.0 ;
      RECT  129150.0 1656150.0 130050.0 1657050.0 ;
      RECT  129150.0 1654950.0 130050.0 1655850.0 ;
      RECT  129150.0 1655850.0 130050.0 1656600.0 ;
      RECT  129600.0 1656150.0 136200.0 1657050.0 ;
      RECT  136200.0 1656150.0 137400.0 1657050.0 ;
      RECT  145650.0 1656150.0 146550.0 1657050.0 ;
      RECT  145650.0 1654950.0 146550.0 1655850.0 ;
      RECT  141600.0 1656150.0 146100.0 1657050.0 ;
      RECT  145650.0 1655400.0 146550.0 1656600.0 ;
      RECT  146100.0 1654950.0 150600.0 1655850.0 ;
      RECT  121050.0 1669350.0 126600.0 1670250.0 ;
      RECT  129150.0 1668150.0 130050.0 1669050.0 ;
      RECT  129150.0 1669350.0 130050.0 1670250.0 ;
      RECT  129150.0 1668600.0 130050.0 1670250.0 ;
      RECT  129600.0 1668150.0 136200.0 1669050.0 ;
      RECT  136200.0 1668150.0 137400.0 1669050.0 ;
      RECT  145650.0 1668150.0 146550.0 1669050.0 ;
      RECT  145650.0 1669350.0 146550.0 1670250.0 ;
      RECT  141600.0 1668150.0 146100.0 1669050.0 ;
      RECT  145650.0 1668600.0 146550.0 1669800.0 ;
      RECT  146100.0 1669350.0 150600.0 1670250.0 ;
      RECT  121050.0 1682550.0 126600.0 1683450.0 ;
      RECT  129150.0 1683750.0 130050.0 1684650.0 ;
      RECT  129150.0 1682550.0 130050.0 1683450.0 ;
      RECT  129150.0 1683450.0 130050.0 1684200.0 ;
      RECT  129600.0 1683750.0 136200.0 1684650.0 ;
      RECT  136200.0 1683750.0 137400.0 1684650.0 ;
      RECT  145650.0 1683750.0 146550.0 1684650.0 ;
      RECT  145650.0 1682550.0 146550.0 1683450.0 ;
      RECT  141600.0 1683750.0 146100.0 1684650.0 ;
      RECT  145650.0 1683000.0 146550.0 1684200.0 ;
      RECT  146100.0 1682550.0 150600.0 1683450.0 ;
      RECT  121050.0 1696950.0 126600.0 1697850.0 ;
      RECT  129150.0 1695750.0 130050.0 1696650.0 ;
      RECT  129150.0 1696950.0 130050.0 1697850.0 ;
      RECT  129150.0 1696200.0 130050.0 1697850.0 ;
      RECT  129600.0 1695750.0 136200.0 1696650.0 ;
      RECT  136200.0 1695750.0 137400.0 1696650.0 ;
      RECT  145650.0 1695750.0 146550.0 1696650.0 ;
      RECT  145650.0 1696950.0 146550.0 1697850.0 ;
      RECT  141600.0 1695750.0 146100.0 1696650.0 ;
      RECT  145650.0 1696200.0 146550.0 1697400.0 ;
      RECT  146100.0 1696950.0 150600.0 1697850.0 ;
      RECT  121050.0 1710150.0 126600.0 1711050.0 ;
      RECT  129150.0 1711350.0 130050.0 1712250.0 ;
      RECT  129150.0 1710150.0 130050.0 1711050.0 ;
      RECT  129150.0 1711050.0 130050.0 1711800.0 ;
      RECT  129600.0 1711350.0 136200.0 1712250.0 ;
      RECT  136200.0 1711350.0 137400.0 1712250.0 ;
      RECT  145650.0 1711350.0 146550.0 1712250.0 ;
      RECT  145650.0 1710150.0 146550.0 1711050.0 ;
      RECT  141600.0 1711350.0 146100.0 1712250.0 ;
      RECT  145650.0 1710600.0 146550.0 1711800.0 ;
      RECT  146100.0 1710150.0 150600.0 1711050.0 ;
      RECT  121050.0 1724550.0 126600.0 1725450.0 ;
      RECT  129150.0 1723350.0 130050.0 1724250.0 ;
      RECT  129150.0 1724550.0 130050.0 1725450.0 ;
      RECT  129150.0 1723800.0 130050.0 1725450.0 ;
      RECT  129600.0 1723350.0 136200.0 1724250.0 ;
      RECT  136200.0 1723350.0 137400.0 1724250.0 ;
      RECT  145650.0 1723350.0 146550.0 1724250.0 ;
      RECT  145650.0 1724550.0 146550.0 1725450.0 ;
      RECT  141600.0 1723350.0 146100.0 1724250.0 ;
      RECT  145650.0 1723800.0 146550.0 1725000.0 ;
      RECT  146100.0 1724550.0 150600.0 1725450.0 ;
      RECT  121050.0 1737750.0 126600.0 1738650.0 ;
      RECT  129150.0 1738950.0 130050.0 1739850.0 ;
      RECT  129150.0 1737750.0 130050.0 1738650.0 ;
      RECT  129150.0 1738650.0 130050.0 1739400.0 ;
      RECT  129600.0 1738950.0 136200.0 1739850.0 ;
      RECT  136200.0 1738950.0 137400.0 1739850.0 ;
      RECT  145650.0 1738950.0 146550.0 1739850.0 ;
      RECT  145650.0 1737750.0 146550.0 1738650.0 ;
      RECT  141600.0 1738950.0 146100.0 1739850.0 ;
      RECT  145650.0 1738200.0 146550.0 1739400.0 ;
      RECT  146100.0 1737750.0 150600.0 1738650.0 ;
      RECT  121050.0 1752150.0 126600.0 1753050.0 ;
      RECT  129150.0 1750950.0 130050.0 1751850.0 ;
      RECT  129150.0 1752150.0 130050.0 1753050.0 ;
      RECT  129150.0 1751400.0 130050.0 1753050.0 ;
      RECT  129600.0 1750950.0 136200.0 1751850.0 ;
      RECT  136200.0 1750950.0 137400.0 1751850.0 ;
      RECT  145650.0 1750950.0 146550.0 1751850.0 ;
      RECT  145650.0 1752150.0 146550.0 1753050.0 ;
      RECT  141600.0 1750950.0 146100.0 1751850.0 ;
      RECT  145650.0 1751400.0 146550.0 1752600.0 ;
      RECT  146100.0 1752150.0 150600.0 1753050.0 ;
      RECT  121050.0 1765350.0 126600.0 1766250.0 ;
      RECT  129150.0 1766550.0 130050.0 1767450.0 ;
      RECT  129150.0 1765350.0 130050.0 1766250.0 ;
      RECT  129150.0 1766250.0 130050.0 1767000.0 ;
      RECT  129600.0 1766550.0 136200.0 1767450.0 ;
      RECT  136200.0 1766550.0 137400.0 1767450.0 ;
      RECT  145650.0 1766550.0 146550.0 1767450.0 ;
      RECT  145650.0 1765350.0 146550.0 1766250.0 ;
      RECT  141600.0 1766550.0 146100.0 1767450.0 ;
      RECT  145650.0 1765800.0 146550.0 1767000.0 ;
      RECT  146100.0 1765350.0 150600.0 1766250.0 ;
      RECT  121050.0 1779750.0 126600.0 1780650.0 ;
      RECT  129150.0 1778550.0 130050.0 1779450.0 ;
      RECT  129150.0 1779750.0 130050.0 1780650.0 ;
      RECT  129150.0 1779000.0 130050.0 1780650.0 ;
      RECT  129600.0 1778550.0 136200.0 1779450.0 ;
      RECT  136200.0 1778550.0 137400.0 1779450.0 ;
      RECT  145650.0 1778550.0 146550.0 1779450.0 ;
      RECT  145650.0 1779750.0 146550.0 1780650.0 ;
      RECT  141600.0 1778550.0 146100.0 1779450.0 ;
      RECT  145650.0 1779000.0 146550.0 1780200.0 ;
      RECT  146100.0 1779750.0 150600.0 1780650.0 ;
      RECT  121050.0 1792950.0 126600.0 1793850.0 ;
      RECT  129150.0 1794150.0 130050.0 1795050.0 ;
      RECT  129150.0 1792950.0 130050.0 1793850.0 ;
      RECT  129150.0 1793850.0 130050.0 1794600.0 ;
      RECT  129600.0 1794150.0 136200.0 1795050.0 ;
      RECT  136200.0 1794150.0 137400.0 1795050.0 ;
      RECT  145650.0 1794150.0 146550.0 1795050.0 ;
      RECT  145650.0 1792950.0 146550.0 1793850.0 ;
      RECT  141600.0 1794150.0 146100.0 1795050.0 ;
      RECT  145650.0 1793400.0 146550.0 1794600.0 ;
      RECT  146100.0 1792950.0 150600.0 1793850.0 ;
      RECT  121050.0 1807350.0 126600.0 1808250.0 ;
      RECT  129150.0 1806150.0 130050.0 1807050.0 ;
      RECT  129150.0 1807350.0 130050.0 1808250.0 ;
      RECT  129150.0 1806600.0 130050.0 1808250.0 ;
      RECT  129600.0 1806150.0 136200.0 1807050.0 ;
      RECT  136200.0 1806150.0 137400.0 1807050.0 ;
      RECT  145650.0 1806150.0 146550.0 1807050.0 ;
      RECT  145650.0 1807350.0 146550.0 1808250.0 ;
      RECT  141600.0 1806150.0 146100.0 1807050.0 ;
      RECT  145650.0 1806600.0 146550.0 1807800.0 ;
      RECT  146100.0 1807350.0 150600.0 1808250.0 ;
      RECT  121050.0 1820550.0 126600.0 1821450.0 ;
      RECT  129150.0 1821750.0 130050.0 1822650.0 ;
      RECT  129150.0 1820550.0 130050.0 1821450.0 ;
      RECT  129150.0 1821450.0 130050.0 1822200.0 ;
      RECT  129600.0 1821750.0 136200.0 1822650.0 ;
      RECT  136200.0 1821750.0 137400.0 1822650.0 ;
      RECT  145650.0 1821750.0 146550.0 1822650.0 ;
      RECT  145650.0 1820550.0 146550.0 1821450.0 ;
      RECT  141600.0 1821750.0 146100.0 1822650.0 ;
      RECT  145650.0 1821000.0 146550.0 1822200.0 ;
      RECT  146100.0 1820550.0 150600.0 1821450.0 ;
      RECT  121050.0 1834950.0 126600.0 1835850.0 ;
      RECT  129150.0 1833750.0 130050.0 1834650.0 ;
      RECT  129150.0 1834950.0 130050.0 1835850.0 ;
      RECT  129150.0 1834200.0 130050.0 1835850.0 ;
      RECT  129600.0 1833750.0 136200.0 1834650.0 ;
      RECT  136200.0 1833750.0 137400.0 1834650.0 ;
      RECT  145650.0 1833750.0 146550.0 1834650.0 ;
      RECT  145650.0 1834950.0 146550.0 1835850.0 ;
      RECT  141600.0 1833750.0 146100.0 1834650.0 ;
      RECT  145650.0 1834200.0 146550.0 1835400.0 ;
      RECT  146100.0 1834950.0 150600.0 1835850.0 ;
      RECT  121050.0 1848150.0 126600.0 1849050.0 ;
      RECT  129150.0 1849350.0 130050.0 1850250.0 ;
      RECT  129150.0 1848150.0 130050.0 1849050.0 ;
      RECT  129150.0 1849050.0 130050.0 1849800.0 ;
      RECT  129600.0 1849350.0 136200.0 1850250.0 ;
      RECT  136200.0 1849350.0 137400.0 1850250.0 ;
      RECT  145650.0 1849350.0 146550.0 1850250.0 ;
      RECT  145650.0 1848150.0 146550.0 1849050.0 ;
      RECT  141600.0 1849350.0 146100.0 1850250.0 ;
      RECT  145650.0 1848600.0 146550.0 1849800.0 ;
      RECT  146100.0 1848150.0 150600.0 1849050.0 ;
      RECT  121050.0 1862550.0 126600.0 1863450.0 ;
      RECT  129150.0 1861350.0 130050.0 1862250.0 ;
      RECT  129150.0 1862550.0 130050.0 1863450.0 ;
      RECT  129150.0 1861800.0 130050.0 1863450.0 ;
      RECT  129600.0 1861350.0 136200.0 1862250.0 ;
      RECT  136200.0 1861350.0 137400.0 1862250.0 ;
      RECT  145650.0 1861350.0 146550.0 1862250.0 ;
      RECT  145650.0 1862550.0 146550.0 1863450.0 ;
      RECT  141600.0 1861350.0 146100.0 1862250.0 ;
      RECT  145650.0 1861800.0 146550.0 1863000.0 ;
      RECT  146100.0 1862550.0 150600.0 1863450.0 ;
      RECT  121050.0 1875750.0 126600.0 1876650.0 ;
      RECT  129150.0 1876950.0 130050.0 1877850.0 ;
      RECT  129150.0 1875750.0 130050.0 1876650.0 ;
      RECT  129150.0 1876650.0 130050.0 1877400.0 ;
      RECT  129600.0 1876950.0 136200.0 1877850.0 ;
      RECT  136200.0 1876950.0 137400.0 1877850.0 ;
      RECT  145650.0 1876950.0 146550.0 1877850.0 ;
      RECT  145650.0 1875750.0 146550.0 1876650.0 ;
      RECT  141600.0 1876950.0 146100.0 1877850.0 ;
      RECT  145650.0 1876200.0 146550.0 1877400.0 ;
      RECT  146100.0 1875750.0 150600.0 1876650.0 ;
      RECT  121050.0 1890150.0 126600.0 1891050.0 ;
      RECT  129150.0 1888950.0 130050.0 1889850.0 ;
      RECT  129150.0 1890150.0 130050.0 1891050.0 ;
      RECT  129150.0 1889400.0 130050.0 1891050.0 ;
      RECT  129600.0 1888950.0 136200.0 1889850.0 ;
      RECT  136200.0 1888950.0 137400.0 1889850.0 ;
      RECT  145650.0 1888950.0 146550.0 1889850.0 ;
      RECT  145650.0 1890150.0 146550.0 1891050.0 ;
      RECT  141600.0 1888950.0 146100.0 1889850.0 ;
      RECT  145650.0 1889400.0 146550.0 1890600.0 ;
      RECT  146100.0 1890150.0 150600.0 1891050.0 ;
      RECT  121050.0 1903350.0 126600.0 1904250.0 ;
      RECT  129150.0 1904550.0 130050.0 1905450.0 ;
      RECT  129150.0 1903350.0 130050.0 1904250.0 ;
      RECT  129150.0 1904250.0 130050.0 1905000.0 ;
      RECT  129600.0 1904550.0 136200.0 1905450.0 ;
      RECT  136200.0 1904550.0 137400.0 1905450.0 ;
      RECT  145650.0 1904550.0 146550.0 1905450.0 ;
      RECT  145650.0 1903350.0 146550.0 1904250.0 ;
      RECT  141600.0 1904550.0 146100.0 1905450.0 ;
      RECT  145650.0 1903800.0 146550.0 1905000.0 ;
      RECT  146100.0 1903350.0 150600.0 1904250.0 ;
      RECT  121050.0 1917750.0 126600.0 1918650.0 ;
      RECT  129150.0 1916550.0 130050.0 1917450.0 ;
      RECT  129150.0 1917750.0 130050.0 1918650.0 ;
      RECT  129150.0 1917000.0 130050.0 1918650.0 ;
      RECT  129600.0 1916550.0 136200.0 1917450.0 ;
      RECT  136200.0 1916550.0 137400.0 1917450.0 ;
      RECT  145650.0 1916550.0 146550.0 1917450.0 ;
      RECT  145650.0 1917750.0 146550.0 1918650.0 ;
      RECT  141600.0 1916550.0 146100.0 1917450.0 ;
      RECT  145650.0 1917000.0 146550.0 1918200.0 ;
      RECT  146100.0 1917750.0 150600.0 1918650.0 ;
      RECT  121050.0 1930950.0 126600.0 1931850.0 ;
      RECT  129150.0 1932150.0 130050.0 1933050.0 ;
      RECT  129150.0 1930950.0 130050.0 1931850.0 ;
      RECT  129150.0 1931850.0 130050.0 1932600.0 ;
      RECT  129600.0 1932150.0 136200.0 1933050.0 ;
      RECT  136200.0 1932150.0 137400.0 1933050.0 ;
      RECT  145650.0 1932150.0 146550.0 1933050.0 ;
      RECT  145650.0 1930950.0 146550.0 1931850.0 ;
      RECT  141600.0 1932150.0 146100.0 1933050.0 ;
      RECT  145650.0 1931400.0 146550.0 1932600.0 ;
      RECT  146100.0 1930950.0 150600.0 1931850.0 ;
      RECT  121050.0 1945350.0 126600.0 1946250.0 ;
      RECT  129150.0 1944150.0 130050.0 1945050.0 ;
      RECT  129150.0 1945350.0 130050.0 1946250.0 ;
      RECT  129150.0 1944600.0 130050.0 1946250.0 ;
      RECT  129600.0 1944150.0 136200.0 1945050.0 ;
      RECT  136200.0 1944150.0 137400.0 1945050.0 ;
      RECT  145650.0 1944150.0 146550.0 1945050.0 ;
      RECT  145650.0 1945350.0 146550.0 1946250.0 ;
      RECT  141600.0 1944150.0 146100.0 1945050.0 ;
      RECT  145650.0 1944600.0 146550.0 1945800.0 ;
      RECT  146100.0 1945350.0 150600.0 1946250.0 ;
      RECT  121050.0 1958550.0 126600.0 1959450.0 ;
      RECT  129150.0 1959750.0 130050.0 1960650.0 ;
      RECT  129150.0 1958550.0 130050.0 1959450.0 ;
      RECT  129150.0 1959450.0 130050.0 1960200.0 ;
      RECT  129600.0 1959750.0 136200.0 1960650.0 ;
      RECT  136200.0 1959750.0 137400.0 1960650.0 ;
      RECT  145650.0 1959750.0 146550.0 1960650.0 ;
      RECT  145650.0 1958550.0 146550.0 1959450.0 ;
      RECT  141600.0 1959750.0 146100.0 1960650.0 ;
      RECT  145650.0 1959000.0 146550.0 1960200.0 ;
      RECT  146100.0 1958550.0 150600.0 1959450.0 ;
      RECT  121050.0 1972950.0 126600.0 1973850.0 ;
      RECT  129150.0 1971750.0 130050.0 1972650.0 ;
      RECT  129150.0 1972950.0 130050.0 1973850.0 ;
      RECT  129150.0 1972200.0 130050.0 1973850.0 ;
      RECT  129600.0 1971750.0 136200.0 1972650.0 ;
      RECT  136200.0 1971750.0 137400.0 1972650.0 ;
      RECT  145650.0 1971750.0 146550.0 1972650.0 ;
      RECT  145650.0 1972950.0 146550.0 1973850.0 ;
      RECT  141600.0 1971750.0 146100.0 1972650.0 ;
      RECT  145650.0 1972200.0 146550.0 1973400.0 ;
      RECT  146100.0 1972950.0 150600.0 1973850.0 ;
      RECT  121050.0 1986150.0 126600.0 1987050.0 ;
      RECT  129150.0 1987350.0 130050.0 1988250.0 ;
      RECT  129150.0 1986150.0 130050.0 1987050.0 ;
      RECT  129150.0 1987050.0 130050.0 1987800.0 ;
      RECT  129600.0 1987350.0 136200.0 1988250.0 ;
      RECT  136200.0 1987350.0 137400.0 1988250.0 ;
      RECT  145650.0 1987350.0 146550.0 1988250.0 ;
      RECT  145650.0 1986150.0 146550.0 1987050.0 ;
      RECT  141600.0 1987350.0 146100.0 1988250.0 ;
      RECT  145650.0 1986600.0 146550.0 1987800.0 ;
      RECT  146100.0 1986150.0 150600.0 1987050.0 ;
      RECT  121050.0 2000550.0 126600.0 2001450.0 ;
      RECT  129150.0 1999350.0 130050.0 2000250.0 ;
      RECT  129150.0 2000550.0 130050.0 2001450.0 ;
      RECT  129150.0 1999800.0 130050.0 2001450.0 ;
      RECT  129600.0 1999350.0 136200.0 2000250.0 ;
      RECT  136200.0 1999350.0 137400.0 2000250.0 ;
      RECT  145650.0 1999350.0 146550.0 2000250.0 ;
      RECT  145650.0 2000550.0 146550.0 2001450.0 ;
      RECT  141600.0 1999350.0 146100.0 2000250.0 ;
      RECT  145650.0 1999800.0 146550.0 2001000.0 ;
      RECT  146100.0 2000550.0 150600.0 2001450.0 ;
      RECT  121050.0 2013750.0 126600.0 2014650.0 ;
      RECT  129150.0 2014950.0 130050.0 2015850.0 ;
      RECT  129150.0 2013750.0 130050.0 2014650.0 ;
      RECT  129150.0 2014650.0 130050.0 2015400.0 ;
      RECT  129600.0 2014950.0 136200.0 2015850.0 ;
      RECT  136200.0 2014950.0 137400.0 2015850.0 ;
      RECT  145650.0 2014950.0 146550.0 2015850.0 ;
      RECT  145650.0 2013750.0 146550.0 2014650.0 ;
      RECT  141600.0 2014950.0 146100.0 2015850.0 ;
      RECT  145650.0 2014200.0 146550.0 2015400.0 ;
      RECT  146100.0 2013750.0 150600.0 2014650.0 ;
      RECT  121050.0 2028150.0 126600.0 2029050.0 ;
      RECT  129150.0 2026950.0 130050.0 2027850.0 ;
      RECT  129150.0 2028150.0 130050.0 2029050.0 ;
      RECT  129150.0 2027400.0 130050.0 2029050.0 ;
      RECT  129600.0 2026950.0 136200.0 2027850.0 ;
      RECT  136200.0 2026950.0 137400.0 2027850.0 ;
      RECT  145650.0 2026950.0 146550.0 2027850.0 ;
      RECT  145650.0 2028150.0 146550.0 2029050.0 ;
      RECT  141600.0 2026950.0 146100.0 2027850.0 ;
      RECT  145650.0 2027400.0 146550.0 2028600.0 ;
      RECT  146100.0 2028150.0 150600.0 2029050.0 ;
      RECT  121050.0 2041350.0 126600.0 2042250.0 ;
      RECT  129150.0 2042550.0 130050.0 2043450.0 ;
      RECT  129150.0 2041350.0 130050.0 2042250.0 ;
      RECT  129150.0 2042250.0 130050.0 2043000.0 ;
      RECT  129600.0 2042550.0 136200.0 2043450.0 ;
      RECT  136200.0 2042550.0 137400.0 2043450.0 ;
      RECT  145650.0 2042550.0 146550.0 2043450.0 ;
      RECT  145650.0 2041350.0 146550.0 2042250.0 ;
      RECT  141600.0 2042550.0 146100.0 2043450.0 ;
      RECT  145650.0 2041800.0 146550.0 2043000.0 ;
      RECT  146100.0 2041350.0 150600.0 2042250.0 ;
      RECT  121050.0 2055750.0 126600.0 2056650.0 ;
      RECT  129150.0 2054550.0 130050.0 2055450.0 ;
      RECT  129150.0 2055750.0 130050.0 2056650.0 ;
      RECT  129150.0 2055000.0 130050.0 2056650.0 ;
      RECT  129600.0 2054550.0 136200.0 2055450.0 ;
      RECT  136200.0 2054550.0 137400.0 2055450.0 ;
      RECT  145650.0 2054550.0 146550.0 2055450.0 ;
      RECT  145650.0 2055750.0 146550.0 2056650.0 ;
      RECT  141600.0 2054550.0 146100.0 2055450.0 ;
      RECT  145650.0 2055000.0 146550.0 2056200.0 ;
      RECT  146100.0 2055750.0 150600.0 2056650.0 ;
      RECT  121050.0 2068950.0 126600.0 2069850.0 ;
      RECT  129150.0 2070150.0 130050.0 2071050.0 ;
      RECT  129150.0 2068950.0 130050.0 2069850.0 ;
      RECT  129150.0 2069850.0 130050.0 2070600.0 ;
      RECT  129600.0 2070150.0 136200.0 2071050.0 ;
      RECT  136200.0 2070150.0 137400.0 2071050.0 ;
      RECT  145650.0 2070150.0 146550.0 2071050.0 ;
      RECT  145650.0 2068950.0 146550.0 2069850.0 ;
      RECT  141600.0 2070150.0 146100.0 2071050.0 ;
      RECT  145650.0 2069400.0 146550.0 2070600.0 ;
      RECT  146100.0 2068950.0 150600.0 2069850.0 ;
      RECT  121050.0 2083350.0 126600.0 2084250.0 ;
      RECT  129150.0 2082150.0 130050.0 2083050.0 ;
      RECT  129150.0 2083350.0 130050.0 2084250.0 ;
      RECT  129150.0 2082600.0 130050.0 2084250.0 ;
      RECT  129600.0 2082150.0 136200.0 2083050.0 ;
      RECT  136200.0 2082150.0 137400.0 2083050.0 ;
      RECT  145650.0 2082150.0 146550.0 2083050.0 ;
      RECT  145650.0 2083350.0 146550.0 2084250.0 ;
      RECT  141600.0 2082150.0 146100.0 2083050.0 ;
      RECT  145650.0 2082600.0 146550.0 2083800.0 ;
      RECT  146100.0 2083350.0 150600.0 2084250.0 ;
      RECT  121050.0 2096550.0 126600.0 2097450.0 ;
      RECT  129150.0 2097750.0 130050.0 2098650.0 ;
      RECT  129150.0 2096550.0 130050.0 2097450.0 ;
      RECT  129150.0 2097450.0 130050.0 2098200.0 ;
      RECT  129600.0 2097750.0 136200.0 2098650.0 ;
      RECT  136200.0 2097750.0 137400.0 2098650.0 ;
      RECT  145650.0 2097750.0 146550.0 2098650.0 ;
      RECT  145650.0 2096550.0 146550.0 2097450.0 ;
      RECT  141600.0 2097750.0 146100.0 2098650.0 ;
      RECT  145650.0 2097000.0 146550.0 2098200.0 ;
      RECT  146100.0 2096550.0 150600.0 2097450.0 ;
      RECT  121050.0 2110950.0 126600.0 2111850.0 ;
      RECT  129150.0 2109750.0 130050.0 2110650.0 ;
      RECT  129150.0 2110950.0 130050.0 2111850.0 ;
      RECT  129150.0 2110200.0 130050.0 2111850.0 ;
      RECT  129600.0 2109750.0 136200.0 2110650.0 ;
      RECT  136200.0 2109750.0 137400.0 2110650.0 ;
      RECT  145650.0 2109750.0 146550.0 2110650.0 ;
      RECT  145650.0 2110950.0 146550.0 2111850.0 ;
      RECT  141600.0 2109750.0 146100.0 2110650.0 ;
      RECT  145650.0 2110200.0 146550.0 2111400.0 ;
      RECT  146100.0 2110950.0 150600.0 2111850.0 ;
      RECT  121050.0 2124150.0 126600.0 2125050.0 ;
      RECT  129150.0 2125350.0 130050.0 2126250.0 ;
      RECT  129150.0 2124150.0 130050.0 2125050.0 ;
      RECT  129150.0 2125050.0 130050.0 2125800.0 ;
      RECT  129600.0 2125350.0 136200.0 2126250.0 ;
      RECT  136200.0 2125350.0 137400.0 2126250.0 ;
      RECT  145650.0 2125350.0 146550.0 2126250.0 ;
      RECT  145650.0 2124150.0 146550.0 2125050.0 ;
      RECT  141600.0 2125350.0 146100.0 2126250.0 ;
      RECT  145650.0 2124600.0 146550.0 2125800.0 ;
      RECT  146100.0 2124150.0 150600.0 2125050.0 ;
      RECT  121050.0 2138550.0 126600.0 2139450.0 ;
      RECT  129150.0 2137350.0 130050.0 2138250.0 ;
      RECT  129150.0 2138550.0 130050.0 2139450.0 ;
      RECT  129150.0 2137800.0 130050.0 2139450.0 ;
      RECT  129600.0 2137350.0 136200.0 2138250.0 ;
      RECT  136200.0 2137350.0 137400.0 2138250.0 ;
      RECT  145650.0 2137350.0 146550.0 2138250.0 ;
      RECT  145650.0 2138550.0 146550.0 2139450.0 ;
      RECT  141600.0 2137350.0 146100.0 2138250.0 ;
      RECT  145650.0 2137800.0 146550.0 2139000.0 ;
      RECT  146100.0 2138550.0 150600.0 2139450.0 ;
      RECT  130800.0 391050.0 132000.0 393000.0 ;
      RECT  130800.0 379200.0 132000.0 381150.0 ;
      RECT  126000.0 380550.0 127200.0 378750.0 ;
      RECT  126000.0 389850.0 127200.0 393450.0 ;
      RECT  128700.0 380550.0 129600.0 389850.0 ;
      RECT  126000.0 389850.0 127200.0 391050.0 ;
      RECT  128400.0 389850.0 129600.0 391050.0 ;
      RECT  128400.0 389850.0 129600.0 391050.0 ;
      RECT  126000.0 389850.0 127200.0 391050.0 ;
      RECT  126000.0 380550.0 127200.0 381750.0 ;
      RECT  128400.0 380550.0 129600.0 381750.0 ;
      RECT  128400.0 380550.0 129600.0 381750.0 ;
      RECT  126000.0 380550.0 127200.0 381750.0 ;
      RECT  130800.0 390450.0 132000.0 391650.0 ;
      RECT  130800.0 380550.0 132000.0 381750.0 ;
      RECT  126600.0 385200.0 127800.0 386400.0 ;
      RECT  126600.0 385200.0 127800.0 386400.0 ;
      RECT  129150.0 385350.0 130050.0 386250.0 ;
      RECT  124200.0 392550.0 133800.0 393450.0 ;
      RECT  124200.0 378750.0 133800.0 379650.0 ;
      RECT  135600.0 381150.0 136800.0 378750.0 ;
      RECT  135600.0 389850.0 136800.0 393450.0 ;
      RECT  140400.0 389850.0 141600.0 393450.0 ;
      RECT  142800.0 391050.0 144000.0 393000.0 ;
      RECT  142800.0 379200.0 144000.0 381150.0 ;
      RECT  135600.0 389850.0 136800.0 391050.0 ;
      RECT  138000.0 389850.0 139200.0 391050.0 ;
      RECT  138000.0 389850.0 139200.0 391050.0 ;
      RECT  135600.0 389850.0 136800.0 391050.0 ;
      RECT  138000.0 389850.0 139200.0 391050.0 ;
      RECT  140400.0 389850.0 141600.0 391050.0 ;
      RECT  140400.0 389850.0 141600.0 391050.0 ;
      RECT  138000.0 389850.0 139200.0 391050.0 ;
      RECT  135600.0 381150.0 136800.0 382350.0 ;
      RECT  138000.0 381150.0 139200.0 382350.0 ;
      RECT  138000.0 381150.0 139200.0 382350.0 ;
      RECT  135600.0 381150.0 136800.0 382350.0 ;
      RECT  138000.0 381150.0 139200.0 382350.0 ;
      RECT  140400.0 381150.0 141600.0 382350.0 ;
      RECT  140400.0 381150.0 141600.0 382350.0 ;
      RECT  138000.0 381150.0 139200.0 382350.0 ;
      RECT  142800.0 390450.0 144000.0 391650.0 ;
      RECT  142800.0 380550.0 144000.0 381750.0 ;
      RECT  140400.0 383700.0 139200.0 384900.0 ;
      RECT  137400.0 386400.0 136200.0 387600.0 ;
      RECT  138000.0 389850.0 139200.0 391050.0 ;
      RECT  140400.0 381150.0 141600.0 382350.0 ;
      RECT  141600.0 386400.0 140400.0 387600.0 ;
      RECT  136200.0 386400.0 137400.0 387600.0 ;
      RECT  139200.0 383700.0 140400.0 384900.0 ;
      RECT  140400.0 386400.0 141600.0 387600.0 ;
      RECT  133800.0 392550.0 148200.0 393450.0 ;
      RECT  133800.0 378750.0 148200.0 379650.0 ;
      RECT  154800.0 391050.0 156000.0 393000.0 ;
      RECT  154800.0 379200.0 156000.0 381150.0 ;
      RECT  150000.0 380550.0 151200.0 378750.0 ;
      RECT  150000.0 389850.0 151200.0 393450.0 ;
      RECT  152700.0 380550.0 153600.0 389850.0 ;
      RECT  150000.0 389850.0 151200.0 391050.0 ;
      RECT  152400.0 389850.0 153600.0 391050.0 ;
      RECT  152400.0 389850.0 153600.0 391050.0 ;
      RECT  150000.0 389850.0 151200.0 391050.0 ;
      RECT  150000.0 380550.0 151200.0 381750.0 ;
      RECT  152400.0 380550.0 153600.0 381750.0 ;
      RECT  152400.0 380550.0 153600.0 381750.0 ;
      RECT  150000.0 380550.0 151200.0 381750.0 ;
      RECT  154800.0 390450.0 156000.0 391650.0 ;
      RECT  154800.0 380550.0 156000.0 381750.0 ;
      RECT  150600.0 385200.0 151800.0 386400.0 ;
      RECT  150600.0 385200.0 151800.0 386400.0 ;
      RECT  153150.0 385350.0 154050.0 386250.0 ;
      RECT  148200.0 392550.0 157800.0 393450.0 ;
      RECT  148200.0 378750.0 157800.0 379650.0 ;
      RECT  120450.0 385200.0 121650.0 386400.0 ;
      RECT  122400.0 382800.0 123600.0 384000.0 ;
      RECT  139200.0 383700.0 138000.0 384900.0 ;
      RECT  130800.0 394950.0 132000.0 393000.0 ;
      RECT  130800.0 406800.0 132000.0 404850.0 ;
      RECT  126000.0 405450.0 127200.0 407250.0 ;
      RECT  126000.0 396150.0 127200.0 392550.0 ;
      RECT  128700.0 405450.0 129600.0 396150.0 ;
      RECT  126000.0 396150.0 127200.0 394950.0 ;
      RECT  128400.0 396150.0 129600.0 394950.0 ;
      RECT  128400.0 396150.0 129600.0 394950.0 ;
      RECT  126000.0 396150.0 127200.0 394950.0 ;
      RECT  126000.0 405450.0 127200.0 404250.0 ;
      RECT  128400.0 405450.0 129600.0 404250.0 ;
      RECT  128400.0 405450.0 129600.0 404250.0 ;
      RECT  126000.0 405450.0 127200.0 404250.0 ;
      RECT  130800.0 395550.0 132000.0 394350.0 ;
      RECT  130800.0 405450.0 132000.0 404250.0 ;
      RECT  126600.0 400800.0 127800.0 399600.0 ;
      RECT  126600.0 400800.0 127800.0 399600.0 ;
      RECT  129150.0 400650.0 130050.0 399750.0 ;
      RECT  124200.0 393450.0 133800.0 392550.0 ;
      RECT  124200.0 407250.0 133800.0 406350.0 ;
      RECT  135600.0 404850.0 136800.0 407250.0 ;
      RECT  135600.0 396150.0 136800.0 392550.0 ;
      RECT  140400.0 396150.0 141600.0 392550.0 ;
      RECT  142800.0 394950.0 144000.0 393000.0 ;
      RECT  142800.0 406800.0 144000.0 404850.0 ;
      RECT  135600.0 396150.0 136800.0 394950.0 ;
      RECT  138000.0 396150.0 139200.0 394950.0 ;
      RECT  138000.0 396150.0 139200.0 394950.0 ;
      RECT  135600.0 396150.0 136800.0 394950.0 ;
      RECT  138000.0 396150.0 139200.0 394950.0 ;
      RECT  140400.0 396150.0 141600.0 394950.0 ;
      RECT  140400.0 396150.0 141600.0 394950.0 ;
      RECT  138000.0 396150.0 139200.0 394950.0 ;
      RECT  135600.0 404850.0 136800.0 403650.0 ;
      RECT  138000.0 404850.0 139200.0 403650.0 ;
      RECT  138000.0 404850.0 139200.0 403650.0 ;
      RECT  135600.0 404850.0 136800.0 403650.0 ;
      RECT  138000.0 404850.0 139200.0 403650.0 ;
      RECT  140400.0 404850.0 141600.0 403650.0 ;
      RECT  140400.0 404850.0 141600.0 403650.0 ;
      RECT  138000.0 404850.0 139200.0 403650.0 ;
      RECT  142800.0 395550.0 144000.0 394350.0 ;
      RECT  142800.0 405450.0 144000.0 404250.0 ;
      RECT  140400.0 402300.0 139200.0 401100.0 ;
      RECT  137400.0 399600.0 136200.0 398400.0 ;
      RECT  138000.0 396150.0 139200.0 394950.0 ;
      RECT  140400.0 404850.0 141600.0 403650.0 ;
      RECT  141600.0 399600.0 140400.0 398400.0 ;
      RECT  136200.0 399600.0 137400.0 398400.0 ;
      RECT  139200.0 402300.0 140400.0 401100.0 ;
      RECT  140400.0 399600.0 141600.0 398400.0 ;
      RECT  133800.0 393450.0 148200.0 392550.0 ;
      RECT  133800.0 407250.0 148200.0 406350.0 ;
      RECT  154800.0 394950.0 156000.0 393000.0 ;
      RECT  154800.0 406800.0 156000.0 404850.0 ;
      RECT  150000.0 405450.0 151200.0 407250.0 ;
      RECT  150000.0 396150.0 151200.0 392550.0 ;
      RECT  152700.0 405450.0 153600.0 396150.0 ;
      RECT  150000.0 396150.0 151200.0 394950.0 ;
      RECT  152400.0 396150.0 153600.0 394950.0 ;
      RECT  152400.0 396150.0 153600.0 394950.0 ;
      RECT  150000.0 396150.0 151200.0 394950.0 ;
      RECT  150000.0 405450.0 151200.0 404250.0 ;
      RECT  152400.0 405450.0 153600.0 404250.0 ;
      RECT  152400.0 405450.0 153600.0 404250.0 ;
      RECT  150000.0 405450.0 151200.0 404250.0 ;
      RECT  154800.0 395550.0 156000.0 394350.0 ;
      RECT  154800.0 405450.0 156000.0 404250.0 ;
      RECT  150600.0 400800.0 151800.0 399600.0 ;
      RECT  150600.0 400800.0 151800.0 399600.0 ;
      RECT  153150.0 400650.0 154050.0 399750.0 ;
      RECT  148200.0 393450.0 157800.0 392550.0 ;
      RECT  148200.0 407250.0 157800.0 406350.0 ;
      RECT  120450.0 399600.0 121650.0 400800.0 ;
      RECT  122400.0 402000.0 123600.0 403200.0 ;
      RECT  139200.0 401100.0 138000.0 402300.0 ;
      RECT  130800.0 418650.0 132000.0 420600.0 ;
      RECT  130800.0 406800.0 132000.0 408750.0 ;
      RECT  126000.0 408150.0 127200.0 406350.0 ;
      RECT  126000.0 417450.0 127200.0 421050.0 ;
      RECT  128700.0 408150.0 129600.0 417450.0 ;
      RECT  126000.0 417450.0 127200.0 418650.0 ;
      RECT  128400.0 417450.0 129600.0 418650.0 ;
      RECT  128400.0 417450.0 129600.0 418650.0 ;
      RECT  126000.0 417450.0 127200.0 418650.0 ;
      RECT  126000.0 408150.0 127200.0 409350.0 ;
      RECT  128400.0 408150.0 129600.0 409350.0 ;
      RECT  128400.0 408150.0 129600.0 409350.0 ;
      RECT  126000.0 408150.0 127200.0 409350.0 ;
      RECT  130800.0 418050.0 132000.0 419250.0 ;
      RECT  130800.0 408150.0 132000.0 409350.0 ;
      RECT  126600.0 412800.0 127800.0 414000.0 ;
      RECT  126600.0 412800.0 127800.0 414000.0 ;
      RECT  129150.0 412950.0 130050.0 413850.0 ;
      RECT  124200.0 420150.0 133800.0 421050.0 ;
      RECT  124200.0 406350.0 133800.0 407250.0 ;
      RECT  135600.0 408750.0 136800.0 406350.0 ;
      RECT  135600.0 417450.0 136800.0 421050.0 ;
      RECT  140400.0 417450.0 141600.0 421050.0 ;
      RECT  142800.0 418650.0 144000.0 420600.0 ;
      RECT  142800.0 406800.0 144000.0 408750.0 ;
      RECT  135600.0 417450.0 136800.0 418650.0 ;
      RECT  138000.0 417450.0 139200.0 418650.0 ;
      RECT  138000.0 417450.0 139200.0 418650.0 ;
      RECT  135600.0 417450.0 136800.0 418650.0 ;
      RECT  138000.0 417450.0 139200.0 418650.0 ;
      RECT  140400.0 417450.0 141600.0 418650.0 ;
      RECT  140400.0 417450.0 141600.0 418650.0 ;
      RECT  138000.0 417450.0 139200.0 418650.0 ;
      RECT  135600.0 408750.0 136800.0 409950.0 ;
      RECT  138000.0 408750.0 139200.0 409950.0 ;
      RECT  138000.0 408750.0 139200.0 409950.0 ;
      RECT  135600.0 408750.0 136800.0 409950.0 ;
      RECT  138000.0 408750.0 139200.0 409950.0 ;
      RECT  140400.0 408750.0 141600.0 409950.0 ;
      RECT  140400.0 408750.0 141600.0 409950.0 ;
      RECT  138000.0 408750.0 139200.0 409950.0 ;
      RECT  142800.0 418050.0 144000.0 419250.0 ;
      RECT  142800.0 408150.0 144000.0 409350.0 ;
      RECT  140400.0 411300.0 139200.0 412500.0 ;
      RECT  137400.0 414000.0 136200.0 415200.0 ;
      RECT  138000.0 417450.0 139200.0 418650.0 ;
      RECT  140400.0 408750.0 141600.0 409950.0 ;
      RECT  141600.0 414000.0 140400.0 415200.0 ;
      RECT  136200.0 414000.0 137400.0 415200.0 ;
      RECT  139200.0 411300.0 140400.0 412500.0 ;
      RECT  140400.0 414000.0 141600.0 415200.0 ;
      RECT  133800.0 420150.0 148200.0 421050.0 ;
      RECT  133800.0 406350.0 148200.0 407250.0 ;
      RECT  154800.0 418650.0 156000.0 420600.0 ;
      RECT  154800.0 406800.0 156000.0 408750.0 ;
      RECT  150000.0 408150.0 151200.0 406350.0 ;
      RECT  150000.0 417450.0 151200.0 421050.0 ;
      RECT  152700.0 408150.0 153600.0 417450.0 ;
      RECT  150000.0 417450.0 151200.0 418650.0 ;
      RECT  152400.0 417450.0 153600.0 418650.0 ;
      RECT  152400.0 417450.0 153600.0 418650.0 ;
      RECT  150000.0 417450.0 151200.0 418650.0 ;
      RECT  150000.0 408150.0 151200.0 409350.0 ;
      RECT  152400.0 408150.0 153600.0 409350.0 ;
      RECT  152400.0 408150.0 153600.0 409350.0 ;
      RECT  150000.0 408150.0 151200.0 409350.0 ;
      RECT  154800.0 418050.0 156000.0 419250.0 ;
      RECT  154800.0 408150.0 156000.0 409350.0 ;
      RECT  150600.0 412800.0 151800.0 414000.0 ;
      RECT  150600.0 412800.0 151800.0 414000.0 ;
      RECT  153150.0 412950.0 154050.0 413850.0 ;
      RECT  148200.0 420150.0 157800.0 421050.0 ;
      RECT  148200.0 406350.0 157800.0 407250.0 ;
      RECT  120450.0 412800.0 121650.0 414000.0 ;
      RECT  122400.0 410400.0 123600.0 411600.0 ;
      RECT  139200.0 411300.0 138000.0 412500.0 ;
      RECT  130800.0 422550.0 132000.0 420600.0 ;
      RECT  130800.0 434400.0 132000.0 432450.0 ;
      RECT  126000.0 433050.0 127200.0 434850.0 ;
      RECT  126000.0 423750.0 127200.0 420150.0 ;
      RECT  128700.0 433050.0 129600.0 423750.0 ;
      RECT  126000.0 423750.0 127200.0 422550.0 ;
      RECT  128400.0 423750.0 129600.0 422550.0 ;
      RECT  128400.0 423750.0 129600.0 422550.0 ;
      RECT  126000.0 423750.0 127200.0 422550.0 ;
      RECT  126000.0 433050.0 127200.0 431850.0 ;
      RECT  128400.0 433050.0 129600.0 431850.0 ;
      RECT  128400.0 433050.0 129600.0 431850.0 ;
      RECT  126000.0 433050.0 127200.0 431850.0 ;
      RECT  130800.0 423150.0 132000.0 421950.0 ;
      RECT  130800.0 433050.0 132000.0 431850.0 ;
      RECT  126600.0 428400.0 127800.0 427200.0 ;
      RECT  126600.0 428400.0 127800.0 427200.0 ;
      RECT  129150.0 428250.0 130050.0 427350.0 ;
      RECT  124200.0 421050.0 133800.0 420150.0 ;
      RECT  124200.0 434850.0 133800.0 433950.0 ;
      RECT  135600.0 432450.0 136800.0 434850.0 ;
      RECT  135600.0 423750.0 136800.0 420150.0 ;
      RECT  140400.0 423750.0 141600.0 420150.0 ;
      RECT  142800.0 422550.0 144000.0 420600.0 ;
      RECT  142800.0 434400.0 144000.0 432450.0 ;
      RECT  135600.0 423750.0 136800.0 422550.0 ;
      RECT  138000.0 423750.0 139200.0 422550.0 ;
      RECT  138000.0 423750.0 139200.0 422550.0 ;
      RECT  135600.0 423750.0 136800.0 422550.0 ;
      RECT  138000.0 423750.0 139200.0 422550.0 ;
      RECT  140400.0 423750.0 141600.0 422550.0 ;
      RECT  140400.0 423750.0 141600.0 422550.0 ;
      RECT  138000.0 423750.0 139200.0 422550.0 ;
      RECT  135600.0 432450.0 136800.0 431250.0 ;
      RECT  138000.0 432450.0 139200.0 431250.0 ;
      RECT  138000.0 432450.0 139200.0 431250.0 ;
      RECT  135600.0 432450.0 136800.0 431250.0 ;
      RECT  138000.0 432450.0 139200.0 431250.0 ;
      RECT  140400.0 432450.0 141600.0 431250.0 ;
      RECT  140400.0 432450.0 141600.0 431250.0 ;
      RECT  138000.0 432450.0 139200.0 431250.0 ;
      RECT  142800.0 423150.0 144000.0 421950.0 ;
      RECT  142800.0 433050.0 144000.0 431850.0 ;
      RECT  140400.0 429900.0 139200.0 428700.0 ;
      RECT  137400.0 427200.0 136200.0 426000.0 ;
      RECT  138000.0 423750.0 139200.0 422550.0 ;
      RECT  140400.0 432450.0 141600.0 431250.0 ;
      RECT  141600.0 427200.0 140400.0 426000.0 ;
      RECT  136200.0 427200.0 137400.0 426000.0 ;
      RECT  139200.0 429900.0 140400.0 428700.0 ;
      RECT  140400.0 427200.0 141600.0 426000.0 ;
      RECT  133800.0 421050.0 148200.0 420150.0 ;
      RECT  133800.0 434850.0 148200.0 433950.0 ;
      RECT  154800.0 422550.0 156000.0 420600.0 ;
      RECT  154800.0 434400.0 156000.0 432450.0 ;
      RECT  150000.0 433050.0 151200.0 434850.0 ;
      RECT  150000.0 423750.0 151200.0 420150.0 ;
      RECT  152700.0 433050.0 153600.0 423750.0 ;
      RECT  150000.0 423750.0 151200.0 422550.0 ;
      RECT  152400.0 423750.0 153600.0 422550.0 ;
      RECT  152400.0 423750.0 153600.0 422550.0 ;
      RECT  150000.0 423750.0 151200.0 422550.0 ;
      RECT  150000.0 433050.0 151200.0 431850.0 ;
      RECT  152400.0 433050.0 153600.0 431850.0 ;
      RECT  152400.0 433050.0 153600.0 431850.0 ;
      RECT  150000.0 433050.0 151200.0 431850.0 ;
      RECT  154800.0 423150.0 156000.0 421950.0 ;
      RECT  154800.0 433050.0 156000.0 431850.0 ;
      RECT  150600.0 428400.0 151800.0 427200.0 ;
      RECT  150600.0 428400.0 151800.0 427200.0 ;
      RECT  153150.0 428250.0 154050.0 427350.0 ;
      RECT  148200.0 421050.0 157800.0 420150.0 ;
      RECT  148200.0 434850.0 157800.0 433950.0 ;
      RECT  120450.0 427200.0 121650.0 428400.0 ;
      RECT  122400.0 429600.0 123600.0 430800.0 ;
      RECT  139200.0 428700.0 138000.0 429900.0 ;
      RECT  130800.0 446250.0 132000.0 448200.0 ;
      RECT  130800.0 434400.0 132000.0 436350.0 ;
      RECT  126000.0 435750.0 127200.0 433950.0 ;
      RECT  126000.0 445050.0 127200.0 448650.0 ;
      RECT  128700.0 435750.0 129600.0 445050.0 ;
      RECT  126000.0 445050.0 127200.0 446250.0 ;
      RECT  128400.0 445050.0 129600.0 446250.0 ;
      RECT  128400.0 445050.0 129600.0 446250.0 ;
      RECT  126000.0 445050.0 127200.0 446250.0 ;
      RECT  126000.0 435750.0 127200.0 436950.0 ;
      RECT  128400.0 435750.0 129600.0 436950.0 ;
      RECT  128400.0 435750.0 129600.0 436950.0 ;
      RECT  126000.0 435750.0 127200.0 436950.0 ;
      RECT  130800.0 445650.0 132000.0 446850.0 ;
      RECT  130800.0 435750.0 132000.0 436950.0 ;
      RECT  126600.0 440400.0 127800.0 441600.0 ;
      RECT  126600.0 440400.0 127800.0 441600.0 ;
      RECT  129150.0 440550.0 130050.0 441450.0 ;
      RECT  124200.0 447750.0 133800.0 448650.0 ;
      RECT  124200.0 433950.0 133800.0 434850.0 ;
      RECT  135600.0 436350.0 136800.0 433950.0 ;
      RECT  135600.0 445050.0 136800.0 448650.0 ;
      RECT  140400.0 445050.0 141600.0 448650.0 ;
      RECT  142800.0 446250.0 144000.0 448200.0 ;
      RECT  142800.0 434400.0 144000.0 436350.0 ;
      RECT  135600.0 445050.0 136800.0 446250.0 ;
      RECT  138000.0 445050.0 139200.0 446250.0 ;
      RECT  138000.0 445050.0 139200.0 446250.0 ;
      RECT  135600.0 445050.0 136800.0 446250.0 ;
      RECT  138000.0 445050.0 139200.0 446250.0 ;
      RECT  140400.0 445050.0 141600.0 446250.0 ;
      RECT  140400.0 445050.0 141600.0 446250.0 ;
      RECT  138000.0 445050.0 139200.0 446250.0 ;
      RECT  135600.0 436350.0 136800.0 437550.0 ;
      RECT  138000.0 436350.0 139200.0 437550.0 ;
      RECT  138000.0 436350.0 139200.0 437550.0 ;
      RECT  135600.0 436350.0 136800.0 437550.0 ;
      RECT  138000.0 436350.0 139200.0 437550.0 ;
      RECT  140400.0 436350.0 141600.0 437550.0 ;
      RECT  140400.0 436350.0 141600.0 437550.0 ;
      RECT  138000.0 436350.0 139200.0 437550.0 ;
      RECT  142800.0 445650.0 144000.0 446850.0 ;
      RECT  142800.0 435750.0 144000.0 436950.0 ;
      RECT  140400.0 438900.0 139200.0 440100.0 ;
      RECT  137400.0 441600.0 136200.0 442800.0 ;
      RECT  138000.0 445050.0 139200.0 446250.0 ;
      RECT  140400.0 436350.0 141600.0 437550.0 ;
      RECT  141600.0 441600.0 140400.0 442800.0 ;
      RECT  136200.0 441600.0 137400.0 442800.0 ;
      RECT  139200.0 438900.0 140400.0 440100.0 ;
      RECT  140400.0 441600.0 141600.0 442800.0 ;
      RECT  133800.0 447750.0 148200.0 448650.0 ;
      RECT  133800.0 433950.0 148200.0 434850.0 ;
      RECT  154800.0 446250.0 156000.0 448200.0 ;
      RECT  154800.0 434400.0 156000.0 436350.0 ;
      RECT  150000.0 435750.0 151200.0 433950.0 ;
      RECT  150000.0 445050.0 151200.0 448650.0 ;
      RECT  152700.0 435750.0 153600.0 445050.0 ;
      RECT  150000.0 445050.0 151200.0 446250.0 ;
      RECT  152400.0 445050.0 153600.0 446250.0 ;
      RECT  152400.0 445050.0 153600.0 446250.0 ;
      RECT  150000.0 445050.0 151200.0 446250.0 ;
      RECT  150000.0 435750.0 151200.0 436950.0 ;
      RECT  152400.0 435750.0 153600.0 436950.0 ;
      RECT  152400.0 435750.0 153600.0 436950.0 ;
      RECT  150000.0 435750.0 151200.0 436950.0 ;
      RECT  154800.0 445650.0 156000.0 446850.0 ;
      RECT  154800.0 435750.0 156000.0 436950.0 ;
      RECT  150600.0 440400.0 151800.0 441600.0 ;
      RECT  150600.0 440400.0 151800.0 441600.0 ;
      RECT  153150.0 440550.0 154050.0 441450.0 ;
      RECT  148200.0 447750.0 157800.0 448650.0 ;
      RECT  148200.0 433950.0 157800.0 434850.0 ;
      RECT  120450.0 440400.0 121650.0 441600.0 ;
      RECT  122400.0 438000.0 123600.0 439200.0 ;
      RECT  139200.0 438900.0 138000.0 440100.0 ;
      RECT  130800.0 450150.0 132000.0 448200.0 ;
      RECT  130800.0 462000.0 132000.0 460050.0 ;
      RECT  126000.0 460650.0 127200.0 462450.0 ;
      RECT  126000.0 451350.0 127200.0 447750.0 ;
      RECT  128700.0 460650.0 129600.0 451350.0 ;
      RECT  126000.0 451350.0 127200.0 450150.0 ;
      RECT  128400.0 451350.0 129600.0 450150.0 ;
      RECT  128400.0 451350.0 129600.0 450150.0 ;
      RECT  126000.0 451350.0 127200.0 450150.0 ;
      RECT  126000.0 460650.0 127200.0 459450.0 ;
      RECT  128400.0 460650.0 129600.0 459450.0 ;
      RECT  128400.0 460650.0 129600.0 459450.0 ;
      RECT  126000.0 460650.0 127200.0 459450.0 ;
      RECT  130800.0 450750.0 132000.0 449550.0 ;
      RECT  130800.0 460650.0 132000.0 459450.0 ;
      RECT  126600.0 456000.0 127800.0 454800.0 ;
      RECT  126600.0 456000.0 127800.0 454800.0 ;
      RECT  129150.0 455850.0 130050.0 454950.0 ;
      RECT  124200.0 448650.0 133800.0 447750.0 ;
      RECT  124200.0 462450.0 133800.0 461550.0 ;
      RECT  135600.0 460050.0 136800.0 462450.0 ;
      RECT  135600.0 451350.0 136800.0 447750.0 ;
      RECT  140400.0 451350.0 141600.0 447750.0 ;
      RECT  142800.0 450150.0 144000.0 448200.0 ;
      RECT  142800.0 462000.0 144000.0 460050.0 ;
      RECT  135600.0 451350.0 136800.0 450150.0 ;
      RECT  138000.0 451350.0 139200.0 450150.0 ;
      RECT  138000.0 451350.0 139200.0 450150.0 ;
      RECT  135600.0 451350.0 136800.0 450150.0 ;
      RECT  138000.0 451350.0 139200.0 450150.0 ;
      RECT  140400.0 451350.0 141600.0 450150.0 ;
      RECT  140400.0 451350.0 141600.0 450150.0 ;
      RECT  138000.0 451350.0 139200.0 450150.0 ;
      RECT  135600.0 460050.0 136800.0 458850.0 ;
      RECT  138000.0 460050.0 139200.0 458850.0 ;
      RECT  138000.0 460050.0 139200.0 458850.0 ;
      RECT  135600.0 460050.0 136800.0 458850.0 ;
      RECT  138000.0 460050.0 139200.0 458850.0 ;
      RECT  140400.0 460050.0 141600.0 458850.0 ;
      RECT  140400.0 460050.0 141600.0 458850.0 ;
      RECT  138000.0 460050.0 139200.0 458850.0 ;
      RECT  142800.0 450750.0 144000.0 449550.0 ;
      RECT  142800.0 460650.0 144000.0 459450.0 ;
      RECT  140400.0 457500.0 139200.0 456300.0 ;
      RECT  137400.0 454800.0 136200.0 453600.0 ;
      RECT  138000.0 451350.0 139200.0 450150.0 ;
      RECT  140400.0 460050.0 141600.0 458850.0 ;
      RECT  141600.0 454800.0 140400.0 453600.0 ;
      RECT  136200.0 454800.0 137400.0 453600.0 ;
      RECT  139200.0 457500.0 140400.0 456300.0 ;
      RECT  140400.0 454800.0 141600.0 453600.0 ;
      RECT  133800.0 448650.0 148200.0 447750.0 ;
      RECT  133800.0 462450.0 148200.0 461550.0 ;
      RECT  154800.0 450150.0 156000.0 448200.0 ;
      RECT  154800.0 462000.0 156000.0 460050.0 ;
      RECT  150000.0 460650.0 151200.0 462450.0 ;
      RECT  150000.0 451350.0 151200.0 447750.0 ;
      RECT  152700.0 460650.0 153600.0 451350.0 ;
      RECT  150000.0 451350.0 151200.0 450150.0 ;
      RECT  152400.0 451350.0 153600.0 450150.0 ;
      RECT  152400.0 451350.0 153600.0 450150.0 ;
      RECT  150000.0 451350.0 151200.0 450150.0 ;
      RECT  150000.0 460650.0 151200.0 459450.0 ;
      RECT  152400.0 460650.0 153600.0 459450.0 ;
      RECT  152400.0 460650.0 153600.0 459450.0 ;
      RECT  150000.0 460650.0 151200.0 459450.0 ;
      RECT  154800.0 450750.0 156000.0 449550.0 ;
      RECT  154800.0 460650.0 156000.0 459450.0 ;
      RECT  150600.0 456000.0 151800.0 454800.0 ;
      RECT  150600.0 456000.0 151800.0 454800.0 ;
      RECT  153150.0 455850.0 154050.0 454950.0 ;
      RECT  148200.0 448650.0 157800.0 447750.0 ;
      RECT  148200.0 462450.0 157800.0 461550.0 ;
      RECT  120450.0 454800.0 121650.0 456000.0 ;
      RECT  122400.0 457200.0 123600.0 458400.0 ;
      RECT  139200.0 456300.0 138000.0 457500.0 ;
      RECT  130800.0 473850.0 132000.0 475800.0 ;
      RECT  130800.0 462000.0 132000.0 463950.0 ;
      RECT  126000.0 463350.0 127200.0 461550.0 ;
      RECT  126000.0 472650.0 127200.0 476250.0 ;
      RECT  128700.0 463350.0 129600.0 472650.0 ;
      RECT  126000.0 472650.0 127200.0 473850.0 ;
      RECT  128400.0 472650.0 129600.0 473850.0 ;
      RECT  128400.0 472650.0 129600.0 473850.0 ;
      RECT  126000.0 472650.0 127200.0 473850.0 ;
      RECT  126000.0 463350.0 127200.0 464550.0 ;
      RECT  128400.0 463350.0 129600.0 464550.0 ;
      RECT  128400.0 463350.0 129600.0 464550.0 ;
      RECT  126000.0 463350.0 127200.0 464550.0 ;
      RECT  130800.0 473250.0 132000.0 474450.0 ;
      RECT  130800.0 463350.0 132000.0 464550.0 ;
      RECT  126600.0 468000.0 127800.0 469200.0 ;
      RECT  126600.0 468000.0 127800.0 469200.0 ;
      RECT  129150.0 468150.0 130050.0 469050.0 ;
      RECT  124200.0 475350.0 133800.0 476250.0 ;
      RECT  124200.0 461550.0 133800.0 462450.0 ;
      RECT  135600.0 463950.0 136800.0 461550.0 ;
      RECT  135600.0 472650.0 136800.0 476250.0 ;
      RECT  140400.0 472650.0 141600.0 476250.0 ;
      RECT  142800.0 473850.0 144000.0 475800.0 ;
      RECT  142800.0 462000.0 144000.0 463950.0 ;
      RECT  135600.0 472650.0 136800.0 473850.0 ;
      RECT  138000.0 472650.0 139200.0 473850.0 ;
      RECT  138000.0 472650.0 139200.0 473850.0 ;
      RECT  135600.0 472650.0 136800.0 473850.0 ;
      RECT  138000.0 472650.0 139200.0 473850.0 ;
      RECT  140400.0 472650.0 141600.0 473850.0 ;
      RECT  140400.0 472650.0 141600.0 473850.0 ;
      RECT  138000.0 472650.0 139200.0 473850.0 ;
      RECT  135600.0 463950.0 136800.0 465150.0 ;
      RECT  138000.0 463950.0 139200.0 465150.0 ;
      RECT  138000.0 463950.0 139200.0 465150.0 ;
      RECT  135600.0 463950.0 136800.0 465150.0 ;
      RECT  138000.0 463950.0 139200.0 465150.0 ;
      RECT  140400.0 463950.0 141600.0 465150.0 ;
      RECT  140400.0 463950.0 141600.0 465150.0 ;
      RECT  138000.0 463950.0 139200.0 465150.0 ;
      RECT  142800.0 473250.0 144000.0 474450.0 ;
      RECT  142800.0 463350.0 144000.0 464550.0 ;
      RECT  140400.0 466500.0 139200.0 467700.0 ;
      RECT  137400.0 469200.0 136200.0 470400.0 ;
      RECT  138000.0 472650.0 139200.0 473850.0 ;
      RECT  140400.0 463950.0 141600.0 465150.0 ;
      RECT  141600.0 469200.0 140400.0 470400.0 ;
      RECT  136200.0 469200.0 137400.0 470400.0 ;
      RECT  139200.0 466500.0 140400.0 467700.0 ;
      RECT  140400.0 469200.0 141600.0 470400.0 ;
      RECT  133800.0 475350.0 148200.0 476250.0 ;
      RECT  133800.0 461550.0 148200.0 462450.0 ;
      RECT  154800.0 473850.0 156000.0 475800.0 ;
      RECT  154800.0 462000.0 156000.0 463950.0 ;
      RECT  150000.0 463350.0 151200.0 461550.0 ;
      RECT  150000.0 472650.0 151200.0 476250.0 ;
      RECT  152700.0 463350.0 153600.0 472650.0 ;
      RECT  150000.0 472650.0 151200.0 473850.0 ;
      RECT  152400.0 472650.0 153600.0 473850.0 ;
      RECT  152400.0 472650.0 153600.0 473850.0 ;
      RECT  150000.0 472650.0 151200.0 473850.0 ;
      RECT  150000.0 463350.0 151200.0 464550.0 ;
      RECT  152400.0 463350.0 153600.0 464550.0 ;
      RECT  152400.0 463350.0 153600.0 464550.0 ;
      RECT  150000.0 463350.0 151200.0 464550.0 ;
      RECT  154800.0 473250.0 156000.0 474450.0 ;
      RECT  154800.0 463350.0 156000.0 464550.0 ;
      RECT  150600.0 468000.0 151800.0 469200.0 ;
      RECT  150600.0 468000.0 151800.0 469200.0 ;
      RECT  153150.0 468150.0 154050.0 469050.0 ;
      RECT  148200.0 475350.0 157800.0 476250.0 ;
      RECT  148200.0 461550.0 157800.0 462450.0 ;
      RECT  120450.0 468000.0 121650.0 469200.0 ;
      RECT  122400.0 465600.0 123600.0 466800.0 ;
      RECT  139200.0 466500.0 138000.0 467700.0 ;
      RECT  130800.0 477750.0 132000.0 475800.0 ;
      RECT  130800.0 489600.0 132000.0 487650.0 ;
      RECT  126000.0 488250.0 127200.0 490050.0 ;
      RECT  126000.0 478950.0 127200.0 475350.0 ;
      RECT  128700.0 488250.0 129600.0 478950.0 ;
      RECT  126000.0 478950.0 127200.0 477750.0 ;
      RECT  128400.0 478950.0 129600.0 477750.0 ;
      RECT  128400.0 478950.0 129600.0 477750.0 ;
      RECT  126000.0 478950.0 127200.0 477750.0 ;
      RECT  126000.0 488250.0 127200.0 487050.0 ;
      RECT  128400.0 488250.0 129600.0 487050.0 ;
      RECT  128400.0 488250.0 129600.0 487050.0 ;
      RECT  126000.0 488250.0 127200.0 487050.0 ;
      RECT  130800.0 478350.0 132000.0 477150.0 ;
      RECT  130800.0 488250.0 132000.0 487050.0 ;
      RECT  126600.0 483600.0 127800.0 482400.0 ;
      RECT  126600.0 483600.0 127800.0 482400.0 ;
      RECT  129150.0 483450.0 130050.0 482550.0 ;
      RECT  124200.0 476250.0 133800.0 475350.0 ;
      RECT  124200.0 490050.0 133800.0 489150.0 ;
      RECT  135600.0 487650.0 136800.0 490050.0 ;
      RECT  135600.0 478950.0 136800.0 475350.0 ;
      RECT  140400.0 478950.0 141600.0 475350.0 ;
      RECT  142800.0 477750.0 144000.0 475800.0 ;
      RECT  142800.0 489600.0 144000.0 487650.0 ;
      RECT  135600.0 478950.0 136800.0 477750.0 ;
      RECT  138000.0 478950.0 139200.0 477750.0 ;
      RECT  138000.0 478950.0 139200.0 477750.0 ;
      RECT  135600.0 478950.0 136800.0 477750.0 ;
      RECT  138000.0 478950.0 139200.0 477750.0 ;
      RECT  140400.0 478950.0 141600.0 477750.0 ;
      RECT  140400.0 478950.0 141600.0 477750.0 ;
      RECT  138000.0 478950.0 139200.0 477750.0 ;
      RECT  135600.0 487650.0 136800.0 486450.0 ;
      RECT  138000.0 487650.0 139200.0 486450.0 ;
      RECT  138000.0 487650.0 139200.0 486450.0 ;
      RECT  135600.0 487650.0 136800.0 486450.0 ;
      RECT  138000.0 487650.0 139200.0 486450.0 ;
      RECT  140400.0 487650.0 141600.0 486450.0 ;
      RECT  140400.0 487650.0 141600.0 486450.0 ;
      RECT  138000.0 487650.0 139200.0 486450.0 ;
      RECT  142800.0 478350.0 144000.0 477150.0 ;
      RECT  142800.0 488250.0 144000.0 487050.0 ;
      RECT  140400.0 485100.0 139200.0 483900.0 ;
      RECT  137400.0 482400.0 136200.0 481200.0 ;
      RECT  138000.0 478950.0 139200.0 477750.0 ;
      RECT  140400.0 487650.0 141600.0 486450.0 ;
      RECT  141600.0 482400.0 140400.0 481200.0 ;
      RECT  136200.0 482400.0 137400.0 481200.0 ;
      RECT  139200.0 485100.0 140400.0 483900.0 ;
      RECT  140400.0 482400.0 141600.0 481200.0 ;
      RECT  133800.0 476250.0 148200.0 475350.0 ;
      RECT  133800.0 490050.0 148200.0 489150.0 ;
      RECT  154800.0 477750.0 156000.0 475800.0 ;
      RECT  154800.0 489600.0 156000.0 487650.0 ;
      RECT  150000.0 488250.0 151200.0 490050.0 ;
      RECT  150000.0 478950.0 151200.0 475350.0 ;
      RECT  152700.0 488250.0 153600.0 478950.0 ;
      RECT  150000.0 478950.0 151200.0 477750.0 ;
      RECT  152400.0 478950.0 153600.0 477750.0 ;
      RECT  152400.0 478950.0 153600.0 477750.0 ;
      RECT  150000.0 478950.0 151200.0 477750.0 ;
      RECT  150000.0 488250.0 151200.0 487050.0 ;
      RECT  152400.0 488250.0 153600.0 487050.0 ;
      RECT  152400.0 488250.0 153600.0 487050.0 ;
      RECT  150000.0 488250.0 151200.0 487050.0 ;
      RECT  154800.0 478350.0 156000.0 477150.0 ;
      RECT  154800.0 488250.0 156000.0 487050.0 ;
      RECT  150600.0 483600.0 151800.0 482400.0 ;
      RECT  150600.0 483600.0 151800.0 482400.0 ;
      RECT  153150.0 483450.0 154050.0 482550.0 ;
      RECT  148200.0 476250.0 157800.0 475350.0 ;
      RECT  148200.0 490050.0 157800.0 489150.0 ;
      RECT  120450.0 482400.0 121650.0 483600.0 ;
      RECT  122400.0 484800.0 123600.0 486000.0 ;
      RECT  139200.0 483900.0 138000.0 485100.0 ;
      RECT  130800.0 501450.0 132000.0 503400.0 ;
      RECT  130800.0 489600.0 132000.0 491550.0 ;
      RECT  126000.0 490950.0 127200.0 489150.0 ;
      RECT  126000.0 500250.0 127200.0 503850.0 ;
      RECT  128700.0 490950.0 129600.0 500250.0 ;
      RECT  126000.0 500250.0 127200.0 501450.0 ;
      RECT  128400.0 500250.0 129600.0 501450.0 ;
      RECT  128400.0 500250.0 129600.0 501450.0 ;
      RECT  126000.0 500250.0 127200.0 501450.0 ;
      RECT  126000.0 490950.0 127200.0 492150.0 ;
      RECT  128400.0 490950.0 129600.0 492150.0 ;
      RECT  128400.0 490950.0 129600.0 492150.0 ;
      RECT  126000.0 490950.0 127200.0 492150.0 ;
      RECT  130800.0 500850.0 132000.0 502050.0 ;
      RECT  130800.0 490950.0 132000.0 492150.0 ;
      RECT  126600.0 495600.0 127800.0 496800.0 ;
      RECT  126600.0 495600.0 127800.0 496800.0 ;
      RECT  129150.0 495750.0 130050.0 496650.0 ;
      RECT  124200.0 502950.0 133800.0 503850.0 ;
      RECT  124200.0 489150.0 133800.0 490050.0 ;
      RECT  135600.0 491550.0 136800.0 489150.0 ;
      RECT  135600.0 500250.0 136800.0 503850.0 ;
      RECT  140400.0 500250.0 141600.0 503850.0 ;
      RECT  142800.0 501450.0 144000.0 503400.0 ;
      RECT  142800.0 489600.0 144000.0 491550.0 ;
      RECT  135600.0 500250.0 136800.0 501450.0 ;
      RECT  138000.0 500250.0 139200.0 501450.0 ;
      RECT  138000.0 500250.0 139200.0 501450.0 ;
      RECT  135600.0 500250.0 136800.0 501450.0 ;
      RECT  138000.0 500250.0 139200.0 501450.0 ;
      RECT  140400.0 500250.0 141600.0 501450.0 ;
      RECT  140400.0 500250.0 141600.0 501450.0 ;
      RECT  138000.0 500250.0 139200.0 501450.0 ;
      RECT  135600.0 491550.0 136800.0 492750.0 ;
      RECT  138000.0 491550.0 139200.0 492750.0 ;
      RECT  138000.0 491550.0 139200.0 492750.0 ;
      RECT  135600.0 491550.0 136800.0 492750.0 ;
      RECT  138000.0 491550.0 139200.0 492750.0 ;
      RECT  140400.0 491550.0 141600.0 492750.0 ;
      RECT  140400.0 491550.0 141600.0 492750.0 ;
      RECT  138000.0 491550.0 139200.0 492750.0 ;
      RECT  142800.0 500850.0 144000.0 502050.0 ;
      RECT  142800.0 490950.0 144000.0 492150.0 ;
      RECT  140400.0 494100.0 139200.0 495300.0 ;
      RECT  137400.0 496800.0 136200.0 498000.0 ;
      RECT  138000.0 500250.0 139200.0 501450.0 ;
      RECT  140400.0 491550.0 141600.0 492750.0 ;
      RECT  141600.0 496800.0 140400.0 498000.0 ;
      RECT  136200.0 496800.0 137400.0 498000.0 ;
      RECT  139200.0 494100.0 140400.0 495300.0 ;
      RECT  140400.0 496800.0 141600.0 498000.0 ;
      RECT  133800.0 502950.0 148200.0 503850.0 ;
      RECT  133800.0 489150.0 148200.0 490050.0 ;
      RECT  154800.0 501450.0 156000.0 503400.0 ;
      RECT  154800.0 489600.0 156000.0 491550.0 ;
      RECT  150000.0 490950.0 151200.0 489150.0 ;
      RECT  150000.0 500250.0 151200.0 503850.0 ;
      RECT  152700.0 490950.0 153600.0 500250.0 ;
      RECT  150000.0 500250.0 151200.0 501450.0 ;
      RECT  152400.0 500250.0 153600.0 501450.0 ;
      RECT  152400.0 500250.0 153600.0 501450.0 ;
      RECT  150000.0 500250.0 151200.0 501450.0 ;
      RECT  150000.0 490950.0 151200.0 492150.0 ;
      RECT  152400.0 490950.0 153600.0 492150.0 ;
      RECT  152400.0 490950.0 153600.0 492150.0 ;
      RECT  150000.0 490950.0 151200.0 492150.0 ;
      RECT  154800.0 500850.0 156000.0 502050.0 ;
      RECT  154800.0 490950.0 156000.0 492150.0 ;
      RECT  150600.0 495600.0 151800.0 496800.0 ;
      RECT  150600.0 495600.0 151800.0 496800.0 ;
      RECT  153150.0 495750.0 154050.0 496650.0 ;
      RECT  148200.0 502950.0 157800.0 503850.0 ;
      RECT  148200.0 489150.0 157800.0 490050.0 ;
      RECT  120450.0 495600.0 121650.0 496800.0 ;
      RECT  122400.0 493200.0 123600.0 494400.0 ;
      RECT  139200.0 494100.0 138000.0 495300.0 ;
      RECT  130800.0 505350.0 132000.0 503400.0 ;
      RECT  130800.0 517200.0 132000.0 515250.0 ;
      RECT  126000.0 515850.0 127200.0 517650.0 ;
      RECT  126000.0 506550.0 127200.0 502950.0 ;
      RECT  128700.0 515850.0 129600.0 506550.0 ;
      RECT  126000.0 506550.0 127200.0 505350.0 ;
      RECT  128400.0 506550.0 129600.0 505350.0 ;
      RECT  128400.0 506550.0 129600.0 505350.0 ;
      RECT  126000.0 506550.0 127200.0 505350.0 ;
      RECT  126000.0 515850.0 127200.0 514650.0 ;
      RECT  128400.0 515850.0 129600.0 514650.0 ;
      RECT  128400.0 515850.0 129600.0 514650.0 ;
      RECT  126000.0 515850.0 127200.0 514650.0 ;
      RECT  130800.0 505950.0 132000.0 504750.0 ;
      RECT  130800.0 515850.0 132000.0 514650.0 ;
      RECT  126600.0 511200.0 127800.0 510000.0 ;
      RECT  126600.0 511200.0 127800.0 510000.0 ;
      RECT  129150.0 511050.0 130050.0 510150.0 ;
      RECT  124200.0 503850.0 133800.0 502950.0 ;
      RECT  124200.0 517650.0 133800.0 516750.0 ;
      RECT  135600.0 515250.0 136800.0 517650.0 ;
      RECT  135600.0 506550.0 136800.0 502950.0 ;
      RECT  140400.0 506550.0 141600.0 502950.0 ;
      RECT  142800.0 505350.0 144000.0 503400.0 ;
      RECT  142800.0 517200.0 144000.0 515250.0 ;
      RECT  135600.0 506550.0 136800.0 505350.0 ;
      RECT  138000.0 506550.0 139200.0 505350.0 ;
      RECT  138000.0 506550.0 139200.0 505350.0 ;
      RECT  135600.0 506550.0 136800.0 505350.0 ;
      RECT  138000.0 506550.0 139200.0 505350.0 ;
      RECT  140400.0 506550.0 141600.0 505350.0 ;
      RECT  140400.0 506550.0 141600.0 505350.0 ;
      RECT  138000.0 506550.0 139200.0 505350.0 ;
      RECT  135600.0 515250.0 136800.0 514050.0 ;
      RECT  138000.0 515250.0 139200.0 514050.0 ;
      RECT  138000.0 515250.0 139200.0 514050.0 ;
      RECT  135600.0 515250.0 136800.0 514050.0 ;
      RECT  138000.0 515250.0 139200.0 514050.0 ;
      RECT  140400.0 515250.0 141600.0 514050.0 ;
      RECT  140400.0 515250.0 141600.0 514050.0 ;
      RECT  138000.0 515250.0 139200.0 514050.0 ;
      RECT  142800.0 505950.0 144000.0 504750.0 ;
      RECT  142800.0 515850.0 144000.0 514650.0 ;
      RECT  140400.0 512700.0 139200.0 511500.0 ;
      RECT  137400.0 510000.0 136200.0 508800.0 ;
      RECT  138000.0 506550.0 139200.0 505350.0 ;
      RECT  140400.0 515250.0 141600.0 514050.0 ;
      RECT  141600.0 510000.0 140400.0 508800.0 ;
      RECT  136200.0 510000.0 137400.0 508800.0 ;
      RECT  139200.0 512700.0 140400.0 511500.0 ;
      RECT  140400.0 510000.0 141600.0 508800.0 ;
      RECT  133800.0 503850.0 148200.0 502950.0 ;
      RECT  133800.0 517650.0 148200.0 516750.0 ;
      RECT  154800.0 505350.0 156000.0 503400.0 ;
      RECT  154800.0 517200.0 156000.0 515250.0 ;
      RECT  150000.0 515850.0 151200.0 517650.0 ;
      RECT  150000.0 506550.0 151200.0 502950.0 ;
      RECT  152700.0 515850.0 153600.0 506550.0 ;
      RECT  150000.0 506550.0 151200.0 505350.0 ;
      RECT  152400.0 506550.0 153600.0 505350.0 ;
      RECT  152400.0 506550.0 153600.0 505350.0 ;
      RECT  150000.0 506550.0 151200.0 505350.0 ;
      RECT  150000.0 515850.0 151200.0 514650.0 ;
      RECT  152400.0 515850.0 153600.0 514650.0 ;
      RECT  152400.0 515850.0 153600.0 514650.0 ;
      RECT  150000.0 515850.0 151200.0 514650.0 ;
      RECT  154800.0 505950.0 156000.0 504750.0 ;
      RECT  154800.0 515850.0 156000.0 514650.0 ;
      RECT  150600.0 511200.0 151800.0 510000.0 ;
      RECT  150600.0 511200.0 151800.0 510000.0 ;
      RECT  153150.0 511050.0 154050.0 510150.0 ;
      RECT  148200.0 503850.0 157800.0 502950.0 ;
      RECT  148200.0 517650.0 157800.0 516750.0 ;
      RECT  120450.0 510000.0 121650.0 511200.0 ;
      RECT  122400.0 512400.0 123600.0 513600.0 ;
      RECT  139200.0 511500.0 138000.0 512700.0 ;
      RECT  130800.0 529050.0 132000.0 531000.0 ;
      RECT  130800.0 517200.0 132000.0 519150.0 ;
      RECT  126000.0 518550.0 127200.0 516750.0 ;
      RECT  126000.0 527850.0 127200.0 531450.0 ;
      RECT  128700.0 518550.0 129600.0 527850.0 ;
      RECT  126000.0 527850.0 127200.0 529050.0 ;
      RECT  128400.0 527850.0 129600.0 529050.0 ;
      RECT  128400.0 527850.0 129600.0 529050.0 ;
      RECT  126000.0 527850.0 127200.0 529050.0 ;
      RECT  126000.0 518550.0 127200.0 519750.0 ;
      RECT  128400.0 518550.0 129600.0 519750.0 ;
      RECT  128400.0 518550.0 129600.0 519750.0 ;
      RECT  126000.0 518550.0 127200.0 519750.0 ;
      RECT  130800.0 528450.0 132000.0 529650.0 ;
      RECT  130800.0 518550.0 132000.0 519750.0 ;
      RECT  126600.0 523200.0 127800.0 524400.0 ;
      RECT  126600.0 523200.0 127800.0 524400.0 ;
      RECT  129150.0 523350.0 130050.0 524250.0 ;
      RECT  124200.0 530550.0 133800.0 531450.0 ;
      RECT  124200.0 516750.0 133800.0 517650.0 ;
      RECT  135600.0 519150.0 136800.0 516750.0 ;
      RECT  135600.0 527850.0 136800.0 531450.0 ;
      RECT  140400.0 527850.0 141600.0 531450.0 ;
      RECT  142800.0 529050.0 144000.0 531000.0 ;
      RECT  142800.0 517200.0 144000.0 519150.0 ;
      RECT  135600.0 527850.0 136800.0 529050.0 ;
      RECT  138000.0 527850.0 139200.0 529050.0 ;
      RECT  138000.0 527850.0 139200.0 529050.0 ;
      RECT  135600.0 527850.0 136800.0 529050.0 ;
      RECT  138000.0 527850.0 139200.0 529050.0 ;
      RECT  140400.0 527850.0 141600.0 529050.0 ;
      RECT  140400.0 527850.0 141600.0 529050.0 ;
      RECT  138000.0 527850.0 139200.0 529050.0 ;
      RECT  135600.0 519150.0 136800.0 520350.0 ;
      RECT  138000.0 519150.0 139200.0 520350.0 ;
      RECT  138000.0 519150.0 139200.0 520350.0 ;
      RECT  135600.0 519150.0 136800.0 520350.0 ;
      RECT  138000.0 519150.0 139200.0 520350.0 ;
      RECT  140400.0 519150.0 141600.0 520350.0 ;
      RECT  140400.0 519150.0 141600.0 520350.0 ;
      RECT  138000.0 519150.0 139200.0 520350.0 ;
      RECT  142800.0 528450.0 144000.0 529650.0 ;
      RECT  142800.0 518550.0 144000.0 519750.0 ;
      RECT  140400.0 521700.0 139200.0 522900.0 ;
      RECT  137400.0 524400.0 136200.0 525600.0 ;
      RECT  138000.0 527850.0 139200.0 529050.0 ;
      RECT  140400.0 519150.0 141600.0 520350.0 ;
      RECT  141600.0 524400.0 140400.0 525600.0 ;
      RECT  136200.0 524400.0 137400.0 525600.0 ;
      RECT  139200.0 521700.0 140400.0 522900.0 ;
      RECT  140400.0 524400.0 141600.0 525600.0 ;
      RECT  133800.0 530550.0 148200.0 531450.0 ;
      RECT  133800.0 516750.0 148200.0 517650.0 ;
      RECT  154800.0 529050.0 156000.0 531000.0 ;
      RECT  154800.0 517200.0 156000.0 519150.0 ;
      RECT  150000.0 518550.0 151200.0 516750.0 ;
      RECT  150000.0 527850.0 151200.0 531450.0 ;
      RECT  152700.0 518550.0 153600.0 527850.0 ;
      RECT  150000.0 527850.0 151200.0 529050.0 ;
      RECT  152400.0 527850.0 153600.0 529050.0 ;
      RECT  152400.0 527850.0 153600.0 529050.0 ;
      RECT  150000.0 527850.0 151200.0 529050.0 ;
      RECT  150000.0 518550.0 151200.0 519750.0 ;
      RECT  152400.0 518550.0 153600.0 519750.0 ;
      RECT  152400.0 518550.0 153600.0 519750.0 ;
      RECT  150000.0 518550.0 151200.0 519750.0 ;
      RECT  154800.0 528450.0 156000.0 529650.0 ;
      RECT  154800.0 518550.0 156000.0 519750.0 ;
      RECT  150600.0 523200.0 151800.0 524400.0 ;
      RECT  150600.0 523200.0 151800.0 524400.0 ;
      RECT  153150.0 523350.0 154050.0 524250.0 ;
      RECT  148200.0 530550.0 157800.0 531450.0 ;
      RECT  148200.0 516750.0 157800.0 517650.0 ;
      RECT  120450.0 523200.0 121650.0 524400.0 ;
      RECT  122400.0 520800.0 123600.0 522000.0 ;
      RECT  139200.0 521700.0 138000.0 522900.0 ;
      RECT  130800.0 532950.0 132000.0 531000.0 ;
      RECT  130800.0 544800.0 132000.0 542850.0 ;
      RECT  126000.0 543450.0 127200.0 545250.0 ;
      RECT  126000.0 534150.0 127200.0 530550.0 ;
      RECT  128700.0 543450.0 129600.0 534150.0 ;
      RECT  126000.0 534150.0 127200.0 532950.0 ;
      RECT  128400.0 534150.0 129600.0 532950.0 ;
      RECT  128400.0 534150.0 129600.0 532950.0 ;
      RECT  126000.0 534150.0 127200.0 532950.0 ;
      RECT  126000.0 543450.0 127200.0 542250.0 ;
      RECT  128400.0 543450.0 129600.0 542250.0 ;
      RECT  128400.0 543450.0 129600.0 542250.0 ;
      RECT  126000.0 543450.0 127200.0 542250.0 ;
      RECT  130800.0 533550.0 132000.0 532350.0 ;
      RECT  130800.0 543450.0 132000.0 542250.0 ;
      RECT  126600.0 538800.0 127800.0 537600.0 ;
      RECT  126600.0 538800.0 127800.0 537600.0 ;
      RECT  129150.0 538650.0 130050.0 537750.0 ;
      RECT  124200.0 531450.0 133800.0 530550.0 ;
      RECT  124200.0 545250.0 133800.0 544350.0 ;
      RECT  135600.0 542850.0 136800.0 545250.0 ;
      RECT  135600.0 534150.0 136800.0 530550.0 ;
      RECT  140400.0 534150.0 141600.0 530550.0 ;
      RECT  142800.0 532950.0 144000.0 531000.0 ;
      RECT  142800.0 544800.0 144000.0 542850.0 ;
      RECT  135600.0 534150.0 136800.0 532950.0 ;
      RECT  138000.0 534150.0 139200.0 532950.0 ;
      RECT  138000.0 534150.0 139200.0 532950.0 ;
      RECT  135600.0 534150.0 136800.0 532950.0 ;
      RECT  138000.0 534150.0 139200.0 532950.0 ;
      RECT  140400.0 534150.0 141600.0 532950.0 ;
      RECT  140400.0 534150.0 141600.0 532950.0 ;
      RECT  138000.0 534150.0 139200.0 532950.0 ;
      RECT  135600.0 542850.0 136800.0 541650.0 ;
      RECT  138000.0 542850.0 139200.0 541650.0 ;
      RECT  138000.0 542850.0 139200.0 541650.0 ;
      RECT  135600.0 542850.0 136800.0 541650.0 ;
      RECT  138000.0 542850.0 139200.0 541650.0 ;
      RECT  140400.0 542850.0 141600.0 541650.0 ;
      RECT  140400.0 542850.0 141600.0 541650.0 ;
      RECT  138000.0 542850.0 139200.0 541650.0 ;
      RECT  142800.0 533550.0 144000.0 532350.0 ;
      RECT  142800.0 543450.0 144000.0 542250.0 ;
      RECT  140400.0 540300.0 139200.0 539100.0 ;
      RECT  137400.0 537600.0 136200.0 536400.0 ;
      RECT  138000.0 534150.0 139200.0 532950.0 ;
      RECT  140400.0 542850.0 141600.0 541650.0 ;
      RECT  141600.0 537600.0 140400.0 536400.0 ;
      RECT  136200.0 537600.0 137400.0 536400.0 ;
      RECT  139200.0 540300.0 140400.0 539100.0 ;
      RECT  140400.0 537600.0 141600.0 536400.0 ;
      RECT  133800.0 531450.0 148200.0 530550.0 ;
      RECT  133800.0 545250.0 148200.0 544350.0 ;
      RECT  154800.0 532950.0 156000.0 531000.0 ;
      RECT  154800.0 544800.0 156000.0 542850.0 ;
      RECT  150000.0 543450.0 151200.0 545250.0 ;
      RECT  150000.0 534150.0 151200.0 530550.0 ;
      RECT  152700.0 543450.0 153600.0 534150.0 ;
      RECT  150000.0 534150.0 151200.0 532950.0 ;
      RECT  152400.0 534150.0 153600.0 532950.0 ;
      RECT  152400.0 534150.0 153600.0 532950.0 ;
      RECT  150000.0 534150.0 151200.0 532950.0 ;
      RECT  150000.0 543450.0 151200.0 542250.0 ;
      RECT  152400.0 543450.0 153600.0 542250.0 ;
      RECT  152400.0 543450.0 153600.0 542250.0 ;
      RECT  150000.0 543450.0 151200.0 542250.0 ;
      RECT  154800.0 533550.0 156000.0 532350.0 ;
      RECT  154800.0 543450.0 156000.0 542250.0 ;
      RECT  150600.0 538800.0 151800.0 537600.0 ;
      RECT  150600.0 538800.0 151800.0 537600.0 ;
      RECT  153150.0 538650.0 154050.0 537750.0 ;
      RECT  148200.0 531450.0 157800.0 530550.0 ;
      RECT  148200.0 545250.0 157800.0 544350.0 ;
      RECT  120450.0 537600.0 121650.0 538800.0 ;
      RECT  122400.0 540000.0 123600.0 541200.0 ;
      RECT  139200.0 539100.0 138000.0 540300.0 ;
      RECT  130800.0 556650.0 132000.0 558600.0 ;
      RECT  130800.0 544800.0 132000.0 546750.0 ;
      RECT  126000.0 546150.0 127200.0 544350.0 ;
      RECT  126000.0 555450.0 127200.0 559050.0 ;
      RECT  128700.0 546150.0 129600.0 555450.0 ;
      RECT  126000.0 555450.0 127200.0 556650.0 ;
      RECT  128400.0 555450.0 129600.0 556650.0 ;
      RECT  128400.0 555450.0 129600.0 556650.0 ;
      RECT  126000.0 555450.0 127200.0 556650.0 ;
      RECT  126000.0 546150.0 127200.0 547350.0 ;
      RECT  128400.0 546150.0 129600.0 547350.0 ;
      RECT  128400.0 546150.0 129600.0 547350.0 ;
      RECT  126000.0 546150.0 127200.0 547350.0 ;
      RECT  130800.0 556050.0 132000.0 557250.0 ;
      RECT  130800.0 546150.0 132000.0 547350.0 ;
      RECT  126600.0 550800.0 127800.0 552000.0 ;
      RECT  126600.0 550800.0 127800.0 552000.0 ;
      RECT  129150.0 550950.0 130050.0 551850.0 ;
      RECT  124200.0 558150.0 133800.0 559050.0 ;
      RECT  124200.0 544350.0 133800.0 545250.0 ;
      RECT  135600.0 546750.0 136800.0 544350.0 ;
      RECT  135600.0 555450.0 136800.0 559050.0 ;
      RECT  140400.0 555450.0 141600.0 559050.0 ;
      RECT  142800.0 556650.0 144000.0 558600.0 ;
      RECT  142800.0 544800.0 144000.0 546750.0 ;
      RECT  135600.0 555450.0 136800.0 556650.0 ;
      RECT  138000.0 555450.0 139200.0 556650.0 ;
      RECT  138000.0 555450.0 139200.0 556650.0 ;
      RECT  135600.0 555450.0 136800.0 556650.0 ;
      RECT  138000.0 555450.0 139200.0 556650.0 ;
      RECT  140400.0 555450.0 141600.0 556650.0 ;
      RECT  140400.0 555450.0 141600.0 556650.0 ;
      RECT  138000.0 555450.0 139200.0 556650.0 ;
      RECT  135600.0 546750.0 136800.0 547950.0 ;
      RECT  138000.0 546750.0 139200.0 547950.0 ;
      RECT  138000.0 546750.0 139200.0 547950.0 ;
      RECT  135600.0 546750.0 136800.0 547950.0 ;
      RECT  138000.0 546750.0 139200.0 547950.0 ;
      RECT  140400.0 546750.0 141600.0 547950.0 ;
      RECT  140400.0 546750.0 141600.0 547950.0 ;
      RECT  138000.0 546750.0 139200.0 547950.0 ;
      RECT  142800.0 556050.0 144000.0 557250.0 ;
      RECT  142800.0 546150.0 144000.0 547350.0 ;
      RECT  140400.0 549300.0 139200.0 550500.0 ;
      RECT  137400.0 552000.0 136200.0 553200.0 ;
      RECT  138000.0 555450.0 139200.0 556650.0 ;
      RECT  140400.0 546750.0 141600.0 547950.0 ;
      RECT  141600.0 552000.0 140400.0 553200.0 ;
      RECT  136200.0 552000.0 137400.0 553200.0 ;
      RECT  139200.0 549300.0 140400.0 550500.0 ;
      RECT  140400.0 552000.0 141600.0 553200.0 ;
      RECT  133800.0 558150.0 148200.0 559050.0 ;
      RECT  133800.0 544350.0 148200.0 545250.0 ;
      RECT  154800.0 556650.0 156000.0 558600.0 ;
      RECT  154800.0 544800.0 156000.0 546750.0 ;
      RECT  150000.0 546150.0 151200.0 544350.0 ;
      RECT  150000.0 555450.0 151200.0 559050.0 ;
      RECT  152700.0 546150.0 153600.0 555450.0 ;
      RECT  150000.0 555450.0 151200.0 556650.0 ;
      RECT  152400.0 555450.0 153600.0 556650.0 ;
      RECT  152400.0 555450.0 153600.0 556650.0 ;
      RECT  150000.0 555450.0 151200.0 556650.0 ;
      RECT  150000.0 546150.0 151200.0 547350.0 ;
      RECT  152400.0 546150.0 153600.0 547350.0 ;
      RECT  152400.0 546150.0 153600.0 547350.0 ;
      RECT  150000.0 546150.0 151200.0 547350.0 ;
      RECT  154800.0 556050.0 156000.0 557250.0 ;
      RECT  154800.0 546150.0 156000.0 547350.0 ;
      RECT  150600.0 550800.0 151800.0 552000.0 ;
      RECT  150600.0 550800.0 151800.0 552000.0 ;
      RECT  153150.0 550950.0 154050.0 551850.0 ;
      RECT  148200.0 558150.0 157800.0 559050.0 ;
      RECT  148200.0 544350.0 157800.0 545250.0 ;
      RECT  120450.0 550800.0 121650.0 552000.0 ;
      RECT  122400.0 548400.0 123600.0 549600.0 ;
      RECT  139200.0 549300.0 138000.0 550500.0 ;
      RECT  130800.0 560550.0 132000.0 558600.0 ;
      RECT  130800.0 572400.0 132000.0 570450.0 ;
      RECT  126000.0 571050.0 127200.0 572850.0 ;
      RECT  126000.0 561750.0 127200.0 558150.0 ;
      RECT  128700.0 571050.0 129600.0 561750.0 ;
      RECT  126000.0 561750.0 127200.0 560550.0 ;
      RECT  128400.0 561750.0 129600.0 560550.0 ;
      RECT  128400.0 561750.0 129600.0 560550.0 ;
      RECT  126000.0 561750.0 127200.0 560550.0 ;
      RECT  126000.0 571050.0 127200.0 569850.0 ;
      RECT  128400.0 571050.0 129600.0 569850.0 ;
      RECT  128400.0 571050.0 129600.0 569850.0 ;
      RECT  126000.0 571050.0 127200.0 569850.0 ;
      RECT  130800.0 561150.0 132000.0 559950.0 ;
      RECT  130800.0 571050.0 132000.0 569850.0 ;
      RECT  126600.0 566400.0 127800.0 565200.0 ;
      RECT  126600.0 566400.0 127800.0 565200.0 ;
      RECT  129150.0 566250.0 130050.0 565350.0 ;
      RECT  124200.0 559050.0 133800.0 558150.0 ;
      RECT  124200.0 572850.0 133800.0 571950.0 ;
      RECT  135600.0 570450.0 136800.0 572850.0 ;
      RECT  135600.0 561750.0 136800.0 558150.0 ;
      RECT  140400.0 561750.0 141600.0 558150.0 ;
      RECT  142800.0 560550.0 144000.0 558600.0 ;
      RECT  142800.0 572400.0 144000.0 570450.0 ;
      RECT  135600.0 561750.0 136800.0 560550.0 ;
      RECT  138000.0 561750.0 139200.0 560550.0 ;
      RECT  138000.0 561750.0 139200.0 560550.0 ;
      RECT  135600.0 561750.0 136800.0 560550.0 ;
      RECT  138000.0 561750.0 139200.0 560550.0 ;
      RECT  140400.0 561750.0 141600.0 560550.0 ;
      RECT  140400.0 561750.0 141600.0 560550.0 ;
      RECT  138000.0 561750.0 139200.0 560550.0 ;
      RECT  135600.0 570450.0 136800.0 569250.0 ;
      RECT  138000.0 570450.0 139200.0 569250.0 ;
      RECT  138000.0 570450.0 139200.0 569250.0 ;
      RECT  135600.0 570450.0 136800.0 569250.0 ;
      RECT  138000.0 570450.0 139200.0 569250.0 ;
      RECT  140400.0 570450.0 141600.0 569250.0 ;
      RECT  140400.0 570450.0 141600.0 569250.0 ;
      RECT  138000.0 570450.0 139200.0 569250.0 ;
      RECT  142800.0 561150.0 144000.0 559950.0 ;
      RECT  142800.0 571050.0 144000.0 569850.0 ;
      RECT  140400.0 567900.0 139200.0 566700.0 ;
      RECT  137400.0 565200.0 136200.0 564000.0 ;
      RECT  138000.0 561750.0 139200.0 560550.0 ;
      RECT  140400.0 570450.0 141600.0 569250.0 ;
      RECT  141600.0 565200.0 140400.0 564000.0 ;
      RECT  136200.0 565200.0 137400.0 564000.0 ;
      RECT  139200.0 567900.0 140400.0 566700.0 ;
      RECT  140400.0 565200.0 141600.0 564000.0 ;
      RECT  133800.0 559050.0 148200.0 558150.0 ;
      RECT  133800.0 572850.0 148200.0 571950.0 ;
      RECT  154800.0 560550.0 156000.0 558600.0 ;
      RECT  154800.0 572400.0 156000.0 570450.0 ;
      RECT  150000.0 571050.0 151200.0 572850.0 ;
      RECT  150000.0 561750.0 151200.0 558150.0 ;
      RECT  152700.0 571050.0 153600.0 561750.0 ;
      RECT  150000.0 561750.0 151200.0 560550.0 ;
      RECT  152400.0 561750.0 153600.0 560550.0 ;
      RECT  152400.0 561750.0 153600.0 560550.0 ;
      RECT  150000.0 561750.0 151200.0 560550.0 ;
      RECT  150000.0 571050.0 151200.0 569850.0 ;
      RECT  152400.0 571050.0 153600.0 569850.0 ;
      RECT  152400.0 571050.0 153600.0 569850.0 ;
      RECT  150000.0 571050.0 151200.0 569850.0 ;
      RECT  154800.0 561150.0 156000.0 559950.0 ;
      RECT  154800.0 571050.0 156000.0 569850.0 ;
      RECT  150600.0 566400.0 151800.0 565200.0 ;
      RECT  150600.0 566400.0 151800.0 565200.0 ;
      RECT  153150.0 566250.0 154050.0 565350.0 ;
      RECT  148200.0 559050.0 157800.0 558150.0 ;
      RECT  148200.0 572850.0 157800.0 571950.0 ;
      RECT  120450.0 565200.0 121650.0 566400.0 ;
      RECT  122400.0 567600.0 123600.0 568800.0 ;
      RECT  139200.0 566700.0 138000.0 567900.0 ;
      RECT  130800.0 584250.0 132000.0 586200.0 ;
      RECT  130800.0 572400.0 132000.0 574350.0 ;
      RECT  126000.0 573750.0 127200.0 571950.0 ;
      RECT  126000.0 583050.0 127200.0 586650.0 ;
      RECT  128700.0 573750.0 129600.0 583050.0 ;
      RECT  126000.0 583050.0 127200.0 584250.0 ;
      RECT  128400.0 583050.0 129600.0 584250.0 ;
      RECT  128400.0 583050.0 129600.0 584250.0 ;
      RECT  126000.0 583050.0 127200.0 584250.0 ;
      RECT  126000.0 573750.0 127200.0 574950.0 ;
      RECT  128400.0 573750.0 129600.0 574950.0 ;
      RECT  128400.0 573750.0 129600.0 574950.0 ;
      RECT  126000.0 573750.0 127200.0 574950.0 ;
      RECT  130800.0 583650.0 132000.0 584850.0 ;
      RECT  130800.0 573750.0 132000.0 574950.0 ;
      RECT  126600.0 578400.0 127800.0 579600.0 ;
      RECT  126600.0 578400.0 127800.0 579600.0 ;
      RECT  129150.0 578550.0 130050.0 579450.0 ;
      RECT  124200.0 585750.0 133800.0 586650.0 ;
      RECT  124200.0 571950.0 133800.0 572850.0 ;
      RECT  135600.0 574350.0 136800.0 571950.0 ;
      RECT  135600.0 583050.0 136800.0 586650.0 ;
      RECT  140400.0 583050.0 141600.0 586650.0 ;
      RECT  142800.0 584250.0 144000.0 586200.0 ;
      RECT  142800.0 572400.0 144000.0 574350.0 ;
      RECT  135600.0 583050.0 136800.0 584250.0 ;
      RECT  138000.0 583050.0 139200.0 584250.0 ;
      RECT  138000.0 583050.0 139200.0 584250.0 ;
      RECT  135600.0 583050.0 136800.0 584250.0 ;
      RECT  138000.0 583050.0 139200.0 584250.0 ;
      RECT  140400.0 583050.0 141600.0 584250.0 ;
      RECT  140400.0 583050.0 141600.0 584250.0 ;
      RECT  138000.0 583050.0 139200.0 584250.0 ;
      RECT  135600.0 574350.0 136800.0 575550.0 ;
      RECT  138000.0 574350.0 139200.0 575550.0 ;
      RECT  138000.0 574350.0 139200.0 575550.0 ;
      RECT  135600.0 574350.0 136800.0 575550.0 ;
      RECT  138000.0 574350.0 139200.0 575550.0 ;
      RECT  140400.0 574350.0 141600.0 575550.0 ;
      RECT  140400.0 574350.0 141600.0 575550.0 ;
      RECT  138000.0 574350.0 139200.0 575550.0 ;
      RECT  142800.0 583650.0 144000.0 584850.0 ;
      RECT  142800.0 573750.0 144000.0 574950.0 ;
      RECT  140400.0 576900.0 139200.0 578100.0 ;
      RECT  137400.0 579600.0 136200.0 580800.0 ;
      RECT  138000.0 583050.0 139200.0 584250.0 ;
      RECT  140400.0 574350.0 141600.0 575550.0 ;
      RECT  141600.0 579600.0 140400.0 580800.0 ;
      RECT  136200.0 579600.0 137400.0 580800.0 ;
      RECT  139200.0 576900.0 140400.0 578100.0 ;
      RECT  140400.0 579600.0 141600.0 580800.0 ;
      RECT  133800.0 585750.0 148200.0 586650.0 ;
      RECT  133800.0 571950.0 148200.0 572850.0 ;
      RECT  154800.0 584250.0 156000.0 586200.0 ;
      RECT  154800.0 572400.0 156000.0 574350.0 ;
      RECT  150000.0 573750.0 151200.0 571950.0 ;
      RECT  150000.0 583050.0 151200.0 586650.0 ;
      RECT  152700.0 573750.0 153600.0 583050.0 ;
      RECT  150000.0 583050.0 151200.0 584250.0 ;
      RECT  152400.0 583050.0 153600.0 584250.0 ;
      RECT  152400.0 583050.0 153600.0 584250.0 ;
      RECT  150000.0 583050.0 151200.0 584250.0 ;
      RECT  150000.0 573750.0 151200.0 574950.0 ;
      RECT  152400.0 573750.0 153600.0 574950.0 ;
      RECT  152400.0 573750.0 153600.0 574950.0 ;
      RECT  150000.0 573750.0 151200.0 574950.0 ;
      RECT  154800.0 583650.0 156000.0 584850.0 ;
      RECT  154800.0 573750.0 156000.0 574950.0 ;
      RECT  150600.0 578400.0 151800.0 579600.0 ;
      RECT  150600.0 578400.0 151800.0 579600.0 ;
      RECT  153150.0 578550.0 154050.0 579450.0 ;
      RECT  148200.0 585750.0 157800.0 586650.0 ;
      RECT  148200.0 571950.0 157800.0 572850.0 ;
      RECT  120450.0 578400.0 121650.0 579600.0 ;
      RECT  122400.0 576000.0 123600.0 577200.0 ;
      RECT  139200.0 576900.0 138000.0 578100.0 ;
      RECT  130800.0 588150.0 132000.0 586200.0 ;
      RECT  130800.0 600000.0 132000.0 598050.0 ;
      RECT  126000.0 598650.0 127200.0 600450.0 ;
      RECT  126000.0 589350.0 127200.0 585750.0 ;
      RECT  128700.0 598650.0 129600.0 589350.0 ;
      RECT  126000.0 589350.0 127200.0 588150.0 ;
      RECT  128400.0 589350.0 129600.0 588150.0 ;
      RECT  128400.0 589350.0 129600.0 588150.0 ;
      RECT  126000.0 589350.0 127200.0 588150.0 ;
      RECT  126000.0 598650.0 127200.0 597450.0 ;
      RECT  128400.0 598650.0 129600.0 597450.0 ;
      RECT  128400.0 598650.0 129600.0 597450.0 ;
      RECT  126000.0 598650.0 127200.0 597450.0 ;
      RECT  130800.0 588750.0 132000.0 587550.0 ;
      RECT  130800.0 598650.0 132000.0 597450.0 ;
      RECT  126600.0 594000.0 127800.0 592800.0 ;
      RECT  126600.0 594000.0 127800.0 592800.0 ;
      RECT  129150.0 593850.0 130050.0 592950.0 ;
      RECT  124200.0 586650.0 133800.0 585750.0 ;
      RECT  124200.0 600450.0 133800.0 599550.0 ;
      RECT  135600.0 598050.0 136800.0 600450.0 ;
      RECT  135600.0 589350.0 136800.0 585750.0 ;
      RECT  140400.0 589350.0 141600.0 585750.0 ;
      RECT  142800.0 588150.0 144000.0 586200.0 ;
      RECT  142800.0 600000.0 144000.0 598050.0 ;
      RECT  135600.0 589350.0 136800.0 588150.0 ;
      RECT  138000.0 589350.0 139200.0 588150.0 ;
      RECT  138000.0 589350.0 139200.0 588150.0 ;
      RECT  135600.0 589350.0 136800.0 588150.0 ;
      RECT  138000.0 589350.0 139200.0 588150.0 ;
      RECT  140400.0 589350.0 141600.0 588150.0 ;
      RECT  140400.0 589350.0 141600.0 588150.0 ;
      RECT  138000.0 589350.0 139200.0 588150.0 ;
      RECT  135600.0 598050.0 136800.0 596850.0 ;
      RECT  138000.0 598050.0 139200.0 596850.0 ;
      RECT  138000.0 598050.0 139200.0 596850.0 ;
      RECT  135600.0 598050.0 136800.0 596850.0 ;
      RECT  138000.0 598050.0 139200.0 596850.0 ;
      RECT  140400.0 598050.0 141600.0 596850.0 ;
      RECT  140400.0 598050.0 141600.0 596850.0 ;
      RECT  138000.0 598050.0 139200.0 596850.0 ;
      RECT  142800.0 588750.0 144000.0 587550.0 ;
      RECT  142800.0 598650.0 144000.0 597450.0 ;
      RECT  140400.0 595500.0 139200.0 594300.0 ;
      RECT  137400.0 592800.0 136200.0 591600.0 ;
      RECT  138000.0 589350.0 139200.0 588150.0 ;
      RECT  140400.0 598050.0 141600.0 596850.0 ;
      RECT  141600.0 592800.0 140400.0 591600.0 ;
      RECT  136200.0 592800.0 137400.0 591600.0 ;
      RECT  139200.0 595500.0 140400.0 594300.0 ;
      RECT  140400.0 592800.0 141600.0 591600.0 ;
      RECT  133800.0 586650.0 148200.0 585750.0 ;
      RECT  133800.0 600450.0 148200.0 599550.0 ;
      RECT  154800.0 588150.0 156000.0 586200.0 ;
      RECT  154800.0 600000.0 156000.0 598050.0 ;
      RECT  150000.0 598650.0 151200.0 600450.0 ;
      RECT  150000.0 589350.0 151200.0 585750.0 ;
      RECT  152700.0 598650.0 153600.0 589350.0 ;
      RECT  150000.0 589350.0 151200.0 588150.0 ;
      RECT  152400.0 589350.0 153600.0 588150.0 ;
      RECT  152400.0 589350.0 153600.0 588150.0 ;
      RECT  150000.0 589350.0 151200.0 588150.0 ;
      RECT  150000.0 598650.0 151200.0 597450.0 ;
      RECT  152400.0 598650.0 153600.0 597450.0 ;
      RECT  152400.0 598650.0 153600.0 597450.0 ;
      RECT  150000.0 598650.0 151200.0 597450.0 ;
      RECT  154800.0 588750.0 156000.0 587550.0 ;
      RECT  154800.0 598650.0 156000.0 597450.0 ;
      RECT  150600.0 594000.0 151800.0 592800.0 ;
      RECT  150600.0 594000.0 151800.0 592800.0 ;
      RECT  153150.0 593850.0 154050.0 592950.0 ;
      RECT  148200.0 586650.0 157800.0 585750.0 ;
      RECT  148200.0 600450.0 157800.0 599550.0 ;
      RECT  120450.0 592800.0 121650.0 594000.0 ;
      RECT  122400.0 595200.0 123600.0 596400.0 ;
      RECT  139200.0 594300.0 138000.0 595500.0 ;
      RECT  130800.0 611850.0 132000.0 613800.0 ;
      RECT  130800.0 600000.0 132000.0 601950.0 ;
      RECT  126000.0 601350.0 127200.0 599550.0 ;
      RECT  126000.0 610650.0 127200.0 614250.0 ;
      RECT  128700.0 601350.0 129600.0 610650.0 ;
      RECT  126000.0 610650.0 127200.0 611850.0 ;
      RECT  128400.0 610650.0 129600.0 611850.0 ;
      RECT  128400.0 610650.0 129600.0 611850.0 ;
      RECT  126000.0 610650.0 127200.0 611850.0 ;
      RECT  126000.0 601350.0 127200.0 602550.0 ;
      RECT  128400.0 601350.0 129600.0 602550.0 ;
      RECT  128400.0 601350.0 129600.0 602550.0 ;
      RECT  126000.0 601350.0 127200.0 602550.0 ;
      RECT  130800.0 611250.0 132000.0 612450.0 ;
      RECT  130800.0 601350.0 132000.0 602550.0 ;
      RECT  126600.0 606000.0 127800.0 607200.0 ;
      RECT  126600.0 606000.0 127800.0 607200.0 ;
      RECT  129150.0 606150.0 130050.0 607050.0 ;
      RECT  124200.0 613350.0 133800.0 614250.0 ;
      RECT  124200.0 599550.0 133800.0 600450.0 ;
      RECT  135600.0 601950.0 136800.0 599550.0 ;
      RECT  135600.0 610650.0 136800.0 614250.0 ;
      RECT  140400.0 610650.0 141600.0 614250.0 ;
      RECT  142800.0 611850.0 144000.0 613800.0 ;
      RECT  142800.0 600000.0 144000.0 601950.0 ;
      RECT  135600.0 610650.0 136800.0 611850.0 ;
      RECT  138000.0 610650.0 139200.0 611850.0 ;
      RECT  138000.0 610650.0 139200.0 611850.0 ;
      RECT  135600.0 610650.0 136800.0 611850.0 ;
      RECT  138000.0 610650.0 139200.0 611850.0 ;
      RECT  140400.0 610650.0 141600.0 611850.0 ;
      RECT  140400.0 610650.0 141600.0 611850.0 ;
      RECT  138000.0 610650.0 139200.0 611850.0 ;
      RECT  135600.0 601950.0 136800.0 603150.0 ;
      RECT  138000.0 601950.0 139200.0 603150.0 ;
      RECT  138000.0 601950.0 139200.0 603150.0 ;
      RECT  135600.0 601950.0 136800.0 603150.0 ;
      RECT  138000.0 601950.0 139200.0 603150.0 ;
      RECT  140400.0 601950.0 141600.0 603150.0 ;
      RECT  140400.0 601950.0 141600.0 603150.0 ;
      RECT  138000.0 601950.0 139200.0 603150.0 ;
      RECT  142800.0 611250.0 144000.0 612450.0 ;
      RECT  142800.0 601350.0 144000.0 602550.0 ;
      RECT  140400.0 604500.0 139200.0 605700.0 ;
      RECT  137400.0 607200.0 136200.0 608400.0 ;
      RECT  138000.0 610650.0 139200.0 611850.0 ;
      RECT  140400.0 601950.0 141600.0 603150.0 ;
      RECT  141600.0 607200.0 140400.0 608400.0 ;
      RECT  136200.0 607200.0 137400.0 608400.0 ;
      RECT  139200.0 604500.0 140400.0 605700.0 ;
      RECT  140400.0 607200.0 141600.0 608400.0 ;
      RECT  133800.0 613350.0 148200.0 614250.0 ;
      RECT  133800.0 599550.0 148200.0 600450.0 ;
      RECT  154800.0 611850.0 156000.0 613800.0 ;
      RECT  154800.0 600000.0 156000.0 601950.0 ;
      RECT  150000.0 601350.0 151200.0 599550.0 ;
      RECT  150000.0 610650.0 151200.0 614250.0 ;
      RECT  152700.0 601350.0 153600.0 610650.0 ;
      RECT  150000.0 610650.0 151200.0 611850.0 ;
      RECT  152400.0 610650.0 153600.0 611850.0 ;
      RECT  152400.0 610650.0 153600.0 611850.0 ;
      RECT  150000.0 610650.0 151200.0 611850.0 ;
      RECT  150000.0 601350.0 151200.0 602550.0 ;
      RECT  152400.0 601350.0 153600.0 602550.0 ;
      RECT  152400.0 601350.0 153600.0 602550.0 ;
      RECT  150000.0 601350.0 151200.0 602550.0 ;
      RECT  154800.0 611250.0 156000.0 612450.0 ;
      RECT  154800.0 601350.0 156000.0 602550.0 ;
      RECT  150600.0 606000.0 151800.0 607200.0 ;
      RECT  150600.0 606000.0 151800.0 607200.0 ;
      RECT  153150.0 606150.0 154050.0 607050.0 ;
      RECT  148200.0 613350.0 157800.0 614250.0 ;
      RECT  148200.0 599550.0 157800.0 600450.0 ;
      RECT  120450.0 606000.0 121650.0 607200.0 ;
      RECT  122400.0 603600.0 123600.0 604800.0 ;
      RECT  139200.0 604500.0 138000.0 605700.0 ;
      RECT  130800.0 615750.0 132000.0 613800.0 ;
      RECT  130800.0 627600.0 132000.0 625650.0 ;
      RECT  126000.0 626250.0 127200.0 628050.0 ;
      RECT  126000.0 616950.0 127200.0 613350.0 ;
      RECT  128700.0 626250.0 129600.0 616950.0 ;
      RECT  126000.0 616950.0 127200.0 615750.0 ;
      RECT  128400.0 616950.0 129600.0 615750.0 ;
      RECT  128400.0 616950.0 129600.0 615750.0 ;
      RECT  126000.0 616950.0 127200.0 615750.0 ;
      RECT  126000.0 626250.0 127200.0 625050.0 ;
      RECT  128400.0 626250.0 129600.0 625050.0 ;
      RECT  128400.0 626250.0 129600.0 625050.0 ;
      RECT  126000.0 626250.0 127200.0 625050.0 ;
      RECT  130800.0 616350.0 132000.0 615150.0 ;
      RECT  130800.0 626250.0 132000.0 625050.0 ;
      RECT  126600.0 621600.0 127800.0 620400.0 ;
      RECT  126600.0 621600.0 127800.0 620400.0 ;
      RECT  129150.0 621450.0 130050.0 620550.0 ;
      RECT  124200.0 614250.0 133800.0 613350.0 ;
      RECT  124200.0 628050.0 133800.0 627150.0 ;
      RECT  135600.0 625650.0 136800.0 628050.0 ;
      RECT  135600.0 616950.0 136800.0 613350.0 ;
      RECT  140400.0 616950.0 141600.0 613350.0 ;
      RECT  142800.0 615750.0 144000.0 613800.0 ;
      RECT  142800.0 627600.0 144000.0 625650.0 ;
      RECT  135600.0 616950.0 136800.0 615750.0 ;
      RECT  138000.0 616950.0 139200.0 615750.0 ;
      RECT  138000.0 616950.0 139200.0 615750.0 ;
      RECT  135600.0 616950.0 136800.0 615750.0 ;
      RECT  138000.0 616950.0 139200.0 615750.0 ;
      RECT  140400.0 616950.0 141600.0 615750.0 ;
      RECT  140400.0 616950.0 141600.0 615750.0 ;
      RECT  138000.0 616950.0 139200.0 615750.0 ;
      RECT  135600.0 625650.0 136800.0 624450.0 ;
      RECT  138000.0 625650.0 139200.0 624450.0 ;
      RECT  138000.0 625650.0 139200.0 624450.0 ;
      RECT  135600.0 625650.0 136800.0 624450.0 ;
      RECT  138000.0 625650.0 139200.0 624450.0 ;
      RECT  140400.0 625650.0 141600.0 624450.0 ;
      RECT  140400.0 625650.0 141600.0 624450.0 ;
      RECT  138000.0 625650.0 139200.0 624450.0 ;
      RECT  142800.0 616350.0 144000.0 615150.0 ;
      RECT  142800.0 626250.0 144000.0 625050.0 ;
      RECT  140400.0 623100.0 139200.0 621900.0 ;
      RECT  137400.0 620400.0 136200.0 619200.0 ;
      RECT  138000.0 616950.0 139200.0 615750.0 ;
      RECT  140400.0 625650.0 141600.0 624450.0 ;
      RECT  141600.0 620400.0 140400.0 619200.0 ;
      RECT  136200.0 620400.0 137400.0 619200.0 ;
      RECT  139200.0 623100.0 140400.0 621900.0 ;
      RECT  140400.0 620400.0 141600.0 619200.0 ;
      RECT  133800.0 614250.0 148200.0 613350.0 ;
      RECT  133800.0 628050.0 148200.0 627150.0 ;
      RECT  154800.0 615750.0 156000.0 613800.0 ;
      RECT  154800.0 627600.0 156000.0 625650.0 ;
      RECT  150000.0 626250.0 151200.0 628050.0 ;
      RECT  150000.0 616950.0 151200.0 613350.0 ;
      RECT  152700.0 626250.0 153600.0 616950.0 ;
      RECT  150000.0 616950.0 151200.0 615750.0 ;
      RECT  152400.0 616950.0 153600.0 615750.0 ;
      RECT  152400.0 616950.0 153600.0 615750.0 ;
      RECT  150000.0 616950.0 151200.0 615750.0 ;
      RECT  150000.0 626250.0 151200.0 625050.0 ;
      RECT  152400.0 626250.0 153600.0 625050.0 ;
      RECT  152400.0 626250.0 153600.0 625050.0 ;
      RECT  150000.0 626250.0 151200.0 625050.0 ;
      RECT  154800.0 616350.0 156000.0 615150.0 ;
      RECT  154800.0 626250.0 156000.0 625050.0 ;
      RECT  150600.0 621600.0 151800.0 620400.0 ;
      RECT  150600.0 621600.0 151800.0 620400.0 ;
      RECT  153150.0 621450.0 154050.0 620550.0 ;
      RECT  148200.0 614250.0 157800.0 613350.0 ;
      RECT  148200.0 628050.0 157800.0 627150.0 ;
      RECT  120450.0 620400.0 121650.0 621600.0 ;
      RECT  122400.0 622800.0 123600.0 624000.0 ;
      RECT  139200.0 621900.0 138000.0 623100.0 ;
      RECT  130800.0 639450.0 132000.0 641400.0 ;
      RECT  130800.0 627600.0 132000.0 629550.0 ;
      RECT  126000.0 628950.0 127200.0 627150.0 ;
      RECT  126000.0 638250.0 127200.0 641850.0 ;
      RECT  128700.0 628950.0 129600.0 638250.0 ;
      RECT  126000.0 638250.0 127200.0 639450.0 ;
      RECT  128400.0 638250.0 129600.0 639450.0 ;
      RECT  128400.0 638250.0 129600.0 639450.0 ;
      RECT  126000.0 638250.0 127200.0 639450.0 ;
      RECT  126000.0 628950.0 127200.0 630150.0 ;
      RECT  128400.0 628950.0 129600.0 630150.0 ;
      RECT  128400.0 628950.0 129600.0 630150.0 ;
      RECT  126000.0 628950.0 127200.0 630150.0 ;
      RECT  130800.0 638850.0 132000.0 640050.0 ;
      RECT  130800.0 628950.0 132000.0 630150.0 ;
      RECT  126600.0 633600.0 127800.0 634800.0 ;
      RECT  126600.0 633600.0 127800.0 634800.0 ;
      RECT  129150.0 633750.0 130050.0 634650.0 ;
      RECT  124200.0 640950.0 133800.0 641850.0 ;
      RECT  124200.0 627150.0 133800.0 628050.0 ;
      RECT  135600.0 629550.0 136800.0 627150.0 ;
      RECT  135600.0 638250.0 136800.0 641850.0 ;
      RECT  140400.0 638250.0 141600.0 641850.0 ;
      RECT  142800.0 639450.0 144000.0 641400.0 ;
      RECT  142800.0 627600.0 144000.0 629550.0 ;
      RECT  135600.0 638250.0 136800.0 639450.0 ;
      RECT  138000.0 638250.0 139200.0 639450.0 ;
      RECT  138000.0 638250.0 139200.0 639450.0 ;
      RECT  135600.0 638250.0 136800.0 639450.0 ;
      RECT  138000.0 638250.0 139200.0 639450.0 ;
      RECT  140400.0 638250.0 141600.0 639450.0 ;
      RECT  140400.0 638250.0 141600.0 639450.0 ;
      RECT  138000.0 638250.0 139200.0 639450.0 ;
      RECT  135600.0 629550.0 136800.0 630750.0 ;
      RECT  138000.0 629550.0 139200.0 630750.0 ;
      RECT  138000.0 629550.0 139200.0 630750.0 ;
      RECT  135600.0 629550.0 136800.0 630750.0 ;
      RECT  138000.0 629550.0 139200.0 630750.0 ;
      RECT  140400.0 629550.0 141600.0 630750.0 ;
      RECT  140400.0 629550.0 141600.0 630750.0 ;
      RECT  138000.0 629550.0 139200.0 630750.0 ;
      RECT  142800.0 638850.0 144000.0 640050.0 ;
      RECT  142800.0 628950.0 144000.0 630150.0 ;
      RECT  140400.0 632100.0 139200.0 633300.0 ;
      RECT  137400.0 634800.0 136200.0 636000.0 ;
      RECT  138000.0 638250.0 139200.0 639450.0 ;
      RECT  140400.0 629550.0 141600.0 630750.0 ;
      RECT  141600.0 634800.0 140400.0 636000.0 ;
      RECT  136200.0 634800.0 137400.0 636000.0 ;
      RECT  139200.0 632100.0 140400.0 633300.0 ;
      RECT  140400.0 634800.0 141600.0 636000.0 ;
      RECT  133800.0 640950.0 148200.0 641850.0 ;
      RECT  133800.0 627150.0 148200.0 628050.0 ;
      RECT  154800.0 639450.0 156000.0 641400.0 ;
      RECT  154800.0 627600.0 156000.0 629550.0 ;
      RECT  150000.0 628950.0 151200.0 627150.0 ;
      RECT  150000.0 638250.0 151200.0 641850.0 ;
      RECT  152700.0 628950.0 153600.0 638250.0 ;
      RECT  150000.0 638250.0 151200.0 639450.0 ;
      RECT  152400.0 638250.0 153600.0 639450.0 ;
      RECT  152400.0 638250.0 153600.0 639450.0 ;
      RECT  150000.0 638250.0 151200.0 639450.0 ;
      RECT  150000.0 628950.0 151200.0 630150.0 ;
      RECT  152400.0 628950.0 153600.0 630150.0 ;
      RECT  152400.0 628950.0 153600.0 630150.0 ;
      RECT  150000.0 628950.0 151200.0 630150.0 ;
      RECT  154800.0 638850.0 156000.0 640050.0 ;
      RECT  154800.0 628950.0 156000.0 630150.0 ;
      RECT  150600.0 633600.0 151800.0 634800.0 ;
      RECT  150600.0 633600.0 151800.0 634800.0 ;
      RECT  153150.0 633750.0 154050.0 634650.0 ;
      RECT  148200.0 640950.0 157800.0 641850.0 ;
      RECT  148200.0 627150.0 157800.0 628050.0 ;
      RECT  120450.0 633600.0 121650.0 634800.0 ;
      RECT  122400.0 631200.0 123600.0 632400.0 ;
      RECT  139200.0 632100.0 138000.0 633300.0 ;
      RECT  130800.0 643350.0 132000.0 641400.0 ;
      RECT  130800.0 655200.0 132000.0 653250.0 ;
      RECT  126000.0 653850.0 127200.0 655650.0 ;
      RECT  126000.0 644550.0 127200.0 640950.0 ;
      RECT  128700.0 653850.0 129600.0 644550.0 ;
      RECT  126000.0 644550.0 127200.0 643350.0 ;
      RECT  128400.0 644550.0 129600.0 643350.0 ;
      RECT  128400.0 644550.0 129600.0 643350.0 ;
      RECT  126000.0 644550.0 127200.0 643350.0 ;
      RECT  126000.0 653850.0 127200.0 652650.0 ;
      RECT  128400.0 653850.0 129600.0 652650.0 ;
      RECT  128400.0 653850.0 129600.0 652650.0 ;
      RECT  126000.0 653850.0 127200.0 652650.0 ;
      RECT  130800.0 643950.0 132000.0 642750.0 ;
      RECT  130800.0 653850.0 132000.0 652650.0 ;
      RECT  126600.0 649200.0 127800.0 648000.0 ;
      RECT  126600.0 649200.0 127800.0 648000.0 ;
      RECT  129150.0 649050.0 130050.0 648150.0 ;
      RECT  124200.0 641850.0 133800.0 640950.0 ;
      RECT  124200.0 655650.0 133800.0 654750.0 ;
      RECT  135600.0 653250.0 136800.0 655650.0 ;
      RECT  135600.0 644550.0 136800.0 640950.0 ;
      RECT  140400.0 644550.0 141600.0 640950.0 ;
      RECT  142800.0 643350.0 144000.0 641400.0 ;
      RECT  142800.0 655200.0 144000.0 653250.0 ;
      RECT  135600.0 644550.0 136800.0 643350.0 ;
      RECT  138000.0 644550.0 139200.0 643350.0 ;
      RECT  138000.0 644550.0 139200.0 643350.0 ;
      RECT  135600.0 644550.0 136800.0 643350.0 ;
      RECT  138000.0 644550.0 139200.0 643350.0 ;
      RECT  140400.0 644550.0 141600.0 643350.0 ;
      RECT  140400.0 644550.0 141600.0 643350.0 ;
      RECT  138000.0 644550.0 139200.0 643350.0 ;
      RECT  135600.0 653250.0 136800.0 652050.0 ;
      RECT  138000.0 653250.0 139200.0 652050.0 ;
      RECT  138000.0 653250.0 139200.0 652050.0 ;
      RECT  135600.0 653250.0 136800.0 652050.0 ;
      RECT  138000.0 653250.0 139200.0 652050.0 ;
      RECT  140400.0 653250.0 141600.0 652050.0 ;
      RECT  140400.0 653250.0 141600.0 652050.0 ;
      RECT  138000.0 653250.0 139200.0 652050.0 ;
      RECT  142800.0 643950.0 144000.0 642750.0 ;
      RECT  142800.0 653850.0 144000.0 652650.0 ;
      RECT  140400.0 650700.0 139200.0 649500.0 ;
      RECT  137400.0 648000.0 136200.0 646800.0 ;
      RECT  138000.0 644550.0 139200.0 643350.0 ;
      RECT  140400.0 653250.0 141600.0 652050.0 ;
      RECT  141600.0 648000.0 140400.0 646800.0 ;
      RECT  136200.0 648000.0 137400.0 646800.0 ;
      RECT  139200.0 650700.0 140400.0 649500.0 ;
      RECT  140400.0 648000.0 141600.0 646800.0 ;
      RECT  133800.0 641850.0 148200.0 640950.0 ;
      RECT  133800.0 655650.0 148200.0 654750.0 ;
      RECT  154800.0 643350.0 156000.0 641400.0 ;
      RECT  154800.0 655200.0 156000.0 653250.0 ;
      RECT  150000.0 653850.0 151200.0 655650.0 ;
      RECT  150000.0 644550.0 151200.0 640950.0 ;
      RECT  152700.0 653850.0 153600.0 644550.0 ;
      RECT  150000.0 644550.0 151200.0 643350.0 ;
      RECT  152400.0 644550.0 153600.0 643350.0 ;
      RECT  152400.0 644550.0 153600.0 643350.0 ;
      RECT  150000.0 644550.0 151200.0 643350.0 ;
      RECT  150000.0 653850.0 151200.0 652650.0 ;
      RECT  152400.0 653850.0 153600.0 652650.0 ;
      RECT  152400.0 653850.0 153600.0 652650.0 ;
      RECT  150000.0 653850.0 151200.0 652650.0 ;
      RECT  154800.0 643950.0 156000.0 642750.0 ;
      RECT  154800.0 653850.0 156000.0 652650.0 ;
      RECT  150600.0 649200.0 151800.0 648000.0 ;
      RECT  150600.0 649200.0 151800.0 648000.0 ;
      RECT  153150.0 649050.0 154050.0 648150.0 ;
      RECT  148200.0 641850.0 157800.0 640950.0 ;
      RECT  148200.0 655650.0 157800.0 654750.0 ;
      RECT  120450.0 648000.0 121650.0 649200.0 ;
      RECT  122400.0 650400.0 123600.0 651600.0 ;
      RECT  139200.0 649500.0 138000.0 650700.0 ;
      RECT  130800.0 667050.0 132000.0 669000.0 ;
      RECT  130800.0 655200.0 132000.0 657150.0 ;
      RECT  126000.0 656550.0 127200.0 654750.0 ;
      RECT  126000.0 665850.0 127200.0 669450.0 ;
      RECT  128700.0 656550.0 129600.0 665850.0 ;
      RECT  126000.0 665850.0 127200.0 667050.0 ;
      RECT  128400.0 665850.0 129600.0 667050.0 ;
      RECT  128400.0 665850.0 129600.0 667050.0 ;
      RECT  126000.0 665850.0 127200.0 667050.0 ;
      RECT  126000.0 656550.0 127200.0 657750.0 ;
      RECT  128400.0 656550.0 129600.0 657750.0 ;
      RECT  128400.0 656550.0 129600.0 657750.0 ;
      RECT  126000.0 656550.0 127200.0 657750.0 ;
      RECT  130800.0 666450.0 132000.0 667650.0 ;
      RECT  130800.0 656550.0 132000.0 657750.0 ;
      RECT  126600.0 661200.0 127800.0 662400.0 ;
      RECT  126600.0 661200.0 127800.0 662400.0 ;
      RECT  129150.0 661350.0 130050.0 662250.0 ;
      RECT  124200.0 668550.0 133800.0 669450.0 ;
      RECT  124200.0 654750.0 133800.0 655650.0 ;
      RECT  135600.0 657150.0 136800.0 654750.0 ;
      RECT  135600.0 665850.0 136800.0 669450.0 ;
      RECT  140400.0 665850.0 141600.0 669450.0 ;
      RECT  142800.0 667050.0 144000.0 669000.0 ;
      RECT  142800.0 655200.0 144000.0 657150.0 ;
      RECT  135600.0 665850.0 136800.0 667050.0 ;
      RECT  138000.0 665850.0 139200.0 667050.0 ;
      RECT  138000.0 665850.0 139200.0 667050.0 ;
      RECT  135600.0 665850.0 136800.0 667050.0 ;
      RECT  138000.0 665850.0 139200.0 667050.0 ;
      RECT  140400.0 665850.0 141600.0 667050.0 ;
      RECT  140400.0 665850.0 141600.0 667050.0 ;
      RECT  138000.0 665850.0 139200.0 667050.0 ;
      RECT  135600.0 657150.0 136800.0 658350.0 ;
      RECT  138000.0 657150.0 139200.0 658350.0 ;
      RECT  138000.0 657150.0 139200.0 658350.0 ;
      RECT  135600.0 657150.0 136800.0 658350.0 ;
      RECT  138000.0 657150.0 139200.0 658350.0 ;
      RECT  140400.0 657150.0 141600.0 658350.0 ;
      RECT  140400.0 657150.0 141600.0 658350.0 ;
      RECT  138000.0 657150.0 139200.0 658350.0 ;
      RECT  142800.0 666450.0 144000.0 667650.0 ;
      RECT  142800.0 656550.0 144000.0 657750.0 ;
      RECT  140400.0 659700.0 139200.0 660900.0 ;
      RECT  137400.0 662400.0 136200.0 663600.0 ;
      RECT  138000.0 665850.0 139200.0 667050.0 ;
      RECT  140400.0 657150.0 141600.0 658350.0 ;
      RECT  141600.0 662400.0 140400.0 663600.0 ;
      RECT  136200.0 662400.0 137400.0 663600.0 ;
      RECT  139200.0 659700.0 140400.0 660900.0 ;
      RECT  140400.0 662400.0 141600.0 663600.0 ;
      RECT  133800.0 668550.0 148200.0 669450.0 ;
      RECT  133800.0 654750.0 148200.0 655650.0 ;
      RECT  154800.0 667050.0 156000.0 669000.0 ;
      RECT  154800.0 655200.0 156000.0 657150.0 ;
      RECT  150000.0 656550.0 151200.0 654750.0 ;
      RECT  150000.0 665850.0 151200.0 669450.0 ;
      RECT  152700.0 656550.0 153600.0 665850.0 ;
      RECT  150000.0 665850.0 151200.0 667050.0 ;
      RECT  152400.0 665850.0 153600.0 667050.0 ;
      RECT  152400.0 665850.0 153600.0 667050.0 ;
      RECT  150000.0 665850.0 151200.0 667050.0 ;
      RECT  150000.0 656550.0 151200.0 657750.0 ;
      RECT  152400.0 656550.0 153600.0 657750.0 ;
      RECT  152400.0 656550.0 153600.0 657750.0 ;
      RECT  150000.0 656550.0 151200.0 657750.0 ;
      RECT  154800.0 666450.0 156000.0 667650.0 ;
      RECT  154800.0 656550.0 156000.0 657750.0 ;
      RECT  150600.0 661200.0 151800.0 662400.0 ;
      RECT  150600.0 661200.0 151800.0 662400.0 ;
      RECT  153150.0 661350.0 154050.0 662250.0 ;
      RECT  148200.0 668550.0 157800.0 669450.0 ;
      RECT  148200.0 654750.0 157800.0 655650.0 ;
      RECT  120450.0 661200.0 121650.0 662400.0 ;
      RECT  122400.0 658800.0 123600.0 660000.0 ;
      RECT  139200.0 659700.0 138000.0 660900.0 ;
      RECT  130800.0 670950.0 132000.0 669000.0 ;
      RECT  130800.0 682800.0 132000.0 680850.0 ;
      RECT  126000.0 681450.0 127200.0 683250.0 ;
      RECT  126000.0 672150.0 127200.0 668550.0 ;
      RECT  128700.0 681450.0 129600.0 672150.0 ;
      RECT  126000.0 672150.0 127200.0 670950.0 ;
      RECT  128400.0 672150.0 129600.0 670950.0 ;
      RECT  128400.0 672150.0 129600.0 670950.0 ;
      RECT  126000.0 672150.0 127200.0 670950.0 ;
      RECT  126000.0 681450.0 127200.0 680250.0 ;
      RECT  128400.0 681450.0 129600.0 680250.0 ;
      RECT  128400.0 681450.0 129600.0 680250.0 ;
      RECT  126000.0 681450.0 127200.0 680250.0 ;
      RECT  130800.0 671550.0 132000.0 670350.0 ;
      RECT  130800.0 681450.0 132000.0 680250.0 ;
      RECT  126600.0 676800.0 127800.0 675600.0 ;
      RECT  126600.0 676800.0 127800.0 675600.0 ;
      RECT  129150.0 676650.0 130050.0 675750.0 ;
      RECT  124200.0 669450.0 133800.0 668550.0 ;
      RECT  124200.0 683250.0 133800.0 682350.0 ;
      RECT  135600.0 680850.0 136800.0 683250.0 ;
      RECT  135600.0 672150.0 136800.0 668550.0 ;
      RECT  140400.0 672150.0 141600.0 668550.0 ;
      RECT  142800.0 670950.0 144000.0 669000.0 ;
      RECT  142800.0 682800.0 144000.0 680850.0 ;
      RECT  135600.0 672150.0 136800.0 670950.0 ;
      RECT  138000.0 672150.0 139200.0 670950.0 ;
      RECT  138000.0 672150.0 139200.0 670950.0 ;
      RECT  135600.0 672150.0 136800.0 670950.0 ;
      RECT  138000.0 672150.0 139200.0 670950.0 ;
      RECT  140400.0 672150.0 141600.0 670950.0 ;
      RECT  140400.0 672150.0 141600.0 670950.0 ;
      RECT  138000.0 672150.0 139200.0 670950.0 ;
      RECT  135600.0 680850.0 136800.0 679650.0 ;
      RECT  138000.0 680850.0 139200.0 679650.0 ;
      RECT  138000.0 680850.0 139200.0 679650.0 ;
      RECT  135600.0 680850.0 136800.0 679650.0 ;
      RECT  138000.0 680850.0 139200.0 679650.0 ;
      RECT  140400.0 680850.0 141600.0 679650.0 ;
      RECT  140400.0 680850.0 141600.0 679650.0 ;
      RECT  138000.0 680850.0 139200.0 679650.0 ;
      RECT  142800.0 671550.0 144000.0 670350.0 ;
      RECT  142800.0 681450.0 144000.0 680250.0 ;
      RECT  140400.0 678300.0 139200.0 677100.0 ;
      RECT  137400.0 675600.0 136200.0 674400.0 ;
      RECT  138000.0 672150.0 139200.0 670950.0 ;
      RECT  140400.0 680850.0 141600.0 679650.0 ;
      RECT  141600.0 675600.0 140400.0 674400.0 ;
      RECT  136200.0 675600.0 137400.0 674400.0 ;
      RECT  139200.0 678300.0 140400.0 677100.0 ;
      RECT  140400.0 675600.0 141600.0 674400.0 ;
      RECT  133800.0 669450.0 148200.0 668550.0 ;
      RECT  133800.0 683250.0 148200.0 682350.0 ;
      RECT  154800.0 670950.0 156000.0 669000.0 ;
      RECT  154800.0 682800.0 156000.0 680850.0 ;
      RECT  150000.0 681450.0 151200.0 683250.0 ;
      RECT  150000.0 672150.0 151200.0 668550.0 ;
      RECT  152700.0 681450.0 153600.0 672150.0 ;
      RECT  150000.0 672150.0 151200.0 670950.0 ;
      RECT  152400.0 672150.0 153600.0 670950.0 ;
      RECT  152400.0 672150.0 153600.0 670950.0 ;
      RECT  150000.0 672150.0 151200.0 670950.0 ;
      RECT  150000.0 681450.0 151200.0 680250.0 ;
      RECT  152400.0 681450.0 153600.0 680250.0 ;
      RECT  152400.0 681450.0 153600.0 680250.0 ;
      RECT  150000.0 681450.0 151200.0 680250.0 ;
      RECT  154800.0 671550.0 156000.0 670350.0 ;
      RECT  154800.0 681450.0 156000.0 680250.0 ;
      RECT  150600.0 676800.0 151800.0 675600.0 ;
      RECT  150600.0 676800.0 151800.0 675600.0 ;
      RECT  153150.0 676650.0 154050.0 675750.0 ;
      RECT  148200.0 669450.0 157800.0 668550.0 ;
      RECT  148200.0 683250.0 157800.0 682350.0 ;
      RECT  120450.0 675600.0 121650.0 676800.0 ;
      RECT  122400.0 678000.0 123600.0 679200.0 ;
      RECT  139200.0 677100.0 138000.0 678300.0 ;
      RECT  130800.0 694650.0 132000.0 696600.0 ;
      RECT  130800.0 682800.0 132000.0 684750.0 ;
      RECT  126000.0 684150.0 127200.0 682350.0 ;
      RECT  126000.0 693450.0 127200.0 697050.0 ;
      RECT  128700.0 684150.0 129600.0 693450.0 ;
      RECT  126000.0 693450.0 127200.0 694650.0 ;
      RECT  128400.0 693450.0 129600.0 694650.0 ;
      RECT  128400.0 693450.0 129600.0 694650.0 ;
      RECT  126000.0 693450.0 127200.0 694650.0 ;
      RECT  126000.0 684150.0 127200.0 685350.0 ;
      RECT  128400.0 684150.0 129600.0 685350.0 ;
      RECT  128400.0 684150.0 129600.0 685350.0 ;
      RECT  126000.0 684150.0 127200.0 685350.0 ;
      RECT  130800.0 694050.0 132000.0 695250.0 ;
      RECT  130800.0 684150.0 132000.0 685350.0 ;
      RECT  126600.0 688800.0 127800.0 690000.0 ;
      RECT  126600.0 688800.0 127800.0 690000.0 ;
      RECT  129150.0 688950.0 130050.0 689850.0 ;
      RECT  124200.0 696150.0 133800.0 697050.0 ;
      RECT  124200.0 682350.0 133800.0 683250.0 ;
      RECT  135600.0 684750.0 136800.0 682350.0 ;
      RECT  135600.0 693450.0 136800.0 697050.0 ;
      RECT  140400.0 693450.0 141600.0 697050.0 ;
      RECT  142800.0 694650.0 144000.0 696600.0 ;
      RECT  142800.0 682800.0 144000.0 684750.0 ;
      RECT  135600.0 693450.0 136800.0 694650.0 ;
      RECT  138000.0 693450.0 139200.0 694650.0 ;
      RECT  138000.0 693450.0 139200.0 694650.0 ;
      RECT  135600.0 693450.0 136800.0 694650.0 ;
      RECT  138000.0 693450.0 139200.0 694650.0 ;
      RECT  140400.0 693450.0 141600.0 694650.0 ;
      RECT  140400.0 693450.0 141600.0 694650.0 ;
      RECT  138000.0 693450.0 139200.0 694650.0 ;
      RECT  135600.0 684750.0 136800.0 685950.0 ;
      RECT  138000.0 684750.0 139200.0 685950.0 ;
      RECT  138000.0 684750.0 139200.0 685950.0 ;
      RECT  135600.0 684750.0 136800.0 685950.0 ;
      RECT  138000.0 684750.0 139200.0 685950.0 ;
      RECT  140400.0 684750.0 141600.0 685950.0 ;
      RECT  140400.0 684750.0 141600.0 685950.0 ;
      RECT  138000.0 684750.0 139200.0 685950.0 ;
      RECT  142800.0 694050.0 144000.0 695250.0 ;
      RECT  142800.0 684150.0 144000.0 685350.0 ;
      RECT  140400.0 687300.0 139200.0 688500.0 ;
      RECT  137400.0 690000.0 136200.0 691200.0 ;
      RECT  138000.0 693450.0 139200.0 694650.0 ;
      RECT  140400.0 684750.0 141600.0 685950.0 ;
      RECT  141600.0 690000.0 140400.0 691200.0 ;
      RECT  136200.0 690000.0 137400.0 691200.0 ;
      RECT  139200.0 687300.0 140400.0 688500.0 ;
      RECT  140400.0 690000.0 141600.0 691200.0 ;
      RECT  133800.0 696150.0 148200.0 697050.0 ;
      RECT  133800.0 682350.0 148200.0 683250.0 ;
      RECT  154800.0 694650.0 156000.0 696600.0 ;
      RECT  154800.0 682800.0 156000.0 684750.0 ;
      RECT  150000.0 684150.0 151200.0 682350.0 ;
      RECT  150000.0 693450.0 151200.0 697050.0 ;
      RECT  152700.0 684150.0 153600.0 693450.0 ;
      RECT  150000.0 693450.0 151200.0 694650.0 ;
      RECT  152400.0 693450.0 153600.0 694650.0 ;
      RECT  152400.0 693450.0 153600.0 694650.0 ;
      RECT  150000.0 693450.0 151200.0 694650.0 ;
      RECT  150000.0 684150.0 151200.0 685350.0 ;
      RECT  152400.0 684150.0 153600.0 685350.0 ;
      RECT  152400.0 684150.0 153600.0 685350.0 ;
      RECT  150000.0 684150.0 151200.0 685350.0 ;
      RECT  154800.0 694050.0 156000.0 695250.0 ;
      RECT  154800.0 684150.0 156000.0 685350.0 ;
      RECT  150600.0 688800.0 151800.0 690000.0 ;
      RECT  150600.0 688800.0 151800.0 690000.0 ;
      RECT  153150.0 688950.0 154050.0 689850.0 ;
      RECT  148200.0 696150.0 157800.0 697050.0 ;
      RECT  148200.0 682350.0 157800.0 683250.0 ;
      RECT  120450.0 688800.0 121650.0 690000.0 ;
      RECT  122400.0 686400.0 123600.0 687600.0 ;
      RECT  139200.0 687300.0 138000.0 688500.0 ;
      RECT  130800.0 698550.0 132000.0 696600.0 ;
      RECT  130800.0 710400.0 132000.0 708450.0 ;
      RECT  126000.0 709050.0 127200.0 710850.0 ;
      RECT  126000.0 699750.0 127200.0 696150.0 ;
      RECT  128700.0 709050.0 129600.0 699750.0 ;
      RECT  126000.0 699750.0 127200.0 698550.0 ;
      RECT  128400.0 699750.0 129600.0 698550.0 ;
      RECT  128400.0 699750.0 129600.0 698550.0 ;
      RECT  126000.0 699750.0 127200.0 698550.0 ;
      RECT  126000.0 709050.0 127200.0 707850.0 ;
      RECT  128400.0 709050.0 129600.0 707850.0 ;
      RECT  128400.0 709050.0 129600.0 707850.0 ;
      RECT  126000.0 709050.0 127200.0 707850.0 ;
      RECT  130800.0 699150.0 132000.0 697950.0 ;
      RECT  130800.0 709050.0 132000.0 707850.0 ;
      RECT  126600.0 704400.0 127800.0 703200.0 ;
      RECT  126600.0 704400.0 127800.0 703200.0 ;
      RECT  129150.0 704250.0 130050.0 703350.0 ;
      RECT  124200.0 697050.0 133800.0 696150.0 ;
      RECT  124200.0 710850.0 133800.0 709950.0 ;
      RECT  135600.0 708450.0 136800.0 710850.0 ;
      RECT  135600.0 699750.0 136800.0 696150.0 ;
      RECT  140400.0 699750.0 141600.0 696150.0 ;
      RECT  142800.0 698550.0 144000.0 696600.0 ;
      RECT  142800.0 710400.0 144000.0 708450.0 ;
      RECT  135600.0 699750.0 136800.0 698550.0 ;
      RECT  138000.0 699750.0 139200.0 698550.0 ;
      RECT  138000.0 699750.0 139200.0 698550.0 ;
      RECT  135600.0 699750.0 136800.0 698550.0 ;
      RECT  138000.0 699750.0 139200.0 698550.0 ;
      RECT  140400.0 699750.0 141600.0 698550.0 ;
      RECT  140400.0 699750.0 141600.0 698550.0 ;
      RECT  138000.0 699750.0 139200.0 698550.0 ;
      RECT  135600.0 708450.0 136800.0 707250.0 ;
      RECT  138000.0 708450.0 139200.0 707250.0 ;
      RECT  138000.0 708450.0 139200.0 707250.0 ;
      RECT  135600.0 708450.0 136800.0 707250.0 ;
      RECT  138000.0 708450.0 139200.0 707250.0 ;
      RECT  140400.0 708450.0 141600.0 707250.0 ;
      RECT  140400.0 708450.0 141600.0 707250.0 ;
      RECT  138000.0 708450.0 139200.0 707250.0 ;
      RECT  142800.0 699150.0 144000.0 697950.0 ;
      RECT  142800.0 709050.0 144000.0 707850.0 ;
      RECT  140400.0 705900.0 139200.0 704700.0 ;
      RECT  137400.0 703200.0 136200.0 702000.0 ;
      RECT  138000.0 699750.0 139200.0 698550.0 ;
      RECT  140400.0 708450.0 141600.0 707250.0 ;
      RECT  141600.0 703200.0 140400.0 702000.0 ;
      RECT  136200.0 703200.0 137400.0 702000.0 ;
      RECT  139200.0 705900.0 140400.0 704700.0 ;
      RECT  140400.0 703200.0 141600.0 702000.0 ;
      RECT  133800.0 697050.0 148200.0 696150.0 ;
      RECT  133800.0 710850.0 148200.0 709950.0 ;
      RECT  154800.0 698550.0 156000.0 696600.0 ;
      RECT  154800.0 710400.0 156000.0 708450.0 ;
      RECT  150000.0 709050.0 151200.0 710850.0 ;
      RECT  150000.0 699750.0 151200.0 696150.0 ;
      RECT  152700.0 709050.0 153600.0 699750.0 ;
      RECT  150000.0 699750.0 151200.0 698550.0 ;
      RECT  152400.0 699750.0 153600.0 698550.0 ;
      RECT  152400.0 699750.0 153600.0 698550.0 ;
      RECT  150000.0 699750.0 151200.0 698550.0 ;
      RECT  150000.0 709050.0 151200.0 707850.0 ;
      RECT  152400.0 709050.0 153600.0 707850.0 ;
      RECT  152400.0 709050.0 153600.0 707850.0 ;
      RECT  150000.0 709050.0 151200.0 707850.0 ;
      RECT  154800.0 699150.0 156000.0 697950.0 ;
      RECT  154800.0 709050.0 156000.0 707850.0 ;
      RECT  150600.0 704400.0 151800.0 703200.0 ;
      RECT  150600.0 704400.0 151800.0 703200.0 ;
      RECT  153150.0 704250.0 154050.0 703350.0 ;
      RECT  148200.0 697050.0 157800.0 696150.0 ;
      RECT  148200.0 710850.0 157800.0 709950.0 ;
      RECT  120450.0 703200.0 121650.0 704400.0 ;
      RECT  122400.0 705600.0 123600.0 706800.0 ;
      RECT  139200.0 704700.0 138000.0 705900.0 ;
      RECT  130800.0 722250.0 132000.0 724200.0 ;
      RECT  130800.0 710400.0 132000.0 712350.0 ;
      RECT  126000.0 711750.0 127200.0 709950.0 ;
      RECT  126000.0 721050.0 127200.0 724650.0 ;
      RECT  128700.0 711750.0 129600.0 721050.0 ;
      RECT  126000.0 721050.0 127200.0 722250.0 ;
      RECT  128400.0 721050.0 129600.0 722250.0 ;
      RECT  128400.0 721050.0 129600.0 722250.0 ;
      RECT  126000.0 721050.0 127200.0 722250.0 ;
      RECT  126000.0 711750.0 127200.0 712950.0 ;
      RECT  128400.0 711750.0 129600.0 712950.0 ;
      RECT  128400.0 711750.0 129600.0 712950.0 ;
      RECT  126000.0 711750.0 127200.0 712950.0 ;
      RECT  130800.0 721650.0 132000.0 722850.0 ;
      RECT  130800.0 711750.0 132000.0 712950.0 ;
      RECT  126600.0 716400.0 127800.0 717600.0 ;
      RECT  126600.0 716400.0 127800.0 717600.0 ;
      RECT  129150.0 716550.0 130050.0 717450.0 ;
      RECT  124200.0 723750.0 133800.0 724650.0 ;
      RECT  124200.0 709950.0 133800.0 710850.0 ;
      RECT  135600.0 712350.0 136800.0 709950.0 ;
      RECT  135600.0 721050.0 136800.0 724650.0 ;
      RECT  140400.0 721050.0 141600.0 724650.0 ;
      RECT  142800.0 722250.0 144000.0 724200.0 ;
      RECT  142800.0 710400.0 144000.0 712350.0 ;
      RECT  135600.0 721050.0 136800.0 722250.0 ;
      RECT  138000.0 721050.0 139200.0 722250.0 ;
      RECT  138000.0 721050.0 139200.0 722250.0 ;
      RECT  135600.0 721050.0 136800.0 722250.0 ;
      RECT  138000.0 721050.0 139200.0 722250.0 ;
      RECT  140400.0 721050.0 141600.0 722250.0 ;
      RECT  140400.0 721050.0 141600.0 722250.0 ;
      RECT  138000.0 721050.0 139200.0 722250.0 ;
      RECT  135600.0 712350.0 136800.0 713550.0 ;
      RECT  138000.0 712350.0 139200.0 713550.0 ;
      RECT  138000.0 712350.0 139200.0 713550.0 ;
      RECT  135600.0 712350.0 136800.0 713550.0 ;
      RECT  138000.0 712350.0 139200.0 713550.0 ;
      RECT  140400.0 712350.0 141600.0 713550.0 ;
      RECT  140400.0 712350.0 141600.0 713550.0 ;
      RECT  138000.0 712350.0 139200.0 713550.0 ;
      RECT  142800.0 721650.0 144000.0 722850.0 ;
      RECT  142800.0 711750.0 144000.0 712950.0 ;
      RECT  140400.0 714900.0 139200.0 716100.0 ;
      RECT  137400.0 717600.0 136200.0 718800.0 ;
      RECT  138000.0 721050.0 139200.0 722250.0 ;
      RECT  140400.0 712350.0 141600.0 713550.0 ;
      RECT  141600.0 717600.0 140400.0 718800.0 ;
      RECT  136200.0 717600.0 137400.0 718800.0 ;
      RECT  139200.0 714900.0 140400.0 716100.0 ;
      RECT  140400.0 717600.0 141600.0 718800.0 ;
      RECT  133800.0 723750.0 148200.0 724650.0 ;
      RECT  133800.0 709950.0 148200.0 710850.0 ;
      RECT  154800.0 722250.0 156000.0 724200.0 ;
      RECT  154800.0 710400.0 156000.0 712350.0 ;
      RECT  150000.0 711750.0 151200.0 709950.0 ;
      RECT  150000.0 721050.0 151200.0 724650.0 ;
      RECT  152700.0 711750.0 153600.0 721050.0 ;
      RECT  150000.0 721050.0 151200.0 722250.0 ;
      RECT  152400.0 721050.0 153600.0 722250.0 ;
      RECT  152400.0 721050.0 153600.0 722250.0 ;
      RECT  150000.0 721050.0 151200.0 722250.0 ;
      RECT  150000.0 711750.0 151200.0 712950.0 ;
      RECT  152400.0 711750.0 153600.0 712950.0 ;
      RECT  152400.0 711750.0 153600.0 712950.0 ;
      RECT  150000.0 711750.0 151200.0 712950.0 ;
      RECT  154800.0 721650.0 156000.0 722850.0 ;
      RECT  154800.0 711750.0 156000.0 712950.0 ;
      RECT  150600.0 716400.0 151800.0 717600.0 ;
      RECT  150600.0 716400.0 151800.0 717600.0 ;
      RECT  153150.0 716550.0 154050.0 717450.0 ;
      RECT  148200.0 723750.0 157800.0 724650.0 ;
      RECT  148200.0 709950.0 157800.0 710850.0 ;
      RECT  120450.0 716400.0 121650.0 717600.0 ;
      RECT  122400.0 714000.0 123600.0 715200.0 ;
      RECT  139200.0 714900.0 138000.0 716100.0 ;
      RECT  130800.0 726150.0 132000.0 724200.0 ;
      RECT  130800.0 738000.0 132000.0 736050.0 ;
      RECT  126000.0 736650.0 127200.0 738450.0 ;
      RECT  126000.0 727350.0 127200.0 723750.0 ;
      RECT  128700.0 736650.0 129600.0 727350.0 ;
      RECT  126000.0 727350.0 127200.0 726150.0 ;
      RECT  128400.0 727350.0 129600.0 726150.0 ;
      RECT  128400.0 727350.0 129600.0 726150.0 ;
      RECT  126000.0 727350.0 127200.0 726150.0 ;
      RECT  126000.0 736650.0 127200.0 735450.0 ;
      RECT  128400.0 736650.0 129600.0 735450.0 ;
      RECT  128400.0 736650.0 129600.0 735450.0 ;
      RECT  126000.0 736650.0 127200.0 735450.0 ;
      RECT  130800.0 726750.0 132000.0 725550.0 ;
      RECT  130800.0 736650.0 132000.0 735450.0 ;
      RECT  126600.0 732000.0 127800.0 730800.0 ;
      RECT  126600.0 732000.0 127800.0 730800.0 ;
      RECT  129150.0 731850.0 130050.0 730950.0 ;
      RECT  124200.0 724650.0 133800.0 723750.0 ;
      RECT  124200.0 738450.0 133800.0 737550.0 ;
      RECT  135600.0 736050.0 136800.0 738450.0 ;
      RECT  135600.0 727350.0 136800.0 723750.0 ;
      RECT  140400.0 727350.0 141600.0 723750.0 ;
      RECT  142800.0 726150.0 144000.0 724200.0 ;
      RECT  142800.0 738000.0 144000.0 736050.0 ;
      RECT  135600.0 727350.0 136800.0 726150.0 ;
      RECT  138000.0 727350.0 139200.0 726150.0 ;
      RECT  138000.0 727350.0 139200.0 726150.0 ;
      RECT  135600.0 727350.0 136800.0 726150.0 ;
      RECT  138000.0 727350.0 139200.0 726150.0 ;
      RECT  140400.0 727350.0 141600.0 726150.0 ;
      RECT  140400.0 727350.0 141600.0 726150.0 ;
      RECT  138000.0 727350.0 139200.0 726150.0 ;
      RECT  135600.0 736050.0 136800.0 734850.0 ;
      RECT  138000.0 736050.0 139200.0 734850.0 ;
      RECT  138000.0 736050.0 139200.0 734850.0 ;
      RECT  135600.0 736050.0 136800.0 734850.0 ;
      RECT  138000.0 736050.0 139200.0 734850.0 ;
      RECT  140400.0 736050.0 141600.0 734850.0 ;
      RECT  140400.0 736050.0 141600.0 734850.0 ;
      RECT  138000.0 736050.0 139200.0 734850.0 ;
      RECT  142800.0 726750.0 144000.0 725550.0 ;
      RECT  142800.0 736650.0 144000.0 735450.0 ;
      RECT  140400.0 733500.0 139200.0 732300.0 ;
      RECT  137400.0 730800.0 136200.0 729600.0 ;
      RECT  138000.0 727350.0 139200.0 726150.0 ;
      RECT  140400.0 736050.0 141600.0 734850.0 ;
      RECT  141600.0 730800.0 140400.0 729600.0 ;
      RECT  136200.0 730800.0 137400.0 729600.0 ;
      RECT  139200.0 733500.0 140400.0 732300.0 ;
      RECT  140400.0 730800.0 141600.0 729600.0 ;
      RECT  133800.0 724650.0 148200.0 723750.0 ;
      RECT  133800.0 738450.0 148200.0 737550.0 ;
      RECT  154800.0 726150.0 156000.0 724200.0 ;
      RECT  154800.0 738000.0 156000.0 736050.0 ;
      RECT  150000.0 736650.0 151200.0 738450.0 ;
      RECT  150000.0 727350.0 151200.0 723750.0 ;
      RECT  152700.0 736650.0 153600.0 727350.0 ;
      RECT  150000.0 727350.0 151200.0 726150.0 ;
      RECT  152400.0 727350.0 153600.0 726150.0 ;
      RECT  152400.0 727350.0 153600.0 726150.0 ;
      RECT  150000.0 727350.0 151200.0 726150.0 ;
      RECT  150000.0 736650.0 151200.0 735450.0 ;
      RECT  152400.0 736650.0 153600.0 735450.0 ;
      RECT  152400.0 736650.0 153600.0 735450.0 ;
      RECT  150000.0 736650.0 151200.0 735450.0 ;
      RECT  154800.0 726750.0 156000.0 725550.0 ;
      RECT  154800.0 736650.0 156000.0 735450.0 ;
      RECT  150600.0 732000.0 151800.0 730800.0 ;
      RECT  150600.0 732000.0 151800.0 730800.0 ;
      RECT  153150.0 731850.0 154050.0 730950.0 ;
      RECT  148200.0 724650.0 157800.0 723750.0 ;
      RECT  148200.0 738450.0 157800.0 737550.0 ;
      RECT  120450.0 730800.0 121650.0 732000.0 ;
      RECT  122400.0 733200.0 123600.0 734400.0 ;
      RECT  139200.0 732300.0 138000.0 733500.0 ;
      RECT  130800.0 749850.0 132000.0 751800.0 ;
      RECT  130800.0 738000.0 132000.0 739950.0 ;
      RECT  126000.0 739350.0 127200.0 737550.0 ;
      RECT  126000.0 748650.0 127200.0 752250.0 ;
      RECT  128700.0 739350.0 129600.0 748650.0 ;
      RECT  126000.0 748650.0 127200.0 749850.0 ;
      RECT  128400.0 748650.0 129600.0 749850.0 ;
      RECT  128400.0 748650.0 129600.0 749850.0 ;
      RECT  126000.0 748650.0 127200.0 749850.0 ;
      RECT  126000.0 739350.0 127200.0 740550.0 ;
      RECT  128400.0 739350.0 129600.0 740550.0 ;
      RECT  128400.0 739350.0 129600.0 740550.0 ;
      RECT  126000.0 739350.0 127200.0 740550.0 ;
      RECT  130800.0 749250.0 132000.0 750450.0 ;
      RECT  130800.0 739350.0 132000.0 740550.0 ;
      RECT  126600.0 744000.0 127800.0 745200.0 ;
      RECT  126600.0 744000.0 127800.0 745200.0 ;
      RECT  129150.0 744150.0 130050.0 745050.0 ;
      RECT  124200.0 751350.0 133800.0 752250.0 ;
      RECT  124200.0 737550.0 133800.0 738450.0 ;
      RECT  135600.0 739950.0 136800.0 737550.0 ;
      RECT  135600.0 748650.0 136800.0 752250.0 ;
      RECT  140400.0 748650.0 141600.0 752250.0 ;
      RECT  142800.0 749850.0 144000.0 751800.0 ;
      RECT  142800.0 738000.0 144000.0 739950.0 ;
      RECT  135600.0 748650.0 136800.0 749850.0 ;
      RECT  138000.0 748650.0 139200.0 749850.0 ;
      RECT  138000.0 748650.0 139200.0 749850.0 ;
      RECT  135600.0 748650.0 136800.0 749850.0 ;
      RECT  138000.0 748650.0 139200.0 749850.0 ;
      RECT  140400.0 748650.0 141600.0 749850.0 ;
      RECT  140400.0 748650.0 141600.0 749850.0 ;
      RECT  138000.0 748650.0 139200.0 749850.0 ;
      RECT  135600.0 739950.0 136800.0 741150.0 ;
      RECT  138000.0 739950.0 139200.0 741150.0 ;
      RECT  138000.0 739950.0 139200.0 741150.0 ;
      RECT  135600.0 739950.0 136800.0 741150.0 ;
      RECT  138000.0 739950.0 139200.0 741150.0 ;
      RECT  140400.0 739950.0 141600.0 741150.0 ;
      RECT  140400.0 739950.0 141600.0 741150.0 ;
      RECT  138000.0 739950.0 139200.0 741150.0 ;
      RECT  142800.0 749250.0 144000.0 750450.0 ;
      RECT  142800.0 739350.0 144000.0 740550.0 ;
      RECT  140400.0 742500.0 139200.0 743700.0 ;
      RECT  137400.0 745200.0 136200.0 746400.0 ;
      RECT  138000.0 748650.0 139200.0 749850.0 ;
      RECT  140400.0 739950.0 141600.0 741150.0 ;
      RECT  141600.0 745200.0 140400.0 746400.0 ;
      RECT  136200.0 745200.0 137400.0 746400.0 ;
      RECT  139200.0 742500.0 140400.0 743700.0 ;
      RECT  140400.0 745200.0 141600.0 746400.0 ;
      RECT  133800.0 751350.0 148200.0 752250.0 ;
      RECT  133800.0 737550.0 148200.0 738450.0 ;
      RECT  154800.0 749850.0 156000.0 751800.0 ;
      RECT  154800.0 738000.0 156000.0 739950.0 ;
      RECT  150000.0 739350.0 151200.0 737550.0 ;
      RECT  150000.0 748650.0 151200.0 752250.0 ;
      RECT  152700.0 739350.0 153600.0 748650.0 ;
      RECT  150000.0 748650.0 151200.0 749850.0 ;
      RECT  152400.0 748650.0 153600.0 749850.0 ;
      RECT  152400.0 748650.0 153600.0 749850.0 ;
      RECT  150000.0 748650.0 151200.0 749850.0 ;
      RECT  150000.0 739350.0 151200.0 740550.0 ;
      RECT  152400.0 739350.0 153600.0 740550.0 ;
      RECT  152400.0 739350.0 153600.0 740550.0 ;
      RECT  150000.0 739350.0 151200.0 740550.0 ;
      RECT  154800.0 749250.0 156000.0 750450.0 ;
      RECT  154800.0 739350.0 156000.0 740550.0 ;
      RECT  150600.0 744000.0 151800.0 745200.0 ;
      RECT  150600.0 744000.0 151800.0 745200.0 ;
      RECT  153150.0 744150.0 154050.0 745050.0 ;
      RECT  148200.0 751350.0 157800.0 752250.0 ;
      RECT  148200.0 737550.0 157800.0 738450.0 ;
      RECT  120450.0 744000.0 121650.0 745200.0 ;
      RECT  122400.0 741600.0 123600.0 742800.0 ;
      RECT  139200.0 742500.0 138000.0 743700.0 ;
      RECT  130800.0 753750.0 132000.0 751800.0 ;
      RECT  130800.0 765600.0 132000.0 763650.0 ;
      RECT  126000.0 764250.0 127200.0 766050.0 ;
      RECT  126000.0 754950.0 127200.0 751350.0 ;
      RECT  128700.0 764250.0 129600.0 754950.0 ;
      RECT  126000.0 754950.0 127200.0 753750.0 ;
      RECT  128400.0 754950.0 129600.0 753750.0 ;
      RECT  128400.0 754950.0 129600.0 753750.0 ;
      RECT  126000.0 754950.0 127200.0 753750.0 ;
      RECT  126000.0 764250.0 127200.0 763050.0 ;
      RECT  128400.0 764250.0 129600.0 763050.0 ;
      RECT  128400.0 764250.0 129600.0 763050.0 ;
      RECT  126000.0 764250.0 127200.0 763050.0 ;
      RECT  130800.0 754350.0 132000.0 753150.0 ;
      RECT  130800.0 764250.0 132000.0 763050.0 ;
      RECT  126600.0 759600.0 127800.0 758400.0 ;
      RECT  126600.0 759600.0 127800.0 758400.0 ;
      RECT  129150.0 759450.0 130050.0 758550.0 ;
      RECT  124200.0 752250.0 133800.0 751350.0 ;
      RECT  124200.0 766050.0 133800.0 765150.0 ;
      RECT  135600.0 763650.0 136800.0 766050.0 ;
      RECT  135600.0 754950.0 136800.0 751350.0 ;
      RECT  140400.0 754950.0 141600.0 751350.0 ;
      RECT  142800.0 753750.0 144000.0 751800.0 ;
      RECT  142800.0 765600.0 144000.0 763650.0 ;
      RECT  135600.0 754950.0 136800.0 753750.0 ;
      RECT  138000.0 754950.0 139200.0 753750.0 ;
      RECT  138000.0 754950.0 139200.0 753750.0 ;
      RECT  135600.0 754950.0 136800.0 753750.0 ;
      RECT  138000.0 754950.0 139200.0 753750.0 ;
      RECT  140400.0 754950.0 141600.0 753750.0 ;
      RECT  140400.0 754950.0 141600.0 753750.0 ;
      RECT  138000.0 754950.0 139200.0 753750.0 ;
      RECT  135600.0 763650.0 136800.0 762450.0 ;
      RECT  138000.0 763650.0 139200.0 762450.0 ;
      RECT  138000.0 763650.0 139200.0 762450.0 ;
      RECT  135600.0 763650.0 136800.0 762450.0 ;
      RECT  138000.0 763650.0 139200.0 762450.0 ;
      RECT  140400.0 763650.0 141600.0 762450.0 ;
      RECT  140400.0 763650.0 141600.0 762450.0 ;
      RECT  138000.0 763650.0 139200.0 762450.0 ;
      RECT  142800.0 754350.0 144000.0 753150.0 ;
      RECT  142800.0 764250.0 144000.0 763050.0 ;
      RECT  140400.0 761100.0 139200.0 759900.0 ;
      RECT  137400.0 758400.0 136200.0 757200.0 ;
      RECT  138000.0 754950.0 139200.0 753750.0 ;
      RECT  140400.0 763650.0 141600.0 762450.0 ;
      RECT  141600.0 758400.0 140400.0 757200.0 ;
      RECT  136200.0 758400.0 137400.0 757200.0 ;
      RECT  139200.0 761100.0 140400.0 759900.0 ;
      RECT  140400.0 758400.0 141600.0 757200.0 ;
      RECT  133800.0 752250.0 148200.0 751350.0 ;
      RECT  133800.0 766050.0 148200.0 765150.0 ;
      RECT  154800.0 753750.0 156000.0 751800.0 ;
      RECT  154800.0 765600.0 156000.0 763650.0 ;
      RECT  150000.0 764250.0 151200.0 766050.0 ;
      RECT  150000.0 754950.0 151200.0 751350.0 ;
      RECT  152700.0 764250.0 153600.0 754950.0 ;
      RECT  150000.0 754950.0 151200.0 753750.0 ;
      RECT  152400.0 754950.0 153600.0 753750.0 ;
      RECT  152400.0 754950.0 153600.0 753750.0 ;
      RECT  150000.0 754950.0 151200.0 753750.0 ;
      RECT  150000.0 764250.0 151200.0 763050.0 ;
      RECT  152400.0 764250.0 153600.0 763050.0 ;
      RECT  152400.0 764250.0 153600.0 763050.0 ;
      RECT  150000.0 764250.0 151200.0 763050.0 ;
      RECT  154800.0 754350.0 156000.0 753150.0 ;
      RECT  154800.0 764250.0 156000.0 763050.0 ;
      RECT  150600.0 759600.0 151800.0 758400.0 ;
      RECT  150600.0 759600.0 151800.0 758400.0 ;
      RECT  153150.0 759450.0 154050.0 758550.0 ;
      RECT  148200.0 752250.0 157800.0 751350.0 ;
      RECT  148200.0 766050.0 157800.0 765150.0 ;
      RECT  120450.0 758400.0 121650.0 759600.0 ;
      RECT  122400.0 760800.0 123600.0 762000.0 ;
      RECT  139200.0 759900.0 138000.0 761100.0 ;
      RECT  130800.0 777450.0 132000.0 779400.0 ;
      RECT  130800.0 765600.0 132000.0 767550.0 ;
      RECT  126000.0 766950.0 127200.0 765150.0 ;
      RECT  126000.0 776250.0 127200.0 779850.0 ;
      RECT  128700.0 766950.0 129600.0 776250.0 ;
      RECT  126000.0 776250.0 127200.0 777450.0 ;
      RECT  128400.0 776250.0 129600.0 777450.0 ;
      RECT  128400.0 776250.0 129600.0 777450.0 ;
      RECT  126000.0 776250.0 127200.0 777450.0 ;
      RECT  126000.0 766950.0 127200.0 768150.0 ;
      RECT  128400.0 766950.0 129600.0 768150.0 ;
      RECT  128400.0 766950.0 129600.0 768150.0 ;
      RECT  126000.0 766950.0 127200.0 768150.0 ;
      RECT  130800.0 776850.0 132000.0 778050.0 ;
      RECT  130800.0 766950.0 132000.0 768150.0 ;
      RECT  126600.0 771600.0 127800.0 772800.0 ;
      RECT  126600.0 771600.0 127800.0 772800.0 ;
      RECT  129150.0 771750.0 130050.0 772650.0 ;
      RECT  124200.0 778950.0 133800.0 779850.0 ;
      RECT  124200.0 765150.0 133800.0 766050.0 ;
      RECT  135600.0 767550.0 136800.0 765150.0 ;
      RECT  135600.0 776250.0 136800.0 779850.0 ;
      RECT  140400.0 776250.0 141600.0 779850.0 ;
      RECT  142800.0 777450.0 144000.0 779400.0 ;
      RECT  142800.0 765600.0 144000.0 767550.0 ;
      RECT  135600.0 776250.0 136800.0 777450.0 ;
      RECT  138000.0 776250.0 139200.0 777450.0 ;
      RECT  138000.0 776250.0 139200.0 777450.0 ;
      RECT  135600.0 776250.0 136800.0 777450.0 ;
      RECT  138000.0 776250.0 139200.0 777450.0 ;
      RECT  140400.0 776250.0 141600.0 777450.0 ;
      RECT  140400.0 776250.0 141600.0 777450.0 ;
      RECT  138000.0 776250.0 139200.0 777450.0 ;
      RECT  135600.0 767550.0 136800.0 768750.0 ;
      RECT  138000.0 767550.0 139200.0 768750.0 ;
      RECT  138000.0 767550.0 139200.0 768750.0 ;
      RECT  135600.0 767550.0 136800.0 768750.0 ;
      RECT  138000.0 767550.0 139200.0 768750.0 ;
      RECT  140400.0 767550.0 141600.0 768750.0 ;
      RECT  140400.0 767550.0 141600.0 768750.0 ;
      RECT  138000.0 767550.0 139200.0 768750.0 ;
      RECT  142800.0 776850.0 144000.0 778050.0 ;
      RECT  142800.0 766950.0 144000.0 768150.0 ;
      RECT  140400.0 770100.0 139200.0 771300.0 ;
      RECT  137400.0 772800.0 136200.0 774000.0 ;
      RECT  138000.0 776250.0 139200.0 777450.0 ;
      RECT  140400.0 767550.0 141600.0 768750.0 ;
      RECT  141600.0 772800.0 140400.0 774000.0 ;
      RECT  136200.0 772800.0 137400.0 774000.0 ;
      RECT  139200.0 770100.0 140400.0 771300.0 ;
      RECT  140400.0 772800.0 141600.0 774000.0 ;
      RECT  133800.0 778950.0 148200.0 779850.0 ;
      RECT  133800.0 765150.0 148200.0 766050.0 ;
      RECT  154800.0 777450.0 156000.0 779400.0 ;
      RECT  154800.0 765600.0 156000.0 767550.0 ;
      RECT  150000.0 766950.0 151200.0 765150.0 ;
      RECT  150000.0 776250.0 151200.0 779850.0 ;
      RECT  152700.0 766950.0 153600.0 776250.0 ;
      RECT  150000.0 776250.0 151200.0 777450.0 ;
      RECT  152400.0 776250.0 153600.0 777450.0 ;
      RECT  152400.0 776250.0 153600.0 777450.0 ;
      RECT  150000.0 776250.0 151200.0 777450.0 ;
      RECT  150000.0 766950.0 151200.0 768150.0 ;
      RECT  152400.0 766950.0 153600.0 768150.0 ;
      RECT  152400.0 766950.0 153600.0 768150.0 ;
      RECT  150000.0 766950.0 151200.0 768150.0 ;
      RECT  154800.0 776850.0 156000.0 778050.0 ;
      RECT  154800.0 766950.0 156000.0 768150.0 ;
      RECT  150600.0 771600.0 151800.0 772800.0 ;
      RECT  150600.0 771600.0 151800.0 772800.0 ;
      RECT  153150.0 771750.0 154050.0 772650.0 ;
      RECT  148200.0 778950.0 157800.0 779850.0 ;
      RECT  148200.0 765150.0 157800.0 766050.0 ;
      RECT  120450.0 771600.0 121650.0 772800.0 ;
      RECT  122400.0 769200.0 123600.0 770400.0 ;
      RECT  139200.0 770100.0 138000.0 771300.0 ;
      RECT  130800.0 781350.0 132000.0 779400.0 ;
      RECT  130800.0 793200.0 132000.0 791250.0 ;
      RECT  126000.0 791850.0 127200.0 793650.0 ;
      RECT  126000.0 782550.0 127200.0 778950.0 ;
      RECT  128700.0 791850.0 129600.0 782550.0 ;
      RECT  126000.0 782550.0 127200.0 781350.0 ;
      RECT  128400.0 782550.0 129600.0 781350.0 ;
      RECT  128400.0 782550.0 129600.0 781350.0 ;
      RECT  126000.0 782550.0 127200.0 781350.0 ;
      RECT  126000.0 791850.0 127200.0 790650.0 ;
      RECT  128400.0 791850.0 129600.0 790650.0 ;
      RECT  128400.0 791850.0 129600.0 790650.0 ;
      RECT  126000.0 791850.0 127200.0 790650.0 ;
      RECT  130800.0 781950.0 132000.0 780750.0 ;
      RECT  130800.0 791850.0 132000.0 790650.0 ;
      RECT  126600.0 787200.0 127800.0 786000.0 ;
      RECT  126600.0 787200.0 127800.0 786000.0 ;
      RECT  129150.0 787050.0 130050.0 786150.0 ;
      RECT  124200.0 779850.0 133800.0 778950.0 ;
      RECT  124200.0 793650.0 133800.0 792750.0 ;
      RECT  135600.0 791250.0 136800.0 793650.0 ;
      RECT  135600.0 782550.0 136800.0 778950.0 ;
      RECT  140400.0 782550.0 141600.0 778950.0 ;
      RECT  142800.0 781350.0 144000.0 779400.0 ;
      RECT  142800.0 793200.0 144000.0 791250.0 ;
      RECT  135600.0 782550.0 136800.0 781350.0 ;
      RECT  138000.0 782550.0 139200.0 781350.0 ;
      RECT  138000.0 782550.0 139200.0 781350.0 ;
      RECT  135600.0 782550.0 136800.0 781350.0 ;
      RECT  138000.0 782550.0 139200.0 781350.0 ;
      RECT  140400.0 782550.0 141600.0 781350.0 ;
      RECT  140400.0 782550.0 141600.0 781350.0 ;
      RECT  138000.0 782550.0 139200.0 781350.0 ;
      RECT  135600.0 791250.0 136800.0 790050.0 ;
      RECT  138000.0 791250.0 139200.0 790050.0 ;
      RECT  138000.0 791250.0 139200.0 790050.0 ;
      RECT  135600.0 791250.0 136800.0 790050.0 ;
      RECT  138000.0 791250.0 139200.0 790050.0 ;
      RECT  140400.0 791250.0 141600.0 790050.0 ;
      RECT  140400.0 791250.0 141600.0 790050.0 ;
      RECT  138000.0 791250.0 139200.0 790050.0 ;
      RECT  142800.0 781950.0 144000.0 780750.0 ;
      RECT  142800.0 791850.0 144000.0 790650.0 ;
      RECT  140400.0 788700.0 139200.0 787500.0 ;
      RECT  137400.0 786000.0 136200.0 784800.0 ;
      RECT  138000.0 782550.0 139200.0 781350.0 ;
      RECT  140400.0 791250.0 141600.0 790050.0 ;
      RECT  141600.0 786000.0 140400.0 784800.0 ;
      RECT  136200.0 786000.0 137400.0 784800.0 ;
      RECT  139200.0 788700.0 140400.0 787500.0 ;
      RECT  140400.0 786000.0 141600.0 784800.0 ;
      RECT  133800.0 779850.0 148200.0 778950.0 ;
      RECT  133800.0 793650.0 148200.0 792750.0 ;
      RECT  154800.0 781350.0 156000.0 779400.0 ;
      RECT  154800.0 793200.0 156000.0 791250.0 ;
      RECT  150000.0 791850.0 151200.0 793650.0 ;
      RECT  150000.0 782550.0 151200.0 778950.0 ;
      RECT  152700.0 791850.0 153600.0 782550.0 ;
      RECT  150000.0 782550.0 151200.0 781350.0 ;
      RECT  152400.0 782550.0 153600.0 781350.0 ;
      RECT  152400.0 782550.0 153600.0 781350.0 ;
      RECT  150000.0 782550.0 151200.0 781350.0 ;
      RECT  150000.0 791850.0 151200.0 790650.0 ;
      RECT  152400.0 791850.0 153600.0 790650.0 ;
      RECT  152400.0 791850.0 153600.0 790650.0 ;
      RECT  150000.0 791850.0 151200.0 790650.0 ;
      RECT  154800.0 781950.0 156000.0 780750.0 ;
      RECT  154800.0 791850.0 156000.0 790650.0 ;
      RECT  150600.0 787200.0 151800.0 786000.0 ;
      RECT  150600.0 787200.0 151800.0 786000.0 ;
      RECT  153150.0 787050.0 154050.0 786150.0 ;
      RECT  148200.0 779850.0 157800.0 778950.0 ;
      RECT  148200.0 793650.0 157800.0 792750.0 ;
      RECT  120450.0 786000.0 121650.0 787200.0 ;
      RECT  122400.0 788400.0 123600.0 789600.0 ;
      RECT  139200.0 787500.0 138000.0 788700.0 ;
      RECT  130800.0 805050.0 132000.0 807000.0 ;
      RECT  130800.0 793200.0 132000.0 795150.0 ;
      RECT  126000.0 794550.0 127200.0 792750.0 ;
      RECT  126000.0 803850.0 127200.0 807450.0 ;
      RECT  128700.0 794550.0 129600.0 803850.0 ;
      RECT  126000.0 803850.0 127200.0 805050.0 ;
      RECT  128400.0 803850.0 129600.0 805050.0 ;
      RECT  128400.0 803850.0 129600.0 805050.0 ;
      RECT  126000.0 803850.0 127200.0 805050.0 ;
      RECT  126000.0 794550.0 127200.0 795750.0 ;
      RECT  128400.0 794550.0 129600.0 795750.0 ;
      RECT  128400.0 794550.0 129600.0 795750.0 ;
      RECT  126000.0 794550.0 127200.0 795750.0 ;
      RECT  130800.0 804450.0 132000.0 805650.0 ;
      RECT  130800.0 794550.0 132000.0 795750.0 ;
      RECT  126600.0 799200.0 127800.0 800400.0 ;
      RECT  126600.0 799200.0 127800.0 800400.0 ;
      RECT  129150.0 799350.0 130050.0 800250.0 ;
      RECT  124200.0 806550.0 133800.0 807450.0 ;
      RECT  124200.0 792750.0 133800.0 793650.0 ;
      RECT  135600.0 795150.0 136800.0 792750.0 ;
      RECT  135600.0 803850.0 136800.0 807450.0 ;
      RECT  140400.0 803850.0 141600.0 807450.0 ;
      RECT  142800.0 805050.0 144000.0 807000.0 ;
      RECT  142800.0 793200.0 144000.0 795150.0 ;
      RECT  135600.0 803850.0 136800.0 805050.0 ;
      RECT  138000.0 803850.0 139200.0 805050.0 ;
      RECT  138000.0 803850.0 139200.0 805050.0 ;
      RECT  135600.0 803850.0 136800.0 805050.0 ;
      RECT  138000.0 803850.0 139200.0 805050.0 ;
      RECT  140400.0 803850.0 141600.0 805050.0 ;
      RECT  140400.0 803850.0 141600.0 805050.0 ;
      RECT  138000.0 803850.0 139200.0 805050.0 ;
      RECT  135600.0 795150.0 136800.0 796350.0 ;
      RECT  138000.0 795150.0 139200.0 796350.0 ;
      RECT  138000.0 795150.0 139200.0 796350.0 ;
      RECT  135600.0 795150.0 136800.0 796350.0 ;
      RECT  138000.0 795150.0 139200.0 796350.0 ;
      RECT  140400.0 795150.0 141600.0 796350.0 ;
      RECT  140400.0 795150.0 141600.0 796350.0 ;
      RECT  138000.0 795150.0 139200.0 796350.0 ;
      RECT  142800.0 804450.0 144000.0 805650.0 ;
      RECT  142800.0 794550.0 144000.0 795750.0 ;
      RECT  140400.0 797700.0 139200.0 798900.0 ;
      RECT  137400.0 800400.0 136200.0 801600.0 ;
      RECT  138000.0 803850.0 139200.0 805050.0 ;
      RECT  140400.0 795150.0 141600.0 796350.0 ;
      RECT  141600.0 800400.0 140400.0 801600.0 ;
      RECT  136200.0 800400.0 137400.0 801600.0 ;
      RECT  139200.0 797700.0 140400.0 798900.0 ;
      RECT  140400.0 800400.0 141600.0 801600.0 ;
      RECT  133800.0 806550.0 148200.0 807450.0 ;
      RECT  133800.0 792750.0 148200.0 793650.0 ;
      RECT  154800.0 805050.0 156000.0 807000.0 ;
      RECT  154800.0 793200.0 156000.0 795150.0 ;
      RECT  150000.0 794550.0 151200.0 792750.0 ;
      RECT  150000.0 803850.0 151200.0 807450.0 ;
      RECT  152700.0 794550.0 153600.0 803850.0 ;
      RECT  150000.0 803850.0 151200.0 805050.0 ;
      RECT  152400.0 803850.0 153600.0 805050.0 ;
      RECT  152400.0 803850.0 153600.0 805050.0 ;
      RECT  150000.0 803850.0 151200.0 805050.0 ;
      RECT  150000.0 794550.0 151200.0 795750.0 ;
      RECT  152400.0 794550.0 153600.0 795750.0 ;
      RECT  152400.0 794550.0 153600.0 795750.0 ;
      RECT  150000.0 794550.0 151200.0 795750.0 ;
      RECT  154800.0 804450.0 156000.0 805650.0 ;
      RECT  154800.0 794550.0 156000.0 795750.0 ;
      RECT  150600.0 799200.0 151800.0 800400.0 ;
      RECT  150600.0 799200.0 151800.0 800400.0 ;
      RECT  153150.0 799350.0 154050.0 800250.0 ;
      RECT  148200.0 806550.0 157800.0 807450.0 ;
      RECT  148200.0 792750.0 157800.0 793650.0 ;
      RECT  120450.0 799200.0 121650.0 800400.0 ;
      RECT  122400.0 796800.0 123600.0 798000.0 ;
      RECT  139200.0 797700.0 138000.0 798900.0 ;
      RECT  130800.0 808950.0 132000.0 807000.0 ;
      RECT  130800.0 820800.0 132000.0 818850.0 ;
      RECT  126000.0 819450.0 127200.0 821250.0 ;
      RECT  126000.0 810150.0 127200.0 806550.0 ;
      RECT  128700.0 819450.0 129600.0 810150.0 ;
      RECT  126000.0 810150.0 127200.0 808950.0 ;
      RECT  128400.0 810150.0 129600.0 808950.0 ;
      RECT  128400.0 810150.0 129600.0 808950.0 ;
      RECT  126000.0 810150.0 127200.0 808950.0 ;
      RECT  126000.0 819450.0 127200.0 818250.0 ;
      RECT  128400.0 819450.0 129600.0 818250.0 ;
      RECT  128400.0 819450.0 129600.0 818250.0 ;
      RECT  126000.0 819450.0 127200.0 818250.0 ;
      RECT  130800.0 809550.0 132000.0 808350.0 ;
      RECT  130800.0 819450.0 132000.0 818250.0 ;
      RECT  126600.0 814800.0 127800.0 813600.0 ;
      RECT  126600.0 814800.0 127800.0 813600.0 ;
      RECT  129150.0 814650.0 130050.0 813750.0 ;
      RECT  124200.0 807450.0 133800.0 806550.0 ;
      RECT  124200.0 821250.0 133800.0 820350.0 ;
      RECT  135600.0 818850.0 136800.0 821250.0 ;
      RECT  135600.0 810150.0 136800.0 806550.0 ;
      RECT  140400.0 810150.0 141600.0 806550.0 ;
      RECT  142800.0 808950.0 144000.0 807000.0 ;
      RECT  142800.0 820800.0 144000.0 818850.0 ;
      RECT  135600.0 810150.0 136800.0 808950.0 ;
      RECT  138000.0 810150.0 139200.0 808950.0 ;
      RECT  138000.0 810150.0 139200.0 808950.0 ;
      RECT  135600.0 810150.0 136800.0 808950.0 ;
      RECT  138000.0 810150.0 139200.0 808950.0 ;
      RECT  140400.0 810150.0 141600.0 808950.0 ;
      RECT  140400.0 810150.0 141600.0 808950.0 ;
      RECT  138000.0 810150.0 139200.0 808950.0 ;
      RECT  135600.0 818850.0 136800.0 817650.0 ;
      RECT  138000.0 818850.0 139200.0 817650.0 ;
      RECT  138000.0 818850.0 139200.0 817650.0 ;
      RECT  135600.0 818850.0 136800.0 817650.0 ;
      RECT  138000.0 818850.0 139200.0 817650.0 ;
      RECT  140400.0 818850.0 141600.0 817650.0 ;
      RECT  140400.0 818850.0 141600.0 817650.0 ;
      RECT  138000.0 818850.0 139200.0 817650.0 ;
      RECT  142800.0 809550.0 144000.0 808350.0 ;
      RECT  142800.0 819450.0 144000.0 818250.0 ;
      RECT  140400.0 816300.0 139200.0 815100.0 ;
      RECT  137400.0 813600.0 136200.0 812400.0 ;
      RECT  138000.0 810150.0 139200.0 808950.0 ;
      RECT  140400.0 818850.0 141600.0 817650.0 ;
      RECT  141600.0 813600.0 140400.0 812400.0 ;
      RECT  136200.0 813600.0 137400.0 812400.0 ;
      RECT  139200.0 816300.0 140400.0 815100.0 ;
      RECT  140400.0 813600.0 141600.0 812400.0 ;
      RECT  133800.0 807450.0 148200.0 806550.0 ;
      RECT  133800.0 821250.0 148200.0 820350.0 ;
      RECT  154800.0 808950.0 156000.0 807000.0 ;
      RECT  154800.0 820800.0 156000.0 818850.0 ;
      RECT  150000.0 819450.0 151200.0 821250.0 ;
      RECT  150000.0 810150.0 151200.0 806550.0 ;
      RECT  152700.0 819450.0 153600.0 810150.0 ;
      RECT  150000.0 810150.0 151200.0 808950.0 ;
      RECT  152400.0 810150.0 153600.0 808950.0 ;
      RECT  152400.0 810150.0 153600.0 808950.0 ;
      RECT  150000.0 810150.0 151200.0 808950.0 ;
      RECT  150000.0 819450.0 151200.0 818250.0 ;
      RECT  152400.0 819450.0 153600.0 818250.0 ;
      RECT  152400.0 819450.0 153600.0 818250.0 ;
      RECT  150000.0 819450.0 151200.0 818250.0 ;
      RECT  154800.0 809550.0 156000.0 808350.0 ;
      RECT  154800.0 819450.0 156000.0 818250.0 ;
      RECT  150600.0 814800.0 151800.0 813600.0 ;
      RECT  150600.0 814800.0 151800.0 813600.0 ;
      RECT  153150.0 814650.0 154050.0 813750.0 ;
      RECT  148200.0 807450.0 157800.0 806550.0 ;
      RECT  148200.0 821250.0 157800.0 820350.0 ;
      RECT  120450.0 813600.0 121650.0 814800.0 ;
      RECT  122400.0 816000.0 123600.0 817200.0 ;
      RECT  139200.0 815100.0 138000.0 816300.0 ;
      RECT  130800.0 832650.0 132000.0 834600.0 ;
      RECT  130800.0 820800.0 132000.0 822750.0 ;
      RECT  126000.0 822150.0 127200.0 820350.0 ;
      RECT  126000.0 831450.0 127200.0 835050.0 ;
      RECT  128700.0 822150.0 129600.0 831450.0 ;
      RECT  126000.0 831450.0 127200.0 832650.0 ;
      RECT  128400.0 831450.0 129600.0 832650.0 ;
      RECT  128400.0 831450.0 129600.0 832650.0 ;
      RECT  126000.0 831450.0 127200.0 832650.0 ;
      RECT  126000.0 822150.0 127200.0 823350.0 ;
      RECT  128400.0 822150.0 129600.0 823350.0 ;
      RECT  128400.0 822150.0 129600.0 823350.0 ;
      RECT  126000.0 822150.0 127200.0 823350.0 ;
      RECT  130800.0 832050.0 132000.0 833250.0 ;
      RECT  130800.0 822150.0 132000.0 823350.0 ;
      RECT  126600.0 826800.0 127800.0 828000.0 ;
      RECT  126600.0 826800.0 127800.0 828000.0 ;
      RECT  129150.0 826950.0 130050.0 827850.0 ;
      RECT  124200.0 834150.0 133800.0 835050.0 ;
      RECT  124200.0 820350.0 133800.0 821250.0 ;
      RECT  135600.0 822750.0 136800.0 820350.0 ;
      RECT  135600.0 831450.0 136800.0 835050.0 ;
      RECT  140400.0 831450.0 141600.0 835050.0 ;
      RECT  142800.0 832650.0 144000.0 834600.0 ;
      RECT  142800.0 820800.0 144000.0 822750.0 ;
      RECT  135600.0 831450.0 136800.0 832650.0 ;
      RECT  138000.0 831450.0 139200.0 832650.0 ;
      RECT  138000.0 831450.0 139200.0 832650.0 ;
      RECT  135600.0 831450.0 136800.0 832650.0 ;
      RECT  138000.0 831450.0 139200.0 832650.0 ;
      RECT  140400.0 831450.0 141600.0 832650.0 ;
      RECT  140400.0 831450.0 141600.0 832650.0 ;
      RECT  138000.0 831450.0 139200.0 832650.0 ;
      RECT  135600.0 822750.0 136800.0 823950.0 ;
      RECT  138000.0 822750.0 139200.0 823950.0 ;
      RECT  138000.0 822750.0 139200.0 823950.0 ;
      RECT  135600.0 822750.0 136800.0 823950.0 ;
      RECT  138000.0 822750.0 139200.0 823950.0 ;
      RECT  140400.0 822750.0 141600.0 823950.0 ;
      RECT  140400.0 822750.0 141600.0 823950.0 ;
      RECT  138000.0 822750.0 139200.0 823950.0 ;
      RECT  142800.0 832050.0 144000.0 833250.0 ;
      RECT  142800.0 822150.0 144000.0 823350.0 ;
      RECT  140400.0 825300.0 139200.0 826500.0 ;
      RECT  137400.0 828000.0 136200.0 829200.0 ;
      RECT  138000.0 831450.0 139200.0 832650.0 ;
      RECT  140400.0 822750.0 141600.0 823950.0 ;
      RECT  141600.0 828000.0 140400.0 829200.0 ;
      RECT  136200.0 828000.0 137400.0 829200.0 ;
      RECT  139200.0 825300.0 140400.0 826500.0 ;
      RECT  140400.0 828000.0 141600.0 829200.0 ;
      RECT  133800.0 834150.0 148200.0 835050.0 ;
      RECT  133800.0 820350.0 148200.0 821250.0 ;
      RECT  154800.0 832650.0 156000.0 834600.0 ;
      RECT  154800.0 820800.0 156000.0 822750.0 ;
      RECT  150000.0 822150.0 151200.0 820350.0 ;
      RECT  150000.0 831450.0 151200.0 835050.0 ;
      RECT  152700.0 822150.0 153600.0 831450.0 ;
      RECT  150000.0 831450.0 151200.0 832650.0 ;
      RECT  152400.0 831450.0 153600.0 832650.0 ;
      RECT  152400.0 831450.0 153600.0 832650.0 ;
      RECT  150000.0 831450.0 151200.0 832650.0 ;
      RECT  150000.0 822150.0 151200.0 823350.0 ;
      RECT  152400.0 822150.0 153600.0 823350.0 ;
      RECT  152400.0 822150.0 153600.0 823350.0 ;
      RECT  150000.0 822150.0 151200.0 823350.0 ;
      RECT  154800.0 832050.0 156000.0 833250.0 ;
      RECT  154800.0 822150.0 156000.0 823350.0 ;
      RECT  150600.0 826800.0 151800.0 828000.0 ;
      RECT  150600.0 826800.0 151800.0 828000.0 ;
      RECT  153150.0 826950.0 154050.0 827850.0 ;
      RECT  148200.0 834150.0 157800.0 835050.0 ;
      RECT  148200.0 820350.0 157800.0 821250.0 ;
      RECT  120450.0 826800.0 121650.0 828000.0 ;
      RECT  122400.0 824400.0 123600.0 825600.0 ;
      RECT  139200.0 825300.0 138000.0 826500.0 ;
      RECT  130800.0 836550.0 132000.0 834600.0 ;
      RECT  130800.0 848400.0 132000.0 846450.0 ;
      RECT  126000.0 847050.0 127200.0 848850.0 ;
      RECT  126000.0 837750.0 127200.0 834150.0 ;
      RECT  128700.0 847050.0 129600.0 837750.0 ;
      RECT  126000.0 837750.0 127200.0 836550.0 ;
      RECT  128400.0 837750.0 129600.0 836550.0 ;
      RECT  128400.0 837750.0 129600.0 836550.0 ;
      RECT  126000.0 837750.0 127200.0 836550.0 ;
      RECT  126000.0 847050.0 127200.0 845850.0 ;
      RECT  128400.0 847050.0 129600.0 845850.0 ;
      RECT  128400.0 847050.0 129600.0 845850.0 ;
      RECT  126000.0 847050.0 127200.0 845850.0 ;
      RECT  130800.0 837150.0 132000.0 835950.0 ;
      RECT  130800.0 847050.0 132000.0 845850.0 ;
      RECT  126600.0 842400.0 127800.0 841200.0 ;
      RECT  126600.0 842400.0 127800.0 841200.0 ;
      RECT  129150.0 842250.0 130050.0 841350.0 ;
      RECT  124200.0 835050.0 133800.0 834150.0 ;
      RECT  124200.0 848850.0 133800.0 847950.0 ;
      RECT  135600.0 846450.0 136800.0 848850.0 ;
      RECT  135600.0 837750.0 136800.0 834150.0 ;
      RECT  140400.0 837750.0 141600.0 834150.0 ;
      RECT  142800.0 836550.0 144000.0 834600.0 ;
      RECT  142800.0 848400.0 144000.0 846450.0 ;
      RECT  135600.0 837750.0 136800.0 836550.0 ;
      RECT  138000.0 837750.0 139200.0 836550.0 ;
      RECT  138000.0 837750.0 139200.0 836550.0 ;
      RECT  135600.0 837750.0 136800.0 836550.0 ;
      RECT  138000.0 837750.0 139200.0 836550.0 ;
      RECT  140400.0 837750.0 141600.0 836550.0 ;
      RECT  140400.0 837750.0 141600.0 836550.0 ;
      RECT  138000.0 837750.0 139200.0 836550.0 ;
      RECT  135600.0 846450.0 136800.0 845250.0 ;
      RECT  138000.0 846450.0 139200.0 845250.0 ;
      RECT  138000.0 846450.0 139200.0 845250.0 ;
      RECT  135600.0 846450.0 136800.0 845250.0 ;
      RECT  138000.0 846450.0 139200.0 845250.0 ;
      RECT  140400.0 846450.0 141600.0 845250.0 ;
      RECT  140400.0 846450.0 141600.0 845250.0 ;
      RECT  138000.0 846450.0 139200.0 845250.0 ;
      RECT  142800.0 837150.0 144000.0 835950.0 ;
      RECT  142800.0 847050.0 144000.0 845850.0 ;
      RECT  140400.0 843900.0 139200.0 842700.0 ;
      RECT  137400.0 841200.0 136200.0 840000.0 ;
      RECT  138000.0 837750.0 139200.0 836550.0 ;
      RECT  140400.0 846450.0 141600.0 845250.0 ;
      RECT  141600.0 841200.0 140400.0 840000.0 ;
      RECT  136200.0 841200.0 137400.0 840000.0 ;
      RECT  139200.0 843900.0 140400.0 842700.0 ;
      RECT  140400.0 841200.0 141600.0 840000.0 ;
      RECT  133800.0 835050.0 148200.0 834150.0 ;
      RECT  133800.0 848850.0 148200.0 847950.0 ;
      RECT  154800.0 836550.0 156000.0 834600.0 ;
      RECT  154800.0 848400.0 156000.0 846450.0 ;
      RECT  150000.0 847050.0 151200.0 848850.0 ;
      RECT  150000.0 837750.0 151200.0 834150.0 ;
      RECT  152700.0 847050.0 153600.0 837750.0 ;
      RECT  150000.0 837750.0 151200.0 836550.0 ;
      RECT  152400.0 837750.0 153600.0 836550.0 ;
      RECT  152400.0 837750.0 153600.0 836550.0 ;
      RECT  150000.0 837750.0 151200.0 836550.0 ;
      RECT  150000.0 847050.0 151200.0 845850.0 ;
      RECT  152400.0 847050.0 153600.0 845850.0 ;
      RECT  152400.0 847050.0 153600.0 845850.0 ;
      RECT  150000.0 847050.0 151200.0 845850.0 ;
      RECT  154800.0 837150.0 156000.0 835950.0 ;
      RECT  154800.0 847050.0 156000.0 845850.0 ;
      RECT  150600.0 842400.0 151800.0 841200.0 ;
      RECT  150600.0 842400.0 151800.0 841200.0 ;
      RECT  153150.0 842250.0 154050.0 841350.0 ;
      RECT  148200.0 835050.0 157800.0 834150.0 ;
      RECT  148200.0 848850.0 157800.0 847950.0 ;
      RECT  120450.0 841200.0 121650.0 842400.0 ;
      RECT  122400.0 843600.0 123600.0 844800.0 ;
      RECT  139200.0 842700.0 138000.0 843900.0 ;
      RECT  130800.0 860250.0 132000.0 862200.0 ;
      RECT  130800.0 848400.0 132000.0 850350.0 ;
      RECT  126000.0 849750.0 127200.0 847950.0 ;
      RECT  126000.0 859050.0 127200.0 862650.0 ;
      RECT  128700.0 849750.0 129600.0 859050.0 ;
      RECT  126000.0 859050.0 127200.0 860250.0 ;
      RECT  128400.0 859050.0 129600.0 860250.0 ;
      RECT  128400.0 859050.0 129600.0 860250.0 ;
      RECT  126000.0 859050.0 127200.0 860250.0 ;
      RECT  126000.0 849750.0 127200.0 850950.0 ;
      RECT  128400.0 849750.0 129600.0 850950.0 ;
      RECT  128400.0 849750.0 129600.0 850950.0 ;
      RECT  126000.0 849750.0 127200.0 850950.0 ;
      RECT  130800.0 859650.0 132000.0 860850.0 ;
      RECT  130800.0 849750.0 132000.0 850950.0 ;
      RECT  126600.0 854400.0 127800.0 855600.0 ;
      RECT  126600.0 854400.0 127800.0 855600.0 ;
      RECT  129150.0 854550.0 130050.0 855450.0 ;
      RECT  124200.0 861750.0 133800.0 862650.0 ;
      RECT  124200.0 847950.0 133800.0 848850.0 ;
      RECT  135600.0 850350.0 136800.0 847950.0 ;
      RECT  135600.0 859050.0 136800.0 862650.0 ;
      RECT  140400.0 859050.0 141600.0 862650.0 ;
      RECT  142800.0 860250.0 144000.0 862200.0 ;
      RECT  142800.0 848400.0 144000.0 850350.0 ;
      RECT  135600.0 859050.0 136800.0 860250.0 ;
      RECT  138000.0 859050.0 139200.0 860250.0 ;
      RECT  138000.0 859050.0 139200.0 860250.0 ;
      RECT  135600.0 859050.0 136800.0 860250.0 ;
      RECT  138000.0 859050.0 139200.0 860250.0 ;
      RECT  140400.0 859050.0 141600.0 860250.0 ;
      RECT  140400.0 859050.0 141600.0 860250.0 ;
      RECT  138000.0 859050.0 139200.0 860250.0 ;
      RECT  135600.0 850350.0 136800.0 851550.0 ;
      RECT  138000.0 850350.0 139200.0 851550.0 ;
      RECT  138000.0 850350.0 139200.0 851550.0 ;
      RECT  135600.0 850350.0 136800.0 851550.0 ;
      RECT  138000.0 850350.0 139200.0 851550.0 ;
      RECT  140400.0 850350.0 141600.0 851550.0 ;
      RECT  140400.0 850350.0 141600.0 851550.0 ;
      RECT  138000.0 850350.0 139200.0 851550.0 ;
      RECT  142800.0 859650.0 144000.0 860850.0 ;
      RECT  142800.0 849750.0 144000.0 850950.0 ;
      RECT  140400.0 852900.0 139200.0 854100.0 ;
      RECT  137400.0 855600.0 136200.0 856800.0 ;
      RECT  138000.0 859050.0 139200.0 860250.0 ;
      RECT  140400.0 850350.0 141600.0 851550.0 ;
      RECT  141600.0 855600.0 140400.0 856800.0 ;
      RECT  136200.0 855600.0 137400.0 856800.0 ;
      RECT  139200.0 852900.0 140400.0 854100.0 ;
      RECT  140400.0 855600.0 141600.0 856800.0 ;
      RECT  133800.0 861750.0 148200.0 862650.0 ;
      RECT  133800.0 847950.0 148200.0 848850.0 ;
      RECT  154800.0 860250.0 156000.0 862200.0 ;
      RECT  154800.0 848400.0 156000.0 850350.0 ;
      RECT  150000.0 849750.0 151200.0 847950.0 ;
      RECT  150000.0 859050.0 151200.0 862650.0 ;
      RECT  152700.0 849750.0 153600.0 859050.0 ;
      RECT  150000.0 859050.0 151200.0 860250.0 ;
      RECT  152400.0 859050.0 153600.0 860250.0 ;
      RECT  152400.0 859050.0 153600.0 860250.0 ;
      RECT  150000.0 859050.0 151200.0 860250.0 ;
      RECT  150000.0 849750.0 151200.0 850950.0 ;
      RECT  152400.0 849750.0 153600.0 850950.0 ;
      RECT  152400.0 849750.0 153600.0 850950.0 ;
      RECT  150000.0 849750.0 151200.0 850950.0 ;
      RECT  154800.0 859650.0 156000.0 860850.0 ;
      RECT  154800.0 849750.0 156000.0 850950.0 ;
      RECT  150600.0 854400.0 151800.0 855600.0 ;
      RECT  150600.0 854400.0 151800.0 855600.0 ;
      RECT  153150.0 854550.0 154050.0 855450.0 ;
      RECT  148200.0 861750.0 157800.0 862650.0 ;
      RECT  148200.0 847950.0 157800.0 848850.0 ;
      RECT  120450.0 854400.0 121650.0 855600.0 ;
      RECT  122400.0 852000.0 123600.0 853200.0 ;
      RECT  139200.0 852900.0 138000.0 854100.0 ;
      RECT  130800.0 864150.0 132000.0 862200.0 ;
      RECT  130800.0 876000.0 132000.0 874050.0 ;
      RECT  126000.0 874650.0 127200.0 876450.0 ;
      RECT  126000.0 865350.0 127200.0 861750.0 ;
      RECT  128700.0 874650.0 129600.0 865350.0 ;
      RECT  126000.0 865350.0 127200.0 864150.0 ;
      RECT  128400.0 865350.0 129600.0 864150.0 ;
      RECT  128400.0 865350.0 129600.0 864150.0 ;
      RECT  126000.0 865350.0 127200.0 864150.0 ;
      RECT  126000.0 874650.0 127200.0 873450.0 ;
      RECT  128400.0 874650.0 129600.0 873450.0 ;
      RECT  128400.0 874650.0 129600.0 873450.0 ;
      RECT  126000.0 874650.0 127200.0 873450.0 ;
      RECT  130800.0 864750.0 132000.0 863550.0 ;
      RECT  130800.0 874650.0 132000.0 873450.0 ;
      RECT  126600.0 870000.0 127800.0 868800.0 ;
      RECT  126600.0 870000.0 127800.0 868800.0 ;
      RECT  129150.0 869850.0 130050.0 868950.0 ;
      RECT  124200.0 862650.0 133800.0 861750.0 ;
      RECT  124200.0 876450.0 133800.0 875550.0 ;
      RECT  135600.0 874050.0 136800.0 876450.0 ;
      RECT  135600.0 865350.0 136800.0 861750.0 ;
      RECT  140400.0 865350.0 141600.0 861750.0 ;
      RECT  142800.0 864150.0 144000.0 862200.0 ;
      RECT  142800.0 876000.0 144000.0 874050.0 ;
      RECT  135600.0 865350.0 136800.0 864150.0 ;
      RECT  138000.0 865350.0 139200.0 864150.0 ;
      RECT  138000.0 865350.0 139200.0 864150.0 ;
      RECT  135600.0 865350.0 136800.0 864150.0 ;
      RECT  138000.0 865350.0 139200.0 864150.0 ;
      RECT  140400.0 865350.0 141600.0 864150.0 ;
      RECT  140400.0 865350.0 141600.0 864150.0 ;
      RECT  138000.0 865350.0 139200.0 864150.0 ;
      RECT  135600.0 874050.0 136800.0 872850.0 ;
      RECT  138000.0 874050.0 139200.0 872850.0 ;
      RECT  138000.0 874050.0 139200.0 872850.0 ;
      RECT  135600.0 874050.0 136800.0 872850.0 ;
      RECT  138000.0 874050.0 139200.0 872850.0 ;
      RECT  140400.0 874050.0 141600.0 872850.0 ;
      RECT  140400.0 874050.0 141600.0 872850.0 ;
      RECT  138000.0 874050.0 139200.0 872850.0 ;
      RECT  142800.0 864750.0 144000.0 863550.0 ;
      RECT  142800.0 874650.0 144000.0 873450.0 ;
      RECT  140400.0 871500.0 139200.0 870300.0 ;
      RECT  137400.0 868800.0 136200.0 867600.0 ;
      RECT  138000.0 865350.0 139200.0 864150.0 ;
      RECT  140400.0 874050.0 141600.0 872850.0 ;
      RECT  141600.0 868800.0 140400.0 867600.0 ;
      RECT  136200.0 868800.0 137400.0 867600.0 ;
      RECT  139200.0 871500.0 140400.0 870300.0 ;
      RECT  140400.0 868800.0 141600.0 867600.0 ;
      RECT  133800.0 862650.0 148200.0 861750.0 ;
      RECT  133800.0 876450.0 148200.0 875550.0 ;
      RECT  154800.0 864150.0 156000.0 862200.0 ;
      RECT  154800.0 876000.0 156000.0 874050.0 ;
      RECT  150000.0 874650.0 151200.0 876450.0 ;
      RECT  150000.0 865350.0 151200.0 861750.0 ;
      RECT  152700.0 874650.0 153600.0 865350.0 ;
      RECT  150000.0 865350.0 151200.0 864150.0 ;
      RECT  152400.0 865350.0 153600.0 864150.0 ;
      RECT  152400.0 865350.0 153600.0 864150.0 ;
      RECT  150000.0 865350.0 151200.0 864150.0 ;
      RECT  150000.0 874650.0 151200.0 873450.0 ;
      RECT  152400.0 874650.0 153600.0 873450.0 ;
      RECT  152400.0 874650.0 153600.0 873450.0 ;
      RECT  150000.0 874650.0 151200.0 873450.0 ;
      RECT  154800.0 864750.0 156000.0 863550.0 ;
      RECT  154800.0 874650.0 156000.0 873450.0 ;
      RECT  150600.0 870000.0 151800.0 868800.0 ;
      RECT  150600.0 870000.0 151800.0 868800.0 ;
      RECT  153150.0 869850.0 154050.0 868950.0 ;
      RECT  148200.0 862650.0 157800.0 861750.0 ;
      RECT  148200.0 876450.0 157800.0 875550.0 ;
      RECT  120450.0 868800.0 121650.0 870000.0 ;
      RECT  122400.0 871200.0 123600.0 872400.0 ;
      RECT  139200.0 870300.0 138000.0 871500.0 ;
      RECT  130800.0 887850.0 132000.0 889800.0 ;
      RECT  130800.0 876000.0 132000.0 877950.0 ;
      RECT  126000.0 877350.0 127200.0 875550.0 ;
      RECT  126000.0 886650.0 127200.0 890250.0 ;
      RECT  128700.0 877350.0 129600.0 886650.0 ;
      RECT  126000.0 886650.0 127200.0 887850.0 ;
      RECT  128400.0 886650.0 129600.0 887850.0 ;
      RECT  128400.0 886650.0 129600.0 887850.0 ;
      RECT  126000.0 886650.0 127200.0 887850.0 ;
      RECT  126000.0 877350.0 127200.0 878550.0 ;
      RECT  128400.0 877350.0 129600.0 878550.0 ;
      RECT  128400.0 877350.0 129600.0 878550.0 ;
      RECT  126000.0 877350.0 127200.0 878550.0 ;
      RECT  130800.0 887250.0 132000.0 888450.0 ;
      RECT  130800.0 877350.0 132000.0 878550.0 ;
      RECT  126600.0 882000.0 127800.0 883200.0 ;
      RECT  126600.0 882000.0 127800.0 883200.0 ;
      RECT  129150.0 882150.0 130050.0 883050.0 ;
      RECT  124200.0 889350.0 133800.0 890250.0 ;
      RECT  124200.0 875550.0 133800.0 876450.0 ;
      RECT  135600.0 877950.0 136800.0 875550.0 ;
      RECT  135600.0 886650.0 136800.0 890250.0 ;
      RECT  140400.0 886650.0 141600.0 890250.0 ;
      RECT  142800.0 887850.0 144000.0 889800.0 ;
      RECT  142800.0 876000.0 144000.0 877950.0 ;
      RECT  135600.0 886650.0 136800.0 887850.0 ;
      RECT  138000.0 886650.0 139200.0 887850.0 ;
      RECT  138000.0 886650.0 139200.0 887850.0 ;
      RECT  135600.0 886650.0 136800.0 887850.0 ;
      RECT  138000.0 886650.0 139200.0 887850.0 ;
      RECT  140400.0 886650.0 141600.0 887850.0 ;
      RECT  140400.0 886650.0 141600.0 887850.0 ;
      RECT  138000.0 886650.0 139200.0 887850.0 ;
      RECT  135600.0 877950.0 136800.0 879150.0 ;
      RECT  138000.0 877950.0 139200.0 879150.0 ;
      RECT  138000.0 877950.0 139200.0 879150.0 ;
      RECT  135600.0 877950.0 136800.0 879150.0 ;
      RECT  138000.0 877950.0 139200.0 879150.0 ;
      RECT  140400.0 877950.0 141600.0 879150.0 ;
      RECT  140400.0 877950.0 141600.0 879150.0 ;
      RECT  138000.0 877950.0 139200.0 879150.0 ;
      RECT  142800.0 887250.0 144000.0 888450.0 ;
      RECT  142800.0 877350.0 144000.0 878550.0 ;
      RECT  140400.0 880500.0 139200.0 881700.0 ;
      RECT  137400.0 883200.0 136200.0 884400.0 ;
      RECT  138000.0 886650.0 139200.0 887850.0 ;
      RECT  140400.0 877950.0 141600.0 879150.0 ;
      RECT  141600.0 883200.0 140400.0 884400.0 ;
      RECT  136200.0 883200.0 137400.0 884400.0 ;
      RECT  139200.0 880500.0 140400.0 881700.0 ;
      RECT  140400.0 883200.0 141600.0 884400.0 ;
      RECT  133800.0 889350.0 148200.0 890250.0 ;
      RECT  133800.0 875550.0 148200.0 876450.0 ;
      RECT  154800.0 887850.0 156000.0 889800.0 ;
      RECT  154800.0 876000.0 156000.0 877950.0 ;
      RECT  150000.0 877350.0 151200.0 875550.0 ;
      RECT  150000.0 886650.0 151200.0 890250.0 ;
      RECT  152700.0 877350.0 153600.0 886650.0 ;
      RECT  150000.0 886650.0 151200.0 887850.0 ;
      RECT  152400.0 886650.0 153600.0 887850.0 ;
      RECT  152400.0 886650.0 153600.0 887850.0 ;
      RECT  150000.0 886650.0 151200.0 887850.0 ;
      RECT  150000.0 877350.0 151200.0 878550.0 ;
      RECT  152400.0 877350.0 153600.0 878550.0 ;
      RECT  152400.0 877350.0 153600.0 878550.0 ;
      RECT  150000.0 877350.0 151200.0 878550.0 ;
      RECT  154800.0 887250.0 156000.0 888450.0 ;
      RECT  154800.0 877350.0 156000.0 878550.0 ;
      RECT  150600.0 882000.0 151800.0 883200.0 ;
      RECT  150600.0 882000.0 151800.0 883200.0 ;
      RECT  153150.0 882150.0 154050.0 883050.0 ;
      RECT  148200.0 889350.0 157800.0 890250.0 ;
      RECT  148200.0 875550.0 157800.0 876450.0 ;
      RECT  120450.0 882000.0 121650.0 883200.0 ;
      RECT  122400.0 879600.0 123600.0 880800.0 ;
      RECT  139200.0 880500.0 138000.0 881700.0 ;
      RECT  130800.0 891750.0 132000.0 889800.0 ;
      RECT  130800.0 903600.0 132000.0 901650.0 ;
      RECT  126000.0 902250.0 127200.0 904050.0 ;
      RECT  126000.0 892950.0 127200.0 889350.0 ;
      RECT  128700.0 902250.0 129600.0 892950.0 ;
      RECT  126000.0 892950.0 127200.0 891750.0 ;
      RECT  128400.0 892950.0 129600.0 891750.0 ;
      RECT  128400.0 892950.0 129600.0 891750.0 ;
      RECT  126000.0 892950.0 127200.0 891750.0 ;
      RECT  126000.0 902250.0 127200.0 901050.0 ;
      RECT  128400.0 902250.0 129600.0 901050.0 ;
      RECT  128400.0 902250.0 129600.0 901050.0 ;
      RECT  126000.0 902250.0 127200.0 901050.0 ;
      RECT  130800.0 892350.0 132000.0 891150.0 ;
      RECT  130800.0 902250.0 132000.0 901050.0 ;
      RECT  126600.0 897600.0 127800.0 896400.0 ;
      RECT  126600.0 897600.0 127800.0 896400.0 ;
      RECT  129150.0 897450.0 130050.0 896550.0 ;
      RECT  124200.0 890250.0 133800.0 889350.0 ;
      RECT  124200.0 904050.0 133800.0 903150.0 ;
      RECT  135600.0 901650.0 136800.0 904050.0 ;
      RECT  135600.0 892950.0 136800.0 889350.0 ;
      RECT  140400.0 892950.0 141600.0 889350.0 ;
      RECT  142800.0 891750.0 144000.0 889800.0 ;
      RECT  142800.0 903600.0 144000.0 901650.0 ;
      RECT  135600.0 892950.0 136800.0 891750.0 ;
      RECT  138000.0 892950.0 139200.0 891750.0 ;
      RECT  138000.0 892950.0 139200.0 891750.0 ;
      RECT  135600.0 892950.0 136800.0 891750.0 ;
      RECT  138000.0 892950.0 139200.0 891750.0 ;
      RECT  140400.0 892950.0 141600.0 891750.0 ;
      RECT  140400.0 892950.0 141600.0 891750.0 ;
      RECT  138000.0 892950.0 139200.0 891750.0 ;
      RECT  135600.0 901650.0 136800.0 900450.0 ;
      RECT  138000.0 901650.0 139200.0 900450.0 ;
      RECT  138000.0 901650.0 139200.0 900450.0 ;
      RECT  135600.0 901650.0 136800.0 900450.0 ;
      RECT  138000.0 901650.0 139200.0 900450.0 ;
      RECT  140400.0 901650.0 141600.0 900450.0 ;
      RECT  140400.0 901650.0 141600.0 900450.0 ;
      RECT  138000.0 901650.0 139200.0 900450.0 ;
      RECT  142800.0 892350.0 144000.0 891150.0 ;
      RECT  142800.0 902250.0 144000.0 901050.0 ;
      RECT  140400.0 899100.0 139200.0 897900.0 ;
      RECT  137400.0 896400.0 136200.0 895200.0 ;
      RECT  138000.0 892950.0 139200.0 891750.0 ;
      RECT  140400.0 901650.0 141600.0 900450.0 ;
      RECT  141600.0 896400.0 140400.0 895200.0 ;
      RECT  136200.0 896400.0 137400.0 895200.0 ;
      RECT  139200.0 899100.0 140400.0 897900.0 ;
      RECT  140400.0 896400.0 141600.0 895200.0 ;
      RECT  133800.0 890250.0 148200.0 889350.0 ;
      RECT  133800.0 904050.0 148200.0 903150.0 ;
      RECT  154800.0 891750.0 156000.0 889800.0 ;
      RECT  154800.0 903600.0 156000.0 901650.0 ;
      RECT  150000.0 902250.0 151200.0 904050.0 ;
      RECT  150000.0 892950.0 151200.0 889350.0 ;
      RECT  152700.0 902250.0 153600.0 892950.0 ;
      RECT  150000.0 892950.0 151200.0 891750.0 ;
      RECT  152400.0 892950.0 153600.0 891750.0 ;
      RECT  152400.0 892950.0 153600.0 891750.0 ;
      RECT  150000.0 892950.0 151200.0 891750.0 ;
      RECT  150000.0 902250.0 151200.0 901050.0 ;
      RECT  152400.0 902250.0 153600.0 901050.0 ;
      RECT  152400.0 902250.0 153600.0 901050.0 ;
      RECT  150000.0 902250.0 151200.0 901050.0 ;
      RECT  154800.0 892350.0 156000.0 891150.0 ;
      RECT  154800.0 902250.0 156000.0 901050.0 ;
      RECT  150600.0 897600.0 151800.0 896400.0 ;
      RECT  150600.0 897600.0 151800.0 896400.0 ;
      RECT  153150.0 897450.0 154050.0 896550.0 ;
      RECT  148200.0 890250.0 157800.0 889350.0 ;
      RECT  148200.0 904050.0 157800.0 903150.0 ;
      RECT  120450.0 896400.0 121650.0 897600.0 ;
      RECT  122400.0 898800.0 123600.0 900000.0 ;
      RECT  139200.0 897900.0 138000.0 899100.0 ;
      RECT  130800.0 915450.0 132000.0 917400.0 ;
      RECT  130800.0 903600.0 132000.0 905550.0 ;
      RECT  126000.0 904950.0 127200.0 903150.0 ;
      RECT  126000.0 914250.0 127200.0 917850.0 ;
      RECT  128700.0 904950.0 129600.0 914250.0 ;
      RECT  126000.0 914250.0 127200.0 915450.0 ;
      RECT  128400.0 914250.0 129600.0 915450.0 ;
      RECT  128400.0 914250.0 129600.0 915450.0 ;
      RECT  126000.0 914250.0 127200.0 915450.0 ;
      RECT  126000.0 904950.0 127200.0 906150.0 ;
      RECT  128400.0 904950.0 129600.0 906150.0 ;
      RECT  128400.0 904950.0 129600.0 906150.0 ;
      RECT  126000.0 904950.0 127200.0 906150.0 ;
      RECT  130800.0 914850.0 132000.0 916050.0 ;
      RECT  130800.0 904950.0 132000.0 906150.0 ;
      RECT  126600.0 909600.0 127800.0 910800.0 ;
      RECT  126600.0 909600.0 127800.0 910800.0 ;
      RECT  129150.0 909750.0 130050.0 910650.0 ;
      RECT  124200.0 916950.0 133800.0 917850.0 ;
      RECT  124200.0 903150.0 133800.0 904050.0 ;
      RECT  135600.0 905550.0 136800.0 903150.0 ;
      RECT  135600.0 914250.0 136800.0 917850.0 ;
      RECT  140400.0 914250.0 141600.0 917850.0 ;
      RECT  142800.0 915450.0 144000.0 917400.0 ;
      RECT  142800.0 903600.0 144000.0 905550.0 ;
      RECT  135600.0 914250.0 136800.0 915450.0 ;
      RECT  138000.0 914250.0 139200.0 915450.0 ;
      RECT  138000.0 914250.0 139200.0 915450.0 ;
      RECT  135600.0 914250.0 136800.0 915450.0 ;
      RECT  138000.0 914250.0 139200.0 915450.0 ;
      RECT  140400.0 914250.0 141600.0 915450.0 ;
      RECT  140400.0 914250.0 141600.0 915450.0 ;
      RECT  138000.0 914250.0 139200.0 915450.0 ;
      RECT  135600.0 905550.0 136800.0 906750.0 ;
      RECT  138000.0 905550.0 139200.0 906750.0 ;
      RECT  138000.0 905550.0 139200.0 906750.0 ;
      RECT  135600.0 905550.0 136800.0 906750.0 ;
      RECT  138000.0 905550.0 139200.0 906750.0 ;
      RECT  140400.0 905550.0 141600.0 906750.0 ;
      RECT  140400.0 905550.0 141600.0 906750.0 ;
      RECT  138000.0 905550.0 139200.0 906750.0 ;
      RECT  142800.0 914850.0 144000.0 916050.0 ;
      RECT  142800.0 904950.0 144000.0 906150.0 ;
      RECT  140400.0 908100.0 139200.0 909300.0 ;
      RECT  137400.0 910800.0 136200.0 912000.0 ;
      RECT  138000.0 914250.0 139200.0 915450.0 ;
      RECT  140400.0 905550.0 141600.0 906750.0 ;
      RECT  141600.0 910800.0 140400.0 912000.0 ;
      RECT  136200.0 910800.0 137400.0 912000.0 ;
      RECT  139200.0 908100.0 140400.0 909300.0 ;
      RECT  140400.0 910800.0 141600.0 912000.0 ;
      RECT  133800.0 916950.0 148200.0 917850.0 ;
      RECT  133800.0 903150.0 148200.0 904050.0 ;
      RECT  154800.0 915450.0 156000.0 917400.0 ;
      RECT  154800.0 903600.0 156000.0 905550.0 ;
      RECT  150000.0 904950.0 151200.0 903150.0 ;
      RECT  150000.0 914250.0 151200.0 917850.0 ;
      RECT  152700.0 904950.0 153600.0 914250.0 ;
      RECT  150000.0 914250.0 151200.0 915450.0 ;
      RECT  152400.0 914250.0 153600.0 915450.0 ;
      RECT  152400.0 914250.0 153600.0 915450.0 ;
      RECT  150000.0 914250.0 151200.0 915450.0 ;
      RECT  150000.0 904950.0 151200.0 906150.0 ;
      RECT  152400.0 904950.0 153600.0 906150.0 ;
      RECT  152400.0 904950.0 153600.0 906150.0 ;
      RECT  150000.0 904950.0 151200.0 906150.0 ;
      RECT  154800.0 914850.0 156000.0 916050.0 ;
      RECT  154800.0 904950.0 156000.0 906150.0 ;
      RECT  150600.0 909600.0 151800.0 910800.0 ;
      RECT  150600.0 909600.0 151800.0 910800.0 ;
      RECT  153150.0 909750.0 154050.0 910650.0 ;
      RECT  148200.0 916950.0 157800.0 917850.0 ;
      RECT  148200.0 903150.0 157800.0 904050.0 ;
      RECT  120450.0 909600.0 121650.0 910800.0 ;
      RECT  122400.0 907200.0 123600.0 908400.0 ;
      RECT  139200.0 908100.0 138000.0 909300.0 ;
      RECT  130800.0 919350.0 132000.0 917400.0 ;
      RECT  130800.0 931200.0 132000.0 929250.0 ;
      RECT  126000.0 929850.0 127200.0 931650.0 ;
      RECT  126000.0 920550.0 127200.0 916950.0 ;
      RECT  128700.0 929850.0 129600.0 920550.0 ;
      RECT  126000.0 920550.0 127200.0 919350.0 ;
      RECT  128400.0 920550.0 129600.0 919350.0 ;
      RECT  128400.0 920550.0 129600.0 919350.0 ;
      RECT  126000.0 920550.0 127200.0 919350.0 ;
      RECT  126000.0 929850.0 127200.0 928650.0 ;
      RECT  128400.0 929850.0 129600.0 928650.0 ;
      RECT  128400.0 929850.0 129600.0 928650.0 ;
      RECT  126000.0 929850.0 127200.0 928650.0 ;
      RECT  130800.0 919950.0 132000.0 918750.0 ;
      RECT  130800.0 929850.0 132000.0 928650.0 ;
      RECT  126600.0 925200.0 127800.0 924000.0 ;
      RECT  126600.0 925200.0 127800.0 924000.0 ;
      RECT  129150.0 925050.0 130050.0 924150.0 ;
      RECT  124200.0 917850.0 133800.0 916950.0 ;
      RECT  124200.0 931650.0 133800.0 930750.0 ;
      RECT  135600.0 929250.0 136800.0 931650.0 ;
      RECT  135600.0 920550.0 136800.0 916950.0 ;
      RECT  140400.0 920550.0 141600.0 916950.0 ;
      RECT  142800.0 919350.0 144000.0 917400.0 ;
      RECT  142800.0 931200.0 144000.0 929250.0 ;
      RECT  135600.0 920550.0 136800.0 919350.0 ;
      RECT  138000.0 920550.0 139200.0 919350.0 ;
      RECT  138000.0 920550.0 139200.0 919350.0 ;
      RECT  135600.0 920550.0 136800.0 919350.0 ;
      RECT  138000.0 920550.0 139200.0 919350.0 ;
      RECT  140400.0 920550.0 141600.0 919350.0 ;
      RECT  140400.0 920550.0 141600.0 919350.0 ;
      RECT  138000.0 920550.0 139200.0 919350.0 ;
      RECT  135600.0 929250.0 136800.0 928050.0 ;
      RECT  138000.0 929250.0 139200.0 928050.0 ;
      RECT  138000.0 929250.0 139200.0 928050.0 ;
      RECT  135600.0 929250.0 136800.0 928050.0 ;
      RECT  138000.0 929250.0 139200.0 928050.0 ;
      RECT  140400.0 929250.0 141600.0 928050.0 ;
      RECT  140400.0 929250.0 141600.0 928050.0 ;
      RECT  138000.0 929250.0 139200.0 928050.0 ;
      RECT  142800.0 919950.0 144000.0 918750.0 ;
      RECT  142800.0 929850.0 144000.0 928650.0 ;
      RECT  140400.0 926700.0 139200.0 925500.0 ;
      RECT  137400.0 924000.0 136200.0 922800.0 ;
      RECT  138000.0 920550.0 139200.0 919350.0 ;
      RECT  140400.0 929250.0 141600.0 928050.0 ;
      RECT  141600.0 924000.0 140400.0 922800.0 ;
      RECT  136200.0 924000.0 137400.0 922800.0 ;
      RECT  139200.0 926700.0 140400.0 925500.0 ;
      RECT  140400.0 924000.0 141600.0 922800.0 ;
      RECT  133800.0 917850.0 148200.0 916950.0 ;
      RECT  133800.0 931650.0 148200.0 930750.0 ;
      RECT  154800.0 919350.0 156000.0 917400.0 ;
      RECT  154800.0 931200.0 156000.0 929250.0 ;
      RECT  150000.0 929850.0 151200.0 931650.0 ;
      RECT  150000.0 920550.0 151200.0 916950.0 ;
      RECT  152700.0 929850.0 153600.0 920550.0 ;
      RECT  150000.0 920550.0 151200.0 919350.0 ;
      RECT  152400.0 920550.0 153600.0 919350.0 ;
      RECT  152400.0 920550.0 153600.0 919350.0 ;
      RECT  150000.0 920550.0 151200.0 919350.0 ;
      RECT  150000.0 929850.0 151200.0 928650.0 ;
      RECT  152400.0 929850.0 153600.0 928650.0 ;
      RECT  152400.0 929850.0 153600.0 928650.0 ;
      RECT  150000.0 929850.0 151200.0 928650.0 ;
      RECT  154800.0 919950.0 156000.0 918750.0 ;
      RECT  154800.0 929850.0 156000.0 928650.0 ;
      RECT  150600.0 925200.0 151800.0 924000.0 ;
      RECT  150600.0 925200.0 151800.0 924000.0 ;
      RECT  153150.0 925050.0 154050.0 924150.0 ;
      RECT  148200.0 917850.0 157800.0 916950.0 ;
      RECT  148200.0 931650.0 157800.0 930750.0 ;
      RECT  120450.0 924000.0 121650.0 925200.0 ;
      RECT  122400.0 926400.0 123600.0 927600.0 ;
      RECT  139200.0 925500.0 138000.0 926700.0 ;
      RECT  130800.0 943050.0 132000.0 945000.0 ;
      RECT  130800.0 931200.0 132000.0 933150.0 ;
      RECT  126000.0 932550.0 127200.0 930750.0 ;
      RECT  126000.0 941850.0 127200.0 945450.0 ;
      RECT  128700.0 932550.0 129600.0 941850.0 ;
      RECT  126000.0 941850.0 127200.0 943050.0 ;
      RECT  128400.0 941850.0 129600.0 943050.0 ;
      RECT  128400.0 941850.0 129600.0 943050.0 ;
      RECT  126000.0 941850.0 127200.0 943050.0 ;
      RECT  126000.0 932550.0 127200.0 933750.0 ;
      RECT  128400.0 932550.0 129600.0 933750.0 ;
      RECT  128400.0 932550.0 129600.0 933750.0 ;
      RECT  126000.0 932550.0 127200.0 933750.0 ;
      RECT  130800.0 942450.0 132000.0 943650.0 ;
      RECT  130800.0 932550.0 132000.0 933750.0 ;
      RECT  126600.0 937200.0 127800.0 938400.0 ;
      RECT  126600.0 937200.0 127800.0 938400.0 ;
      RECT  129150.0 937350.0 130050.0 938250.0 ;
      RECT  124200.0 944550.0 133800.0 945450.0 ;
      RECT  124200.0 930750.0 133800.0 931650.0 ;
      RECT  135600.0 933150.0 136800.0 930750.0 ;
      RECT  135600.0 941850.0 136800.0 945450.0 ;
      RECT  140400.0 941850.0 141600.0 945450.0 ;
      RECT  142800.0 943050.0 144000.0 945000.0 ;
      RECT  142800.0 931200.0 144000.0 933150.0 ;
      RECT  135600.0 941850.0 136800.0 943050.0 ;
      RECT  138000.0 941850.0 139200.0 943050.0 ;
      RECT  138000.0 941850.0 139200.0 943050.0 ;
      RECT  135600.0 941850.0 136800.0 943050.0 ;
      RECT  138000.0 941850.0 139200.0 943050.0 ;
      RECT  140400.0 941850.0 141600.0 943050.0 ;
      RECT  140400.0 941850.0 141600.0 943050.0 ;
      RECT  138000.0 941850.0 139200.0 943050.0 ;
      RECT  135600.0 933150.0 136800.0 934350.0 ;
      RECT  138000.0 933150.0 139200.0 934350.0 ;
      RECT  138000.0 933150.0 139200.0 934350.0 ;
      RECT  135600.0 933150.0 136800.0 934350.0 ;
      RECT  138000.0 933150.0 139200.0 934350.0 ;
      RECT  140400.0 933150.0 141600.0 934350.0 ;
      RECT  140400.0 933150.0 141600.0 934350.0 ;
      RECT  138000.0 933150.0 139200.0 934350.0 ;
      RECT  142800.0 942450.0 144000.0 943650.0 ;
      RECT  142800.0 932550.0 144000.0 933750.0 ;
      RECT  140400.0 935700.0 139200.0 936900.0 ;
      RECT  137400.0 938400.0 136200.0 939600.0 ;
      RECT  138000.0 941850.0 139200.0 943050.0 ;
      RECT  140400.0 933150.0 141600.0 934350.0 ;
      RECT  141600.0 938400.0 140400.0 939600.0 ;
      RECT  136200.0 938400.0 137400.0 939600.0 ;
      RECT  139200.0 935700.0 140400.0 936900.0 ;
      RECT  140400.0 938400.0 141600.0 939600.0 ;
      RECT  133800.0 944550.0 148200.0 945450.0 ;
      RECT  133800.0 930750.0 148200.0 931650.0 ;
      RECT  154800.0 943050.0 156000.0 945000.0 ;
      RECT  154800.0 931200.0 156000.0 933150.0 ;
      RECT  150000.0 932550.0 151200.0 930750.0 ;
      RECT  150000.0 941850.0 151200.0 945450.0 ;
      RECT  152700.0 932550.0 153600.0 941850.0 ;
      RECT  150000.0 941850.0 151200.0 943050.0 ;
      RECT  152400.0 941850.0 153600.0 943050.0 ;
      RECT  152400.0 941850.0 153600.0 943050.0 ;
      RECT  150000.0 941850.0 151200.0 943050.0 ;
      RECT  150000.0 932550.0 151200.0 933750.0 ;
      RECT  152400.0 932550.0 153600.0 933750.0 ;
      RECT  152400.0 932550.0 153600.0 933750.0 ;
      RECT  150000.0 932550.0 151200.0 933750.0 ;
      RECT  154800.0 942450.0 156000.0 943650.0 ;
      RECT  154800.0 932550.0 156000.0 933750.0 ;
      RECT  150600.0 937200.0 151800.0 938400.0 ;
      RECT  150600.0 937200.0 151800.0 938400.0 ;
      RECT  153150.0 937350.0 154050.0 938250.0 ;
      RECT  148200.0 944550.0 157800.0 945450.0 ;
      RECT  148200.0 930750.0 157800.0 931650.0 ;
      RECT  120450.0 937200.0 121650.0 938400.0 ;
      RECT  122400.0 934800.0 123600.0 936000.0 ;
      RECT  139200.0 935700.0 138000.0 936900.0 ;
      RECT  130800.0 946950.0 132000.0 945000.0 ;
      RECT  130800.0 958800.0 132000.0 956850.0 ;
      RECT  126000.0 957450.0 127200.0 959250.0 ;
      RECT  126000.0 948150.0 127200.0 944550.0 ;
      RECT  128700.0 957450.0 129600.0 948150.0 ;
      RECT  126000.0 948150.0 127200.0 946950.0 ;
      RECT  128400.0 948150.0 129600.0 946950.0 ;
      RECT  128400.0 948150.0 129600.0 946950.0 ;
      RECT  126000.0 948150.0 127200.0 946950.0 ;
      RECT  126000.0 957450.0 127200.0 956250.0 ;
      RECT  128400.0 957450.0 129600.0 956250.0 ;
      RECT  128400.0 957450.0 129600.0 956250.0 ;
      RECT  126000.0 957450.0 127200.0 956250.0 ;
      RECT  130800.0 947550.0 132000.0 946350.0 ;
      RECT  130800.0 957450.0 132000.0 956250.0 ;
      RECT  126600.0 952800.0 127800.0 951600.0 ;
      RECT  126600.0 952800.0 127800.0 951600.0 ;
      RECT  129150.0 952650.0 130050.0 951750.0 ;
      RECT  124200.0 945450.0 133800.0 944550.0 ;
      RECT  124200.0 959250.0 133800.0 958350.0 ;
      RECT  135600.0 956850.0 136800.0 959250.0 ;
      RECT  135600.0 948150.0 136800.0 944550.0 ;
      RECT  140400.0 948150.0 141600.0 944550.0 ;
      RECT  142800.0 946950.0 144000.0 945000.0 ;
      RECT  142800.0 958800.0 144000.0 956850.0 ;
      RECT  135600.0 948150.0 136800.0 946950.0 ;
      RECT  138000.0 948150.0 139200.0 946950.0 ;
      RECT  138000.0 948150.0 139200.0 946950.0 ;
      RECT  135600.0 948150.0 136800.0 946950.0 ;
      RECT  138000.0 948150.0 139200.0 946950.0 ;
      RECT  140400.0 948150.0 141600.0 946950.0 ;
      RECT  140400.0 948150.0 141600.0 946950.0 ;
      RECT  138000.0 948150.0 139200.0 946950.0 ;
      RECT  135600.0 956850.0 136800.0 955650.0 ;
      RECT  138000.0 956850.0 139200.0 955650.0 ;
      RECT  138000.0 956850.0 139200.0 955650.0 ;
      RECT  135600.0 956850.0 136800.0 955650.0 ;
      RECT  138000.0 956850.0 139200.0 955650.0 ;
      RECT  140400.0 956850.0 141600.0 955650.0 ;
      RECT  140400.0 956850.0 141600.0 955650.0 ;
      RECT  138000.0 956850.0 139200.0 955650.0 ;
      RECT  142800.0 947550.0 144000.0 946350.0 ;
      RECT  142800.0 957450.0 144000.0 956250.0 ;
      RECT  140400.0 954300.0 139200.0 953100.0 ;
      RECT  137400.0 951600.0 136200.0 950400.0 ;
      RECT  138000.0 948150.0 139200.0 946950.0 ;
      RECT  140400.0 956850.0 141600.0 955650.0 ;
      RECT  141600.0 951600.0 140400.0 950400.0 ;
      RECT  136200.0 951600.0 137400.0 950400.0 ;
      RECT  139200.0 954300.0 140400.0 953100.0 ;
      RECT  140400.0 951600.0 141600.0 950400.0 ;
      RECT  133800.0 945450.0 148200.0 944550.0 ;
      RECT  133800.0 959250.0 148200.0 958350.0 ;
      RECT  154800.0 946950.0 156000.0 945000.0 ;
      RECT  154800.0 958800.0 156000.0 956850.0 ;
      RECT  150000.0 957450.0 151200.0 959250.0 ;
      RECT  150000.0 948150.0 151200.0 944550.0 ;
      RECT  152700.0 957450.0 153600.0 948150.0 ;
      RECT  150000.0 948150.0 151200.0 946950.0 ;
      RECT  152400.0 948150.0 153600.0 946950.0 ;
      RECT  152400.0 948150.0 153600.0 946950.0 ;
      RECT  150000.0 948150.0 151200.0 946950.0 ;
      RECT  150000.0 957450.0 151200.0 956250.0 ;
      RECT  152400.0 957450.0 153600.0 956250.0 ;
      RECT  152400.0 957450.0 153600.0 956250.0 ;
      RECT  150000.0 957450.0 151200.0 956250.0 ;
      RECT  154800.0 947550.0 156000.0 946350.0 ;
      RECT  154800.0 957450.0 156000.0 956250.0 ;
      RECT  150600.0 952800.0 151800.0 951600.0 ;
      RECT  150600.0 952800.0 151800.0 951600.0 ;
      RECT  153150.0 952650.0 154050.0 951750.0 ;
      RECT  148200.0 945450.0 157800.0 944550.0 ;
      RECT  148200.0 959250.0 157800.0 958350.0 ;
      RECT  120450.0 951600.0 121650.0 952800.0 ;
      RECT  122400.0 954000.0 123600.0 955200.0 ;
      RECT  139200.0 953100.0 138000.0 954300.0 ;
      RECT  130800.0 970650.0 132000.0 972600.0 ;
      RECT  130800.0 958800.0 132000.0 960750.0 ;
      RECT  126000.0 960150.0 127200.0 958350.0 ;
      RECT  126000.0 969450.0 127200.0 973050.0 ;
      RECT  128700.0 960150.0 129600.0 969450.0 ;
      RECT  126000.0 969450.0 127200.0 970650.0 ;
      RECT  128400.0 969450.0 129600.0 970650.0 ;
      RECT  128400.0 969450.0 129600.0 970650.0 ;
      RECT  126000.0 969450.0 127200.0 970650.0 ;
      RECT  126000.0 960150.0 127200.0 961350.0 ;
      RECT  128400.0 960150.0 129600.0 961350.0 ;
      RECT  128400.0 960150.0 129600.0 961350.0 ;
      RECT  126000.0 960150.0 127200.0 961350.0 ;
      RECT  130800.0 970050.0 132000.0 971250.0 ;
      RECT  130800.0 960150.0 132000.0 961350.0 ;
      RECT  126600.0 964800.0 127800.0 966000.0 ;
      RECT  126600.0 964800.0 127800.0 966000.0 ;
      RECT  129150.0 964950.0 130050.0 965850.0 ;
      RECT  124200.0 972150.0 133800.0 973050.0 ;
      RECT  124200.0 958350.0 133800.0 959250.0 ;
      RECT  135600.0 960750.0 136800.0 958350.0 ;
      RECT  135600.0 969450.0 136800.0 973050.0 ;
      RECT  140400.0 969450.0 141600.0 973050.0 ;
      RECT  142800.0 970650.0 144000.0 972600.0 ;
      RECT  142800.0 958800.0 144000.0 960750.0 ;
      RECT  135600.0 969450.0 136800.0 970650.0 ;
      RECT  138000.0 969450.0 139200.0 970650.0 ;
      RECT  138000.0 969450.0 139200.0 970650.0 ;
      RECT  135600.0 969450.0 136800.0 970650.0 ;
      RECT  138000.0 969450.0 139200.0 970650.0 ;
      RECT  140400.0 969450.0 141600.0 970650.0 ;
      RECT  140400.0 969450.0 141600.0 970650.0 ;
      RECT  138000.0 969450.0 139200.0 970650.0 ;
      RECT  135600.0 960750.0 136800.0 961950.0 ;
      RECT  138000.0 960750.0 139200.0 961950.0 ;
      RECT  138000.0 960750.0 139200.0 961950.0 ;
      RECT  135600.0 960750.0 136800.0 961950.0 ;
      RECT  138000.0 960750.0 139200.0 961950.0 ;
      RECT  140400.0 960750.0 141600.0 961950.0 ;
      RECT  140400.0 960750.0 141600.0 961950.0 ;
      RECT  138000.0 960750.0 139200.0 961950.0 ;
      RECT  142800.0 970050.0 144000.0 971250.0 ;
      RECT  142800.0 960150.0 144000.0 961350.0 ;
      RECT  140400.0 963300.0 139200.0 964500.0 ;
      RECT  137400.0 966000.0 136200.0 967200.0 ;
      RECT  138000.0 969450.0 139200.0 970650.0 ;
      RECT  140400.0 960750.0 141600.0 961950.0 ;
      RECT  141600.0 966000.0 140400.0 967200.0 ;
      RECT  136200.0 966000.0 137400.0 967200.0 ;
      RECT  139200.0 963300.0 140400.0 964500.0 ;
      RECT  140400.0 966000.0 141600.0 967200.0 ;
      RECT  133800.0 972150.0 148200.0 973050.0 ;
      RECT  133800.0 958350.0 148200.0 959250.0 ;
      RECT  154800.0 970650.0 156000.0 972600.0 ;
      RECT  154800.0 958800.0 156000.0 960750.0 ;
      RECT  150000.0 960150.0 151200.0 958350.0 ;
      RECT  150000.0 969450.0 151200.0 973050.0 ;
      RECT  152700.0 960150.0 153600.0 969450.0 ;
      RECT  150000.0 969450.0 151200.0 970650.0 ;
      RECT  152400.0 969450.0 153600.0 970650.0 ;
      RECT  152400.0 969450.0 153600.0 970650.0 ;
      RECT  150000.0 969450.0 151200.0 970650.0 ;
      RECT  150000.0 960150.0 151200.0 961350.0 ;
      RECT  152400.0 960150.0 153600.0 961350.0 ;
      RECT  152400.0 960150.0 153600.0 961350.0 ;
      RECT  150000.0 960150.0 151200.0 961350.0 ;
      RECT  154800.0 970050.0 156000.0 971250.0 ;
      RECT  154800.0 960150.0 156000.0 961350.0 ;
      RECT  150600.0 964800.0 151800.0 966000.0 ;
      RECT  150600.0 964800.0 151800.0 966000.0 ;
      RECT  153150.0 964950.0 154050.0 965850.0 ;
      RECT  148200.0 972150.0 157800.0 973050.0 ;
      RECT  148200.0 958350.0 157800.0 959250.0 ;
      RECT  120450.0 964800.0 121650.0 966000.0 ;
      RECT  122400.0 962400.0 123600.0 963600.0 ;
      RECT  139200.0 963300.0 138000.0 964500.0 ;
      RECT  130800.0 974550.0 132000.0 972600.0 ;
      RECT  130800.0 986400.0 132000.0 984450.0 ;
      RECT  126000.0 985050.0 127200.0 986850.0 ;
      RECT  126000.0 975750.0 127200.0 972150.0 ;
      RECT  128700.0 985050.0 129600.0 975750.0 ;
      RECT  126000.0 975750.0 127200.0 974550.0 ;
      RECT  128400.0 975750.0 129600.0 974550.0 ;
      RECT  128400.0 975750.0 129600.0 974550.0 ;
      RECT  126000.0 975750.0 127200.0 974550.0 ;
      RECT  126000.0 985050.0 127200.0 983850.0 ;
      RECT  128400.0 985050.0 129600.0 983850.0 ;
      RECT  128400.0 985050.0 129600.0 983850.0 ;
      RECT  126000.0 985050.0 127200.0 983850.0 ;
      RECT  130800.0 975150.0 132000.0 973950.0 ;
      RECT  130800.0 985050.0 132000.0 983850.0 ;
      RECT  126600.0 980400.0 127800.0 979200.0 ;
      RECT  126600.0 980400.0 127800.0 979200.0 ;
      RECT  129150.0 980250.0 130050.0 979350.0 ;
      RECT  124200.0 973050.0 133800.0 972150.0 ;
      RECT  124200.0 986850.0 133800.0 985950.0 ;
      RECT  135600.0 984450.0 136800.0 986850.0 ;
      RECT  135600.0 975750.0 136800.0 972150.0 ;
      RECT  140400.0 975750.0 141600.0 972150.0 ;
      RECT  142800.0 974550.0 144000.0 972600.0 ;
      RECT  142800.0 986400.0 144000.0 984450.0 ;
      RECT  135600.0 975750.0 136800.0 974550.0 ;
      RECT  138000.0 975750.0 139200.0 974550.0 ;
      RECT  138000.0 975750.0 139200.0 974550.0 ;
      RECT  135600.0 975750.0 136800.0 974550.0 ;
      RECT  138000.0 975750.0 139200.0 974550.0 ;
      RECT  140400.0 975750.0 141600.0 974550.0 ;
      RECT  140400.0 975750.0 141600.0 974550.0 ;
      RECT  138000.0 975750.0 139200.0 974550.0 ;
      RECT  135600.0 984450.0 136800.0 983250.0 ;
      RECT  138000.0 984450.0 139200.0 983250.0 ;
      RECT  138000.0 984450.0 139200.0 983250.0 ;
      RECT  135600.0 984450.0 136800.0 983250.0 ;
      RECT  138000.0 984450.0 139200.0 983250.0 ;
      RECT  140400.0 984450.0 141600.0 983250.0 ;
      RECT  140400.0 984450.0 141600.0 983250.0 ;
      RECT  138000.0 984450.0 139200.0 983250.0 ;
      RECT  142800.0 975150.0 144000.0 973950.0 ;
      RECT  142800.0 985050.0 144000.0 983850.0 ;
      RECT  140400.0 981900.0 139200.0 980700.0 ;
      RECT  137400.0 979200.0 136200.0 978000.0 ;
      RECT  138000.0 975750.0 139200.0 974550.0 ;
      RECT  140400.0 984450.0 141600.0 983250.0 ;
      RECT  141600.0 979200.0 140400.0 978000.0 ;
      RECT  136200.0 979200.0 137400.0 978000.0 ;
      RECT  139200.0 981900.0 140400.0 980700.0 ;
      RECT  140400.0 979200.0 141600.0 978000.0 ;
      RECT  133800.0 973050.0 148200.0 972150.0 ;
      RECT  133800.0 986850.0 148200.0 985950.0 ;
      RECT  154800.0 974550.0 156000.0 972600.0 ;
      RECT  154800.0 986400.0 156000.0 984450.0 ;
      RECT  150000.0 985050.0 151200.0 986850.0 ;
      RECT  150000.0 975750.0 151200.0 972150.0 ;
      RECT  152700.0 985050.0 153600.0 975750.0 ;
      RECT  150000.0 975750.0 151200.0 974550.0 ;
      RECT  152400.0 975750.0 153600.0 974550.0 ;
      RECT  152400.0 975750.0 153600.0 974550.0 ;
      RECT  150000.0 975750.0 151200.0 974550.0 ;
      RECT  150000.0 985050.0 151200.0 983850.0 ;
      RECT  152400.0 985050.0 153600.0 983850.0 ;
      RECT  152400.0 985050.0 153600.0 983850.0 ;
      RECT  150000.0 985050.0 151200.0 983850.0 ;
      RECT  154800.0 975150.0 156000.0 973950.0 ;
      RECT  154800.0 985050.0 156000.0 983850.0 ;
      RECT  150600.0 980400.0 151800.0 979200.0 ;
      RECT  150600.0 980400.0 151800.0 979200.0 ;
      RECT  153150.0 980250.0 154050.0 979350.0 ;
      RECT  148200.0 973050.0 157800.0 972150.0 ;
      RECT  148200.0 986850.0 157800.0 985950.0 ;
      RECT  120450.0 979200.0 121650.0 980400.0 ;
      RECT  122400.0 981600.0 123600.0 982800.0 ;
      RECT  139200.0 980700.0 138000.0 981900.0 ;
      RECT  130800.0 998250.0 132000.0 1000200.0 ;
      RECT  130800.0 986400.0 132000.0 988350.0 ;
      RECT  126000.0 987750.0 127200.0 985950.0 ;
      RECT  126000.0 997050.0 127200.0 1000650.0 ;
      RECT  128700.0 987750.0 129600.0 997050.0 ;
      RECT  126000.0 997050.0 127200.0 998250.0 ;
      RECT  128400.0 997050.0 129600.0 998250.0 ;
      RECT  128400.0 997050.0 129600.0 998250.0 ;
      RECT  126000.0 997050.0 127200.0 998250.0 ;
      RECT  126000.0 987750.0 127200.0 988950.0 ;
      RECT  128400.0 987750.0 129600.0 988950.0 ;
      RECT  128400.0 987750.0 129600.0 988950.0 ;
      RECT  126000.0 987750.0 127200.0 988950.0 ;
      RECT  130800.0 997650.0 132000.0 998850.0 ;
      RECT  130800.0 987750.0 132000.0 988950.0 ;
      RECT  126600.0 992400.0 127800.0 993600.0 ;
      RECT  126600.0 992400.0 127800.0 993600.0 ;
      RECT  129150.0 992550.0 130050.0 993450.0 ;
      RECT  124200.0 999750.0 133800.0 1000650.0 ;
      RECT  124200.0 985950.0 133800.0 986850.0 ;
      RECT  135600.0 988350.0 136800.0 985950.0 ;
      RECT  135600.0 997050.0 136800.0 1000650.0 ;
      RECT  140400.0 997050.0 141600.0 1000650.0 ;
      RECT  142800.0 998250.0 144000.0 1000200.0 ;
      RECT  142800.0 986400.0 144000.0 988350.0 ;
      RECT  135600.0 997050.0 136800.0 998250.0 ;
      RECT  138000.0 997050.0 139200.0 998250.0 ;
      RECT  138000.0 997050.0 139200.0 998250.0 ;
      RECT  135600.0 997050.0 136800.0 998250.0 ;
      RECT  138000.0 997050.0 139200.0 998250.0 ;
      RECT  140400.0 997050.0 141600.0 998250.0 ;
      RECT  140400.0 997050.0 141600.0 998250.0 ;
      RECT  138000.0 997050.0 139200.0 998250.0 ;
      RECT  135600.0 988350.0 136800.0 989550.0 ;
      RECT  138000.0 988350.0 139200.0 989550.0 ;
      RECT  138000.0 988350.0 139200.0 989550.0 ;
      RECT  135600.0 988350.0 136800.0 989550.0 ;
      RECT  138000.0 988350.0 139200.0 989550.0 ;
      RECT  140400.0 988350.0 141600.0 989550.0 ;
      RECT  140400.0 988350.0 141600.0 989550.0 ;
      RECT  138000.0 988350.0 139200.0 989550.0 ;
      RECT  142800.0 997650.0 144000.0 998850.0 ;
      RECT  142800.0 987750.0 144000.0 988950.0 ;
      RECT  140400.0 990900.0 139200.0 992100.0 ;
      RECT  137400.0 993600.0 136200.0 994800.0 ;
      RECT  138000.0 997050.0 139200.0 998250.0 ;
      RECT  140400.0 988350.0 141600.0 989550.0 ;
      RECT  141600.0 993600.0 140400.0 994800.0 ;
      RECT  136200.0 993600.0 137400.0 994800.0 ;
      RECT  139200.0 990900.0 140400.0 992100.0 ;
      RECT  140400.0 993600.0 141600.0 994800.0 ;
      RECT  133800.0 999750.0 148200.0 1000650.0 ;
      RECT  133800.0 985950.0 148200.0 986850.0 ;
      RECT  154800.0 998250.0 156000.0 1000200.0 ;
      RECT  154800.0 986400.0 156000.0 988350.0 ;
      RECT  150000.0 987750.0 151200.0 985950.0 ;
      RECT  150000.0 997050.0 151200.0 1000650.0 ;
      RECT  152700.0 987750.0 153600.0 997050.0 ;
      RECT  150000.0 997050.0 151200.0 998250.0 ;
      RECT  152400.0 997050.0 153600.0 998250.0 ;
      RECT  152400.0 997050.0 153600.0 998250.0 ;
      RECT  150000.0 997050.0 151200.0 998250.0 ;
      RECT  150000.0 987750.0 151200.0 988950.0 ;
      RECT  152400.0 987750.0 153600.0 988950.0 ;
      RECT  152400.0 987750.0 153600.0 988950.0 ;
      RECT  150000.0 987750.0 151200.0 988950.0 ;
      RECT  154800.0 997650.0 156000.0 998850.0 ;
      RECT  154800.0 987750.0 156000.0 988950.0 ;
      RECT  150600.0 992400.0 151800.0 993600.0 ;
      RECT  150600.0 992400.0 151800.0 993600.0 ;
      RECT  153150.0 992550.0 154050.0 993450.0 ;
      RECT  148200.0 999750.0 157800.0 1000650.0 ;
      RECT  148200.0 985950.0 157800.0 986850.0 ;
      RECT  120450.0 992400.0 121650.0 993600.0 ;
      RECT  122400.0 990000.0 123600.0 991200.0 ;
      RECT  139200.0 990900.0 138000.0 992100.0 ;
      RECT  130800.0 1002150.0 132000.0 1000200.0 ;
      RECT  130800.0 1014000.0 132000.0 1012050.0 ;
      RECT  126000.0 1012650.0 127200.0 1014450.0 ;
      RECT  126000.0 1003350.0 127200.0 999750.0 ;
      RECT  128700.0 1012650.0 129600.0 1003350.0 ;
      RECT  126000.0 1003350.0 127200.0 1002150.0 ;
      RECT  128400.0 1003350.0 129600.0 1002150.0 ;
      RECT  128400.0 1003350.0 129600.0 1002150.0 ;
      RECT  126000.0 1003350.0 127200.0 1002150.0 ;
      RECT  126000.0 1012650.0 127200.0 1011450.0 ;
      RECT  128400.0 1012650.0 129600.0 1011450.0 ;
      RECT  128400.0 1012650.0 129600.0 1011450.0 ;
      RECT  126000.0 1012650.0 127200.0 1011450.0 ;
      RECT  130800.0 1002750.0 132000.0 1001550.0 ;
      RECT  130800.0 1012650.0 132000.0 1011450.0 ;
      RECT  126600.0 1008000.0 127800.0 1006800.0 ;
      RECT  126600.0 1008000.0 127800.0 1006800.0 ;
      RECT  129150.0 1007850.0 130050.0 1006950.0 ;
      RECT  124200.0 1000650.0 133800.0 999750.0 ;
      RECT  124200.0 1014450.0 133800.0 1013550.0 ;
      RECT  135600.0 1012050.0 136800.0 1014450.0 ;
      RECT  135600.0 1003350.0 136800.0 999750.0 ;
      RECT  140400.0 1003350.0 141600.0 999750.0 ;
      RECT  142800.0 1002150.0 144000.0 1000200.0 ;
      RECT  142800.0 1014000.0 144000.0 1012050.0 ;
      RECT  135600.0 1003350.0 136800.0 1002150.0 ;
      RECT  138000.0 1003350.0 139200.0 1002150.0 ;
      RECT  138000.0 1003350.0 139200.0 1002150.0 ;
      RECT  135600.0 1003350.0 136800.0 1002150.0 ;
      RECT  138000.0 1003350.0 139200.0 1002150.0 ;
      RECT  140400.0 1003350.0 141600.0 1002150.0 ;
      RECT  140400.0 1003350.0 141600.0 1002150.0 ;
      RECT  138000.0 1003350.0 139200.0 1002150.0 ;
      RECT  135600.0 1012050.0 136800.0 1010850.0 ;
      RECT  138000.0 1012050.0 139200.0 1010850.0 ;
      RECT  138000.0 1012050.0 139200.0 1010850.0 ;
      RECT  135600.0 1012050.0 136800.0 1010850.0 ;
      RECT  138000.0 1012050.0 139200.0 1010850.0 ;
      RECT  140400.0 1012050.0 141600.0 1010850.0 ;
      RECT  140400.0 1012050.0 141600.0 1010850.0 ;
      RECT  138000.0 1012050.0 139200.0 1010850.0 ;
      RECT  142800.0 1002750.0 144000.0 1001550.0 ;
      RECT  142800.0 1012650.0 144000.0 1011450.0 ;
      RECT  140400.0 1009500.0 139200.0 1008300.0 ;
      RECT  137400.0 1006800.0 136200.0 1005600.0 ;
      RECT  138000.0 1003350.0 139200.0 1002150.0 ;
      RECT  140400.0 1012050.0 141600.0 1010850.0 ;
      RECT  141600.0 1006800.0 140400.0 1005600.0 ;
      RECT  136200.0 1006800.0 137400.0 1005600.0 ;
      RECT  139200.0 1009500.0 140400.0 1008300.0 ;
      RECT  140400.0 1006800.0 141600.0 1005600.0 ;
      RECT  133800.0 1000650.0 148200.0 999750.0 ;
      RECT  133800.0 1014450.0 148200.0 1013550.0 ;
      RECT  154800.0 1002150.0 156000.0 1000200.0 ;
      RECT  154800.0 1014000.0 156000.0 1012050.0 ;
      RECT  150000.0 1012650.0 151200.0 1014450.0 ;
      RECT  150000.0 1003350.0 151200.0 999750.0 ;
      RECT  152700.0 1012650.0 153600.0 1003350.0 ;
      RECT  150000.0 1003350.0 151200.0 1002150.0 ;
      RECT  152400.0 1003350.0 153600.0 1002150.0 ;
      RECT  152400.0 1003350.0 153600.0 1002150.0 ;
      RECT  150000.0 1003350.0 151200.0 1002150.0 ;
      RECT  150000.0 1012650.0 151200.0 1011450.0 ;
      RECT  152400.0 1012650.0 153600.0 1011450.0 ;
      RECT  152400.0 1012650.0 153600.0 1011450.0 ;
      RECT  150000.0 1012650.0 151200.0 1011450.0 ;
      RECT  154800.0 1002750.0 156000.0 1001550.0 ;
      RECT  154800.0 1012650.0 156000.0 1011450.0 ;
      RECT  150600.0 1008000.0 151800.0 1006800.0 ;
      RECT  150600.0 1008000.0 151800.0 1006800.0 ;
      RECT  153150.0 1007850.0 154050.0 1006950.0 ;
      RECT  148200.0 1000650.0 157800.0 999750.0 ;
      RECT  148200.0 1014450.0 157800.0 1013550.0 ;
      RECT  120450.0 1006800.0 121650.0 1008000.0 ;
      RECT  122400.0 1009200.0 123600.0 1010400.0 ;
      RECT  139200.0 1008300.0 138000.0 1009500.0 ;
      RECT  130800.0 1025850.0 132000.0 1027800.0 ;
      RECT  130800.0 1014000.0 132000.0 1015950.0 ;
      RECT  126000.0 1015350.0 127200.0 1013550.0 ;
      RECT  126000.0 1024650.0 127200.0 1028250.0 ;
      RECT  128700.0 1015350.0 129600.0 1024650.0 ;
      RECT  126000.0 1024650.0 127200.0 1025850.0 ;
      RECT  128400.0 1024650.0 129600.0 1025850.0 ;
      RECT  128400.0 1024650.0 129600.0 1025850.0 ;
      RECT  126000.0 1024650.0 127200.0 1025850.0 ;
      RECT  126000.0 1015350.0 127200.0 1016550.0 ;
      RECT  128400.0 1015350.0 129600.0 1016550.0 ;
      RECT  128400.0 1015350.0 129600.0 1016550.0 ;
      RECT  126000.0 1015350.0 127200.0 1016550.0 ;
      RECT  130800.0 1025250.0 132000.0 1026450.0 ;
      RECT  130800.0 1015350.0 132000.0 1016550.0 ;
      RECT  126600.0 1020000.0 127800.0 1021200.0 ;
      RECT  126600.0 1020000.0 127800.0 1021200.0 ;
      RECT  129150.0 1020150.0 130050.0 1021050.0 ;
      RECT  124200.0 1027350.0 133800.0 1028250.0 ;
      RECT  124200.0 1013550.0 133800.0 1014450.0 ;
      RECT  135600.0 1015950.0 136800.0 1013550.0 ;
      RECT  135600.0 1024650.0 136800.0 1028250.0 ;
      RECT  140400.0 1024650.0 141600.0 1028250.0 ;
      RECT  142800.0 1025850.0 144000.0 1027800.0 ;
      RECT  142800.0 1014000.0 144000.0 1015950.0 ;
      RECT  135600.0 1024650.0 136800.0 1025850.0 ;
      RECT  138000.0 1024650.0 139200.0 1025850.0 ;
      RECT  138000.0 1024650.0 139200.0 1025850.0 ;
      RECT  135600.0 1024650.0 136800.0 1025850.0 ;
      RECT  138000.0 1024650.0 139200.0 1025850.0 ;
      RECT  140400.0 1024650.0 141600.0 1025850.0 ;
      RECT  140400.0 1024650.0 141600.0 1025850.0 ;
      RECT  138000.0 1024650.0 139200.0 1025850.0 ;
      RECT  135600.0 1015950.0 136800.0 1017150.0 ;
      RECT  138000.0 1015950.0 139200.0 1017150.0 ;
      RECT  138000.0 1015950.0 139200.0 1017150.0 ;
      RECT  135600.0 1015950.0 136800.0 1017150.0 ;
      RECT  138000.0 1015950.0 139200.0 1017150.0 ;
      RECT  140400.0 1015950.0 141600.0 1017150.0 ;
      RECT  140400.0 1015950.0 141600.0 1017150.0 ;
      RECT  138000.0 1015950.0 139200.0 1017150.0 ;
      RECT  142800.0 1025250.0 144000.0 1026450.0 ;
      RECT  142800.0 1015350.0 144000.0 1016550.0 ;
      RECT  140400.0 1018500.0 139200.0 1019700.0 ;
      RECT  137400.0 1021200.0 136200.0 1022400.0 ;
      RECT  138000.0 1024650.0 139200.0 1025850.0 ;
      RECT  140400.0 1015950.0 141600.0 1017150.0 ;
      RECT  141600.0 1021200.0 140400.0 1022400.0 ;
      RECT  136200.0 1021200.0 137400.0 1022400.0 ;
      RECT  139200.0 1018500.0 140400.0 1019700.0 ;
      RECT  140400.0 1021200.0 141600.0 1022400.0 ;
      RECT  133800.0 1027350.0 148200.0 1028250.0 ;
      RECT  133800.0 1013550.0 148200.0 1014450.0 ;
      RECT  154800.0 1025850.0 156000.0 1027800.0 ;
      RECT  154800.0 1014000.0 156000.0 1015950.0 ;
      RECT  150000.0 1015350.0 151200.0 1013550.0 ;
      RECT  150000.0 1024650.0 151200.0 1028250.0 ;
      RECT  152700.0 1015350.0 153600.0 1024650.0 ;
      RECT  150000.0 1024650.0 151200.0 1025850.0 ;
      RECT  152400.0 1024650.0 153600.0 1025850.0 ;
      RECT  152400.0 1024650.0 153600.0 1025850.0 ;
      RECT  150000.0 1024650.0 151200.0 1025850.0 ;
      RECT  150000.0 1015350.0 151200.0 1016550.0 ;
      RECT  152400.0 1015350.0 153600.0 1016550.0 ;
      RECT  152400.0 1015350.0 153600.0 1016550.0 ;
      RECT  150000.0 1015350.0 151200.0 1016550.0 ;
      RECT  154800.0 1025250.0 156000.0 1026450.0 ;
      RECT  154800.0 1015350.0 156000.0 1016550.0 ;
      RECT  150600.0 1020000.0 151800.0 1021200.0 ;
      RECT  150600.0 1020000.0 151800.0 1021200.0 ;
      RECT  153150.0 1020150.0 154050.0 1021050.0 ;
      RECT  148200.0 1027350.0 157800.0 1028250.0 ;
      RECT  148200.0 1013550.0 157800.0 1014450.0 ;
      RECT  120450.0 1020000.0 121650.0 1021200.0 ;
      RECT  122400.0 1017600.0 123600.0 1018800.0 ;
      RECT  139200.0 1018500.0 138000.0 1019700.0 ;
      RECT  130800.0 1029750.0 132000.0 1027800.0 ;
      RECT  130800.0 1041600.0 132000.0 1039650.0 ;
      RECT  126000.0 1040250.0 127200.0 1042050.0 ;
      RECT  126000.0 1030950.0 127200.0 1027350.0 ;
      RECT  128700.0 1040250.0 129600.0 1030950.0 ;
      RECT  126000.0 1030950.0 127200.0 1029750.0 ;
      RECT  128400.0 1030950.0 129600.0 1029750.0 ;
      RECT  128400.0 1030950.0 129600.0 1029750.0 ;
      RECT  126000.0 1030950.0 127200.0 1029750.0 ;
      RECT  126000.0 1040250.0 127200.0 1039050.0 ;
      RECT  128400.0 1040250.0 129600.0 1039050.0 ;
      RECT  128400.0 1040250.0 129600.0 1039050.0 ;
      RECT  126000.0 1040250.0 127200.0 1039050.0 ;
      RECT  130800.0 1030350.0 132000.0 1029150.0 ;
      RECT  130800.0 1040250.0 132000.0 1039050.0 ;
      RECT  126600.0 1035600.0 127800.0 1034400.0 ;
      RECT  126600.0 1035600.0 127800.0 1034400.0 ;
      RECT  129150.0 1035450.0 130050.0 1034550.0 ;
      RECT  124200.0 1028250.0 133800.0 1027350.0 ;
      RECT  124200.0 1042050.0 133800.0 1041150.0 ;
      RECT  135600.0 1039650.0 136800.0 1042050.0 ;
      RECT  135600.0 1030950.0 136800.0 1027350.0 ;
      RECT  140400.0 1030950.0 141600.0 1027350.0 ;
      RECT  142800.0 1029750.0 144000.0 1027800.0 ;
      RECT  142800.0 1041600.0 144000.0 1039650.0 ;
      RECT  135600.0 1030950.0 136800.0 1029750.0 ;
      RECT  138000.0 1030950.0 139200.0 1029750.0 ;
      RECT  138000.0 1030950.0 139200.0 1029750.0 ;
      RECT  135600.0 1030950.0 136800.0 1029750.0 ;
      RECT  138000.0 1030950.0 139200.0 1029750.0 ;
      RECT  140400.0 1030950.0 141600.0 1029750.0 ;
      RECT  140400.0 1030950.0 141600.0 1029750.0 ;
      RECT  138000.0 1030950.0 139200.0 1029750.0 ;
      RECT  135600.0 1039650.0 136800.0 1038450.0 ;
      RECT  138000.0 1039650.0 139200.0 1038450.0 ;
      RECT  138000.0 1039650.0 139200.0 1038450.0 ;
      RECT  135600.0 1039650.0 136800.0 1038450.0 ;
      RECT  138000.0 1039650.0 139200.0 1038450.0 ;
      RECT  140400.0 1039650.0 141600.0 1038450.0 ;
      RECT  140400.0 1039650.0 141600.0 1038450.0 ;
      RECT  138000.0 1039650.0 139200.0 1038450.0 ;
      RECT  142800.0 1030350.0 144000.0 1029150.0 ;
      RECT  142800.0 1040250.0 144000.0 1039050.0 ;
      RECT  140400.0 1037100.0 139200.0 1035900.0 ;
      RECT  137400.0 1034400.0 136200.0 1033200.0 ;
      RECT  138000.0 1030950.0 139200.0 1029750.0 ;
      RECT  140400.0 1039650.0 141600.0 1038450.0 ;
      RECT  141600.0 1034400.0 140400.0 1033200.0 ;
      RECT  136200.0 1034400.0 137400.0 1033200.0 ;
      RECT  139200.0 1037100.0 140400.0 1035900.0 ;
      RECT  140400.0 1034400.0 141600.0 1033200.0 ;
      RECT  133800.0 1028250.0 148200.0 1027350.0 ;
      RECT  133800.0 1042050.0 148200.0 1041150.0 ;
      RECT  154800.0 1029750.0 156000.0 1027800.0 ;
      RECT  154800.0 1041600.0 156000.0 1039650.0 ;
      RECT  150000.0 1040250.0 151200.0 1042050.0 ;
      RECT  150000.0 1030950.0 151200.0 1027350.0 ;
      RECT  152700.0 1040250.0 153600.0 1030950.0 ;
      RECT  150000.0 1030950.0 151200.0 1029750.0 ;
      RECT  152400.0 1030950.0 153600.0 1029750.0 ;
      RECT  152400.0 1030950.0 153600.0 1029750.0 ;
      RECT  150000.0 1030950.0 151200.0 1029750.0 ;
      RECT  150000.0 1040250.0 151200.0 1039050.0 ;
      RECT  152400.0 1040250.0 153600.0 1039050.0 ;
      RECT  152400.0 1040250.0 153600.0 1039050.0 ;
      RECT  150000.0 1040250.0 151200.0 1039050.0 ;
      RECT  154800.0 1030350.0 156000.0 1029150.0 ;
      RECT  154800.0 1040250.0 156000.0 1039050.0 ;
      RECT  150600.0 1035600.0 151800.0 1034400.0 ;
      RECT  150600.0 1035600.0 151800.0 1034400.0 ;
      RECT  153150.0 1035450.0 154050.0 1034550.0 ;
      RECT  148200.0 1028250.0 157800.0 1027350.0 ;
      RECT  148200.0 1042050.0 157800.0 1041150.0 ;
      RECT  120450.0 1034400.0 121650.0 1035600.0 ;
      RECT  122400.0 1036800.0 123600.0 1038000.0 ;
      RECT  139200.0 1035900.0 138000.0 1037100.0 ;
      RECT  130800.0 1053450.0 132000.0 1055400.0 ;
      RECT  130800.0 1041600.0 132000.0 1043550.0 ;
      RECT  126000.0 1042950.0 127200.0 1041150.0 ;
      RECT  126000.0 1052250.0 127200.0 1055850.0 ;
      RECT  128700.0 1042950.0 129600.0 1052250.0 ;
      RECT  126000.0 1052250.0 127200.0 1053450.0 ;
      RECT  128400.0 1052250.0 129600.0 1053450.0 ;
      RECT  128400.0 1052250.0 129600.0 1053450.0 ;
      RECT  126000.0 1052250.0 127200.0 1053450.0 ;
      RECT  126000.0 1042950.0 127200.0 1044150.0 ;
      RECT  128400.0 1042950.0 129600.0 1044150.0 ;
      RECT  128400.0 1042950.0 129600.0 1044150.0 ;
      RECT  126000.0 1042950.0 127200.0 1044150.0 ;
      RECT  130800.0 1052850.0 132000.0 1054050.0 ;
      RECT  130800.0 1042950.0 132000.0 1044150.0 ;
      RECT  126600.0 1047600.0 127800.0 1048800.0 ;
      RECT  126600.0 1047600.0 127800.0 1048800.0 ;
      RECT  129150.0 1047750.0 130050.0 1048650.0 ;
      RECT  124200.0 1054950.0 133800.0 1055850.0 ;
      RECT  124200.0 1041150.0 133800.0 1042050.0 ;
      RECT  135600.0 1043550.0 136800.0 1041150.0 ;
      RECT  135600.0 1052250.0 136800.0 1055850.0 ;
      RECT  140400.0 1052250.0 141600.0 1055850.0 ;
      RECT  142800.0 1053450.0 144000.0 1055400.0 ;
      RECT  142800.0 1041600.0 144000.0 1043550.0 ;
      RECT  135600.0 1052250.0 136800.0 1053450.0 ;
      RECT  138000.0 1052250.0 139200.0 1053450.0 ;
      RECT  138000.0 1052250.0 139200.0 1053450.0 ;
      RECT  135600.0 1052250.0 136800.0 1053450.0 ;
      RECT  138000.0 1052250.0 139200.0 1053450.0 ;
      RECT  140400.0 1052250.0 141600.0 1053450.0 ;
      RECT  140400.0 1052250.0 141600.0 1053450.0 ;
      RECT  138000.0 1052250.0 139200.0 1053450.0 ;
      RECT  135600.0 1043550.0 136800.0 1044750.0 ;
      RECT  138000.0 1043550.0 139200.0 1044750.0 ;
      RECT  138000.0 1043550.0 139200.0 1044750.0 ;
      RECT  135600.0 1043550.0 136800.0 1044750.0 ;
      RECT  138000.0 1043550.0 139200.0 1044750.0 ;
      RECT  140400.0 1043550.0 141600.0 1044750.0 ;
      RECT  140400.0 1043550.0 141600.0 1044750.0 ;
      RECT  138000.0 1043550.0 139200.0 1044750.0 ;
      RECT  142800.0 1052850.0 144000.0 1054050.0 ;
      RECT  142800.0 1042950.0 144000.0 1044150.0 ;
      RECT  140400.0 1046100.0 139200.0 1047300.0 ;
      RECT  137400.0 1048800.0 136200.0 1050000.0 ;
      RECT  138000.0 1052250.0 139200.0 1053450.0 ;
      RECT  140400.0 1043550.0 141600.0 1044750.0 ;
      RECT  141600.0 1048800.0 140400.0 1050000.0 ;
      RECT  136200.0 1048800.0 137400.0 1050000.0 ;
      RECT  139200.0 1046100.0 140400.0 1047300.0 ;
      RECT  140400.0 1048800.0 141600.0 1050000.0 ;
      RECT  133800.0 1054950.0 148200.0 1055850.0 ;
      RECT  133800.0 1041150.0 148200.0 1042050.0 ;
      RECT  154800.0 1053450.0 156000.0 1055400.0 ;
      RECT  154800.0 1041600.0 156000.0 1043550.0 ;
      RECT  150000.0 1042950.0 151200.0 1041150.0 ;
      RECT  150000.0 1052250.0 151200.0 1055850.0 ;
      RECT  152700.0 1042950.0 153600.0 1052250.0 ;
      RECT  150000.0 1052250.0 151200.0 1053450.0 ;
      RECT  152400.0 1052250.0 153600.0 1053450.0 ;
      RECT  152400.0 1052250.0 153600.0 1053450.0 ;
      RECT  150000.0 1052250.0 151200.0 1053450.0 ;
      RECT  150000.0 1042950.0 151200.0 1044150.0 ;
      RECT  152400.0 1042950.0 153600.0 1044150.0 ;
      RECT  152400.0 1042950.0 153600.0 1044150.0 ;
      RECT  150000.0 1042950.0 151200.0 1044150.0 ;
      RECT  154800.0 1052850.0 156000.0 1054050.0 ;
      RECT  154800.0 1042950.0 156000.0 1044150.0 ;
      RECT  150600.0 1047600.0 151800.0 1048800.0 ;
      RECT  150600.0 1047600.0 151800.0 1048800.0 ;
      RECT  153150.0 1047750.0 154050.0 1048650.0 ;
      RECT  148200.0 1054950.0 157800.0 1055850.0 ;
      RECT  148200.0 1041150.0 157800.0 1042050.0 ;
      RECT  120450.0 1047600.0 121650.0 1048800.0 ;
      RECT  122400.0 1045200.0 123600.0 1046400.0 ;
      RECT  139200.0 1046100.0 138000.0 1047300.0 ;
      RECT  130800.0 1057350.0 132000.0 1055400.0 ;
      RECT  130800.0 1069200.0 132000.0 1067250.0 ;
      RECT  126000.0 1067850.0 127200.0 1069650.0 ;
      RECT  126000.0 1058550.0 127200.0 1054950.0 ;
      RECT  128700.0 1067850.0 129600.0 1058550.0 ;
      RECT  126000.0 1058550.0 127200.0 1057350.0 ;
      RECT  128400.0 1058550.0 129600.0 1057350.0 ;
      RECT  128400.0 1058550.0 129600.0 1057350.0 ;
      RECT  126000.0 1058550.0 127200.0 1057350.0 ;
      RECT  126000.0 1067850.0 127200.0 1066650.0 ;
      RECT  128400.0 1067850.0 129600.0 1066650.0 ;
      RECT  128400.0 1067850.0 129600.0 1066650.0 ;
      RECT  126000.0 1067850.0 127200.0 1066650.0 ;
      RECT  130800.0 1057950.0 132000.0 1056750.0 ;
      RECT  130800.0 1067850.0 132000.0 1066650.0 ;
      RECT  126600.0 1063200.0 127800.0 1062000.0 ;
      RECT  126600.0 1063200.0 127800.0 1062000.0 ;
      RECT  129150.0 1063050.0 130050.0 1062150.0 ;
      RECT  124200.0 1055850.0 133800.0 1054950.0 ;
      RECT  124200.0 1069650.0 133800.0 1068750.0 ;
      RECT  135600.0 1067250.0 136800.0 1069650.0 ;
      RECT  135600.0 1058550.0 136800.0 1054950.0 ;
      RECT  140400.0 1058550.0 141600.0 1054950.0 ;
      RECT  142800.0 1057350.0 144000.0 1055400.0 ;
      RECT  142800.0 1069200.0 144000.0 1067250.0 ;
      RECT  135600.0 1058550.0 136800.0 1057350.0 ;
      RECT  138000.0 1058550.0 139200.0 1057350.0 ;
      RECT  138000.0 1058550.0 139200.0 1057350.0 ;
      RECT  135600.0 1058550.0 136800.0 1057350.0 ;
      RECT  138000.0 1058550.0 139200.0 1057350.0 ;
      RECT  140400.0 1058550.0 141600.0 1057350.0 ;
      RECT  140400.0 1058550.0 141600.0 1057350.0 ;
      RECT  138000.0 1058550.0 139200.0 1057350.0 ;
      RECT  135600.0 1067250.0 136800.0 1066050.0 ;
      RECT  138000.0 1067250.0 139200.0 1066050.0 ;
      RECT  138000.0 1067250.0 139200.0 1066050.0 ;
      RECT  135600.0 1067250.0 136800.0 1066050.0 ;
      RECT  138000.0 1067250.0 139200.0 1066050.0 ;
      RECT  140400.0 1067250.0 141600.0 1066050.0 ;
      RECT  140400.0 1067250.0 141600.0 1066050.0 ;
      RECT  138000.0 1067250.0 139200.0 1066050.0 ;
      RECT  142800.0 1057950.0 144000.0 1056750.0 ;
      RECT  142800.0 1067850.0 144000.0 1066650.0 ;
      RECT  140400.0 1064700.0 139200.0 1063500.0 ;
      RECT  137400.0 1062000.0 136200.0 1060800.0 ;
      RECT  138000.0 1058550.0 139200.0 1057350.0 ;
      RECT  140400.0 1067250.0 141600.0 1066050.0 ;
      RECT  141600.0 1062000.0 140400.0 1060800.0 ;
      RECT  136200.0 1062000.0 137400.0 1060800.0 ;
      RECT  139200.0 1064700.0 140400.0 1063500.0 ;
      RECT  140400.0 1062000.0 141600.0 1060800.0 ;
      RECT  133800.0 1055850.0 148200.0 1054950.0 ;
      RECT  133800.0 1069650.0 148200.0 1068750.0 ;
      RECT  154800.0 1057350.0 156000.0 1055400.0 ;
      RECT  154800.0 1069200.0 156000.0 1067250.0 ;
      RECT  150000.0 1067850.0 151200.0 1069650.0 ;
      RECT  150000.0 1058550.0 151200.0 1054950.0 ;
      RECT  152700.0 1067850.0 153600.0 1058550.0 ;
      RECT  150000.0 1058550.0 151200.0 1057350.0 ;
      RECT  152400.0 1058550.0 153600.0 1057350.0 ;
      RECT  152400.0 1058550.0 153600.0 1057350.0 ;
      RECT  150000.0 1058550.0 151200.0 1057350.0 ;
      RECT  150000.0 1067850.0 151200.0 1066650.0 ;
      RECT  152400.0 1067850.0 153600.0 1066650.0 ;
      RECT  152400.0 1067850.0 153600.0 1066650.0 ;
      RECT  150000.0 1067850.0 151200.0 1066650.0 ;
      RECT  154800.0 1057950.0 156000.0 1056750.0 ;
      RECT  154800.0 1067850.0 156000.0 1066650.0 ;
      RECT  150600.0 1063200.0 151800.0 1062000.0 ;
      RECT  150600.0 1063200.0 151800.0 1062000.0 ;
      RECT  153150.0 1063050.0 154050.0 1062150.0 ;
      RECT  148200.0 1055850.0 157800.0 1054950.0 ;
      RECT  148200.0 1069650.0 157800.0 1068750.0 ;
      RECT  120450.0 1062000.0 121650.0 1063200.0 ;
      RECT  122400.0 1064400.0 123600.0 1065600.0 ;
      RECT  139200.0 1063500.0 138000.0 1064700.0 ;
      RECT  130800.0 1081050.0 132000.0 1083000.0 ;
      RECT  130800.0 1069200.0 132000.0 1071150.0 ;
      RECT  126000.0 1070550.0 127200.0 1068750.0 ;
      RECT  126000.0 1079850.0 127200.0 1083450.0 ;
      RECT  128700.0 1070550.0 129600.0 1079850.0 ;
      RECT  126000.0 1079850.0 127200.0 1081050.0 ;
      RECT  128400.0 1079850.0 129600.0 1081050.0 ;
      RECT  128400.0 1079850.0 129600.0 1081050.0 ;
      RECT  126000.0 1079850.0 127200.0 1081050.0 ;
      RECT  126000.0 1070550.0 127200.0 1071750.0 ;
      RECT  128400.0 1070550.0 129600.0 1071750.0 ;
      RECT  128400.0 1070550.0 129600.0 1071750.0 ;
      RECT  126000.0 1070550.0 127200.0 1071750.0 ;
      RECT  130800.0 1080450.0 132000.0 1081650.0 ;
      RECT  130800.0 1070550.0 132000.0 1071750.0 ;
      RECT  126600.0 1075200.0 127800.0 1076400.0 ;
      RECT  126600.0 1075200.0 127800.0 1076400.0 ;
      RECT  129150.0 1075350.0 130050.0 1076250.0 ;
      RECT  124200.0 1082550.0 133800.0 1083450.0 ;
      RECT  124200.0 1068750.0 133800.0 1069650.0 ;
      RECT  135600.0 1071150.0 136800.0 1068750.0 ;
      RECT  135600.0 1079850.0 136800.0 1083450.0 ;
      RECT  140400.0 1079850.0 141600.0 1083450.0 ;
      RECT  142800.0 1081050.0 144000.0 1083000.0 ;
      RECT  142800.0 1069200.0 144000.0 1071150.0 ;
      RECT  135600.0 1079850.0 136800.0 1081050.0 ;
      RECT  138000.0 1079850.0 139200.0 1081050.0 ;
      RECT  138000.0 1079850.0 139200.0 1081050.0 ;
      RECT  135600.0 1079850.0 136800.0 1081050.0 ;
      RECT  138000.0 1079850.0 139200.0 1081050.0 ;
      RECT  140400.0 1079850.0 141600.0 1081050.0 ;
      RECT  140400.0 1079850.0 141600.0 1081050.0 ;
      RECT  138000.0 1079850.0 139200.0 1081050.0 ;
      RECT  135600.0 1071150.0 136800.0 1072350.0 ;
      RECT  138000.0 1071150.0 139200.0 1072350.0 ;
      RECT  138000.0 1071150.0 139200.0 1072350.0 ;
      RECT  135600.0 1071150.0 136800.0 1072350.0 ;
      RECT  138000.0 1071150.0 139200.0 1072350.0 ;
      RECT  140400.0 1071150.0 141600.0 1072350.0 ;
      RECT  140400.0 1071150.0 141600.0 1072350.0 ;
      RECT  138000.0 1071150.0 139200.0 1072350.0 ;
      RECT  142800.0 1080450.0 144000.0 1081650.0 ;
      RECT  142800.0 1070550.0 144000.0 1071750.0 ;
      RECT  140400.0 1073700.0 139200.0 1074900.0 ;
      RECT  137400.0 1076400.0 136200.0 1077600.0 ;
      RECT  138000.0 1079850.0 139200.0 1081050.0 ;
      RECT  140400.0 1071150.0 141600.0 1072350.0 ;
      RECT  141600.0 1076400.0 140400.0 1077600.0 ;
      RECT  136200.0 1076400.0 137400.0 1077600.0 ;
      RECT  139200.0 1073700.0 140400.0 1074900.0 ;
      RECT  140400.0 1076400.0 141600.0 1077600.0 ;
      RECT  133800.0 1082550.0 148200.0 1083450.0 ;
      RECT  133800.0 1068750.0 148200.0 1069650.0 ;
      RECT  154800.0 1081050.0 156000.0 1083000.0 ;
      RECT  154800.0 1069200.0 156000.0 1071150.0 ;
      RECT  150000.0 1070550.0 151200.0 1068750.0 ;
      RECT  150000.0 1079850.0 151200.0 1083450.0 ;
      RECT  152700.0 1070550.0 153600.0 1079850.0 ;
      RECT  150000.0 1079850.0 151200.0 1081050.0 ;
      RECT  152400.0 1079850.0 153600.0 1081050.0 ;
      RECT  152400.0 1079850.0 153600.0 1081050.0 ;
      RECT  150000.0 1079850.0 151200.0 1081050.0 ;
      RECT  150000.0 1070550.0 151200.0 1071750.0 ;
      RECT  152400.0 1070550.0 153600.0 1071750.0 ;
      RECT  152400.0 1070550.0 153600.0 1071750.0 ;
      RECT  150000.0 1070550.0 151200.0 1071750.0 ;
      RECT  154800.0 1080450.0 156000.0 1081650.0 ;
      RECT  154800.0 1070550.0 156000.0 1071750.0 ;
      RECT  150600.0 1075200.0 151800.0 1076400.0 ;
      RECT  150600.0 1075200.0 151800.0 1076400.0 ;
      RECT  153150.0 1075350.0 154050.0 1076250.0 ;
      RECT  148200.0 1082550.0 157800.0 1083450.0 ;
      RECT  148200.0 1068750.0 157800.0 1069650.0 ;
      RECT  120450.0 1075200.0 121650.0 1076400.0 ;
      RECT  122400.0 1072800.0 123600.0 1074000.0 ;
      RECT  139200.0 1073700.0 138000.0 1074900.0 ;
      RECT  130800.0 1084950.0 132000.0 1083000.0 ;
      RECT  130800.0 1096800.0 132000.0 1094850.0 ;
      RECT  126000.0 1095450.0 127200.0 1097250.0 ;
      RECT  126000.0 1086150.0 127200.0 1082550.0 ;
      RECT  128700.0 1095450.0 129600.0 1086150.0 ;
      RECT  126000.0 1086150.0 127200.0 1084950.0 ;
      RECT  128400.0 1086150.0 129600.0 1084950.0 ;
      RECT  128400.0 1086150.0 129600.0 1084950.0 ;
      RECT  126000.0 1086150.0 127200.0 1084950.0 ;
      RECT  126000.0 1095450.0 127200.0 1094250.0 ;
      RECT  128400.0 1095450.0 129600.0 1094250.0 ;
      RECT  128400.0 1095450.0 129600.0 1094250.0 ;
      RECT  126000.0 1095450.0 127200.0 1094250.0 ;
      RECT  130800.0 1085550.0 132000.0 1084350.0 ;
      RECT  130800.0 1095450.0 132000.0 1094250.0 ;
      RECT  126600.0 1090800.0 127800.0 1089600.0 ;
      RECT  126600.0 1090800.0 127800.0 1089600.0 ;
      RECT  129150.0 1090650.0 130050.0 1089750.0 ;
      RECT  124200.0 1083450.0 133800.0 1082550.0 ;
      RECT  124200.0 1097250.0 133800.0 1096350.0 ;
      RECT  135600.0 1094850.0 136800.0 1097250.0 ;
      RECT  135600.0 1086150.0 136800.0 1082550.0 ;
      RECT  140400.0 1086150.0 141600.0 1082550.0 ;
      RECT  142800.0 1084950.0 144000.0 1083000.0 ;
      RECT  142800.0 1096800.0 144000.0 1094850.0 ;
      RECT  135600.0 1086150.0 136800.0 1084950.0 ;
      RECT  138000.0 1086150.0 139200.0 1084950.0 ;
      RECT  138000.0 1086150.0 139200.0 1084950.0 ;
      RECT  135600.0 1086150.0 136800.0 1084950.0 ;
      RECT  138000.0 1086150.0 139200.0 1084950.0 ;
      RECT  140400.0 1086150.0 141600.0 1084950.0 ;
      RECT  140400.0 1086150.0 141600.0 1084950.0 ;
      RECT  138000.0 1086150.0 139200.0 1084950.0 ;
      RECT  135600.0 1094850.0 136800.0 1093650.0 ;
      RECT  138000.0 1094850.0 139200.0 1093650.0 ;
      RECT  138000.0 1094850.0 139200.0 1093650.0 ;
      RECT  135600.0 1094850.0 136800.0 1093650.0 ;
      RECT  138000.0 1094850.0 139200.0 1093650.0 ;
      RECT  140400.0 1094850.0 141600.0 1093650.0 ;
      RECT  140400.0 1094850.0 141600.0 1093650.0 ;
      RECT  138000.0 1094850.0 139200.0 1093650.0 ;
      RECT  142800.0 1085550.0 144000.0 1084350.0 ;
      RECT  142800.0 1095450.0 144000.0 1094250.0 ;
      RECT  140400.0 1092300.0 139200.0 1091100.0 ;
      RECT  137400.0 1089600.0 136200.0 1088400.0 ;
      RECT  138000.0 1086150.0 139200.0 1084950.0 ;
      RECT  140400.0 1094850.0 141600.0 1093650.0 ;
      RECT  141600.0 1089600.0 140400.0 1088400.0 ;
      RECT  136200.0 1089600.0 137400.0 1088400.0 ;
      RECT  139200.0 1092300.0 140400.0 1091100.0 ;
      RECT  140400.0 1089600.0 141600.0 1088400.0 ;
      RECT  133800.0 1083450.0 148200.0 1082550.0 ;
      RECT  133800.0 1097250.0 148200.0 1096350.0 ;
      RECT  154800.0 1084950.0 156000.0 1083000.0 ;
      RECT  154800.0 1096800.0 156000.0 1094850.0 ;
      RECT  150000.0 1095450.0 151200.0 1097250.0 ;
      RECT  150000.0 1086150.0 151200.0 1082550.0 ;
      RECT  152700.0 1095450.0 153600.0 1086150.0 ;
      RECT  150000.0 1086150.0 151200.0 1084950.0 ;
      RECT  152400.0 1086150.0 153600.0 1084950.0 ;
      RECT  152400.0 1086150.0 153600.0 1084950.0 ;
      RECT  150000.0 1086150.0 151200.0 1084950.0 ;
      RECT  150000.0 1095450.0 151200.0 1094250.0 ;
      RECT  152400.0 1095450.0 153600.0 1094250.0 ;
      RECT  152400.0 1095450.0 153600.0 1094250.0 ;
      RECT  150000.0 1095450.0 151200.0 1094250.0 ;
      RECT  154800.0 1085550.0 156000.0 1084350.0 ;
      RECT  154800.0 1095450.0 156000.0 1094250.0 ;
      RECT  150600.0 1090800.0 151800.0 1089600.0 ;
      RECT  150600.0 1090800.0 151800.0 1089600.0 ;
      RECT  153150.0 1090650.0 154050.0 1089750.0 ;
      RECT  148200.0 1083450.0 157800.0 1082550.0 ;
      RECT  148200.0 1097250.0 157800.0 1096350.0 ;
      RECT  120450.0 1089600.0 121650.0 1090800.0 ;
      RECT  122400.0 1092000.0 123600.0 1093200.0 ;
      RECT  139200.0 1091100.0 138000.0 1092300.0 ;
      RECT  130800.0 1108650.0 132000.0 1110600.0 ;
      RECT  130800.0 1096800.0 132000.0 1098750.0 ;
      RECT  126000.0 1098150.0 127200.0 1096350.0 ;
      RECT  126000.0 1107450.0 127200.0 1111050.0 ;
      RECT  128700.0 1098150.0 129600.0 1107450.0 ;
      RECT  126000.0 1107450.0 127200.0 1108650.0 ;
      RECT  128400.0 1107450.0 129600.0 1108650.0 ;
      RECT  128400.0 1107450.0 129600.0 1108650.0 ;
      RECT  126000.0 1107450.0 127200.0 1108650.0 ;
      RECT  126000.0 1098150.0 127200.0 1099350.0 ;
      RECT  128400.0 1098150.0 129600.0 1099350.0 ;
      RECT  128400.0 1098150.0 129600.0 1099350.0 ;
      RECT  126000.0 1098150.0 127200.0 1099350.0 ;
      RECT  130800.0 1108050.0 132000.0 1109250.0 ;
      RECT  130800.0 1098150.0 132000.0 1099350.0 ;
      RECT  126600.0 1102800.0 127800.0 1104000.0 ;
      RECT  126600.0 1102800.0 127800.0 1104000.0 ;
      RECT  129150.0 1102950.0 130050.0 1103850.0 ;
      RECT  124200.0 1110150.0 133800.0 1111050.0 ;
      RECT  124200.0 1096350.0 133800.0 1097250.0 ;
      RECT  135600.0 1098750.0 136800.0 1096350.0 ;
      RECT  135600.0 1107450.0 136800.0 1111050.0 ;
      RECT  140400.0 1107450.0 141600.0 1111050.0 ;
      RECT  142800.0 1108650.0 144000.0 1110600.0 ;
      RECT  142800.0 1096800.0 144000.0 1098750.0 ;
      RECT  135600.0 1107450.0 136800.0 1108650.0 ;
      RECT  138000.0 1107450.0 139200.0 1108650.0 ;
      RECT  138000.0 1107450.0 139200.0 1108650.0 ;
      RECT  135600.0 1107450.0 136800.0 1108650.0 ;
      RECT  138000.0 1107450.0 139200.0 1108650.0 ;
      RECT  140400.0 1107450.0 141600.0 1108650.0 ;
      RECT  140400.0 1107450.0 141600.0 1108650.0 ;
      RECT  138000.0 1107450.0 139200.0 1108650.0 ;
      RECT  135600.0 1098750.0 136800.0 1099950.0 ;
      RECT  138000.0 1098750.0 139200.0 1099950.0 ;
      RECT  138000.0 1098750.0 139200.0 1099950.0 ;
      RECT  135600.0 1098750.0 136800.0 1099950.0 ;
      RECT  138000.0 1098750.0 139200.0 1099950.0 ;
      RECT  140400.0 1098750.0 141600.0 1099950.0 ;
      RECT  140400.0 1098750.0 141600.0 1099950.0 ;
      RECT  138000.0 1098750.0 139200.0 1099950.0 ;
      RECT  142800.0 1108050.0 144000.0 1109250.0 ;
      RECT  142800.0 1098150.0 144000.0 1099350.0 ;
      RECT  140400.0 1101300.0 139200.0 1102500.0 ;
      RECT  137400.0 1104000.0 136200.0 1105200.0 ;
      RECT  138000.0 1107450.0 139200.0 1108650.0 ;
      RECT  140400.0 1098750.0 141600.0 1099950.0 ;
      RECT  141600.0 1104000.0 140400.0 1105200.0 ;
      RECT  136200.0 1104000.0 137400.0 1105200.0 ;
      RECT  139200.0 1101300.0 140400.0 1102500.0 ;
      RECT  140400.0 1104000.0 141600.0 1105200.0 ;
      RECT  133800.0 1110150.0 148200.0 1111050.0 ;
      RECT  133800.0 1096350.0 148200.0 1097250.0 ;
      RECT  154800.0 1108650.0 156000.0 1110600.0 ;
      RECT  154800.0 1096800.0 156000.0 1098750.0 ;
      RECT  150000.0 1098150.0 151200.0 1096350.0 ;
      RECT  150000.0 1107450.0 151200.0 1111050.0 ;
      RECT  152700.0 1098150.0 153600.0 1107450.0 ;
      RECT  150000.0 1107450.0 151200.0 1108650.0 ;
      RECT  152400.0 1107450.0 153600.0 1108650.0 ;
      RECT  152400.0 1107450.0 153600.0 1108650.0 ;
      RECT  150000.0 1107450.0 151200.0 1108650.0 ;
      RECT  150000.0 1098150.0 151200.0 1099350.0 ;
      RECT  152400.0 1098150.0 153600.0 1099350.0 ;
      RECT  152400.0 1098150.0 153600.0 1099350.0 ;
      RECT  150000.0 1098150.0 151200.0 1099350.0 ;
      RECT  154800.0 1108050.0 156000.0 1109250.0 ;
      RECT  154800.0 1098150.0 156000.0 1099350.0 ;
      RECT  150600.0 1102800.0 151800.0 1104000.0 ;
      RECT  150600.0 1102800.0 151800.0 1104000.0 ;
      RECT  153150.0 1102950.0 154050.0 1103850.0 ;
      RECT  148200.0 1110150.0 157800.0 1111050.0 ;
      RECT  148200.0 1096350.0 157800.0 1097250.0 ;
      RECT  120450.0 1102800.0 121650.0 1104000.0 ;
      RECT  122400.0 1100400.0 123600.0 1101600.0 ;
      RECT  139200.0 1101300.0 138000.0 1102500.0 ;
      RECT  130800.0 1112550.0 132000.0 1110600.0 ;
      RECT  130800.0 1124400.0 132000.0 1122450.0 ;
      RECT  126000.0 1123050.0 127200.0 1124850.0 ;
      RECT  126000.0 1113750.0 127200.0 1110150.0 ;
      RECT  128700.0 1123050.0 129600.0 1113750.0 ;
      RECT  126000.0 1113750.0 127200.0 1112550.0 ;
      RECT  128400.0 1113750.0 129600.0 1112550.0 ;
      RECT  128400.0 1113750.0 129600.0 1112550.0 ;
      RECT  126000.0 1113750.0 127200.0 1112550.0 ;
      RECT  126000.0 1123050.0 127200.0 1121850.0 ;
      RECT  128400.0 1123050.0 129600.0 1121850.0 ;
      RECT  128400.0 1123050.0 129600.0 1121850.0 ;
      RECT  126000.0 1123050.0 127200.0 1121850.0 ;
      RECT  130800.0 1113150.0 132000.0 1111950.0 ;
      RECT  130800.0 1123050.0 132000.0 1121850.0 ;
      RECT  126600.0 1118400.0 127800.0 1117200.0 ;
      RECT  126600.0 1118400.0 127800.0 1117200.0 ;
      RECT  129150.0 1118250.0 130050.0 1117350.0 ;
      RECT  124200.0 1111050.0 133800.0 1110150.0 ;
      RECT  124200.0 1124850.0 133800.0 1123950.0 ;
      RECT  135600.0 1122450.0 136800.0 1124850.0 ;
      RECT  135600.0 1113750.0 136800.0 1110150.0 ;
      RECT  140400.0 1113750.0 141600.0 1110150.0 ;
      RECT  142800.0 1112550.0 144000.0 1110600.0 ;
      RECT  142800.0 1124400.0 144000.0 1122450.0 ;
      RECT  135600.0 1113750.0 136800.0 1112550.0 ;
      RECT  138000.0 1113750.0 139200.0 1112550.0 ;
      RECT  138000.0 1113750.0 139200.0 1112550.0 ;
      RECT  135600.0 1113750.0 136800.0 1112550.0 ;
      RECT  138000.0 1113750.0 139200.0 1112550.0 ;
      RECT  140400.0 1113750.0 141600.0 1112550.0 ;
      RECT  140400.0 1113750.0 141600.0 1112550.0 ;
      RECT  138000.0 1113750.0 139200.0 1112550.0 ;
      RECT  135600.0 1122450.0 136800.0 1121250.0 ;
      RECT  138000.0 1122450.0 139200.0 1121250.0 ;
      RECT  138000.0 1122450.0 139200.0 1121250.0 ;
      RECT  135600.0 1122450.0 136800.0 1121250.0 ;
      RECT  138000.0 1122450.0 139200.0 1121250.0 ;
      RECT  140400.0 1122450.0 141600.0 1121250.0 ;
      RECT  140400.0 1122450.0 141600.0 1121250.0 ;
      RECT  138000.0 1122450.0 139200.0 1121250.0 ;
      RECT  142800.0 1113150.0 144000.0 1111950.0 ;
      RECT  142800.0 1123050.0 144000.0 1121850.0 ;
      RECT  140400.0 1119900.0 139200.0 1118700.0 ;
      RECT  137400.0 1117200.0 136200.0 1116000.0 ;
      RECT  138000.0 1113750.0 139200.0 1112550.0 ;
      RECT  140400.0 1122450.0 141600.0 1121250.0 ;
      RECT  141600.0 1117200.0 140400.0 1116000.0 ;
      RECT  136200.0 1117200.0 137400.0 1116000.0 ;
      RECT  139200.0 1119900.0 140400.0 1118700.0 ;
      RECT  140400.0 1117200.0 141600.0 1116000.0 ;
      RECT  133800.0 1111050.0 148200.0 1110150.0 ;
      RECT  133800.0 1124850.0 148200.0 1123950.0 ;
      RECT  154800.0 1112550.0 156000.0 1110600.0 ;
      RECT  154800.0 1124400.0 156000.0 1122450.0 ;
      RECT  150000.0 1123050.0 151200.0 1124850.0 ;
      RECT  150000.0 1113750.0 151200.0 1110150.0 ;
      RECT  152700.0 1123050.0 153600.0 1113750.0 ;
      RECT  150000.0 1113750.0 151200.0 1112550.0 ;
      RECT  152400.0 1113750.0 153600.0 1112550.0 ;
      RECT  152400.0 1113750.0 153600.0 1112550.0 ;
      RECT  150000.0 1113750.0 151200.0 1112550.0 ;
      RECT  150000.0 1123050.0 151200.0 1121850.0 ;
      RECT  152400.0 1123050.0 153600.0 1121850.0 ;
      RECT  152400.0 1123050.0 153600.0 1121850.0 ;
      RECT  150000.0 1123050.0 151200.0 1121850.0 ;
      RECT  154800.0 1113150.0 156000.0 1111950.0 ;
      RECT  154800.0 1123050.0 156000.0 1121850.0 ;
      RECT  150600.0 1118400.0 151800.0 1117200.0 ;
      RECT  150600.0 1118400.0 151800.0 1117200.0 ;
      RECT  153150.0 1118250.0 154050.0 1117350.0 ;
      RECT  148200.0 1111050.0 157800.0 1110150.0 ;
      RECT  148200.0 1124850.0 157800.0 1123950.0 ;
      RECT  120450.0 1117200.0 121650.0 1118400.0 ;
      RECT  122400.0 1119600.0 123600.0 1120800.0 ;
      RECT  139200.0 1118700.0 138000.0 1119900.0 ;
      RECT  130800.0 1136250.0 132000.0 1138200.0 ;
      RECT  130800.0 1124400.0 132000.0 1126350.0 ;
      RECT  126000.0 1125750.0 127200.0 1123950.0 ;
      RECT  126000.0 1135050.0 127200.0 1138650.0 ;
      RECT  128700.0 1125750.0 129600.0 1135050.0 ;
      RECT  126000.0 1135050.0 127200.0 1136250.0 ;
      RECT  128400.0 1135050.0 129600.0 1136250.0 ;
      RECT  128400.0 1135050.0 129600.0 1136250.0 ;
      RECT  126000.0 1135050.0 127200.0 1136250.0 ;
      RECT  126000.0 1125750.0 127200.0 1126950.0 ;
      RECT  128400.0 1125750.0 129600.0 1126950.0 ;
      RECT  128400.0 1125750.0 129600.0 1126950.0 ;
      RECT  126000.0 1125750.0 127200.0 1126950.0 ;
      RECT  130800.0 1135650.0 132000.0 1136850.0 ;
      RECT  130800.0 1125750.0 132000.0 1126950.0 ;
      RECT  126600.0 1130400.0 127800.0 1131600.0 ;
      RECT  126600.0 1130400.0 127800.0 1131600.0 ;
      RECT  129150.0 1130550.0 130050.0 1131450.0 ;
      RECT  124200.0 1137750.0 133800.0 1138650.0 ;
      RECT  124200.0 1123950.0 133800.0 1124850.0 ;
      RECT  135600.0 1126350.0 136800.0 1123950.0 ;
      RECT  135600.0 1135050.0 136800.0 1138650.0 ;
      RECT  140400.0 1135050.0 141600.0 1138650.0 ;
      RECT  142800.0 1136250.0 144000.0 1138200.0 ;
      RECT  142800.0 1124400.0 144000.0 1126350.0 ;
      RECT  135600.0 1135050.0 136800.0 1136250.0 ;
      RECT  138000.0 1135050.0 139200.0 1136250.0 ;
      RECT  138000.0 1135050.0 139200.0 1136250.0 ;
      RECT  135600.0 1135050.0 136800.0 1136250.0 ;
      RECT  138000.0 1135050.0 139200.0 1136250.0 ;
      RECT  140400.0 1135050.0 141600.0 1136250.0 ;
      RECT  140400.0 1135050.0 141600.0 1136250.0 ;
      RECT  138000.0 1135050.0 139200.0 1136250.0 ;
      RECT  135600.0 1126350.0 136800.0 1127550.0 ;
      RECT  138000.0 1126350.0 139200.0 1127550.0 ;
      RECT  138000.0 1126350.0 139200.0 1127550.0 ;
      RECT  135600.0 1126350.0 136800.0 1127550.0 ;
      RECT  138000.0 1126350.0 139200.0 1127550.0 ;
      RECT  140400.0 1126350.0 141600.0 1127550.0 ;
      RECT  140400.0 1126350.0 141600.0 1127550.0 ;
      RECT  138000.0 1126350.0 139200.0 1127550.0 ;
      RECT  142800.0 1135650.0 144000.0 1136850.0 ;
      RECT  142800.0 1125750.0 144000.0 1126950.0 ;
      RECT  140400.0 1128900.0 139200.0 1130100.0 ;
      RECT  137400.0 1131600.0 136200.0 1132800.0 ;
      RECT  138000.0 1135050.0 139200.0 1136250.0 ;
      RECT  140400.0 1126350.0 141600.0 1127550.0 ;
      RECT  141600.0 1131600.0 140400.0 1132800.0 ;
      RECT  136200.0 1131600.0 137400.0 1132800.0 ;
      RECT  139200.0 1128900.0 140400.0 1130100.0 ;
      RECT  140400.0 1131600.0 141600.0 1132800.0 ;
      RECT  133800.0 1137750.0 148200.0 1138650.0 ;
      RECT  133800.0 1123950.0 148200.0 1124850.0 ;
      RECT  154800.0 1136250.0 156000.0 1138200.0 ;
      RECT  154800.0 1124400.0 156000.0 1126350.0 ;
      RECT  150000.0 1125750.0 151200.0 1123950.0 ;
      RECT  150000.0 1135050.0 151200.0 1138650.0 ;
      RECT  152700.0 1125750.0 153600.0 1135050.0 ;
      RECT  150000.0 1135050.0 151200.0 1136250.0 ;
      RECT  152400.0 1135050.0 153600.0 1136250.0 ;
      RECT  152400.0 1135050.0 153600.0 1136250.0 ;
      RECT  150000.0 1135050.0 151200.0 1136250.0 ;
      RECT  150000.0 1125750.0 151200.0 1126950.0 ;
      RECT  152400.0 1125750.0 153600.0 1126950.0 ;
      RECT  152400.0 1125750.0 153600.0 1126950.0 ;
      RECT  150000.0 1125750.0 151200.0 1126950.0 ;
      RECT  154800.0 1135650.0 156000.0 1136850.0 ;
      RECT  154800.0 1125750.0 156000.0 1126950.0 ;
      RECT  150600.0 1130400.0 151800.0 1131600.0 ;
      RECT  150600.0 1130400.0 151800.0 1131600.0 ;
      RECT  153150.0 1130550.0 154050.0 1131450.0 ;
      RECT  148200.0 1137750.0 157800.0 1138650.0 ;
      RECT  148200.0 1123950.0 157800.0 1124850.0 ;
      RECT  120450.0 1130400.0 121650.0 1131600.0 ;
      RECT  122400.0 1128000.0 123600.0 1129200.0 ;
      RECT  139200.0 1128900.0 138000.0 1130100.0 ;
      RECT  130800.0 1140150.0 132000.0 1138200.0 ;
      RECT  130800.0 1152000.0 132000.0 1150050.0 ;
      RECT  126000.0 1150650.0 127200.0 1152450.0 ;
      RECT  126000.0 1141350.0 127200.0 1137750.0 ;
      RECT  128700.0 1150650.0 129600.0 1141350.0 ;
      RECT  126000.0 1141350.0 127200.0 1140150.0 ;
      RECT  128400.0 1141350.0 129600.0 1140150.0 ;
      RECT  128400.0 1141350.0 129600.0 1140150.0 ;
      RECT  126000.0 1141350.0 127200.0 1140150.0 ;
      RECT  126000.0 1150650.0 127200.0 1149450.0 ;
      RECT  128400.0 1150650.0 129600.0 1149450.0 ;
      RECT  128400.0 1150650.0 129600.0 1149450.0 ;
      RECT  126000.0 1150650.0 127200.0 1149450.0 ;
      RECT  130800.0 1140750.0 132000.0 1139550.0 ;
      RECT  130800.0 1150650.0 132000.0 1149450.0 ;
      RECT  126600.0 1146000.0 127800.0 1144800.0 ;
      RECT  126600.0 1146000.0 127800.0 1144800.0 ;
      RECT  129150.0 1145850.0 130050.0 1144950.0 ;
      RECT  124200.0 1138650.0 133800.0 1137750.0 ;
      RECT  124200.0 1152450.0 133800.0 1151550.0 ;
      RECT  135600.0 1150050.0 136800.0 1152450.0 ;
      RECT  135600.0 1141350.0 136800.0 1137750.0 ;
      RECT  140400.0 1141350.0 141600.0 1137750.0 ;
      RECT  142800.0 1140150.0 144000.0 1138200.0 ;
      RECT  142800.0 1152000.0 144000.0 1150050.0 ;
      RECT  135600.0 1141350.0 136800.0 1140150.0 ;
      RECT  138000.0 1141350.0 139200.0 1140150.0 ;
      RECT  138000.0 1141350.0 139200.0 1140150.0 ;
      RECT  135600.0 1141350.0 136800.0 1140150.0 ;
      RECT  138000.0 1141350.0 139200.0 1140150.0 ;
      RECT  140400.0 1141350.0 141600.0 1140150.0 ;
      RECT  140400.0 1141350.0 141600.0 1140150.0 ;
      RECT  138000.0 1141350.0 139200.0 1140150.0 ;
      RECT  135600.0 1150050.0 136800.0 1148850.0 ;
      RECT  138000.0 1150050.0 139200.0 1148850.0 ;
      RECT  138000.0 1150050.0 139200.0 1148850.0 ;
      RECT  135600.0 1150050.0 136800.0 1148850.0 ;
      RECT  138000.0 1150050.0 139200.0 1148850.0 ;
      RECT  140400.0 1150050.0 141600.0 1148850.0 ;
      RECT  140400.0 1150050.0 141600.0 1148850.0 ;
      RECT  138000.0 1150050.0 139200.0 1148850.0 ;
      RECT  142800.0 1140750.0 144000.0 1139550.0 ;
      RECT  142800.0 1150650.0 144000.0 1149450.0 ;
      RECT  140400.0 1147500.0 139200.0 1146300.0 ;
      RECT  137400.0 1144800.0 136200.0 1143600.0 ;
      RECT  138000.0 1141350.0 139200.0 1140150.0 ;
      RECT  140400.0 1150050.0 141600.0 1148850.0 ;
      RECT  141600.0 1144800.0 140400.0 1143600.0 ;
      RECT  136200.0 1144800.0 137400.0 1143600.0 ;
      RECT  139200.0 1147500.0 140400.0 1146300.0 ;
      RECT  140400.0 1144800.0 141600.0 1143600.0 ;
      RECT  133800.0 1138650.0 148200.0 1137750.0 ;
      RECT  133800.0 1152450.0 148200.0 1151550.0 ;
      RECT  154800.0 1140150.0 156000.0 1138200.0 ;
      RECT  154800.0 1152000.0 156000.0 1150050.0 ;
      RECT  150000.0 1150650.0 151200.0 1152450.0 ;
      RECT  150000.0 1141350.0 151200.0 1137750.0 ;
      RECT  152700.0 1150650.0 153600.0 1141350.0 ;
      RECT  150000.0 1141350.0 151200.0 1140150.0 ;
      RECT  152400.0 1141350.0 153600.0 1140150.0 ;
      RECT  152400.0 1141350.0 153600.0 1140150.0 ;
      RECT  150000.0 1141350.0 151200.0 1140150.0 ;
      RECT  150000.0 1150650.0 151200.0 1149450.0 ;
      RECT  152400.0 1150650.0 153600.0 1149450.0 ;
      RECT  152400.0 1150650.0 153600.0 1149450.0 ;
      RECT  150000.0 1150650.0 151200.0 1149450.0 ;
      RECT  154800.0 1140750.0 156000.0 1139550.0 ;
      RECT  154800.0 1150650.0 156000.0 1149450.0 ;
      RECT  150600.0 1146000.0 151800.0 1144800.0 ;
      RECT  150600.0 1146000.0 151800.0 1144800.0 ;
      RECT  153150.0 1145850.0 154050.0 1144950.0 ;
      RECT  148200.0 1138650.0 157800.0 1137750.0 ;
      RECT  148200.0 1152450.0 157800.0 1151550.0 ;
      RECT  120450.0 1144800.0 121650.0 1146000.0 ;
      RECT  122400.0 1147200.0 123600.0 1148400.0 ;
      RECT  139200.0 1146300.0 138000.0 1147500.0 ;
      RECT  130800.0 1163850.0 132000.0 1165800.0 ;
      RECT  130800.0 1152000.0 132000.0 1153950.0 ;
      RECT  126000.0 1153350.0 127200.0 1151550.0 ;
      RECT  126000.0 1162650.0 127200.0 1166250.0 ;
      RECT  128700.0 1153350.0 129600.0 1162650.0 ;
      RECT  126000.0 1162650.0 127200.0 1163850.0 ;
      RECT  128400.0 1162650.0 129600.0 1163850.0 ;
      RECT  128400.0 1162650.0 129600.0 1163850.0 ;
      RECT  126000.0 1162650.0 127200.0 1163850.0 ;
      RECT  126000.0 1153350.0 127200.0 1154550.0 ;
      RECT  128400.0 1153350.0 129600.0 1154550.0 ;
      RECT  128400.0 1153350.0 129600.0 1154550.0 ;
      RECT  126000.0 1153350.0 127200.0 1154550.0 ;
      RECT  130800.0 1163250.0 132000.0 1164450.0 ;
      RECT  130800.0 1153350.0 132000.0 1154550.0 ;
      RECT  126600.0 1158000.0 127800.0 1159200.0 ;
      RECT  126600.0 1158000.0 127800.0 1159200.0 ;
      RECT  129150.0 1158150.0 130050.0 1159050.0 ;
      RECT  124200.0 1165350.0 133800.0 1166250.0 ;
      RECT  124200.0 1151550.0 133800.0 1152450.0 ;
      RECT  135600.0 1153950.0 136800.0 1151550.0 ;
      RECT  135600.0 1162650.0 136800.0 1166250.0 ;
      RECT  140400.0 1162650.0 141600.0 1166250.0 ;
      RECT  142800.0 1163850.0 144000.0 1165800.0 ;
      RECT  142800.0 1152000.0 144000.0 1153950.0 ;
      RECT  135600.0 1162650.0 136800.0 1163850.0 ;
      RECT  138000.0 1162650.0 139200.0 1163850.0 ;
      RECT  138000.0 1162650.0 139200.0 1163850.0 ;
      RECT  135600.0 1162650.0 136800.0 1163850.0 ;
      RECT  138000.0 1162650.0 139200.0 1163850.0 ;
      RECT  140400.0 1162650.0 141600.0 1163850.0 ;
      RECT  140400.0 1162650.0 141600.0 1163850.0 ;
      RECT  138000.0 1162650.0 139200.0 1163850.0 ;
      RECT  135600.0 1153950.0 136800.0 1155150.0 ;
      RECT  138000.0 1153950.0 139200.0 1155150.0 ;
      RECT  138000.0 1153950.0 139200.0 1155150.0 ;
      RECT  135600.0 1153950.0 136800.0 1155150.0 ;
      RECT  138000.0 1153950.0 139200.0 1155150.0 ;
      RECT  140400.0 1153950.0 141600.0 1155150.0 ;
      RECT  140400.0 1153950.0 141600.0 1155150.0 ;
      RECT  138000.0 1153950.0 139200.0 1155150.0 ;
      RECT  142800.0 1163250.0 144000.0 1164450.0 ;
      RECT  142800.0 1153350.0 144000.0 1154550.0 ;
      RECT  140400.0 1156500.0 139200.0 1157700.0 ;
      RECT  137400.0 1159200.0 136200.0 1160400.0 ;
      RECT  138000.0 1162650.0 139200.0 1163850.0 ;
      RECT  140400.0 1153950.0 141600.0 1155150.0 ;
      RECT  141600.0 1159200.0 140400.0 1160400.0 ;
      RECT  136200.0 1159200.0 137400.0 1160400.0 ;
      RECT  139200.0 1156500.0 140400.0 1157700.0 ;
      RECT  140400.0 1159200.0 141600.0 1160400.0 ;
      RECT  133800.0 1165350.0 148200.0 1166250.0 ;
      RECT  133800.0 1151550.0 148200.0 1152450.0 ;
      RECT  154800.0 1163850.0 156000.0 1165800.0 ;
      RECT  154800.0 1152000.0 156000.0 1153950.0 ;
      RECT  150000.0 1153350.0 151200.0 1151550.0 ;
      RECT  150000.0 1162650.0 151200.0 1166250.0 ;
      RECT  152700.0 1153350.0 153600.0 1162650.0 ;
      RECT  150000.0 1162650.0 151200.0 1163850.0 ;
      RECT  152400.0 1162650.0 153600.0 1163850.0 ;
      RECT  152400.0 1162650.0 153600.0 1163850.0 ;
      RECT  150000.0 1162650.0 151200.0 1163850.0 ;
      RECT  150000.0 1153350.0 151200.0 1154550.0 ;
      RECT  152400.0 1153350.0 153600.0 1154550.0 ;
      RECT  152400.0 1153350.0 153600.0 1154550.0 ;
      RECT  150000.0 1153350.0 151200.0 1154550.0 ;
      RECT  154800.0 1163250.0 156000.0 1164450.0 ;
      RECT  154800.0 1153350.0 156000.0 1154550.0 ;
      RECT  150600.0 1158000.0 151800.0 1159200.0 ;
      RECT  150600.0 1158000.0 151800.0 1159200.0 ;
      RECT  153150.0 1158150.0 154050.0 1159050.0 ;
      RECT  148200.0 1165350.0 157800.0 1166250.0 ;
      RECT  148200.0 1151550.0 157800.0 1152450.0 ;
      RECT  120450.0 1158000.0 121650.0 1159200.0 ;
      RECT  122400.0 1155600.0 123600.0 1156800.0 ;
      RECT  139200.0 1156500.0 138000.0 1157700.0 ;
      RECT  130800.0 1167750.0 132000.0 1165800.0 ;
      RECT  130800.0 1179600.0 132000.0 1177650.0 ;
      RECT  126000.0 1178250.0 127200.0 1180050.0 ;
      RECT  126000.0 1168950.0 127200.0 1165350.0 ;
      RECT  128700.0 1178250.0 129600.0 1168950.0 ;
      RECT  126000.0 1168950.0 127200.0 1167750.0 ;
      RECT  128400.0 1168950.0 129600.0 1167750.0 ;
      RECT  128400.0 1168950.0 129600.0 1167750.0 ;
      RECT  126000.0 1168950.0 127200.0 1167750.0 ;
      RECT  126000.0 1178250.0 127200.0 1177050.0 ;
      RECT  128400.0 1178250.0 129600.0 1177050.0 ;
      RECT  128400.0 1178250.0 129600.0 1177050.0 ;
      RECT  126000.0 1178250.0 127200.0 1177050.0 ;
      RECT  130800.0 1168350.0 132000.0 1167150.0 ;
      RECT  130800.0 1178250.0 132000.0 1177050.0 ;
      RECT  126600.0 1173600.0 127800.0 1172400.0 ;
      RECT  126600.0 1173600.0 127800.0 1172400.0 ;
      RECT  129150.0 1173450.0 130050.0 1172550.0 ;
      RECT  124200.0 1166250.0 133800.0 1165350.0 ;
      RECT  124200.0 1180050.0 133800.0 1179150.0 ;
      RECT  135600.0 1177650.0 136800.0 1180050.0 ;
      RECT  135600.0 1168950.0 136800.0 1165350.0 ;
      RECT  140400.0 1168950.0 141600.0 1165350.0 ;
      RECT  142800.0 1167750.0 144000.0 1165800.0 ;
      RECT  142800.0 1179600.0 144000.0 1177650.0 ;
      RECT  135600.0 1168950.0 136800.0 1167750.0 ;
      RECT  138000.0 1168950.0 139200.0 1167750.0 ;
      RECT  138000.0 1168950.0 139200.0 1167750.0 ;
      RECT  135600.0 1168950.0 136800.0 1167750.0 ;
      RECT  138000.0 1168950.0 139200.0 1167750.0 ;
      RECT  140400.0 1168950.0 141600.0 1167750.0 ;
      RECT  140400.0 1168950.0 141600.0 1167750.0 ;
      RECT  138000.0 1168950.0 139200.0 1167750.0 ;
      RECT  135600.0 1177650.0 136800.0 1176450.0 ;
      RECT  138000.0 1177650.0 139200.0 1176450.0 ;
      RECT  138000.0 1177650.0 139200.0 1176450.0 ;
      RECT  135600.0 1177650.0 136800.0 1176450.0 ;
      RECT  138000.0 1177650.0 139200.0 1176450.0 ;
      RECT  140400.0 1177650.0 141600.0 1176450.0 ;
      RECT  140400.0 1177650.0 141600.0 1176450.0 ;
      RECT  138000.0 1177650.0 139200.0 1176450.0 ;
      RECT  142800.0 1168350.0 144000.0 1167150.0 ;
      RECT  142800.0 1178250.0 144000.0 1177050.0 ;
      RECT  140400.0 1175100.0 139200.0 1173900.0 ;
      RECT  137400.0 1172400.0 136200.0 1171200.0 ;
      RECT  138000.0 1168950.0 139200.0 1167750.0 ;
      RECT  140400.0 1177650.0 141600.0 1176450.0 ;
      RECT  141600.0 1172400.0 140400.0 1171200.0 ;
      RECT  136200.0 1172400.0 137400.0 1171200.0 ;
      RECT  139200.0 1175100.0 140400.0 1173900.0 ;
      RECT  140400.0 1172400.0 141600.0 1171200.0 ;
      RECT  133800.0 1166250.0 148200.0 1165350.0 ;
      RECT  133800.0 1180050.0 148200.0 1179150.0 ;
      RECT  154800.0 1167750.0 156000.0 1165800.0 ;
      RECT  154800.0 1179600.0 156000.0 1177650.0 ;
      RECT  150000.0 1178250.0 151200.0 1180050.0 ;
      RECT  150000.0 1168950.0 151200.0 1165350.0 ;
      RECT  152700.0 1178250.0 153600.0 1168950.0 ;
      RECT  150000.0 1168950.0 151200.0 1167750.0 ;
      RECT  152400.0 1168950.0 153600.0 1167750.0 ;
      RECT  152400.0 1168950.0 153600.0 1167750.0 ;
      RECT  150000.0 1168950.0 151200.0 1167750.0 ;
      RECT  150000.0 1178250.0 151200.0 1177050.0 ;
      RECT  152400.0 1178250.0 153600.0 1177050.0 ;
      RECT  152400.0 1178250.0 153600.0 1177050.0 ;
      RECT  150000.0 1178250.0 151200.0 1177050.0 ;
      RECT  154800.0 1168350.0 156000.0 1167150.0 ;
      RECT  154800.0 1178250.0 156000.0 1177050.0 ;
      RECT  150600.0 1173600.0 151800.0 1172400.0 ;
      RECT  150600.0 1173600.0 151800.0 1172400.0 ;
      RECT  153150.0 1173450.0 154050.0 1172550.0 ;
      RECT  148200.0 1166250.0 157800.0 1165350.0 ;
      RECT  148200.0 1180050.0 157800.0 1179150.0 ;
      RECT  120450.0 1172400.0 121650.0 1173600.0 ;
      RECT  122400.0 1174800.0 123600.0 1176000.0 ;
      RECT  139200.0 1173900.0 138000.0 1175100.0 ;
      RECT  130800.0 1191450.0 132000.0 1193400.0 ;
      RECT  130800.0 1179600.0 132000.0 1181550.0 ;
      RECT  126000.0 1180950.0 127200.0 1179150.0 ;
      RECT  126000.0 1190250.0 127200.0 1193850.0 ;
      RECT  128700.0 1180950.0 129600.0 1190250.0 ;
      RECT  126000.0 1190250.0 127200.0 1191450.0 ;
      RECT  128400.0 1190250.0 129600.0 1191450.0 ;
      RECT  128400.0 1190250.0 129600.0 1191450.0 ;
      RECT  126000.0 1190250.0 127200.0 1191450.0 ;
      RECT  126000.0 1180950.0 127200.0 1182150.0 ;
      RECT  128400.0 1180950.0 129600.0 1182150.0 ;
      RECT  128400.0 1180950.0 129600.0 1182150.0 ;
      RECT  126000.0 1180950.0 127200.0 1182150.0 ;
      RECT  130800.0 1190850.0 132000.0 1192050.0 ;
      RECT  130800.0 1180950.0 132000.0 1182150.0 ;
      RECT  126600.0 1185600.0 127800.0 1186800.0 ;
      RECT  126600.0 1185600.0 127800.0 1186800.0 ;
      RECT  129150.0 1185750.0 130050.0 1186650.0 ;
      RECT  124200.0 1192950.0 133800.0 1193850.0 ;
      RECT  124200.0 1179150.0 133800.0 1180050.0 ;
      RECT  135600.0 1181550.0 136800.0 1179150.0 ;
      RECT  135600.0 1190250.0 136800.0 1193850.0 ;
      RECT  140400.0 1190250.0 141600.0 1193850.0 ;
      RECT  142800.0 1191450.0 144000.0 1193400.0 ;
      RECT  142800.0 1179600.0 144000.0 1181550.0 ;
      RECT  135600.0 1190250.0 136800.0 1191450.0 ;
      RECT  138000.0 1190250.0 139200.0 1191450.0 ;
      RECT  138000.0 1190250.0 139200.0 1191450.0 ;
      RECT  135600.0 1190250.0 136800.0 1191450.0 ;
      RECT  138000.0 1190250.0 139200.0 1191450.0 ;
      RECT  140400.0 1190250.0 141600.0 1191450.0 ;
      RECT  140400.0 1190250.0 141600.0 1191450.0 ;
      RECT  138000.0 1190250.0 139200.0 1191450.0 ;
      RECT  135600.0 1181550.0 136800.0 1182750.0 ;
      RECT  138000.0 1181550.0 139200.0 1182750.0 ;
      RECT  138000.0 1181550.0 139200.0 1182750.0 ;
      RECT  135600.0 1181550.0 136800.0 1182750.0 ;
      RECT  138000.0 1181550.0 139200.0 1182750.0 ;
      RECT  140400.0 1181550.0 141600.0 1182750.0 ;
      RECT  140400.0 1181550.0 141600.0 1182750.0 ;
      RECT  138000.0 1181550.0 139200.0 1182750.0 ;
      RECT  142800.0 1190850.0 144000.0 1192050.0 ;
      RECT  142800.0 1180950.0 144000.0 1182150.0 ;
      RECT  140400.0 1184100.0 139200.0 1185300.0 ;
      RECT  137400.0 1186800.0 136200.0 1188000.0 ;
      RECT  138000.0 1190250.0 139200.0 1191450.0 ;
      RECT  140400.0 1181550.0 141600.0 1182750.0 ;
      RECT  141600.0 1186800.0 140400.0 1188000.0 ;
      RECT  136200.0 1186800.0 137400.0 1188000.0 ;
      RECT  139200.0 1184100.0 140400.0 1185300.0 ;
      RECT  140400.0 1186800.0 141600.0 1188000.0 ;
      RECT  133800.0 1192950.0 148200.0 1193850.0 ;
      RECT  133800.0 1179150.0 148200.0 1180050.0 ;
      RECT  154800.0 1191450.0 156000.0 1193400.0 ;
      RECT  154800.0 1179600.0 156000.0 1181550.0 ;
      RECT  150000.0 1180950.0 151200.0 1179150.0 ;
      RECT  150000.0 1190250.0 151200.0 1193850.0 ;
      RECT  152700.0 1180950.0 153600.0 1190250.0 ;
      RECT  150000.0 1190250.0 151200.0 1191450.0 ;
      RECT  152400.0 1190250.0 153600.0 1191450.0 ;
      RECT  152400.0 1190250.0 153600.0 1191450.0 ;
      RECT  150000.0 1190250.0 151200.0 1191450.0 ;
      RECT  150000.0 1180950.0 151200.0 1182150.0 ;
      RECT  152400.0 1180950.0 153600.0 1182150.0 ;
      RECT  152400.0 1180950.0 153600.0 1182150.0 ;
      RECT  150000.0 1180950.0 151200.0 1182150.0 ;
      RECT  154800.0 1190850.0 156000.0 1192050.0 ;
      RECT  154800.0 1180950.0 156000.0 1182150.0 ;
      RECT  150600.0 1185600.0 151800.0 1186800.0 ;
      RECT  150600.0 1185600.0 151800.0 1186800.0 ;
      RECT  153150.0 1185750.0 154050.0 1186650.0 ;
      RECT  148200.0 1192950.0 157800.0 1193850.0 ;
      RECT  148200.0 1179150.0 157800.0 1180050.0 ;
      RECT  120450.0 1185600.0 121650.0 1186800.0 ;
      RECT  122400.0 1183200.0 123600.0 1184400.0 ;
      RECT  139200.0 1184100.0 138000.0 1185300.0 ;
      RECT  130800.0 1195350.0 132000.0 1193400.0 ;
      RECT  130800.0 1207200.0 132000.0 1205250.0 ;
      RECT  126000.0 1205850.0 127200.0 1207650.0 ;
      RECT  126000.0 1196550.0 127200.0 1192950.0 ;
      RECT  128700.0 1205850.0 129600.0 1196550.0 ;
      RECT  126000.0 1196550.0 127200.0 1195350.0 ;
      RECT  128400.0 1196550.0 129600.0 1195350.0 ;
      RECT  128400.0 1196550.0 129600.0 1195350.0 ;
      RECT  126000.0 1196550.0 127200.0 1195350.0 ;
      RECT  126000.0 1205850.0 127200.0 1204650.0 ;
      RECT  128400.0 1205850.0 129600.0 1204650.0 ;
      RECT  128400.0 1205850.0 129600.0 1204650.0 ;
      RECT  126000.0 1205850.0 127200.0 1204650.0 ;
      RECT  130800.0 1195950.0 132000.0 1194750.0 ;
      RECT  130800.0 1205850.0 132000.0 1204650.0 ;
      RECT  126600.0 1201200.0 127800.0 1200000.0 ;
      RECT  126600.0 1201200.0 127800.0 1200000.0 ;
      RECT  129150.0 1201050.0 130050.0 1200150.0 ;
      RECT  124200.0 1193850.0 133800.0 1192950.0 ;
      RECT  124200.0 1207650.0 133800.0 1206750.0 ;
      RECT  135600.0 1205250.0 136800.0 1207650.0 ;
      RECT  135600.0 1196550.0 136800.0 1192950.0 ;
      RECT  140400.0 1196550.0 141600.0 1192950.0 ;
      RECT  142800.0 1195350.0 144000.0 1193400.0 ;
      RECT  142800.0 1207200.0 144000.0 1205250.0 ;
      RECT  135600.0 1196550.0 136800.0 1195350.0 ;
      RECT  138000.0 1196550.0 139200.0 1195350.0 ;
      RECT  138000.0 1196550.0 139200.0 1195350.0 ;
      RECT  135600.0 1196550.0 136800.0 1195350.0 ;
      RECT  138000.0 1196550.0 139200.0 1195350.0 ;
      RECT  140400.0 1196550.0 141600.0 1195350.0 ;
      RECT  140400.0 1196550.0 141600.0 1195350.0 ;
      RECT  138000.0 1196550.0 139200.0 1195350.0 ;
      RECT  135600.0 1205250.0 136800.0 1204050.0 ;
      RECT  138000.0 1205250.0 139200.0 1204050.0 ;
      RECT  138000.0 1205250.0 139200.0 1204050.0 ;
      RECT  135600.0 1205250.0 136800.0 1204050.0 ;
      RECT  138000.0 1205250.0 139200.0 1204050.0 ;
      RECT  140400.0 1205250.0 141600.0 1204050.0 ;
      RECT  140400.0 1205250.0 141600.0 1204050.0 ;
      RECT  138000.0 1205250.0 139200.0 1204050.0 ;
      RECT  142800.0 1195950.0 144000.0 1194750.0 ;
      RECT  142800.0 1205850.0 144000.0 1204650.0 ;
      RECT  140400.0 1202700.0 139200.0 1201500.0 ;
      RECT  137400.0 1200000.0 136200.0 1198800.0 ;
      RECT  138000.0 1196550.0 139200.0 1195350.0 ;
      RECT  140400.0 1205250.0 141600.0 1204050.0 ;
      RECT  141600.0 1200000.0 140400.0 1198800.0 ;
      RECT  136200.0 1200000.0 137400.0 1198800.0 ;
      RECT  139200.0 1202700.0 140400.0 1201500.0 ;
      RECT  140400.0 1200000.0 141600.0 1198800.0 ;
      RECT  133800.0 1193850.0 148200.0 1192950.0 ;
      RECT  133800.0 1207650.0 148200.0 1206750.0 ;
      RECT  154800.0 1195350.0 156000.0 1193400.0 ;
      RECT  154800.0 1207200.0 156000.0 1205250.0 ;
      RECT  150000.0 1205850.0 151200.0 1207650.0 ;
      RECT  150000.0 1196550.0 151200.0 1192950.0 ;
      RECT  152700.0 1205850.0 153600.0 1196550.0 ;
      RECT  150000.0 1196550.0 151200.0 1195350.0 ;
      RECT  152400.0 1196550.0 153600.0 1195350.0 ;
      RECT  152400.0 1196550.0 153600.0 1195350.0 ;
      RECT  150000.0 1196550.0 151200.0 1195350.0 ;
      RECT  150000.0 1205850.0 151200.0 1204650.0 ;
      RECT  152400.0 1205850.0 153600.0 1204650.0 ;
      RECT  152400.0 1205850.0 153600.0 1204650.0 ;
      RECT  150000.0 1205850.0 151200.0 1204650.0 ;
      RECT  154800.0 1195950.0 156000.0 1194750.0 ;
      RECT  154800.0 1205850.0 156000.0 1204650.0 ;
      RECT  150600.0 1201200.0 151800.0 1200000.0 ;
      RECT  150600.0 1201200.0 151800.0 1200000.0 ;
      RECT  153150.0 1201050.0 154050.0 1200150.0 ;
      RECT  148200.0 1193850.0 157800.0 1192950.0 ;
      RECT  148200.0 1207650.0 157800.0 1206750.0 ;
      RECT  120450.0 1200000.0 121650.0 1201200.0 ;
      RECT  122400.0 1202400.0 123600.0 1203600.0 ;
      RECT  139200.0 1201500.0 138000.0 1202700.0 ;
      RECT  130800.0 1219050.0 132000.0 1221000.0 ;
      RECT  130800.0 1207200.0 132000.0 1209150.0 ;
      RECT  126000.0 1208550.0 127200.0 1206750.0 ;
      RECT  126000.0 1217850.0 127200.0 1221450.0 ;
      RECT  128700.0 1208550.0 129600.0 1217850.0 ;
      RECT  126000.0 1217850.0 127200.0 1219050.0 ;
      RECT  128400.0 1217850.0 129600.0 1219050.0 ;
      RECT  128400.0 1217850.0 129600.0 1219050.0 ;
      RECT  126000.0 1217850.0 127200.0 1219050.0 ;
      RECT  126000.0 1208550.0 127200.0 1209750.0 ;
      RECT  128400.0 1208550.0 129600.0 1209750.0 ;
      RECT  128400.0 1208550.0 129600.0 1209750.0 ;
      RECT  126000.0 1208550.0 127200.0 1209750.0 ;
      RECT  130800.0 1218450.0 132000.0 1219650.0 ;
      RECT  130800.0 1208550.0 132000.0 1209750.0 ;
      RECT  126600.0 1213200.0 127800.0 1214400.0 ;
      RECT  126600.0 1213200.0 127800.0 1214400.0 ;
      RECT  129150.0 1213350.0 130050.0 1214250.0 ;
      RECT  124200.0 1220550.0 133800.0 1221450.0 ;
      RECT  124200.0 1206750.0 133800.0 1207650.0 ;
      RECT  135600.0 1209150.0 136800.0 1206750.0 ;
      RECT  135600.0 1217850.0 136800.0 1221450.0 ;
      RECT  140400.0 1217850.0 141600.0 1221450.0 ;
      RECT  142800.0 1219050.0 144000.0 1221000.0 ;
      RECT  142800.0 1207200.0 144000.0 1209150.0 ;
      RECT  135600.0 1217850.0 136800.0 1219050.0 ;
      RECT  138000.0 1217850.0 139200.0 1219050.0 ;
      RECT  138000.0 1217850.0 139200.0 1219050.0 ;
      RECT  135600.0 1217850.0 136800.0 1219050.0 ;
      RECT  138000.0 1217850.0 139200.0 1219050.0 ;
      RECT  140400.0 1217850.0 141600.0 1219050.0 ;
      RECT  140400.0 1217850.0 141600.0 1219050.0 ;
      RECT  138000.0 1217850.0 139200.0 1219050.0 ;
      RECT  135600.0 1209150.0 136800.0 1210350.0 ;
      RECT  138000.0 1209150.0 139200.0 1210350.0 ;
      RECT  138000.0 1209150.0 139200.0 1210350.0 ;
      RECT  135600.0 1209150.0 136800.0 1210350.0 ;
      RECT  138000.0 1209150.0 139200.0 1210350.0 ;
      RECT  140400.0 1209150.0 141600.0 1210350.0 ;
      RECT  140400.0 1209150.0 141600.0 1210350.0 ;
      RECT  138000.0 1209150.0 139200.0 1210350.0 ;
      RECT  142800.0 1218450.0 144000.0 1219650.0 ;
      RECT  142800.0 1208550.0 144000.0 1209750.0 ;
      RECT  140400.0 1211700.0 139200.0 1212900.0 ;
      RECT  137400.0 1214400.0 136200.0 1215600.0 ;
      RECT  138000.0 1217850.0 139200.0 1219050.0 ;
      RECT  140400.0 1209150.0 141600.0 1210350.0 ;
      RECT  141600.0 1214400.0 140400.0 1215600.0 ;
      RECT  136200.0 1214400.0 137400.0 1215600.0 ;
      RECT  139200.0 1211700.0 140400.0 1212900.0 ;
      RECT  140400.0 1214400.0 141600.0 1215600.0 ;
      RECT  133800.0 1220550.0 148200.0 1221450.0 ;
      RECT  133800.0 1206750.0 148200.0 1207650.0 ;
      RECT  154800.0 1219050.0 156000.0 1221000.0 ;
      RECT  154800.0 1207200.0 156000.0 1209150.0 ;
      RECT  150000.0 1208550.0 151200.0 1206750.0 ;
      RECT  150000.0 1217850.0 151200.0 1221450.0 ;
      RECT  152700.0 1208550.0 153600.0 1217850.0 ;
      RECT  150000.0 1217850.0 151200.0 1219050.0 ;
      RECT  152400.0 1217850.0 153600.0 1219050.0 ;
      RECT  152400.0 1217850.0 153600.0 1219050.0 ;
      RECT  150000.0 1217850.0 151200.0 1219050.0 ;
      RECT  150000.0 1208550.0 151200.0 1209750.0 ;
      RECT  152400.0 1208550.0 153600.0 1209750.0 ;
      RECT  152400.0 1208550.0 153600.0 1209750.0 ;
      RECT  150000.0 1208550.0 151200.0 1209750.0 ;
      RECT  154800.0 1218450.0 156000.0 1219650.0 ;
      RECT  154800.0 1208550.0 156000.0 1209750.0 ;
      RECT  150600.0 1213200.0 151800.0 1214400.0 ;
      RECT  150600.0 1213200.0 151800.0 1214400.0 ;
      RECT  153150.0 1213350.0 154050.0 1214250.0 ;
      RECT  148200.0 1220550.0 157800.0 1221450.0 ;
      RECT  148200.0 1206750.0 157800.0 1207650.0 ;
      RECT  120450.0 1213200.0 121650.0 1214400.0 ;
      RECT  122400.0 1210800.0 123600.0 1212000.0 ;
      RECT  139200.0 1211700.0 138000.0 1212900.0 ;
      RECT  130800.0 1222950.0 132000.0 1221000.0 ;
      RECT  130800.0 1234800.0 132000.0 1232850.0 ;
      RECT  126000.0 1233450.0 127200.0 1235250.0 ;
      RECT  126000.0 1224150.0 127200.0 1220550.0 ;
      RECT  128700.0 1233450.0 129600.0 1224150.0 ;
      RECT  126000.0 1224150.0 127200.0 1222950.0 ;
      RECT  128400.0 1224150.0 129600.0 1222950.0 ;
      RECT  128400.0 1224150.0 129600.0 1222950.0 ;
      RECT  126000.0 1224150.0 127200.0 1222950.0 ;
      RECT  126000.0 1233450.0 127200.0 1232250.0 ;
      RECT  128400.0 1233450.0 129600.0 1232250.0 ;
      RECT  128400.0 1233450.0 129600.0 1232250.0 ;
      RECT  126000.0 1233450.0 127200.0 1232250.0 ;
      RECT  130800.0 1223550.0 132000.0 1222350.0 ;
      RECT  130800.0 1233450.0 132000.0 1232250.0 ;
      RECT  126600.0 1228800.0 127800.0 1227600.0 ;
      RECT  126600.0 1228800.0 127800.0 1227600.0 ;
      RECT  129150.0 1228650.0 130050.0 1227750.0 ;
      RECT  124200.0 1221450.0 133800.0 1220550.0 ;
      RECT  124200.0 1235250.0 133800.0 1234350.0 ;
      RECT  135600.0 1232850.0 136800.0 1235250.0 ;
      RECT  135600.0 1224150.0 136800.0 1220550.0 ;
      RECT  140400.0 1224150.0 141600.0 1220550.0 ;
      RECT  142800.0 1222950.0 144000.0 1221000.0 ;
      RECT  142800.0 1234800.0 144000.0 1232850.0 ;
      RECT  135600.0 1224150.0 136800.0 1222950.0 ;
      RECT  138000.0 1224150.0 139200.0 1222950.0 ;
      RECT  138000.0 1224150.0 139200.0 1222950.0 ;
      RECT  135600.0 1224150.0 136800.0 1222950.0 ;
      RECT  138000.0 1224150.0 139200.0 1222950.0 ;
      RECT  140400.0 1224150.0 141600.0 1222950.0 ;
      RECT  140400.0 1224150.0 141600.0 1222950.0 ;
      RECT  138000.0 1224150.0 139200.0 1222950.0 ;
      RECT  135600.0 1232850.0 136800.0 1231650.0 ;
      RECT  138000.0 1232850.0 139200.0 1231650.0 ;
      RECT  138000.0 1232850.0 139200.0 1231650.0 ;
      RECT  135600.0 1232850.0 136800.0 1231650.0 ;
      RECT  138000.0 1232850.0 139200.0 1231650.0 ;
      RECT  140400.0 1232850.0 141600.0 1231650.0 ;
      RECT  140400.0 1232850.0 141600.0 1231650.0 ;
      RECT  138000.0 1232850.0 139200.0 1231650.0 ;
      RECT  142800.0 1223550.0 144000.0 1222350.0 ;
      RECT  142800.0 1233450.0 144000.0 1232250.0 ;
      RECT  140400.0 1230300.0 139200.0 1229100.0 ;
      RECT  137400.0 1227600.0 136200.0 1226400.0 ;
      RECT  138000.0 1224150.0 139200.0 1222950.0 ;
      RECT  140400.0 1232850.0 141600.0 1231650.0 ;
      RECT  141600.0 1227600.0 140400.0 1226400.0 ;
      RECT  136200.0 1227600.0 137400.0 1226400.0 ;
      RECT  139200.0 1230300.0 140400.0 1229100.0 ;
      RECT  140400.0 1227600.0 141600.0 1226400.0 ;
      RECT  133800.0 1221450.0 148200.0 1220550.0 ;
      RECT  133800.0 1235250.0 148200.0 1234350.0 ;
      RECT  154800.0 1222950.0 156000.0 1221000.0 ;
      RECT  154800.0 1234800.0 156000.0 1232850.0 ;
      RECT  150000.0 1233450.0 151200.0 1235250.0 ;
      RECT  150000.0 1224150.0 151200.0 1220550.0 ;
      RECT  152700.0 1233450.0 153600.0 1224150.0 ;
      RECT  150000.0 1224150.0 151200.0 1222950.0 ;
      RECT  152400.0 1224150.0 153600.0 1222950.0 ;
      RECT  152400.0 1224150.0 153600.0 1222950.0 ;
      RECT  150000.0 1224150.0 151200.0 1222950.0 ;
      RECT  150000.0 1233450.0 151200.0 1232250.0 ;
      RECT  152400.0 1233450.0 153600.0 1232250.0 ;
      RECT  152400.0 1233450.0 153600.0 1232250.0 ;
      RECT  150000.0 1233450.0 151200.0 1232250.0 ;
      RECT  154800.0 1223550.0 156000.0 1222350.0 ;
      RECT  154800.0 1233450.0 156000.0 1232250.0 ;
      RECT  150600.0 1228800.0 151800.0 1227600.0 ;
      RECT  150600.0 1228800.0 151800.0 1227600.0 ;
      RECT  153150.0 1228650.0 154050.0 1227750.0 ;
      RECT  148200.0 1221450.0 157800.0 1220550.0 ;
      RECT  148200.0 1235250.0 157800.0 1234350.0 ;
      RECT  120450.0 1227600.0 121650.0 1228800.0 ;
      RECT  122400.0 1230000.0 123600.0 1231200.0 ;
      RECT  139200.0 1229100.0 138000.0 1230300.0 ;
      RECT  130800.0 1246650.0 132000.0 1248600.0 ;
      RECT  130800.0 1234800.0 132000.0 1236750.0 ;
      RECT  126000.0 1236150.0 127200.0 1234350.0 ;
      RECT  126000.0 1245450.0 127200.0 1249050.0 ;
      RECT  128700.0 1236150.0 129600.0 1245450.0 ;
      RECT  126000.0 1245450.0 127200.0 1246650.0 ;
      RECT  128400.0 1245450.0 129600.0 1246650.0 ;
      RECT  128400.0 1245450.0 129600.0 1246650.0 ;
      RECT  126000.0 1245450.0 127200.0 1246650.0 ;
      RECT  126000.0 1236150.0 127200.0 1237350.0 ;
      RECT  128400.0 1236150.0 129600.0 1237350.0 ;
      RECT  128400.0 1236150.0 129600.0 1237350.0 ;
      RECT  126000.0 1236150.0 127200.0 1237350.0 ;
      RECT  130800.0 1246050.0 132000.0 1247250.0 ;
      RECT  130800.0 1236150.0 132000.0 1237350.0 ;
      RECT  126600.0 1240800.0 127800.0 1242000.0 ;
      RECT  126600.0 1240800.0 127800.0 1242000.0 ;
      RECT  129150.0 1240950.0 130050.0 1241850.0 ;
      RECT  124200.0 1248150.0 133800.0 1249050.0 ;
      RECT  124200.0 1234350.0 133800.0 1235250.0 ;
      RECT  135600.0 1236750.0 136800.0 1234350.0 ;
      RECT  135600.0 1245450.0 136800.0 1249050.0 ;
      RECT  140400.0 1245450.0 141600.0 1249050.0 ;
      RECT  142800.0 1246650.0 144000.0 1248600.0 ;
      RECT  142800.0 1234800.0 144000.0 1236750.0 ;
      RECT  135600.0 1245450.0 136800.0 1246650.0 ;
      RECT  138000.0 1245450.0 139200.0 1246650.0 ;
      RECT  138000.0 1245450.0 139200.0 1246650.0 ;
      RECT  135600.0 1245450.0 136800.0 1246650.0 ;
      RECT  138000.0 1245450.0 139200.0 1246650.0 ;
      RECT  140400.0 1245450.0 141600.0 1246650.0 ;
      RECT  140400.0 1245450.0 141600.0 1246650.0 ;
      RECT  138000.0 1245450.0 139200.0 1246650.0 ;
      RECT  135600.0 1236750.0 136800.0 1237950.0 ;
      RECT  138000.0 1236750.0 139200.0 1237950.0 ;
      RECT  138000.0 1236750.0 139200.0 1237950.0 ;
      RECT  135600.0 1236750.0 136800.0 1237950.0 ;
      RECT  138000.0 1236750.0 139200.0 1237950.0 ;
      RECT  140400.0 1236750.0 141600.0 1237950.0 ;
      RECT  140400.0 1236750.0 141600.0 1237950.0 ;
      RECT  138000.0 1236750.0 139200.0 1237950.0 ;
      RECT  142800.0 1246050.0 144000.0 1247250.0 ;
      RECT  142800.0 1236150.0 144000.0 1237350.0 ;
      RECT  140400.0 1239300.0 139200.0 1240500.0 ;
      RECT  137400.0 1242000.0 136200.0 1243200.0 ;
      RECT  138000.0 1245450.0 139200.0 1246650.0 ;
      RECT  140400.0 1236750.0 141600.0 1237950.0 ;
      RECT  141600.0 1242000.0 140400.0 1243200.0 ;
      RECT  136200.0 1242000.0 137400.0 1243200.0 ;
      RECT  139200.0 1239300.0 140400.0 1240500.0 ;
      RECT  140400.0 1242000.0 141600.0 1243200.0 ;
      RECT  133800.0 1248150.0 148200.0 1249050.0 ;
      RECT  133800.0 1234350.0 148200.0 1235250.0 ;
      RECT  154800.0 1246650.0 156000.0 1248600.0 ;
      RECT  154800.0 1234800.0 156000.0 1236750.0 ;
      RECT  150000.0 1236150.0 151200.0 1234350.0 ;
      RECT  150000.0 1245450.0 151200.0 1249050.0 ;
      RECT  152700.0 1236150.0 153600.0 1245450.0 ;
      RECT  150000.0 1245450.0 151200.0 1246650.0 ;
      RECT  152400.0 1245450.0 153600.0 1246650.0 ;
      RECT  152400.0 1245450.0 153600.0 1246650.0 ;
      RECT  150000.0 1245450.0 151200.0 1246650.0 ;
      RECT  150000.0 1236150.0 151200.0 1237350.0 ;
      RECT  152400.0 1236150.0 153600.0 1237350.0 ;
      RECT  152400.0 1236150.0 153600.0 1237350.0 ;
      RECT  150000.0 1236150.0 151200.0 1237350.0 ;
      RECT  154800.0 1246050.0 156000.0 1247250.0 ;
      RECT  154800.0 1236150.0 156000.0 1237350.0 ;
      RECT  150600.0 1240800.0 151800.0 1242000.0 ;
      RECT  150600.0 1240800.0 151800.0 1242000.0 ;
      RECT  153150.0 1240950.0 154050.0 1241850.0 ;
      RECT  148200.0 1248150.0 157800.0 1249050.0 ;
      RECT  148200.0 1234350.0 157800.0 1235250.0 ;
      RECT  120450.0 1240800.0 121650.0 1242000.0 ;
      RECT  122400.0 1238400.0 123600.0 1239600.0 ;
      RECT  139200.0 1239300.0 138000.0 1240500.0 ;
      RECT  130800.0 1250550.0 132000.0 1248600.0 ;
      RECT  130800.0 1262400.0 132000.0 1260450.0 ;
      RECT  126000.0 1261050.0 127200.0 1262850.0 ;
      RECT  126000.0 1251750.0 127200.0 1248150.0 ;
      RECT  128700.0 1261050.0 129600.0 1251750.0 ;
      RECT  126000.0 1251750.0 127200.0 1250550.0 ;
      RECT  128400.0 1251750.0 129600.0 1250550.0 ;
      RECT  128400.0 1251750.0 129600.0 1250550.0 ;
      RECT  126000.0 1251750.0 127200.0 1250550.0 ;
      RECT  126000.0 1261050.0 127200.0 1259850.0 ;
      RECT  128400.0 1261050.0 129600.0 1259850.0 ;
      RECT  128400.0 1261050.0 129600.0 1259850.0 ;
      RECT  126000.0 1261050.0 127200.0 1259850.0 ;
      RECT  130800.0 1251150.0 132000.0 1249950.0 ;
      RECT  130800.0 1261050.0 132000.0 1259850.0 ;
      RECT  126600.0 1256400.0 127800.0 1255200.0 ;
      RECT  126600.0 1256400.0 127800.0 1255200.0 ;
      RECT  129150.0 1256250.0 130050.0 1255350.0 ;
      RECT  124200.0 1249050.0 133800.0 1248150.0 ;
      RECT  124200.0 1262850.0 133800.0 1261950.0 ;
      RECT  135600.0 1260450.0 136800.0 1262850.0 ;
      RECT  135600.0 1251750.0 136800.0 1248150.0 ;
      RECT  140400.0 1251750.0 141600.0 1248150.0 ;
      RECT  142800.0 1250550.0 144000.0 1248600.0 ;
      RECT  142800.0 1262400.0 144000.0 1260450.0 ;
      RECT  135600.0 1251750.0 136800.0 1250550.0 ;
      RECT  138000.0 1251750.0 139200.0 1250550.0 ;
      RECT  138000.0 1251750.0 139200.0 1250550.0 ;
      RECT  135600.0 1251750.0 136800.0 1250550.0 ;
      RECT  138000.0 1251750.0 139200.0 1250550.0 ;
      RECT  140400.0 1251750.0 141600.0 1250550.0 ;
      RECT  140400.0 1251750.0 141600.0 1250550.0 ;
      RECT  138000.0 1251750.0 139200.0 1250550.0 ;
      RECT  135600.0 1260450.0 136800.0 1259250.0 ;
      RECT  138000.0 1260450.0 139200.0 1259250.0 ;
      RECT  138000.0 1260450.0 139200.0 1259250.0 ;
      RECT  135600.0 1260450.0 136800.0 1259250.0 ;
      RECT  138000.0 1260450.0 139200.0 1259250.0 ;
      RECT  140400.0 1260450.0 141600.0 1259250.0 ;
      RECT  140400.0 1260450.0 141600.0 1259250.0 ;
      RECT  138000.0 1260450.0 139200.0 1259250.0 ;
      RECT  142800.0 1251150.0 144000.0 1249950.0 ;
      RECT  142800.0 1261050.0 144000.0 1259850.0 ;
      RECT  140400.0 1257900.0 139200.0 1256700.0 ;
      RECT  137400.0 1255200.0 136200.0 1254000.0 ;
      RECT  138000.0 1251750.0 139200.0 1250550.0 ;
      RECT  140400.0 1260450.0 141600.0 1259250.0 ;
      RECT  141600.0 1255200.0 140400.0 1254000.0 ;
      RECT  136200.0 1255200.0 137400.0 1254000.0 ;
      RECT  139200.0 1257900.0 140400.0 1256700.0 ;
      RECT  140400.0 1255200.0 141600.0 1254000.0 ;
      RECT  133800.0 1249050.0 148200.0 1248150.0 ;
      RECT  133800.0 1262850.0 148200.0 1261950.0 ;
      RECT  154800.0 1250550.0 156000.0 1248600.0 ;
      RECT  154800.0 1262400.0 156000.0 1260450.0 ;
      RECT  150000.0 1261050.0 151200.0 1262850.0 ;
      RECT  150000.0 1251750.0 151200.0 1248150.0 ;
      RECT  152700.0 1261050.0 153600.0 1251750.0 ;
      RECT  150000.0 1251750.0 151200.0 1250550.0 ;
      RECT  152400.0 1251750.0 153600.0 1250550.0 ;
      RECT  152400.0 1251750.0 153600.0 1250550.0 ;
      RECT  150000.0 1251750.0 151200.0 1250550.0 ;
      RECT  150000.0 1261050.0 151200.0 1259850.0 ;
      RECT  152400.0 1261050.0 153600.0 1259850.0 ;
      RECT  152400.0 1261050.0 153600.0 1259850.0 ;
      RECT  150000.0 1261050.0 151200.0 1259850.0 ;
      RECT  154800.0 1251150.0 156000.0 1249950.0 ;
      RECT  154800.0 1261050.0 156000.0 1259850.0 ;
      RECT  150600.0 1256400.0 151800.0 1255200.0 ;
      RECT  150600.0 1256400.0 151800.0 1255200.0 ;
      RECT  153150.0 1256250.0 154050.0 1255350.0 ;
      RECT  148200.0 1249050.0 157800.0 1248150.0 ;
      RECT  148200.0 1262850.0 157800.0 1261950.0 ;
      RECT  120450.0 1255200.0 121650.0 1256400.0 ;
      RECT  122400.0 1257600.0 123600.0 1258800.0 ;
      RECT  139200.0 1256700.0 138000.0 1257900.0 ;
      RECT  130800.0 1274250.0 132000.0 1276200.0 ;
      RECT  130800.0 1262400.0 132000.0 1264350.0 ;
      RECT  126000.0 1263750.0 127200.0 1261950.0 ;
      RECT  126000.0 1273050.0 127200.0 1276650.0 ;
      RECT  128700.0 1263750.0 129600.0 1273050.0 ;
      RECT  126000.0 1273050.0 127200.0 1274250.0 ;
      RECT  128400.0 1273050.0 129600.0 1274250.0 ;
      RECT  128400.0 1273050.0 129600.0 1274250.0 ;
      RECT  126000.0 1273050.0 127200.0 1274250.0 ;
      RECT  126000.0 1263750.0 127200.0 1264950.0 ;
      RECT  128400.0 1263750.0 129600.0 1264950.0 ;
      RECT  128400.0 1263750.0 129600.0 1264950.0 ;
      RECT  126000.0 1263750.0 127200.0 1264950.0 ;
      RECT  130800.0 1273650.0 132000.0 1274850.0 ;
      RECT  130800.0 1263750.0 132000.0 1264950.0 ;
      RECT  126600.0 1268400.0 127800.0 1269600.0 ;
      RECT  126600.0 1268400.0 127800.0 1269600.0 ;
      RECT  129150.0 1268550.0 130050.0 1269450.0 ;
      RECT  124200.0 1275750.0 133800.0 1276650.0 ;
      RECT  124200.0 1261950.0 133800.0 1262850.0 ;
      RECT  135600.0 1264350.0 136800.0 1261950.0 ;
      RECT  135600.0 1273050.0 136800.0 1276650.0 ;
      RECT  140400.0 1273050.0 141600.0 1276650.0 ;
      RECT  142800.0 1274250.0 144000.0 1276200.0 ;
      RECT  142800.0 1262400.0 144000.0 1264350.0 ;
      RECT  135600.0 1273050.0 136800.0 1274250.0 ;
      RECT  138000.0 1273050.0 139200.0 1274250.0 ;
      RECT  138000.0 1273050.0 139200.0 1274250.0 ;
      RECT  135600.0 1273050.0 136800.0 1274250.0 ;
      RECT  138000.0 1273050.0 139200.0 1274250.0 ;
      RECT  140400.0 1273050.0 141600.0 1274250.0 ;
      RECT  140400.0 1273050.0 141600.0 1274250.0 ;
      RECT  138000.0 1273050.0 139200.0 1274250.0 ;
      RECT  135600.0 1264350.0 136800.0 1265550.0 ;
      RECT  138000.0 1264350.0 139200.0 1265550.0 ;
      RECT  138000.0 1264350.0 139200.0 1265550.0 ;
      RECT  135600.0 1264350.0 136800.0 1265550.0 ;
      RECT  138000.0 1264350.0 139200.0 1265550.0 ;
      RECT  140400.0 1264350.0 141600.0 1265550.0 ;
      RECT  140400.0 1264350.0 141600.0 1265550.0 ;
      RECT  138000.0 1264350.0 139200.0 1265550.0 ;
      RECT  142800.0 1273650.0 144000.0 1274850.0 ;
      RECT  142800.0 1263750.0 144000.0 1264950.0 ;
      RECT  140400.0 1266900.0 139200.0 1268100.0 ;
      RECT  137400.0 1269600.0 136200.0 1270800.0 ;
      RECT  138000.0 1273050.0 139200.0 1274250.0 ;
      RECT  140400.0 1264350.0 141600.0 1265550.0 ;
      RECT  141600.0 1269600.0 140400.0 1270800.0 ;
      RECT  136200.0 1269600.0 137400.0 1270800.0 ;
      RECT  139200.0 1266900.0 140400.0 1268100.0 ;
      RECT  140400.0 1269600.0 141600.0 1270800.0 ;
      RECT  133800.0 1275750.0 148200.0 1276650.0 ;
      RECT  133800.0 1261950.0 148200.0 1262850.0 ;
      RECT  154800.0 1274250.0 156000.0 1276200.0 ;
      RECT  154800.0 1262400.0 156000.0 1264350.0 ;
      RECT  150000.0 1263750.0 151200.0 1261950.0 ;
      RECT  150000.0 1273050.0 151200.0 1276650.0 ;
      RECT  152700.0 1263750.0 153600.0 1273050.0 ;
      RECT  150000.0 1273050.0 151200.0 1274250.0 ;
      RECT  152400.0 1273050.0 153600.0 1274250.0 ;
      RECT  152400.0 1273050.0 153600.0 1274250.0 ;
      RECT  150000.0 1273050.0 151200.0 1274250.0 ;
      RECT  150000.0 1263750.0 151200.0 1264950.0 ;
      RECT  152400.0 1263750.0 153600.0 1264950.0 ;
      RECT  152400.0 1263750.0 153600.0 1264950.0 ;
      RECT  150000.0 1263750.0 151200.0 1264950.0 ;
      RECT  154800.0 1273650.0 156000.0 1274850.0 ;
      RECT  154800.0 1263750.0 156000.0 1264950.0 ;
      RECT  150600.0 1268400.0 151800.0 1269600.0 ;
      RECT  150600.0 1268400.0 151800.0 1269600.0 ;
      RECT  153150.0 1268550.0 154050.0 1269450.0 ;
      RECT  148200.0 1275750.0 157800.0 1276650.0 ;
      RECT  148200.0 1261950.0 157800.0 1262850.0 ;
      RECT  120450.0 1268400.0 121650.0 1269600.0 ;
      RECT  122400.0 1266000.0 123600.0 1267200.0 ;
      RECT  139200.0 1266900.0 138000.0 1268100.0 ;
      RECT  130800.0 1278150.0 132000.0 1276200.0 ;
      RECT  130800.0 1290000.0 132000.0 1288050.0 ;
      RECT  126000.0 1288650.0 127200.0 1290450.0 ;
      RECT  126000.0 1279350.0 127200.0 1275750.0 ;
      RECT  128700.0 1288650.0 129600.0 1279350.0 ;
      RECT  126000.0 1279350.0 127200.0 1278150.0 ;
      RECT  128400.0 1279350.0 129600.0 1278150.0 ;
      RECT  128400.0 1279350.0 129600.0 1278150.0 ;
      RECT  126000.0 1279350.0 127200.0 1278150.0 ;
      RECT  126000.0 1288650.0 127200.0 1287450.0 ;
      RECT  128400.0 1288650.0 129600.0 1287450.0 ;
      RECT  128400.0 1288650.0 129600.0 1287450.0 ;
      RECT  126000.0 1288650.0 127200.0 1287450.0 ;
      RECT  130800.0 1278750.0 132000.0 1277550.0 ;
      RECT  130800.0 1288650.0 132000.0 1287450.0 ;
      RECT  126600.0 1284000.0 127800.0 1282800.0 ;
      RECT  126600.0 1284000.0 127800.0 1282800.0 ;
      RECT  129150.0 1283850.0 130050.0 1282950.0 ;
      RECT  124200.0 1276650.0 133800.0 1275750.0 ;
      RECT  124200.0 1290450.0 133800.0 1289550.0 ;
      RECT  135600.0 1288050.0 136800.0 1290450.0 ;
      RECT  135600.0 1279350.0 136800.0 1275750.0 ;
      RECT  140400.0 1279350.0 141600.0 1275750.0 ;
      RECT  142800.0 1278150.0 144000.0 1276200.0 ;
      RECT  142800.0 1290000.0 144000.0 1288050.0 ;
      RECT  135600.0 1279350.0 136800.0 1278150.0 ;
      RECT  138000.0 1279350.0 139200.0 1278150.0 ;
      RECT  138000.0 1279350.0 139200.0 1278150.0 ;
      RECT  135600.0 1279350.0 136800.0 1278150.0 ;
      RECT  138000.0 1279350.0 139200.0 1278150.0 ;
      RECT  140400.0 1279350.0 141600.0 1278150.0 ;
      RECT  140400.0 1279350.0 141600.0 1278150.0 ;
      RECT  138000.0 1279350.0 139200.0 1278150.0 ;
      RECT  135600.0 1288050.0 136800.0 1286850.0 ;
      RECT  138000.0 1288050.0 139200.0 1286850.0 ;
      RECT  138000.0 1288050.0 139200.0 1286850.0 ;
      RECT  135600.0 1288050.0 136800.0 1286850.0 ;
      RECT  138000.0 1288050.0 139200.0 1286850.0 ;
      RECT  140400.0 1288050.0 141600.0 1286850.0 ;
      RECT  140400.0 1288050.0 141600.0 1286850.0 ;
      RECT  138000.0 1288050.0 139200.0 1286850.0 ;
      RECT  142800.0 1278750.0 144000.0 1277550.0 ;
      RECT  142800.0 1288650.0 144000.0 1287450.0 ;
      RECT  140400.0 1285500.0 139200.0 1284300.0 ;
      RECT  137400.0 1282800.0 136200.0 1281600.0 ;
      RECT  138000.0 1279350.0 139200.0 1278150.0 ;
      RECT  140400.0 1288050.0 141600.0 1286850.0 ;
      RECT  141600.0 1282800.0 140400.0 1281600.0 ;
      RECT  136200.0 1282800.0 137400.0 1281600.0 ;
      RECT  139200.0 1285500.0 140400.0 1284300.0 ;
      RECT  140400.0 1282800.0 141600.0 1281600.0 ;
      RECT  133800.0 1276650.0 148200.0 1275750.0 ;
      RECT  133800.0 1290450.0 148200.0 1289550.0 ;
      RECT  154800.0 1278150.0 156000.0 1276200.0 ;
      RECT  154800.0 1290000.0 156000.0 1288050.0 ;
      RECT  150000.0 1288650.0 151200.0 1290450.0 ;
      RECT  150000.0 1279350.0 151200.0 1275750.0 ;
      RECT  152700.0 1288650.0 153600.0 1279350.0 ;
      RECT  150000.0 1279350.0 151200.0 1278150.0 ;
      RECT  152400.0 1279350.0 153600.0 1278150.0 ;
      RECT  152400.0 1279350.0 153600.0 1278150.0 ;
      RECT  150000.0 1279350.0 151200.0 1278150.0 ;
      RECT  150000.0 1288650.0 151200.0 1287450.0 ;
      RECT  152400.0 1288650.0 153600.0 1287450.0 ;
      RECT  152400.0 1288650.0 153600.0 1287450.0 ;
      RECT  150000.0 1288650.0 151200.0 1287450.0 ;
      RECT  154800.0 1278750.0 156000.0 1277550.0 ;
      RECT  154800.0 1288650.0 156000.0 1287450.0 ;
      RECT  150600.0 1284000.0 151800.0 1282800.0 ;
      RECT  150600.0 1284000.0 151800.0 1282800.0 ;
      RECT  153150.0 1283850.0 154050.0 1282950.0 ;
      RECT  148200.0 1276650.0 157800.0 1275750.0 ;
      RECT  148200.0 1290450.0 157800.0 1289550.0 ;
      RECT  120450.0 1282800.0 121650.0 1284000.0 ;
      RECT  122400.0 1285200.0 123600.0 1286400.0 ;
      RECT  139200.0 1284300.0 138000.0 1285500.0 ;
      RECT  130800.0 1301850.0 132000.0 1303800.0 ;
      RECT  130800.0 1290000.0 132000.0 1291950.0 ;
      RECT  126000.0 1291350.0 127200.0 1289550.0 ;
      RECT  126000.0 1300650.0 127200.0 1304250.0 ;
      RECT  128700.0 1291350.0 129600.0 1300650.0 ;
      RECT  126000.0 1300650.0 127200.0 1301850.0 ;
      RECT  128400.0 1300650.0 129600.0 1301850.0 ;
      RECT  128400.0 1300650.0 129600.0 1301850.0 ;
      RECT  126000.0 1300650.0 127200.0 1301850.0 ;
      RECT  126000.0 1291350.0 127200.0 1292550.0 ;
      RECT  128400.0 1291350.0 129600.0 1292550.0 ;
      RECT  128400.0 1291350.0 129600.0 1292550.0 ;
      RECT  126000.0 1291350.0 127200.0 1292550.0 ;
      RECT  130800.0 1301250.0 132000.0 1302450.0 ;
      RECT  130800.0 1291350.0 132000.0 1292550.0 ;
      RECT  126600.0 1296000.0 127800.0 1297200.0 ;
      RECT  126600.0 1296000.0 127800.0 1297200.0 ;
      RECT  129150.0 1296150.0 130050.0 1297050.0 ;
      RECT  124200.0 1303350.0 133800.0 1304250.0 ;
      RECT  124200.0 1289550.0 133800.0 1290450.0 ;
      RECT  135600.0 1291950.0 136800.0 1289550.0 ;
      RECT  135600.0 1300650.0 136800.0 1304250.0 ;
      RECT  140400.0 1300650.0 141600.0 1304250.0 ;
      RECT  142800.0 1301850.0 144000.0 1303800.0 ;
      RECT  142800.0 1290000.0 144000.0 1291950.0 ;
      RECT  135600.0 1300650.0 136800.0 1301850.0 ;
      RECT  138000.0 1300650.0 139200.0 1301850.0 ;
      RECT  138000.0 1300650.0 139200.0 1301850.0 ;
      RECT  135600.0 1300650.0 136800.0 1301850.0 ;
      RECT  138000.0 1300650.0 139200.0 1301850.0 ;
      RECT  140400.0 1300650.0 141600.0 1301850.0 ;
      RECT  140400.0 1300650.0 141600.0 1301850.0 ;
      RECT  138000.0 1300650.0 139200.0 1301850.0 ;
      RECT  135600.0 1291950.0 136800.0 1293150.0 ;
      RECT  138000.0 1291950.0 139200.0 1293150.0 ;
      RECT  138000.0 1291950.0 139200.0 1293150.0 ;
      RECT  135600.0 1291950.0 136800.0 1293150.0 ;
      RECT  138000.0 1291950.0 139200.0 1293150.0 ;
      RECT  140400.0 1291950.0 141600.0 1293150.0 ;
      RECT  140400.0 1291950.0 141600.0 1293150.0 ;
      RECT  138000.0 1291950.0 139200.0 1293150.0 ;
      RECT  142800.0 1301250.0 144000.0 1302450.0 ;
      RECT  142800.0 1291350.0 144000.0 1292550.0 ;
      RECT  140400.0 1294500.0 139200.0 1295700.0 ;
      RECT  137400.0 1297200.0 136200.0 1298400.0 ;
      RECT  138000.0 1300650.0 139200.0 1301850.0 ;
      RECT  140400.0 1291950.0 141600.0 1293150.0 ;
      RECT  141600.0 1297200.0 140400.0 1298400.0 ;
      RECT  136200.0 1297200.0 137400.0 1298400.0 ;
      RECT  139200.0 1294500.0 140400.0 1295700.0 ;
      RECT  140400.0 1297200.0 141600.0 1298400.0 ;
      RECT  133800.0 1303350.0 148200.0 1304250.0 ;
      RECT  133800.0 1289550.0 148200.0 1290450.0 ;
      RECT  154800.0 1301850.0 156000.0 1303800.0 ;
      RECT  154800.0 1290000.0 156000.0 1291950.0 ;
      RECT  150000.0 1291350.0 151200.0 1289550.0 ;
      RECT  150000.0 1300650.0 151200.0 1304250.0 ;
      RECT  152700.0 1291350.0 153600.0 1300650.0 ;
      RECT  150000.0 1300650.0 151200.0 1301850.0 ;
      RECT  152400.0 1300650.0 153600.0 1301850.0 ;
      RECT  152400.0 1300650.0 153600.0 1301850.0 ;
      RECT  150000.0 1300650.0 151200.0 1301850.0 ;
      RECT  150000.0 1291350.0 151200.0 1292550.0 ;
      RECT  152400.0 1291350.0 153600.0 1292550.0 ;
      RECT  152400.0 1291350.0 153600.0 1292550.0 ;
      RECT  150000.0 1291350.0 151200.0 1292550.0 ;
      RECT  154800.0 1301250.0 156000.0 1302450.0 ;
      RECT  154800.0 1291350.0 156000.0 1292550.0 ;
      RECT  150600.0 1296000.0 151800.0 1297200.0 ;
      RECT  150600.0 1296000.0 151800.0 1297200.0 ;
      RECT  153150.0 1296150.0 154050.0 1297050.0 ;
      RECT  148200.0 1303350.0 157800.0 1304250.0 ;
      RECT  148200.0 1289550.0 157800.0 1290450.0 ;
      RECT  120450.0 1296000.0 121650.0 1297200.0 ;
      RECT  122400.0 1293600.0 123600.0 1294800.0 ;
      RECT  139200.0 1294500.0 138000.0 1295700.0 ;
      RECT  130800.0 1305750.0 132000.0 1303800.0 ;
      RECT  130800.0 1317600.0 132000.0 1315650.0 ;
      RECT  126000.0 1316250.0 127200.0 1318050.0 ;
      RECT  126000.0 1306950.0 127200.0 1303350.0 ;
      RECT  128700.0 1316250.0 129600.0 1306950.0 ;
      RECT  126000.0 1306950.0 127200.0 1305750.0 ;
      RECT  128400.0 1306950.0 129600.0 1305750.0 ;
      RECT  128400.0 1306950.0 129600.0 1305750.0 ;
      RECT  126000.0 1306950.0 127200.0 1305750.0 ;
      RECT  126000.0 1316250.0 127200.0 1315050.0 ;
      RECT  128400.0 1316250.0 129600.0 1315050.0 ;
      RECT  128400.0 1316250.0 129600.0 1315050.0 ;
      RECT  126000.0 1316250.0 127200.0 1315050.0 ;
      RECT  130800.0 1306350.0 132000.0 1305150.0 ;
      RECT  130800.0 1316250.0 132000.0 1315050.0 ;
      RECT  126600.0 1311600.0 127800.0 1310400.0 ;
      RECT  126600.0 1311600.0 127800.0 1310400.0 ;
      RECT  129150.0 1311450.0 130050.0 1310550.0 ;
      RECT  124200.0 1304250.0 133800.0 1303350.0 ;
      RECT  124200.0 1318050.0 133800.0 1317150.0 ;
      RECT  135600.0 1315650.0 136800.0 1318050.0 ;
      RECT  135600.0 1306950.0 136800.0 1303350.0 ;
      RECT  140400.0 1306950.0 141600.0 1303350.0 ;
      RECT  142800.0 1305750.0 144000.0 1303800.0 ;
      RECT  142800.0 1317600.0 144000.0 1315650.0 ;
      RECT  135600.0 1306950.0 136800.0 1305750.0 ;
      RECT  138000.0 1306950.0 139200.0 1305750.0 ;
      RECT  138000.0 1306950.0 139200.0 1305750.0 ;
      RECT  135600.0 1306950.0 136800.0 1305750.0 ;
      RECT  138000.0 1306950.0 139200.0 1305750.0 ;
      RECT  140400.0 1306950.0 141600.0 1305750.0 ;
      RECT  140400.0 1306950.0 141600.0 1305750.0 ;
      RECT  138000.0 1306950.0 139200.0 1305750.0 ;
      RECT  135600.0 1315650.0 136800.0 1314450.0 ;
      RECT  138000.0 1315650.0 139200.0 1314450.0 ;
      RECT  138000.0 1315650.0 139200.0 1314450.0 ;
      RECT  135600.0 1315650.0 136800.0 1314450.0 ;
      RECT  138000.0 1315650.0 139200.0 1314450.0 ;
      RECT  140400.0 1315650.0 141600.0 1314450.0 ;
      RECT  140400.0 1315650.0 141600.0 1314450.0 ;
      RECT  138000.0 1315650.0 139200.0 1314450.0 ;
      RECT  142800.0 1306350.0 144000.0 1305150.0 ;
      RECT  142800.0 1316250.0 144000.0 1315050.0 ;
      RECT  140400.0 1313100.0 139200.0 1311900.0 ;
      RECT  137400.0 1310400.0 136200.0 1309200.0 ;
      RECT  138000.0 1306950.0 139200.0 1305750.0 ;
      RECT  140400.0 1315650.0 141600.0 1314450.0 ;
      RECT  141600.0 1310400.0 140400.0 1309200.0 ;
      RECT  136200.0 1310400.0 137400.0 1309200.0 ;
      RECT  139200.0 1313100.0 140400.0 1311900.0 ;
      RECT  140400.0 1310400.0 141600.0 1309200.0 ;
      RECT  133800.0 1304250.0 148200.0 1303350.0 ;
      RECT  133800.0 1318050.0 148200.0 1317150.0 ;
      RECT  154800.0 1305750.0 156000.0 1303800.0 ;
      RECT  154800.0 1317600.0 156000.0 1315650.0 ;
      RECT  150000.0 1316250.0 151200.0 1318050.0 ;
      RECT  150000.0 1306950.0 151200.0 1303350.0 ;
      RECT  152700.0 1316250.0 153600.0 1306950.0 ;
      RECT  150000.0 1306950.0 151200.0 1305750.0 ;
      RECT  152400.0 1306950.0 153600.0 1305750.0 ;
      RECT  152400.0 1306950.0 153600.0 1305750.0 ;
      RECT  150000.0 1306950.0 151200.0 1305750.0 ;
      RECT  150000.0 1316250.0 151200.0 1315050.0 ;
      RECT  152400.0 1316250.0 153600.0 1315050.0 ;
      RECT  152400.0 1316250.0 153600.0 1315050.0 ;
      RECT  150000.0 1316250.0 151200.0 1315050.0 ;
      RECT  154800.0 1306350.0 156000.0 1305150.0 ;
      RECT  154800.0 1316250.0 156000.0 1315050.0 ;
      RECT  150600.0 1311600.0 151800.0 1310400.0 ;
      RECT  150600.0 1311600.0 151800.0 1310400.0 ;
      RECT  153150.0 1311450.0 154050.0 1310550.0 ;
      RECT  148200.0 1304250.0 157800.0 1303350.0 ;
      RECT  148200.0 1318050.0 157800.0 1317150.0 ;
      RECT  120450.0 1310400.0 121650.0 1311600.0 ;
      RECT  122400.0 1312800.0 123600.0 1314000.0 ;
      RECT  139200.0 1311900.0 138000.0 1313100.0 ;
      RECT  130800.0 1329450.0 132000.0 1331400.0 ;
      RECT  130800.0 1317600.0 132000.0 1319550.0 ;
      RECT  126000.0 1318950.0 127200.0 1317150.0 ;
      RECT  126000.0 1328250.0 127200.0 1331850.0 ;
      RECT  128700.0 1318950.0 129600.0 1328250.0 ;
      RECT  126000.0 1328250.0 127200.0 1329450.0 ;
      RECT  128400.0 1328250.0 129600.0 1329450.0 ;
      RECT  128400.0 1328250.0 129600.0 1329450.0 ;
      RECT  126000.0 1328250.0 127200.0 1329450.0 ;
      RECT  126000.0 1318950.0 127200.0 1320150.0 ;
      RECT  128400.0 1318950.0 129600.0 1320150.0 ;
      RECT  128400.0 1318950.0 129600.0 1320150.0 ;
      RECT  126000.0 1318950.0 127200.0 1320150.0 ;
      RECT  130800.0 1328850.0 132000.0 1330050.0 ;
      RECT  130800.0 1318950.0 132000.0 1320150.0 ;
      RECT  126600.0 1323600.0 127800.0 1324800.0 ;
      RECT  126600.0 1323600.0 127800.0 1324800.0 ;
      RECT  129150.0 1323750.0 130050.0 1324650.0 ;
      RECT  124200.0 1330950.0 133800.0 1331850.0 ;
      RECT  124200.0 1317150.0 133800.0 1318050.0 ;
      RECT  135600.0 1319550.0 136800.0 1317150.0 ;
      RECT  135600.0 1328250.0 136800.0 1331850.0 ;
      RECT  140400.0 1328250.0 141600.0 1331850.0 ;
      RECT  142800.0 1329450.0 144000.0 1331400.0 ;
      RECT  142800.0 1317600.0 144000.0 1319550.0 ;
      RECT  135600.0 1328250.0 136800.0 1329450.0 ;
      RECT  138000.0 1328250.0 139200.0 1329450.0 ;
      RECT  138000.0 1328250.0 139200.0 1329450.0 ;
      RECT  135600.0 1328250.0 136800.0 1329450.0 ;
      RECT  138000.0 1328250.0 139200.0 1329450.0 ;
      RECT  140400.0 1328250.0 141600.0 1329450.0 ;
      RECT  140400.0 1328250.0 141600.0 1329450.0 ;
      RECT  138000.0 1328250.0 139200.0 1329450.0 ;
      RECT  135600.0 1319550.0 136800.0 1320750.0 ;
      RECT  138000.0 1319550.0 139200.0 1320750.0 ;
      RECT  138000.0 1319550.0 139200.0 1320750.0 ;
      RECT  135600.0 1319550.0 136800.0 1320750.0 ;
      RECT  138000.0 1319550.0 139200.0 1320750.0 ;
      RECT  140400.0 1319550.0 141600.0 1320750.0 ;
      RECT  140400.0 1319550.0 141600.0 1320750.0 ;
      RECT  138000.0 1319550.0 139200.0 1320750.0 ;
      RECT  142800.0 1328850.0 144000.0 1330050.0 ;
      RECT  142800.0 1318950.0 144000.0 1320150.0 ;
      RECT  140400.0 1322100.0 139200.0 1323300.0 ;
      RECT  137400.0 1324800.0 136200.0 1326000.0 ;
      RECT  138000.0 1328250.0 139200.0 1329450.0 ;
      RECT  140400.0 1319550.0 141600.0 1320750.0 ;
      RECT  141600.0 1324800.0 140400.0 1326000.0 ;
      RECT  136200.0 1324800.0 137400.0 1326000.0 ;
      RECT  139200.0 1322100.0 140400.0 1323300.0 ;
      RECT  140400.0 1324800.0 141600.0 1326000.0 ;
      RECT  133800.0 1330950.0 148200.0 1331850.0 ;
      RECT  133800.0 1317150.0 148200.0 1318050.0 ;
      RECT  154800.0 1329450.0 156000.0 1331400.0 ;
      RECT  154800.0 1317600.0 156000.0 1319550.0 ;
      RECT  150000.0 1318950.0 151200.0 1317150.0 ;
      RECT  150000.0 1328250.0 151200.0 1331850.0 ;
      RECT  152700.0 1318950.0 153600.0 1328250.0 ;
      RECT  150000.0 1328250.0 151200.0 1329450.0 ;
      RECT  152400.0 1328250.0 153600.0 1329450.0 ;
      RECT  152400.0 1328250.0 153600.0 1329450.0 ;
      RECT  150000.0 1328250.0 151200.0 1329450.0 ;
      RECT  150000.0 1318950.0 151200.0 1320150.0 ;
      RECT  152400.0 1318950.0 153600.0 1320150.0 ;
      RECT  152400.0 1318950.0 153600.0 1320150.0 ;
      RECT  150000.0 1318950.0 151200.0 1320150.0 ;
      RECT  154800.0 1328850.0 156000.0 1330050.0 ;
      RECT  154800.0 1318950.0 156000.0 1320150.0 ;
      RECT  150600.0 1323600.0 151800.0 1324800.0 ;
      RECT  150600.0 1323600.0 151800.0 1324800.0 ;
      RECT  153150.0 1323750.0 154050.0 1324650.0 ;
      RECT  148200.0 1330950.0 157800.0 1331850.0 ;
      RECT  148200.0 1317150.0 157800.0 1318050.0 ;
      RECT  120450.0 1323600.0 121650.0 1324800.0 ;
      RECT  122400.0 1321200.0 123600.0 1322400.0 ;
      RECT  139200.0 1322100.0 138000.0 1323300.0 ;
      RECT  130800.0 1333350.0 132000.0 1331400.0 ;
      RECT  130800.0 1345200.0 132000.0 1343250.0 ;
      RECT  126000.0 1343850.0 127200.0 1345650.0 ;
      RECT  126000.0 1334550.0 127200.0 1330950.0 ;
      RECT  128700.0 1343850.0 129600.0 1334550.0 ;
      RECT  126000.0 1334550.0 127200.0 1333350.0 ;
      RECT  128400.0 1334550.0 129600.0 1333350.0 ;
      RECT  128400.0 1334550.0 129600.0 1333350.0 ;
      RECT  126000.0 1334550.0 127200.0 1333350.0 ;
      RECT  126000.0 1343850.0 127200.0 1342650.0 ;
      RECT  128400.0 1343850.0 129600.0 1342650.0 ;
      RECT  128400.0 1343850.0 129600.0 1342650.0 ;
      RECT  126000.0 1343850.0 127200.0 1342650.0 ;
      RECT  130800.0 1333950.0 132000.0 1332750.0 ;
      RECT  130800.0 1343850.0 132000.0 1342650.0 ;
      RECT  126600.0 1339200.0 127800.0 1338000.0 ;
      RECT  126600.0 1339200.0 127800.0 1338000.0 ;
      RECT  129150.0 1339050.0 130050.0 1338150.0 ;
      RECT  124200.0 1331850.0 133800.0 1330950.0 ;
      RECT  124200.0 1345650.0 133800.0 1344750.0 ;
      RECT  135600.0 1343250.0 136800.0 1345650.0 ;
      RECT  135600.0 1334550.0 136800.0 1330950.0 ;
      RECT  140400.0 1334550.0 141600.0 1330950.0 ;
      RECT  142800.0 1333350.0 144000.0 1331400.0 ;
      RECT  142800.0 1345200.0 144000.0 1343250.0 ;
      RECT  135600.0 1334550.0 136800.0 1333350.0 ;
      RECT  138000.0 1334550.0 139200.0 1333350.0 ;
      RECT  138000.0 1334550.0 139200.0 1333350.0 ;
      RECT  135600.0 1334550.0 136800.0 1333350.0 ;
      RECT  138000.0 1334550.0 139200.0 1333350.0 ;
      RECT  140400.0 1334550.0 141600.0 1333350.0 ;
      RECT  140400.0 1334550.0 141600.0 1333350.0 ;
      RECT  138000.0 1334550.0 139200.0 1333350.0 ;
      RECT  135600.0 1343250.0 136800.0 1342050.0 ;
      RECT  138000.0 1343250.0 139200.0 1342050.0 ;
      RECT  138000.0 1343250.0 139200.0 1342050.0 ;
      RECT  135600.0 1343250.0 136800.0 1342050.0 ;
      RECT  138000.0 1343250.0 139200.0 1342050.0 ;
      RECT  140400.0 1343250.0 141600.0 1342050.0 ;
      RECT  140400.0 1343250.0 141600.0 1342050.0 ;
      RECT  138000.0 1343250.0 139200.0 1342050.0 ;
      RECT  142800.0 1333950.0 144000.0 1332750.0 ;
      RECT  142800.0 1343850.0 144000.0 1342650.0 ;
      RECT  140400.0 1340700.0 139200.0 1339500.0 ;
      RECT  137400.0 1338000.0 136200.0 1336800.0 ;
      RECT  138000.0 1334550.0 139200.0 1333350.0 ;
      RECT  140400.0 1343250.0 141600.0 1342050.0 ;
      RECT  141600.0 1338000.0 140400.0 1336800.0 ;
      RECT  136200.0 1338000.0 137400.0 1336800.0 ;
      RECT  139200.0 1340700.0 140400.0 1339500.0 ;
      RECT  140400.0 1338000.0 141600.0 1336800.0 ;
      RECT  133800.0 1331850.0 148200.0 1330950.0 ;
      RECT  133800.0 1345650.0 148200.0 1344750.0 ;
      RECT  154800.0 1333350.0 156000.0 1331400.0 ;
      RECT  154800.0 1345200.0 156000.0 1343250.0 ;
      RECT  150000.0 1343850.0 151200.0 1345650.0 ;
      RECT  150000.0 1334550.0 151200.0 1330950.0 ;
      RECT  152700.0 1343850.0 153600.0 1334550.0 ;
      RECT  150000.0 1334550.0 151200.0 1333350.0 ;
      RECT  152400.0 1334550.0 153600.0 1333350.0 ;
      RECT  152400.0 1334550.0 153600.0 1333350.0 ;
      RECT  150000.0 1334550.0 151200.0 1333350.0 ;
      RECT  150000.0 1343850.0 151200.0 1342650.0 ;
      RECT  152400.0 1343850.0 153600.0 1342650.0 ;
      RECT  152400.0 1343850.0 153600.0 1342650.0 ;
      RECT  150000.0 1343850.0 151200.0 1342650.0 ;
      RECT  154800.0 1333950.0 156000.0 1332750.0 ;
      RECT  154800.0 1343850.0 156000.0 1342650.0 ;
      RECT  150600.0 1339200.0 151800.0 1338000.0 ;
      RECT  150600.0 1339200.0 151800.0 1338000.0 ;
      RECT  153150.0 1339050.0 154050.0 1338150.0 ;
      RECT  148200.0 1331850.0 157800.0 1330950.0 ;
      RECT  148200.0 1345650.0 157800.0 1344750.0 ;
      RECT  120450.0 1338000.0 121650.0 1339200.0 ;
      RECT  122400.0 1340400.0 123600.0 1341600.0 ;
      RECT  139200.0 1339500.0 138000.0 1340700.0 ;
      RECT  130800.0 1357050.0 132000.0 1359000.0 ;
      RECT  130800.0 1345200.0 132000.0 1347150.0 ;
      RECT  126000.0 1346550.0 127200.0 1344750.0 ;
      RECT  126000.0 1355850.0 127200.0 1359450.0 ;
      RECT  128700.0 1346550.0 129600.0 1355850.0 ;
      RECT  126000.0 1355850.0 127200.0 1357050.0 ;
      RECT  128400.0 1355850.0 129600.0 1357050.0 ;
      RECT  128400.0 1355850.0 129600.0 1357050.0 ;
      RECT  126000.0 1355850.0 127200.0 1357050.0 ;
      RECT  126000.0 1346550.0 127200.0 1347750.0 ;
      RECT  128400.0 1346550.0 129600.0 1347750.0 ;
      RECT  128400.0 1346550.0 129600.0 1347750.0 ;
      RECT  126000.0 1346550.0 127200.0 1347750.0 ;
      RECT  130800.0 1356450.0 132000.0 1357650.0 ;
      RECT  130800.0 1346550.0 132000.0 1347750.0 ;
      RECT  126600.0 1351200.0 127800.0 1352400.0 ;
      RECT  126600.0 1351200.0 127800.0 1352400.0 ;
      RECT  129150.0 1351350.0 130050.0 1352250.0 ;
      RECT  124200.0 1358550.0 133800.0 1359450.0 ;
      RECT  124200.0 1344750.0 133800.0 1345650.0 ;
      RECT  135600.0 1347150.0 136800.0 1344750.0 ;
      RECT  135600.0 1355850.0 136800.0 1359450.0 ;
      RECT  140400.0 1355850.0 141600.0 1359450.0 ;
      RECT  142800.0 1357050.0 144000.0 1359000.0 ;
      RECT  142800.0 1345200.0 144000.0 1347150.0 ;
      RECT  135600.0 1355850.0 136800.0 1357050.0 ;
      RECT  138000.0 1355850.0 139200.0 1357050.0 ;
      RECT  138000.0 1355850.0 139200.0 1357050.0 ;
      RECT  135600.0 1355850.0 136800.0 1357050.0 ;
      RECT  138000.0 1355850.0 139200.0 1357050.0 ;
      RECT  140400.0 1355850.0 141600.0 1357050.0 ;
      RECT  140400.0 1355850.0 141600.0 1357050.0 ;
      RECT  138000.0 1355850.0 139200.0 1357050.0 ;
      RECT  135600.0 1347150.0 136800.0 1348350.0 ;
      RECT  138000.0 1347150.0 139200.0 1348350.0 ;
      RECT  138000.0 1347150.0 139200.0 1348350.0 ;
      RECT  135600.0 1347150.0 136800.0 1348350.0 ;
      RECT  138000.0 1347150.0 139200.0 1348350.0 ;
      RECT  140400.0 1347150.0 141600.0 1348350.0 ;
      RECT  140400.0 1347150.0 141600.0 1348350.0 ;
      RECT  138000.0 1347150.0 139200.0 1348350.0 ;
      RECT  142800.0 1356450.0 144000.0 1357650.0 ;
      RECT  142800.0 1346550.0 144000.0 1347750.0 ;
      RECT  140400.0 1349700.0 139200.0 1350900.0 ;
      RECT  137400.0 1352400.0 136200.0 1353600.0 ;
      RECT  138000.0 1355850.0 139200.0 1357050.0 ;
      RECT  140400.0 1347150.0 141600.0 1348350.0 ;
      RECT  141600.0 1352400.0 140400.0 1353600.0 ;
      RECT  136200.0 1352400.0 137400.0 1353600.0 ;
      RECT  139200.0 1349700.0 140400.0 1350900.0 ;
      RECT  140400.0 1352400.0 141600.0 1353600.0 ;
      RECT  133800.0 1358550.0 148200.0 1359450.0 ;
      RECT  133800.0 1344750.0 148200.0 1345650.0 ;
      RECT  154800.0 1357050.0 156000.0 1359000.0 ;
      RECT  154800.0 1345200.0 156000.0 1347150.0 ;
      RECT  150000.0 1346550.0 151200.0 1344750.0 ;
      RECT  150000.0 1355850.0 151200.0 1359450.0 ;
      RECT  152700.0 1346550.0 153600.0 1355850.0 ;
      RECT  150000.0 1355850.0 151200.0 1357050.0 ;
      RECT  152400.0 1355850.0 153600.0 1357050.0 ;
      RECT  152400.0 1355850.0 153600.0 1357050.0 ;
      RECT  150000.0 1355850.0 151200.0 1357050.0 ;
      RECT  150000.0 1346550.0 151200.0 1347750.0 ;
      RECT  152400.0 1346550.0 153600.0 1347750.0 ;
      RECT  152400.0 1346550.0 153600.0 1347750.0 ;
      RECT  150000.0 1346550.0 151200.0 1347750.0 ;
      RECT  154800.0 1356450.0 156000.0 1357650.0 ;
      RECT  154800.0 1346550.0 156000.0 1347750.0 ;
      RECT  150600.0 1351200.0 151800.0 1352400.0 ;
      RECT  150600.0 1351200.0 151800.0 1352400.0 ;
      RECT  153150.0 1351350.0 154050.0 1352250.0 ;
      RECT  148200.0 1358550.0 157800.0 1359450.0 ;
      RECT  148200.0 1344750.0 157800.0 1345650.0 ;
      RECT  120450.0 1351200.0 121650.0 1352400.0 ;
      RECT  122400.0 1348800.0 123600.0 1350000.0 ;
      RECT  139200.0 1349700.0 138000.0 1350900.0 ;
      RECT  130800.0 1360950.0 132000.0 1359000.0 ;
      RECT  130800.0 1372800.0 132000.0 1370850.0 ;
      RECT  126000.0 1371450.0 127200.0 1373250.0 ;
      RECT  126000.0 1362150.0 127200.0 1358550.0 ;
      RECT  128700.0 1371450.0 129600.0 1362150.0 ;
      RECT  126000.0 1362150.0 127200.0 1360950.0 ;
      RECT  128400.0 1362150.0 129600.0 1360950.0 ;
      RECT  128400.0 1362150.0 129600.0 1360950.0 ;
      RECT  126000.0 1362150.0 127200.0 1360950.0 ;
      RECT  126000.0 1371450.0 127200.0 1370250.0 ;
      RECT  128400.0 1371450.0 129600.0 1370250.0 ;
      RECT  128400.0 1371450.0 129600.0 1370250.0 ;
      RECT  126000.0 1371450.0 127200.0 1370250.0 ;
      RECT  130800.0 1361550.0 132000.0 1360350.0 ;
      RECT  130800.0 1371450.0 132000.0 1370250.0 ;
      RECT  126600.0 1366800.0 127800.0 1365600.0 ;
      RECT  126600.0 1366800.0 127800.0 1365600.0 ;
      RECT  129150.0 1366650.0 130050.0 1365750.0 ;
      RECT  124200.0 1359450.0 133800.0 1358550.0 ;
      RECT  124200.0 1373250.0 133800.0 1372350.0 ;
      RECT  135600.0 1370850.0 136800.0 1373250.0 ;
      RECT  135600.0 1362150.0 136800.0 1358550.0 ;
      RECT  140400.0 1362150.0 141600.0 1358550.0 ;
      RECT  142800.0 1360950.0 144000.0 1359000.0 ;
      RECT  142800.0 1372800.0 144000.0 1370850.0 ;
      RECT  135600.0 1362150.0 136800.0 1360950.0 ;
      RECT  138000.0 1362150.0 139200.0 1360950.0 ;
      RECT  138000.0 1362150.0 139200.0 1360950.0 ;
      RECT  135600.0 1362150.0 136800.0 1360950.0 ;
      RECT  138000.0 1362150.0 139200.0 1360950.0 ;
      RECT  140400.0 1362150.0 141600.0 1360950.0 ;
      RECT  140400.0 1362150.0 141600.0 1360950.0 ;
      RECT  138000.0 1362150.0 139200.0 1360950.0 ;
      RECT  135600.0 1370850.0 136800.0 1369650.0 ;
      RECT  138000.0 1370850.0 139200.0 1369650.0 ;
      RECT  138000.0 1370850.0 139200.0 1369650.0 ;
      RECT  135600.0 1370850.0 136800.0 1369650.0 ;
      RECT  138000.0 1370850.0 139200.0 1369650.0 ;
      RECT  140400.0 1370850.0 141600.0 1369650.0 ;
      RECT  140400.0 1370850.0 141600.0 1369650.0 ;
      RECT  138000.0 1370850.0 139200.0 1369650.0 ;
      RECT  142800.0 1361550.0 144000.0 1360350.0 ;
      RECT  142800.0 1371450.0 144000.0 1370250.0 ;
      RECT  140400.0 1368300.0 139200.0 1367100.0 ;
      RECT  137400.0 1365600.0 136200.0 1364400.0 ;
      RECT  138000.0 1362150.0 139200.0 1360950.0 ;
      RECT  140400.0 1370850.0 141600.0 1369650.0 ;
      RECT  141600.0 1365600.0 140400.0 1364400.0 ;
      RECT  136200.0 1365600.0 137400.0 1364400.0 ;
      RECT  139200.0 1368300.0 140400.0 1367100.0 ;
      RECT  140400.0 1365600.0 141600.0 1364400.0 ;
      RECT  133800.0 1359450.0 148200.0 1358550.0 ;
      RECT  133800.0 1373250.0 148200.0 1372350.0 ;
      RECT  154800.0 1360950.0 156000.0 1359000.0 ;
      RECT  154800.0 1372800.0 156000.0 1370850.0 ;
      RECT  150000.0 1371450.0 151200.0 1373250.0 ;
      RECT  150000.0 1362150.0 151200.0 1358550.0 ;
      RECT  152700.0 1371450.0 153600.0 1362150.0 ;
      RECT  150000.0 1362150.0 151200.0 1360950.0 ;
      RECT  152400.0 1362150.0 153600.0 1360950.0 ;
      RECT  152400.0 1362150.0 153600.0 1360950.0 ;
      RECT  150000.0 1362150.0 151200.0 1360950.0 ;
      RECT  150000.0 1371450.0 151200.0 1370250.0 ;
      RECT  152400.0 1371450.0 153600.0 1370250.0 ;
      RECT  152400.0 1371450.0 153600.0 1370250.0 ;
      RECT  150000.0 1371450.0 151200.0 1370250.0 ;
      RECT  154800.0 1361550.0 156000.0 1360350.0 ;
      RECT  154800.0 1371450.0 156000.0 1370250.0 ;
      RECT  150600.0 1366800.0 151800.0 1365600.0 ;
      RECT  150600.0 1366800.0 151800.0 1365600.0 ;
      RECT  153150.0 1366650.0 154050.0 1365750.0 ;
      RECT  148200.0 1359450.0 157800.0 1358550.0 ;
      RECT  148200.0 1373250.0 157800.0 1372350.0 ;
      RECT  120450.0 1365600.0 121650.0 1366800.0 ;
      RECT  122400.0 1368000.0 123600.0 1369200.0 ;
      RECT  139200.0 1367100.0 138000.0 1368300.0 ;
      RECT  130800.0 1384650.0 132000.0 1386600.0 ;
      RECT  130800.0 1372800.0 132000.0 1374750.0 ;
      RECT  126000.0 1374150.0 127200.0 1372350.0 ;
      RECT  126000.0 1383450.0 127200.0 1387050.0 ;
      RECT  128700.0 1374150.0 129600.0 1383450.0 ;
      RECT  126000.0 1383450.0 127200.0 1384650.0 ;
      RECT  128400.0 1383450.0 129600.0 1384650.0 ;
      RECT  128400.0 1383450.0 129600.0 1384650.0 ;
      RECT  126000.0 1383450.0 127200.0 1384650.0 ;
      RECT  126000.0 1374150.0 127200.0 1375350.0 ;
      RECT  128400.0 1374150.0 129600.0 1375350.0 ;
      RECT  128400.0 1374150.0 129600.0 1375350.0 ;
      RECT  126000.0 1374150.0 127200.0 1375350.0 ;
      RECT  130800.0 1384050.0 132000.0 1385250.0 ;
      RECT  130800.0 1374150.0 132000.0 1375350.0 ;
      RECT  126600.0 1378800.0 127800.0 1380000.0 ;
      RECT  126600.0 1378800.0 127800.0 1380000.0 ;
      RECT  129150.0 1378950.0 130050.0 1379850.0 ;
      RECT  124200.0 1386150.0 133800.0 1387050.0 ;
      RECT  124200.0 1372350.0 133800.0 1373250.0 ;
      RECT  135600.0 1374750.0 136800.0 1372350.0 ;
      RECT  135600.0 1383450.0 136800.0 1387050.0 ;
      RECT  140400.0 1383450.0 141600.0 1387050.0 ;
      RECT  142800.0 1384650.0 144000.0 1386600.0 ;
      RECT  142800.0 1372800.0 144000.0 1374750.0 ;
      RECT  135600.0 1383450.0 136800.0 1384650.0 ;
      RECT  138000.0 1383450.0 139200.0 1384650.0 ;
      RECT  138000.0 1383450.0 139200.0 1384650.0 ;
      RECT  135600.0 1383450.0 136800.0 1384650.0 ;
      RECT  138000.0 1383450.0 139200.0 1384650.0 ;
      RECT  140400.0 1383450.0 141600.0 1384650.0 ;
      RECT  140400.0 1383450.0 141600.0 1384650.0 ;
      RECT  138000.0 1383450.0 139200.0 1384650.0 ;
      RECT  135600.0 1374750.0 136800.0 1375950.0 ;
      RECT  138000.0 1374750.0 139200.0 1375950.0 ;
      RECT  138000.0 1374750.0 139200.0 1375950.0 ;
      RECT  135600.0 1374750.0 136800.0 1375950.0 ;
      RECT  138000.0 1374750.0 139200.0 1375950.0 ;
      RECT  140400.0 1374750.0 141600.0 1375950.0 ;
      RECT  140400.0 1374750.0 141600.0 1375950.0 ;
      RECT  138000.0 1374750.0 139200.0 1375950.0 ;
      RECT  142800.0 1384050.0 144000.0 1385250.0 ;
      RECT  142800.0 1374150.0 144000.0 1375350.0 ;
      RECT  140400.0 1377300.0 139200.0 1378500.0 ;
      RECT  137400.0 1380000.0 136200.0 1381200.0 ;
      RECT  138000.0 1383450.0 139200.0 1384650.0 ;
      RECT  140400.0 1374750.0 141600.0 1375950.0 ;
      RECT  141600.0 1380000.0 140400.0 1381200.0 ;
      RECT  136200.0 1380000.0 137400.0 1381200.0 ;
      RECT  139200.0 1377300.0 140400.0 1378500.0 ;
      RECT  140400.0 1380000.0 141600.0 1381200.0 ;
      RECT  133800.0 1386150.0 148200.0 1387050.0 ;
      RECT  133800.0 1372350.0 148200.0 1373250.0 ;
      RECT  154800.0 1384650.0 156000.0 1386600.0 ;
      RECT  154800.0 1372800.0 156000.0 1374750.0 ;
      RECT  150000.0 1374150.0 151200.0 1372350.0 ;
      RECT  150000.0 1383450.0 151200.0 1387050.0 ;
      RECT  152700.0 1374150.0 153600.0 1383450.0 ;
      RECT  150000.0 1383450.0 151200.0 1384650.0 ;
      RECT  152400.0 1383450.0 153600.0 1384650.0 ;
      RECT  152400.0 1383450.0 153600.0 1384650.0 ;
      RECT  150000.0 1383450.0 151200.0 1384650.0 ;
      RECT  150000.0 1374150.0 151200.0 1375350.0 ;
      RECT  152400.0 1374150.0 153600.0 1375350.0 ;
      RECT  152400.0 1374150.0 153600.0 1375350.0 ;
      RECT  150000.0 1374150.0 151200.0 1375350.0 ;
      RECT  154800.0 1384050.0 156000.0 1385250.0 ;
      RECT  154800.0 1374150.0 156000.0 1375350.0 ;
      RECT  150600.0 1378800.0 151800.0 1380000.0 ;
      RECT  150600.0 1378800.0 151800.0 1380000.0 ;
      RECT  153150.0 1378950.0 154050.0 1379850.0 ;
      RECT  148200.0 1386150.0 157800.0 1387050.0 ;
      RECT  148200.0 1372350.0 157800.0 1373250.0 ;
      RECT  120450.0 1378800.0 121650.0 1380000.0 ;
      RECT  122400.0 1376400.0 123600.0 1377600.0 ;
      RECT  139200.0 1377300.0 138000.0 1378500.0 ;
      RECT  130800.0 1388550.0 132000.0 1386600.0 ;
      RECT  130800.0 1400400.0 132000.0 1398450.0 ;
      RECT  126000.0 1399050.0 127200.0 1400850.0 ;
      RECT  126000.0 1389750.0 127200.0 1386150.0 ;
      RECT  128700.0 1399050.0 129600.0 1389750.0 ;
      RECT  126000.0 1389750.0 127200.0 1388550.0 ;
      RECT  128400.0 1389750.0 129600.0 1388550.0 ;
      RECT  128400.0 1389750.0 129600.0 1388550.0 ;
      RECT  126000.0 1389750.0 127200.0 1388550.0 ;
      RECT  126000.0 1399050.0 127200.0 1397850.0 ;
      RECT  128400.0 1399050.0 129600.0 1397850.0 ;
      RECT  128400.0 1399050.0 129600.0 1397850.0 ;
      RECT  126000.0 1399050.0 127200.0 1397850.0 ;
      RECT  130800.0 1389150.0 132000.0 1387950.0 ;
      RECT  130800.0 1399050.0 132000.0 1397850.0 ;
      RECT  126600.0 1394400.0 127800.0 1393200.0 ;
      RECT  126600.0 1394400.0 127800.0 1393200.0 ;
      RECT  129150.0 1394250.0 130050.0 1393350.0 ;
      RECT  124200.0 1387050.0 133800.0 1386150.0 ;
      RECT  124200.0 1400850.0 133800.0 1399950.0 ;
      RECT  135600.0 1398450.0 136800.0 1400850.0 ;
      RECT  135600.0 1389750.0 136800.0 1386150.0 ;
      RECT  140400.0 1389750.0 141600.0 1386150.0 ;
      RECT  142800.0 1388550.0 144000.0 1386600.0 ;
      RECT  142800.0 1400400.0 144000.0 1398450.0 ;
      RECT  135600.0 1389750.0 136800.0 1388550.0 ;
      RECT  138000.0 1389750.0 139200.0 1388550.0 ;
      RECT  138000.0 1389750.0 139200.0 1388550.0 ;
      RECT  135600.0 1389750.0 136800.0 1388550.0 ;
      RECT  138000.0 1389750.0 139200.0 1388550.0 ;
      RECT  140400.0 1389750.0 141600.0 1388550.0 ;
      RECT  140400.0 1389750.0 141600.0 1388550.0 ;
      RECT  138000.0 1389750.0 139200.0 1388550.0 ;
      RECT  135600.0 1398450.0 136800.0 1397250.0 ;
      RECT  138000.0 1398450.0 139200.0 1397250.0 ;
      RECT  138000.0 1398450.0 139200.0 1397250.0 ;
      RECT  135600.0 1398450.0 136800.0 1397250.0 ;
      RECT  138000.0 1398450.0 139200.0 1397250.0 ;
      RECT  140400.0 1398450.0 141600.0 1397250.0 ;
      RECT  140400.0 1398450.0 141600.0 1397250.0 ;
      RECT  138000.0 1398450.0 139200.0 1397250.0 ;
      RECT  142800.0 1389150.0 144000.0 1387950.0 ;
      RECT  142800.0 1399050.0 144000.0 1397850.0 ;
      RECT  140400.0 1395900.0 139200.0 1394700.0 ;
      RECT  137400.0 1393200.0 136200.0 1392000.0 ;
      RECT  138000.0 1389750.0 139200.0 1388550.0 ;
      RECT  140400.0 1398450.0 141600.0 1397250.0 ;
      RECT  141600.0 1393200.0 140400.0 1392000.0 ;
      RECT  136200.0 1393200.0 137400.0 1392000.0 ;
      RECT  139200.0 1395900.0 140400.0 1394700.0 ;
      RECT  140400.0 1393200.0 141600.0 1392000.0 ;
      RECT  133800.0 1387050.0 148200.0 1386150.0 ;
      RECT  133800.0 1400850.0 148200.0 1399950.0 ;
      RECT  154800.0 1388550.0 156000.0 1386600.0 ;
      RECT  154800.0 1400400.0 156000.0 1398450.0 ;
      RECT  150000.0 1399050.0 151200.0 1400850.0 ;
      RECT  150000.0 1389750.0 151200.0 1386150.0 ;
      RECT  152700.0 1399050.0 153600.0 1389750.0 ;
      RECT  150000.0 1389750.0 151200.0 1388550.0 ;
      RECT  152400.0 1389750.0 153600.0 1388550.0 ;
      RECT  152400.0 1389750.0 153600.0 1388550.0 ;
      RECT  150000.0 1389750.0 151200.0 1388550.0 ;
      RECT  150000.0 1399050.0 151200.0 1397850.0 ;
      RECT  152400.0 1399050.0 153600.0 1397850.0 ;
      RECT  152400.0 1399050.0 153600.0 1397850.0 ;
      RECT  150000.0 1399050.0 151200.0 1397850.0 ;
      RECT  154800.0 1389150.0 156000.0 1387950.0 ;
      RECT  154800.0 1399050.0 156000.0 1397850.0 ;
      RECT  150600.0 1394400.0 151800.0 1393200.0 ;
      RECT  150600.0 1394400.0 151800.0 1393200.0 ;
      RECT  153150.0 1394250.0 154050.0 1393350.0 ;
      RECT  148200.0 1387050.0 157800.0 1386150.0 ;
      RECT  148200.0 1400850.0 157800.0 1399950.0 ;
      RECT  120450.0 1393200.0 121650.0 1394400.0 ;
      RECT  122400.0 1395600.0 123600.0 1396800.0 ;
      RECT  139200.0 1394700.0 138000.0 1395900.0 ;
      RECT  130800.0 1412250.0 132000.0 1414200.0 ;
      RECT  130800.0 1400400.0 132000.0 1402350.0 ;
      RECT  126000.0 1401750.0 127200.0 1399950.0 ;
      RECT  126000.0 1411050.0 127200.0 1414650.0 ;
      RECT  128700.0 1401750.0 129600.0 1411050.0 ;
      RECT  126000.0 1411050.0 127200.0 1412250.0 ;
      RECT  128400.0 1411050.0 129600.0 1412250.0 ;
      RECT  128400.0 1411050.0 129600.0 1412250.0 ;
      RECT  126000.0 1411050.0 127200.0 1412250.0 ;
      RECT  126000.0 1401750.0 127200.0 1402950.0 ;
      RECT  128400.0 1401750.0 129600.0 1402950.0 ;
      RECT  128400.0 1401750.0 129600.0 1402950.0 ;
      RECT  126000.0 1401750.0 127200.0 1402950.0 ;
      RECT  130800.0 1411650.0 132000.0 1412850.0 ;
      RECT  130800.0 1401750.0 132000.0 1402950.0 ;
      RECT  126600.0 1406400.0 127800.0 1407600.0 ;
      RECT  126600.0 1406400.0 127800.0 1407600.0 ;
      RECT  129150.0 1406550.0 130050.0 1407450.0 ;
      RECT  124200.0 1413750.0 133800.0 1414650.0 ;
      RECT  124200.0 1399950.0 133800.0 1400850.0 ;
      RECT  135600.0 1402350.0 136800.0 1399950.0 ;
      RECT  135600.0 1411050.0 136800.0 1414650.0 ;
      RECT  140400.0 1411050.0 141600.0 1414650.0 ;
      RECT  142800.0 1412250.0 144000.0 1414200.0 ;
      RECT  142800.0 1400400.0 144000.0 1402350.0 ;
      RECT  135600.0 1411050.0 136800.0 1412250.0 ;
      RECT  138000.0 1411050.0 139200.0 1412250.0 ;
      RECT  138000.0 1411050.0 139200.0 1412250.0 ;
      RECT  135600.0 1411050.0 136800.0 1412250.0 ;
      RECT  138000.0 1411050.0 139200.0 1412250.0 ;
      RECT  140400.0 1411050.0 141600.0 1412250.0 ;
      RECT  140400.0 1411050.0 141600.0 1412250.0 ;
      RECT  138000.0 1411050.0 139200.0 1412250.0 ;
      RECT  135600.0 1402350.0 136800.0 1403550.0 ;
      RECT  138000.0 1402350.0 139200.0 1403550.0 ;
      RECT  138000.0 1402350.0 139200.0 1403550.0 ;
      RECT  135600.0 1402350.0 136800.0 1403550.0 ;
      RECT  138000.0 1402350.0 139200.0 1403550.0 ;
      RECT  140400.0 1402350.0 141600.0 1403550.0 ;
      RECT  140400.0 1402350.0 141600.0 1403550.0 ;
      RECT  138000.0 1402350.0 139200.0 1403550.0 ;
      RECT  142800.0 1411650.0 144000.0 1412850.0 ;
      RECT  142800.0 1401750.0 144000.0 1402950.0 ;
      RECT  140400.0 1404900.0 139200.0 1406100.0 ;
      RECT  137400.0 1407600.0 136200.0 1408800.0 ;
      RECT  138000.0 1411050.0 139200.0 1412250.0 ;
      RECT  140400.0 1402350.0 141600.0 1403550.0 ;
      RECT  141600.0 1407600.0 140400.0 1408800.0 ;
      RECT  136200.0 1407600.0 137400.0 1408800.0 ;
      RECT  139200.0 1404900.0 140400.0 1406100.0 ;
      RECT  140400.0 1407600.0 141600.0 1408800.0 ;
      RECT  133800.0 1413750.0 148200.0 1414650.0 ;
      RECT  133800.0 1399950.0 148200.0 1400850.0 ;
      RECT  154800.0 1412250.0 156000.0 1414200.0 ;
      RECT  154800.0 1400400.0 156000.0 1402350.0 ;
      RECT  150000.0 1401750.0 151200.0 1399950.0 ;
      RECT  150000.0 1411050.0 151200.0 1414650.0 ;
      RECT  152700.0 1401750.0 153600.0 1411050.0 ;
      RECT  150000.0 1411050.0 151200.0 1412250.0 ;
      RECT  152400.0 1411050.0 153600.0 1412250.0 ;
      RECT  152400.0 1411050.0 153600.0 1412250.0 ;
      RECT  150000.0 1411050.0 151200.0 1412250.0 ;
      RECT  150000.0 1401750.0 151200.0 1402950.0 ;
      RECT  152400.0 1401750.0 153600.0 1402950.0 ;
      RECT  152400.0 1401750.0 153600.0 1402950.0 ;
      RECT  150000.0 1401750.0 151200.0 1402950.0 ;
      RECT  154800.0 1411650.0 156000.0 1412850.0 ;
      RECT  154800.0 1401750.0 156000.0 1402950.0 ;
      RECT  150600.0 1406400.0 151800.0 1407600.0 ;
      RECT  150600.0 1406400.0 151800.0 1407600.0 ;
      RECT  153150.0 1406550.0 154050.0 1407450.0 ;
      RECT  148200.0 1413750.0 157800.0 1414650.0 ;
      RECT  148200.0 1399950.0 157800.0 1400850.0 ;
      RECT  120450.0 1406400.0 121650.0 1407600.0 ;
      RECT  122400.0 1404000.0 123600.0 1405200.0 ;
      RECT  139200.0 1404900.0 138000.0 1406100.0 ;
      RECT  130800.0 1416150.0 132000.0 1414200.0 ;
      RECT  130800.0 1428000.0 132000.0 1426050.0 ;
      RECT  126000.0 1426650.0 127200.0 1428450.0 ;
      RECT  126000.0 1417350.0 127200.0 1413750.0 ;
      RECT  128700.0 1426650.0 129600.0 1417350.0 ;
      RECT  126000.0 1417350.0 127200.0 1416150.0 ;
      RECT  128400.0 1417350.0 129600.0 1416150.0 ;
      RECT  128400.0 1417350.0 129600.0 1416150.0 ;
      RECT  126000.0 1417350.0 127200.0 1416150.0 ;
      RECT  126000.0 1426650.0 127200.0 1425450.0 ;
      RECT  128400.0 1426650.0 129600.0 1425450.0 ;
      RECT  128400.0 1426650.0 129600.0 1425450.0 ;
      RECT  126000.0 1426650.0 127200.0 1425450.0 ;
      RECT  130800.0 1416750.0 132000.0 1415550.0 ;
      RECT  130800.0 1426650.0 132000.0 1425450.0 ;
      RECT  126600.0 1422000.0 127800.0 1420800.0 ;
      RECT  126600.0 1422000.0 127800.0 1420800.0 ;
      RECT  129150.0 1421850.0 130050.0 1420950.0 ;
      RECT  124200.0 1414650.0 133800.0 1413750.0 ;
      RECT  124200.0 1428450.0 133800.0 1427550.0 ;
      RECT  135600.0 1426050.0 136800.0 1428450.0 ;
      RECT  135600.0 1417350.0 136800.0 1413750.0 ;
      RECT  140400.0 1417350.0 141600.0 1413750.0 ;
      RECT  142800.0 1416150.0 144000.0 1414200.0 ;
      RECT  142800.0 1428000.0 144000.0 1426050.0 ;
      RECT  135600.0 1417350.0 136800.0 1416150.0 ;
      RECT  138000.0 1417350.0 139200.0 1416150.0 ;
      RECT  138000.0 1417350.0 139200.0 1416150.0 ;
      RECT  135600.0 1417350.0 136800.0 1416150.0 ;
      RECT  138000.0 1417350.0 139200.0 1416150.0 ;
      RECT  140400.0 1417350.0 141600.0 1416150.0 ;
      RECT  140400.0 1417350.0 141600.0 1416150.0 ;
      RECT  138000.0 1417350.0 139200.0 1416150.0 ;
      RECT  135600.0 1426050.0 136800.0 1424850.0 ;
      RECT  138000.0 1426050.0 139200.0 1424850.0 ;
      RECT  138000.0 1426050.0 139200.0 1424850.0 ;
      RECT  135600.0 1426050.0 136800.0 1424850.0 ;
      RECT  138000.0 1426050.0 139200.0 1424850.0 ;
      RECT  140400.0 1426050.0 141600.0 1424850.0 ;
      RECT  140400.0 1426050.0 141600.0 1424850.0 ;
      RECT  138000.0 1426050.0 139200.0 1424850.0 ;
      RECT  142800.0 1416750.0 144000.0 1415550.0 ;
      RECT  142800.0 1426650.0 144000.0 1425450.0 ;
      RECT  140400.0 1423500.0 139200.0 1422300.0 ;
      RECT  137400.0 1420800.0 136200.0 1419600.0 ;
      RECT  138000.0 1417350.0 139200.0 1416150.0 ;
      RECT  140400.0 1426050.0 141600.0 1424850.0 ;
      RECT  141600.0 1420800.0 140400.0 1419600.0 ;
      RECT  136200.0 1420800.0 137400.0 1419600.0 ;
      RECT  139200.0 1423500.0 140400.0 1422300.0 ;
      RECT  140400.0 1420800.0 141600.0 1419600.0 ;
      RECT  133800.0 1414650.0 148200.0 1413750.0 ;
      RECT  133800.0 1428450.0 148200.0 1427550.0 ;
      RECT  154800.0 1416150.0 156000.0 1414200.0 ;
      RECT  154800.0 1428000.0 156000.0 1426050.0 ;
      RECT  150000.0 1426650.0 151200.0 1428450.0 ;
      RECT  150000.0 1417350.0 151200.0 1413750.0 ;
      RECT  152700.0 1426650.0 153600.0 1417350.0 ;
      RECT  150000.0 1417350.0 151200.0 1416150.0 ;
      RECT  152400.0 1417350.0 153600.0 1416150.0 ;
      RECT  152400.0 1417350.0 153600.0 1416150.0 ;
      RECT  150000.0 1417350.0 151200.0 1416150.0 ;
      RECT  150000.0 1426650.0 151200.0 1425450.0 ;
      RECT  152400.0 1426650.0 153600.0 1425450.0 ;
      RECT  152400.0 1426650.0 153600.0 1425450.0 ;
      RECT  150000.0 1426650.0 151200.0 1425450.0 ;
      RECT  154800.0 1416750.0 156000.0 1415550.0 ;
      RECT  154800.0 1426650.0 156000.0 1425450.0 ;
      RECT  150600.0 1422000.0 151800.0 1420800.0 ;
      RECT  150600.0 1422000.0 151800.0 1420800.0 ;
      RECT  153150.0 1421850.0 154050.0 1420950.0 ;
      RECT  148200.0 1414650.0 157800.0 1413750.0 ;
      RECT  148200.0 1428450.0 157800.0 1427550.0 ;
      RECT  120450.0 1420800.0 121650.0 1422000.0 ;
      RECT  122400.0 1423200.0 123600.0 1424400.0 ;
      RECT  139200.0 1422300.0 138000.0 1423500.0 ;
      RECT  130800.0 1439850.0 132000.0 1441800.0 ;
      RECT  130800.0 1428000.0 132000.0 1429950.0 ;
      RECT  126000.0 1429350.0 127200.0 1427550.0 ;
      RECT  126000.0 1438650.0 127200.0 1442250.0 ;
      RECT  128700.0 1429350.0 129600.0 1438650.0 ;
      RECT  126000.0 1438650.0 127200.0 1439850.0 ;
      RECT  128400.0 1438650.0 129600.0 1439850.0 ;
      RECT  128400.0 1438650.0 129600.0 1439850.0 ;
      RECT  126000.0 1438650.0 127200.0 1439850.0 ;
      RECT  126000.0 1429350.0 127200.0 1430550.0 ;
      RECT  128400.0 1429350.0 129600.0 1430550.0 ;
      RECT  128400.0 1429350.0 129600.0 1430550.0 ;
      RECT  126000.0 1429350.0 127200.0 1430550.0 ;
      RECT  130800.0 1439250.0 132000.0 1440450.0 ;
      RECT  130800.0 1429350.0 132000.0 1430550.0 ;
      RECT  126600.0 1434000.0 127800.0 1435200.0 ;
      RECT  126600.0 1434000.0 127800.0 1435200.0 ;
      RECT  129150.0 1434150.0 130050.0 1435050.0 ;
      RECT  124200.0 1441350.0 133800.0 1442250.0 ;
      RECT  124200.0 1427550.0 133800.0 1428450.0 ;
      RECT  135600.0 1429950.0 136800.0 1427550.0 ;
      RECT  135600.0 1438650.0 136800.0 1442250.0 ;
      RECT  140400.0 1438650.0 141600.0 1442250.0 ;
      RECT  142800.0 1439850.0 144000.0 1441800.0 ;
      RECT  142800.0 1428000.0 144000.0 1429950.0 ;
      RECT  135600.0 1438650.0 136800.0 1439850.0 ;
      RECT  138000.0 1438650.0 139200.0 1439850.0 ;
      RECT  138000.0 1438650.0 139200.0 1439850.0 ;
      RECT  135600.0 1438650.0 136800.0 1439850.0 ;
      RECT  138000.0 1438650.0 139200.0 1439850.0 ;
      RECT  140400.0 1438650.0 141600.0 1439850.0 ;
      RECT  140400.0 1438650.0 141600.0 1439850.0 ;
      RECT  138000.0 1438650.0 139200.0 1439850.0 ;
      RECT  135600.0 1429950.0 136800.0 1431150.0 ;
      RECT  138000.0 1429950.0 139200.0 1431150.0 ;
      RECT  138000.0 1429950.0 139200.0 1431150.0 ;
      RECT  135600.0 1429950.0 136800.0 1431150.0 ;
      RECT  138000.0 1429950.0 139200.0 1431150.0 ;
      RECT  140400.0 1429950.0 141600.0 1431150.0 ;
      RECT  140400.0 1429950.0 141600.0 1431150.0 ;
      RECT  138000.0 1429950.0 139200.0 1431150.0 ;
      RECT  142800.0 1439250.0 144000.0 1440450.0 ;
      RECT  142800.0 1429350.0 144000.0 1430550.0 ;
      RECT  140400.0 1432500.0 139200.0 1433700.0 ;
      RECT  137400.0 1435200.0 136200.0 1436400.0 ;
      RECT  138000.0 1438650.0 139200.0 1439850.0 ;
      RECT  140400.0 1429950.0 141600.0 1431150.0 ;
      RECT  141600.0 1435200.0 140400.0 1436400.0 ;
      RECT  136200.0 1435200.0 137400.0 1436400.0 ;
      RECT  139200.0 1432500.0 140400.0 1433700.0 ;
      RECT  140400.0 1435200.0 141600.0 1436400.0 ;
      RECT  133800.0 1441350.0 148200.0 1442250.0 ;
      RECT  133800.0 1427550.0 148200.0 1428450.0 ;
      RECT  154800.0 1439850.0 156000.0 1441800.0 ;
      RECT  154800.0 1428000.0 156000.0 1429950.0 ;
      RECT  150000.0 1429350.0 151200.0 1427550.0 ;
      RECT  150000.0 1438650.0 151200.0 1442250.0 ;
      RECT  152700.0 1429350.0 153600.0 1438650.0 ;
      RECT  150000.0 1438650.0 151200.0 1439850.0 ;
      RECT  152400.0 1438650.0 153600.0 1439850.0 ;
      RECT  152400.0 1438650.0 153600.0 1439850.0 ;
      RECT  150000.0 1438650.0 151200.0 1439850.0 ;
      RECT  150000.0 1429350.0 151200.0 1430550.0 ;
      RECT  152400.0 1429350.0 153600.0 1430550.0 ;
      RECT  152400.0 1429350.0 153600.0 1430550.0 ;
      RECT  150000.0 1429350.0 151200.0 1430550.0 ;
      RECT  154800.0 1439250.0 156000.0 1440450.0 ;
      RECT  154800.0 1429350.0 156000.0 1430550.0 ;
      RECT  150600.0 1434000.0 151800.0 1435200.0 ;
      RECT  150600.0 1434000.0 151800.0 1435200.0 ;
      RECT  153150.0 1434150.0 154050.0 1435050.0 ;
      RECT  148200.0 1441350.0 157800.0 1442250.0 ;
      RECT  148200.0 1427550.0 157800.0 1428450.0 ;
      RECT  120450.0 1434000.0 121650.0 1435200.0 ;
      RECT  122400.0 1431600.0 123600.0 1432800.0 ;
      RECT  139200.0 1432500.0 138000.0 1433700.0 ;
      RECT  130800.0 1443750.0 132000.0 1441800.0 ;
      RECT  130800.0 1455600.0 132000.0 1453650.0 ;
      RECT  126000.0 1454250.0 127200.0 1456050.0 ;
      RECT  126000.0 1444950.0 127200.0 1441350.0 ;
      RECT  128700.0 1454250.0 129600.0 1444950.0 ;
      RECT  126000.0 1444950.0 127200.0 1443750.0 ;
      RECT  128400.0 1444950.0 129600.0 1443750.0 ;
      RECT  128400.0 1444950.0 129600.0 1443750.0 ;
      RECT  126000.0 1444950.0 127200.0 1443750.0 ;
      RECT  126000.0 1454250.0 127200.0 1453050.0 ;
      RECT  128400.0 1454250.0 129600.0 1453050.0 ;
      RECT  128400.0 1454250.0 129600.0 1453050.0 ;
      RECT  126000.0 1454250.0 127200.0 1453050.0 ;
      RECT  130800.0 1444350.0 132000.0 1443150.0 ;
      RECT  130800.0 1454250.0 132000.0 1453050.0 ;
      RECT  126600.0 1449600.0 127800.0 1448400.0 ;
      RECT  126600.0 1449600.0 127800.0 1448400.0 ;
      RECT  129150.0 1449450.0 130050.0 1448550.0 ;
      RECT  124200.0 1442250.0 133800.0 1441350.0 ;
      RECT  124200.0 1456050.0 133800.0 1455150.0 ;
      RECT  135600.0 1453650.0 136800.0 1456050.0 ;
      RECT  135600.0 1444950.0 136800.0 1441350.0 ;
      RECT  140400.0 1444950.0 141600.0 1441350.0 ;
      RECT  142800.0 1443750.0 144000.0 1441800.0 ;
      RECT  142800.0 1455600.0 144000.0 1453650.0 ;
      RECT  135600.0 1444950.0 136800.0 1443750.0 ;
      RECT  138000.0 1444950.0 139200.0 1443750.0 ;
      RECT  138000.0 1444950.0 139200.0 1443750.0 ;
      RECT  135600.0 1444950.0 136800.0 1443750.0 ;
      RECT  138000.0 1444950.0 139200.0 1443750.0 ;
      RECT  140400.0 1444950.0 141600.0 1443750.0 ;
      RECT  140400.0 1444950.0 141600.0 1443750.0 ;
      RECT  138000.0 1444950.0 139200.0 1443750.0 ;
      RECT  135600.0 1453650.0 136800.0 1452450.0 ;
      RECT  138000.0 1453650.0 139200.0 1452450.0 ;
      RECT  138000.0 1453650.0 139200.0 1452450.0 ;
      RECT  135600.0 1453650.0 136800.0 1452450.0 ;
      RECT  138000.0 1453650.0 139200.0 1452450.0 ;
      RECT  140400.0 1453650.0 141600.0 1452450.0 ;
      RECT  140400.0 1453650.0 141600.0 1452450.0 ;
      RECT  138000.0 1453650.0 139200.0 1452450.0 ;
      RECT  142800.0 1444350.0 144000.0 1443150.0 ;
      RECT  142800.0 1454250.0 144000.0 1453050.0 ;
      RECT  140400.0 1451100.0 139200.0 1449900.0 ;
      RECT  137400.0 1448400.0 136200.0 1447200.0 ;
      RECT  138000.0 1444950.0 139200.0 1443750.0 ;
      RECT  140400.0 1453650.0 141600.0 1452450.0 ;
      RECT  141600.0 1448400.0 140400.0 1447200.0 ;
      RECT  136200.0 1448400.0 137400.0 1447200.0 ;
      RECT  139200.0 1451100.0 140400.0 1449900.0 ;
      RECT  140400.0 1448400.0 141600.0 1447200.0 ;
      RECT  133800.0 1442250.0 148200.0 1441350.0 ;
      RECT  133800.0 1456050.0 148200.0 1455150.0 ;
      RECT  154800.0 1443750.0 156000.0 1441800.0 ;
      RECT  154800.0 1455600.0 156000.0 1453650.0 ;
      RECT  150000.0 1454250.0 151200.0 1456050.0 ;
      RECT  150000.0 1444950.0 151200.0 1441350.0 ;
      RECT  152700.0 1454250.0 153600.0 1444950.0 ;
      RECT  150000.0 1444950.0 151200.0 1443750.0 ;
      RECT  152400.0 1444950.0 153600.0 1443750.0 ;
      RECT  152400.0 1444950.0 153600.0 1443750.0 ;
      RECT  150000.0 1444950.0 151200.0 1443750.0 ;
      RECT  150000.0 1454250.0 151200.0 1453050.0 ;
      RECT  152400.0 1454250.0 153600.0 1453050.0 ;
      RECT  152400.0 1454250.0 153600.0 1453050.0 ;
      RECT  150000.0 1454250.0 151200.0 1453050.0 ;
      RECT  154800.0 1444350.0 156000.0 1443150.0 ;
      RECT  154800.0 1454250.0 156000.0 1453050.0 ;
      RECT  150600.0 1449600.0 151800.0 1448400.0 ;
      RECT  150600.0 1449600.0 151800.0 1448400.0 ;
      RECT  153150.0 1449450.0 154050.0 1448550.0 ;
      RECT  148200.0 1442250.0 157800.0 1441350.0 ;
      RECT  148200.0 1456050.0 157800.0 1455150.0 ;
      RECT  120450.0 1448400.0 121650.0 1449600.0 ;
      RECT  122400.0 1450800.0 123600.0 1452000.0 ;
      RECT  139200.0 1449900.0 138000.0 1451100.0 ;
      RECT  130800.0 1467450.0 132000.0 1469400.0 ;
      RECT  130800.0 1455600.0 132000.0 1457550.0 ;
      RECT  126000.0 1456950.0 127200.0 1455150.0 ;
      RECT  126000.0 1466250.0 127200.0 1469850.0 ;
      RECT  128700.0 1456950.0 129600.0 1466250.0 ;
      RECT  126000.0 1466250.0 127200.0 1467450.0 ;
      RECT  128400.0 1466250.0 129600.0 1467450.0 ;
      RECT  128400.0 1466250.0 129600.0 1467450.0 ;
      RECT  126000.0 1466250.0 127200.0 1467450.0 ;
      RECT  126000.0 1456950.0 127200.0 1458150.0 ;
      RECT  128400.0 1456950.0 129600.0 1458150.0 ;
      RECT  128400.0 1456950.0 129600.0 1458150.0 ;
      RECT  126000.0 1456950.0 127200.0 1458150.0 ;
      RECT  130800.0 1466850.0 132000.0 1468050.0 ;
      RECT  130800.0 1456950.0 132000.0 1458150.0 ;
      RECT  126600.0 1461600.0 127800.0 1462800.0 ;
      RECT  126600.0 1461600.0 127800.0 1462800.0 ;
      RECT  129150.0 1461750.0 130050.0 1462650.0 ;
      RECT  124200.0 1468950.0 133800.0 1469850.0 ;
      RECT  124200.0 1455150.0 133800.0 1456050.0 ;
      RECT  135600.0 1457550.0 136800.0 1455150.0 ;
      RECT  135600.0 1466250.0 136800.0 1469850.0 ;
      RECT  140400.0 1466250.0 141600.0 1469850.0 ;
      RECT  142800.0 1467450.0 144000.0 1469400.0 ;
      RECT  142800.0 1455600.0 144000.0 1457550.0 ;
      RECT  135600.0 1466250.0 136800.0 1467450.0 ;
      RECT  138000.0 1466250.0 139200.0 1467450.0 ;
      RECT  138000.0 1466250.0 139200.0 1467450.0 ;
      RECT  135600.0 1466250.0 136800.0 1467450.0 ;
      RECT  138000.0 1466250.0 139200.0 1467450.0 ;
      RECT  140400.0 1466250.0 141600.0 1467450.0 ;
      RECT  140400.0 1466250.0 141600.0 1467450.0 ;
      RECT  138000.0 1466250.0 139200.0 1467450.0 ;
      RECT  135600.0 1457550.0 136800.0 1458750.0 ;
      RECT  138000.0 1457550.0 139200.0 1458750.0 ;
      RECT  138000.0 1457550.0 139200.0 1458750.0 ;
      RECT  135600.0 1457550.0 136800.0 1458750.0 ;
      RECT  138000.0 1457550.0 139200.0 1458750.0 ;
      RECT  140400.0 1457550.0 141600.0 1458750.0 ;
      RECT  140400.0 1457550.0 141600.0 1458750.0 ;
      RECT  138000.0 1457550.0 139200.0 1458750.0 ;
      RECT  142800.0 1466850.0 144000.0 1468050.0 ;
      RECT  142800.0 1456950.0 144000.0 1458150.0 ;
      RECT  140400.0 1460100.0 139200.0 1461300.0 ;
      RECT  137400.0 1462800.0 136200.0 1464000.0 ;
      RECT  138000.0 1466250.0 139200.0 1467450.0 ;
      RECT  140400.0 1457550.0 141600.0 1458750.0 ;
      RECT  141600.0 1462800.0 140400.0 1464000.0 ;
      RECT  136200.0 1462800.0 137400.0 1464000.0 ;
      RECT  139200.0 1460100.0 140400.0 1461300.0 ;
      RECT  140400.0 1462800.0 141600.0 1464000.0 ;
      RECT  133800.0 1468950.0 148200.0 1469850.0 ;
      RECT  133800.0 1455150.0 148200.0 1456050.0 ;
      RECT  154800.0 1467450.0 156000.0 1469400.0 ;
      RECT  154800.0 1455600.0 156000.0 1457550.0 ;
      RECT  150000.0 1456950.0 151200.0 1455150.0 ;
      RECT  150000.0 1466250.0 151200.0 1469850.0 ;
      RECT  152700.0 1456950.0 153600.0 1466250.0 ;
      RECT  150000.0 1466250.0 151200.0 1467450.0 ;
      RECT  152400.0 1466250.0 153600.0 1467450.0 ;
      RECT  152400.0 1466250.0 153600.0 1467450.0 ;
      RECT  150000.0 1466250.0 151200.0 1467450.0 ;
      RECT  150000.0 1456950.0 151200.0 1458150.0 ;
      RECT  152400.0 1456950.0 153600.0 1458150.0 ;
      RECT  152400.0 1456950.0 153600.0 1458150.0 ;
      RECT  150000.0 1456950.0 151200.0 1458150.0 ;
      RECT  154800.0 1466850.0 156000.0 1468050.0 ;
      RECT  154800.0 1456950.0 156000.0 1458150.0 ;
      RECT  150600.0 1461600.0 151800.0 1462800.0 ;
      RECT  150600.0 1461600.0 151800.0 1462800.0 ;
      RECT  153150.0 1461750.0 154050.0 1462650.0 ;
      RECT  148200.0 1468950.0 157800.0 1469850.0 ;
      RECT  148200.0 1455150.0 157800.0 1456050.0 ;
      RECT  120450.0 1461600.0 121650.0 1462800.0 ;
      RECT  122400.0 1459200.0 123600.0 1460400.0 ;
      RECT  139200.0 1460100.0 138000.0 1461300.0 ;
      RECT  130800.0 1471350.0 132000.0 1469400.0 ;
      RECT  130800.0 1483200.0 132000.0 1481250.0 ;
      RECT  126000.0 1481850.0 127200.0 1483650.0 ;
      RECT  126000.0 1472550.0 127200.0 1468950.0 ;
      RECT  128700.0 1481850.0 129600.0 1472550.0 ;
      RECT  126000.0 1472550.0 127200.0 1471350.0 ;
      RECT  128400.0 1472550.0 129600.0 1471350.0 ;
      RECT  128400.0 1472550.0 129600.0 1471350.0 ;
      RECT  126000.0 1472550.0 127200.0 1471350.0 ;
      RECT  126000.0 1481850.0 127200.0 1480650.0 ;
      RECT  128400.0 1481850.0 129600.0 1480650.0 ;
      RECT  128400.0 1481850.0 129600.0 1480650.0 ;
      RECT  126000.0 1481850.0 127200.0 1480650.0 ;
      RECT  130800.0 1471950.0 132000.0 1470750.0 ;
      RECT  130800.0 1481850.0 132000.0 1480650.0 ;
      RECT  126600.0 1477200.0 127800.0 1476000.0 ;
      RECT  126600.0 1477200.0 127800.0 1476000.0 ;
      RECT  129150.0 1477050.0 130050.0 1476150.0 ;
      RECT  124200.0 1469850.0 133800.0 1468950.0 ;
      RECT  124200.0 1483650.0 133800.0 1482750.0 ;
      RECT  135600.0 1481250.0 136800.0 1483650.0 ;
      RECT  135600.0 1472550.0 136800.0 1468950.0 ;
      RECT  140400.0 1472550.0 141600.0 1468950.0 ;
      RECT  142800.0 1471350.0 144000.0 1469400.0 ;
      RECT  142800.0 1483200.0 144000.0 1481250.0 ;
      RECT  135600.0 1472550.0 136800.0 1471350.0 ;
      RECT  138000.0 1472550.0 139200.0 1471350.0 ;
      RECT  138000.0 1472550.0 139200.0 1471350.0 ;
      RECT  135600.0 1472550.0 136800.0 1471350.0 ;
      RECT  138000.0 1472550.0 139200.0 1471350.0 ;
      RECT  140400.0 1472550.0 141600.0 1471350.0 ;
      RECT  140400.0 1472550.0 141600.0 1471350.0 ;
      RECT  138000.0 1472550.0 139200.0 1471350.0 ;
      RECT  135600.0 1481250.0 136800.0 1480050.0 ;
      RECT  138000.0 1481250.0 139200.0 1480050.0 ;
      RECT  138000.0 1481250.0 139200.0 1480050.0 ;
      RECT  135600.0 1481250.0 136800.0 1480050.0 ;
      RECT  138000.0 1481250.0 139200.0 1480050.0 ;
      RECT  140400.0 1481250.0 141600.0 1480050.0 ;
      RECT  140400.0 1481250.0 141600.0 1480050.0 ;
      RECT  138000.0 1481250.0 139200.0 1480050.0 ;
      RECT  142800.0 1471950.0 144000.0 1470750.0 ;
      RECT  142800.0 1481850.0 144000.0 1480650.0 ;
      RECT  140400.0 1478700.0 139200.0 1477500.0 ;
      RECT  137400.0 1476000.0 136200.0 1474800.0 ;
      RECT  138000.0 1472550.0 139200.0 1471350.0 ;
      RECT  140400.0 1481250.0 141600.0 1480050.0 ;
      RECT  141600.0 1476000.0 140400.0 1474800.0 ;
      RECT  136200.0 1476000.0 137400.0 1474800.0 ;
      RECT  139200.0 1478700.0 140400.0 1477500.0 ;
      RECT  140400.0 1476000.0 141600.0 1474800.0 ;
      RECT  133800.0 1469850.0 148200.0 1468950.0 ;
      RECT  133800.0 1483650.0 148200.0 1482750.0 ;
      RECT  154800.0 1471350.0 156000.0 1469400.0 ;
      RECT  154800.0 1483200.0 156000.0 1481250.0 ;
      RECT  150000.0 1481850.0 151200.0 1483650.0 ;
      RECT  150000.0 1472550.0 151200.0 1468950.0 ;
      RECT  152700.0 1481850.0 153600.0 1472550.0 ;
      RECT  150000.0 1472550.0 151200.0 1471350.0 ;
      RECT  152400.0 1472550.0 153600.0 1471350.0 ;
      RECT  152400.0 1472550.0 153600.0 1471350.0 ;
      RECT  150000.0 1472550.0 151200.0 1471350.0 ;
      RECT  150000.0 1481850.0 151200.0 1480650.0 ;
      RECT  152400.0 1481850.0 153600.0 1480650.0 ;
      RECT  152400.0 1481850.0 153600.0 1480650.0 ;
      RECT  150000.0 1481850.0 151200.0 1480650.0 ;
      RECT  154800.0 1471950.0 156000.0 1470750.0 ;
      RECT  154800.0 1481850.0 156000.0 1480650.0 ;
      RECT  150600.0 1477200.0 151800.0 1476000.0 ;
      RECT  150600.0 1477200.0 151800.0 1476000.0 ;
      RECT  153150.0 1477050.0 154050.0 1476150.0 ;
      RECT  148200.0 1469850.0 157800.0 1468950.0 ;
      RECT  148200.0 1483650.0 157800.0 1482750.0 ;
      RECT  120450.0 1476000.0 121650.0 1477200.0 ;
      RECT  122400.0 1478400.0 123600.0 1479600.0 ;
      RECT  139200.0 1477500.0 138000.0 1478700.0 ;
      RECT  130800.0 1495050.0 132000.0 1497000.0 ;
      RECT  130800.0 1483200.0 132000.0 1485150.0 ;
      RECT  126000.0 1484550.0 127200.0 1482750.0 ;
      RECT  126000.0 1493850.0 127200.0 1497450.0 ;
      RECT  128700.0 1484550.0 129600.0 1493850.0 ;
      RECT  126000.0 1493850.0 127200.0 1495050.0 ;
      RECT  128400.0 1493850.0 129600.0 1495050.0 ;
      RECT  128400.0 1493850.0 129600.0 1495050.0 ;
      RECT  126000.0 1493850.0 127200.0 1495050.0 ;
      RECT  126000.0 1484550.0 127200.0 1485750.0 ;
      RECT  128400.0 1484550.0 129600.0 1485750.0 ;
      RECT  128400.0 1484550.0 129600.0 1485750.0 ;
      RECT  126000.0 1484550.0 127200.0 1485750.0 ;
      RECT  130800.0 1494450.0 132000.0 1495650.0 ;
      RECT  130800.0 1484550.0 132000.0 1485750.0 ;
      RECT  126600.0 1489200.0 127800.0 1490400.0 ;
      RECT  126600.0 1489200.0 127800.0 1490400.0 ;
      RECT  129150.0 1489350.0 130050.0 1490250.0 ;
      RECT  124200.0 1496550.0 133800.0 1497450.0 ;
      RECT  124200.0 1482750.0 133800.0 1483650.0 ;
      RECT  135600.0 1485150.0 136800.0 1482750.0 ;
      RECT  135600.0 1493850.0 136800.0 1497450.0 ;
      RECT  140400.0 1493850.0 141600.0 1497450.0 ;
      RECT  142800.0 1495050.0 144000.0 1497000.0 ;
      RECT  142800.0 1483200.0 144000.0 1485150.0 ;
      RECT  135600.0 1493850.0 136800.0 1495050.0 ;
      RECT  138000.0 1493850.0 139200.0 1495050.0 ;
      RECT  138000.0 1493850.0 139200.0 1495050.0 ;
      RECT  135600.0 1493850.0 136800.0 1495050.0 ;
      RECT  138000.0 1493850.0 139200.0 1495050.0 ;
      RECT  140400.0 1493850.0 141600.0 1495050.0 ;
      RECT  140400.0 1493850.0 141600.0 1495050.0 ;
      RECT  138000.0 1493850.0 139200.0 1495050.0 ;
      RECT  135600.0 1485150.0 136800.0 1486350.0 ;
      RECT  138000.0 1485150.0 139200.0 1486350.0 ;
      RECT  138000.0 1485150.0 139200.0 1486350.0 ;
      RECT  135600.0 1485150.0 136800.0 1486350.0 ;
      RECT  138000.0 1485150.0 139200.0 1486350.0 ;
      RECT  140400.0 1485150.0 141600.0 1486350.0 ;
      RECT  140400.0 1485150.0 141600.0 1486350.0 ;
      RECT  138000.0 1485150.0 139200.0 1486350.0 ;
      RECT  142800.0 1494450.0 144000.0 1495650.0 ;
      RECT  142800.0 1484550.0 144000.0 1485750.0 ;
      RECT  140400.0 1487700.0 139200.0 1488900.0 ;
      RECT  137400.0 1490400.0 136200.0 1491600.0 ;
      RECT  138000.0 1493850.0 139200.0 1495050.0 ;
      RECT  140400.0 1485150.0 141600.0 1486350.0 ;
      RECT  141600.0 1490400.0 140400.0 1491600.0 ;
      RECT  136200.0 1490400.0 137400.0 1491600.0 ;
      RECT  139200.0 1487700.0 140400.0 1488900.0 ;
      RECT  140400.0 1490400.0 141600.0 1491600.0 ;
      RECT  133800.0 1496550.0 148200.0 1497450.0 ;
      RECT  133800.0 1482750.0 148200.0 1483650.0 ;
      RECT  154800.0 1495050.0 156000.0 1497000.0 ;
      RECT  154800.0 1483200.0 156000.0 1485150.0 ;
      RECT  150000.0 1484550.0 151200.0 1482750.0 ;
      RECT  150000.0 1493850.0 151200.0 1497450.0 ;
      RECT  152700.0 1484550.0 153600.0 1493850.0 ;
      RECT  150000.0 1493850.0 151200.0 1495050.0 ;
      RECT  152400.0 1493850.0 153600.0 1495050.0 ;
      RECT  152400.0 1493850.0 153600.0 1495050.0 ;
      RECT  150000.0 1493850.0 151200.0 1495050.0 ;
      RECT  150000.0 1484550.0 151200.0 1485750.0 ;
      RECT  152400.0 1484550.0 153600.0 1485750.0 ;
      RECT  152400.0 1484550.0 153600.0 1485750.0 ;
      RECT  150000.0 1484550.0 151200.0 1485750.0 ;
      RECT  154800.0 1494450.0 156000.0 1495650.0 ;
      RECT  154800.0 1484550.0 156000.0 1485750.0 ;
      RECT  150600.0 1489200.0 151800.0 1490400.0 ;
      RECT  150600.0 1489200.0 151800.0 1490400.0 ;
      RECT  153150.0 1489350.0 154050.0 1490250.0 ;
      RECT  148200.0 1496550.0 157800.0 1497450.0 ;
      RECT  148200.0 1482750.0 157800.0 1483650.0 ;
      RECT  120450.0 1489200.0 121650.0 1490400.0 ;
      RECT  122400.0 1486800.0 123600.0 1488000.0 ;
      RECT  139200.0 1487700.0 138000.0 1488900.0 ;
      RECT  130800.0 1498950.0 132000.0 1497000.0 ;
      RECT  130800.0 1510800.0 132000.0 1508850.0 ;
      RECT  126000.0 1509450.0 127200.0 1511250.0 ;
      RECT  126000.0 1500150.0 127200.0 1496550.0 ;
      RECT  128700.0 1509450.0 129600.0 1500150.0 ;
      RECT  126000.0 1500150.0 127200.0 1498950.0 ;
      RECT  128400.0 1500150.0 129600.0 1498950.0 ;
      RECT  128400.0 1500150.0 129600.0 1498950.0 ;
      RECT  126000.0 1500150.0 127200.0 1498950.0 ;
      RECT  126000.0 1509450.0 127200.0 1508250.0 ;
      RECT  128400.0 1509450.0 129600.0 1508250.0 ;
      RECT  128400.0 1509450.0 129600.0 1508250.0 ;
      RECT  126000.0 1509450.0 127200.0 1508250.0 ;
      RECT  130800.0 1499550.0 132000.0 1498350.0 ;
      RECT  130800.0 1509450.0 132000.0 1508250.0 ;
      RECT  126600.0 1504800.0 127800.0 1503600.0 ;
      RECT  126600.0 1504800.0 127800.0 1503600.0 ;
      RECT  129150.0 1504650.0 130050.0 1503750.0 ;
      RECT  124200.0 1497450.0 133800.0 1496550.0 ;
      RECT  124200.0 1511250.0 133800.0 1510350.0 ;
      RECT  135600.0 1508850.0 136800.0 1511250.0 ;
      RECT  135600.0 1500150.0 136800.0 1496550.0 ;
      RECT  140400.0 1500150.0 141600.0 1496550.0 ;
      RECT  142800.0 1498950.0 144000.0 1497000.0 ;
      RECT  142800.0 1510800.0 144000.0 1508850.0 ;
      RECT  135600.0 1500150.0 136800.0 1498950.0 ;
      RECT  138000.0 1500150.0 139200.0 1498950.0 ;
      RECT  138000.0 1500150.0 139200.0 1498950.0 ;
      RECT  135600.0 1500150.0 136800.0 1498950.0 ;
      RECT  138000.0 1500150.0 139200.0 1498950.0 ;
      RECT  140400.0 1500150.0 141600.0 1498950.0 ;
      RECT  140400.0 1500150.0 141600.0 1498950.0 ;
      RECT  138000.0 1500150.0 139200.0 1498950.0 ;
      RECT  135600.0 1508850.0 136800.0 1507650.0 ;
      RECT  138000.0 1508850.0 139200.0 1507650.0 ;
      RECT  138000.0 1508850.0 139200.0 1507650.0 ;
      RECT  135600.0 1508850.0 136800.0 1507650.0 ;
      RECT  138000.0 1508850.0 139200.0 1507650.0 ;
      RECT  140400.0 1508850.0 141600.0 1507650.0 ;
      RECT  140400.0 1508850.0 141600.0 1507650.0 ;
      RECT  138000.0 1508850.0 139200.0 1507650.0 ;
      RECT  142800.0 1499550.0 144000.0 1498350.0 ;
      RECT  142800.0 1509450.0 144000.0 1508250.0 ;
      RECT  140400.0 1506300.0 139200.0 1505100.0 ;
      RECT  137400.0 1503600.0 136200.0 1502400.0 ;
      RECT  138000.0 1500150.0 139200.0 1498950.0 ;
      RECT  140400.0 1508850.0 141600.0 1507650.0 ;
      RECT  141600.0 1503600.0 140400.0 1502400.0 ;
      RECT  136200.0 1503600.0 137400.0 1502400.0 ;
      RECT  139200.0 1506300.0 140400.0 1505100.0 ;
      RECT  140400.0 1503600.0 141600.0 1502400.0 ;
      RECT  133800.0 1497450.0 148200.0 1496550.0 ;
      RECT  133800.0 1511250.0 148200.0 1510350.0 ;
      RECT  154800.0 1498950.0 156000.0 1497000.0 ;
      RECT  154800.0 1510800.0 156000.0 1508850.0 ;
      RECT  150000.0 1509450.0 151200.0 1511250.0 ;
      RECT  150000.0 1500150.0 151200.0 1496550.0 ;
      RECT  152700.0 1509450.0 153600.0 1500150.0 ;
      RECT  150000.0 1500150.0 151200.0 1498950.0 ;
      RECT  152400.0 1500150.0 153600.0 1498950.0 ;
      RECT  152400.0 1500150.0 153600.0 1498950.0 ;
      RECT  150000.0 1500150.0 151200.0 1498950.0 ;
      RECT  150000.0 1509450.0 151200.0 1508250.0 ;
      RECT  152400.0 1509450.0 153600.0 1508250.0 ;
      RECT  152400.0 1509450.0 153600.0 1508250.0 ;
      RECT  150000.0 1509450.0 151200.0 1508250.0 ;
      RECT  154800.0 1499550.0 156000.0 1498350.0 ;
      RECT  154800.0 1509450.0 156000.0 1508250.0 ;
      RECT  150600.0 1504800.0 151800.0 1503600.0 ;
      RECT  150600.0 1504800.0 151800.0 1503600.0 ;
      RECT  153150.0 1504650.0 154050.0 1503750.0 ;
      RECT  148200.0 1497450.0 157800.0 1496550.0 ;
      RECT  148200.0 1511250.0 157800.0 1510350.0 ;
      RECT  120450.0 1503600.0 121650.0 1504800.0 ;
      RECT  122400.0 1506000.0 123600.0 1507200.0 ;
      RECT  139200.0 1505100.0 138000.0 1506300.0 ;
      RECT  130800.0 1522650.0 132000.0 1524600.0 ;
      RECT  130800.0 1510800.0 132000.0 1512750.0 ;
      RECT  126000.0 1512150.0 127200.0 1510350.0 ;
      RECT  126000.0 1521450.0 127200.0 1525050.0 ;
      RECT  128700.0 1512150.0 129600.0 1521450.0 ;
      RECT  126000.0 1521450.0 127200.0 1522650.0 ;
      RECT  128400.0 1521450.0 129600.0 1522650.0 ;
      RECT  128400.0 1521450.0 129600.0 1522650.0 ;
      RECT  126000.0 1521450.0 127200.0 1522650.0 ;
      RECT  126000.0 1512150.0 127200.0 1513350.0 ;
      RECT  128400.0 1512150.0 129600.0 1513350.0 ;
      RECT  128400.0 1512150.0 129600.0 1513350.0 ;
      RECT  126000.0 1512150.0 127200.0 1513350.0 ;
      RECT  130800.0 1522050.0 132000.0 1523250.0 ;
      RECT  130800.0 1512150.0 132000.0 1513350.0 ;
      RECT  126600.0 1516800.0 127800.0 1518000.0 ;
      RECT  126600.0 1516800.0 127800.0 1518000.0 ;
      RECT  129150.0 1516950.0 130050.0 1517850.0 ;
      RECT  124200.0 1524150.0 133800.0 1525050.0 ;
      RECT  124200.0 1510350.0 133800.0 1511250.0 ;
      RECT  135600.0 1512750.0 136800.0 1510350.0 ;
      RECT  135600.0 1521450.0 136800.0 1525050.0 ;
      RECT  140400.0 1521450.0 141600.0 1525050.0 ;
      RECT  142800.0 1522650.0 144000.0 1524600.0 ;
      RECT  142800.0 1510800.0 144000.0 1512750.0 ;
      RECT  135600.0 1521450.0 136800.0 1522650.0 ;
      RECT  138000.0 1521450.0 139200.0 1522650.0 ;
      RECT  138000.0 1521450.0 139200.0 1522650.0 ;
      RECT  135600.0 1521450.0 136800.0 1522650.0 ;
      RECT  138000.0 1521450.0 139200.0 1522650.0 ;
      RECT  140400.0 1521450.0 141600.0 1522650.0 ;
      RECT  140400.0 1521450.0 141600.0 1522650.0 ;
      RECT  138000.0 1521450.0 139200.0 1522650.0 ;
      RECT  135600.0 1512750.0 136800.0 1513950.0 ;
      RECT  138000.0 1512750.0 139200.0 1513950.0 ;
      RECT  138000.0 1512750.0 139200.0 1513950.0 ;
      RECT  135600.0 1512750.0 136800.0 1513950.0 ;
      RECT  138000.0 1512750.0 139200.0 1513950.0 ;
      RECT  140400.0 1512750.0 141600.0 1513950.0 ;
      RECT  140400.0 1512750.0 141600.0 1513950.0 ;
      RECT  138000.0 1512750.0 139200.0 1513950.0 ;
      RECT  142800.0 1522050.0 144000.0 1523250.0 ;
      RECT  142800.0 1512150.0 144000.0 1513350.0 ;
      RECT  140400.0 1515300.0 139200.0 1516500.0 ;
      RECT  137400.0 1518000.0 136200.0 1519200.0 ;
      RECT  138000.0 1521450.0 139200.0 1522650.0 ;
      RECT  140400.0 1512750.0 141600.0 1513950.0 ;
      RECT  141600.0 1518000.0 140400.0 1519200.0 ;
      RECT  136200.0 1518000.0 137400.0 1519200.0 ;
      RECT  139200.0 1515300.0 140400.0 1516500.0 ;
      RECT  140400.0 1518000.0 141600.0 1519200.0 ;
      RECT  133800.0 1524150.0 148200.0 1525050.0 ;
      RECT  133800.0 1510350.0 148200.0 1511250.0 ;
      RECT  154800.0 1522650.0 156000.0 1524600.0 ;
      RECT  154800.0 1510800.0 156000.0 1512750.0 ;
      RECT  150000.0 1512150.0 151200.0 1510350.0 ;
      RECT  150000.0 1521450.0 151200.0 1525050.0 ;
      RECT  152700.0 1512150.0 153600.0 1521450.0 ;
      RECT  150000.0 1521450.0 151200.0 1522650.0 ;
      RECT  152400.0 1521450.0 153600.0 1522650.0 ;
      RECT  152400.0 1521450.0 153600.0 1522650.0 ;
      RECT  150000.0 1521450.0 151200.0 1522650.0 ;
      RECT  150000.0 1512150.0 151200.0 1513350.0 ;
      RECT  152400.0 1512150.0 153600.0 1513350.0 ;
      RECT  152400.0 1512150.0 153600.0 1513350.0 ;
      RECT  150000.0 1512150.0 151200.0 1513350.0 ;
      RECT  154800.0 1522050.0 156000.0 1523250.0 ;
      RECT  154800.0 1512150.0 156000.0 1513350.0 ;
      RECT  150600.0 1516800.0 151800.0 1518000.0 ;
      RECT  150600.0 1516800.0 151800.0 1518000.0 ;
      RECT  153150.0 1516950.0 154050.0 1517850.0 ;
      RECT  148200.0 1524150.0 157800.0 1525050.0 ;
      RECT  148200.0 1510350.0 157800.0 1511250.0 ;
      RECT  120450.0 1516800.0 121650.0 1518000.0 ;
      RECT  122400.0 1514400.0 123600.0 1515600.0 ;
      RECT  139200.0 1515300.0 138000.0 1516500.0 ;
      RECT  130800.0 1526550.0 132000.0 1524600.0 ;
      RECT  130800.0 1538400.0 132000.0 1536450.0 ;
      RECT  126000.0 1537050.0 127200.0 1538850.0 ;
      RECT  126000.0 1527750.0 127200.0 1524150.0 ;
      RECT  128700.0 1537050.0 129600.0 1527750.0 ;
      RECT  126000.0 1527750.0 127200.0 1526550.0 ;
      RECT  128400.0 1527750.0 129600.0 1526550.0 ;
      RECT  128400.0 1527750.0 129600.0 1526550.0 ;
      RECT  126000.0 1527750.0 127200.0 1526550.0 ;
      RECT  126000.0 1537050.0 127200.0 1535850.0 ;
      RECT  128400.0 1537050.0 129600.0 1535850.0 ;
      RECT  128400.0 1537050.0 129600.0 1535850.0 ;
      RECT  126000.0 1537050.0 127200.0 1535850.0 ;
      RECT  130800.0 1527150.0 132000.0 1525950.0 ;
      RECT  130800.0 1537050.0 132000.0 1535850.0 ;
      RECT  126600.0 1532400.0 127800.0 1531200.0 ;
      RECT  126600.0 1532400.0 127800.0 1531200.0 ;
      RECT  129150.0 1532250.0 130050.0 1531350.0 ;
      RECT  124200.0 1525050.0 133800.0 1524150.0 ;
      RECT  124200.0 1538850.0 133800.0 1537950.0 ;
      RECT  135600.0 1536450.0 136800.0 1538850.0 ;
      RECT  135600.0 1527750.0 136800.0 1524150.0 ;
      RECT  140400.0 1527750.0 141600.0 1524150.0 ;
      RECT  142800.0 1526550.0 144000.0 1524600.0 ;
      RECT  142800.0 1538400.0 144000.0 1536450.0 ;
      RECT  135600.0 1527750.0 136800.0 1526550.0 ;
      RECT  138000.0 1527750.0 139200.0 1526550.0 ;
      RECT  138000.0 1527750.0 139200.0 1526550.0 ;
      RECT  135600.0 1527750.0 136800.0 1526550.0 ;
      RECT  138000.0 1527750.0 139200.0 1526550.0 ;
      RECT  140400.0 1527750.0 141600.0 1526550.0 ;
      RECT  140400.0 1527750.0 141600.0 1526550.0 ;
      RECT  138000.0 1527750.0 139200.0 1526550.0 ;
      RECT  135600.0 1536450.0 136800.0 1535250.0 ;
      RECT  138000.0 1536450.0 139200.0 1535250.0 ;
      RECT  138000.0 1536450.0 139200.0 1535250.0 ;
      RECT  135600.0 1536450.0 136800.0 1535250.0 ;
      RECT  138000.0 1536450.0 139200.0 1535250.0 ;
      RECT  140400.0 1536450.0 141600.0 1535250.0 ;
      RECT  140400.0 1536450.0 141600.0 1535250.0 ;
      RECT  138000.0 1536450.0 139200.0 1535250.0 ;
      RECT  142800.0 1527150.0 144000.0 1525950.0 ;
      RECT  142800.0 1537050.0 144000.0 1535850.0 ;
      RECT  140400.0 1533900.0 139200.0 1532700.0 ;
      RECT  137400.0 1531200.0 136200.0 1530000.0 ;
      RECT  138000.0 1527750.0 139200.0 1526550.0 ;
      RECT  140400.0 1536450.0 141600.0 1535250.0 ;
      RECT  141600.0 1531200.0 140400.0 1530000.0 ;
      RECT  136200.0 1531200.0 137400.0 1530000.0 ;
      RECT  139200.0 1533900.0 140400.0 1532700.0 ;
      RECT  140400.0 1531200.0 141600.0 1530000.0 ;
      RECT  133800.0 1525050.0 148200.0 1524150.0 ;
      RECT  133800.0 1538850.0 148200.0 1537950.0 ;
      RECT  154800.0 1526550.0 156000.0 1524600.0 ;
      RECT  154800.0 1538400.0 156000.0 1536450.0 ;
      RECT  150000.0 1537050.0 151200.0 1538850.0 ;
      RECT  150000.0 1527750.0 151200.0 1524150.0 ;
      RECT  152700.0 1537050.0 153600.0 1527750.0 ;
      RECT  150000.0 1527750.0 151200.0 1526550.0 ;
      RECT  152400.0 1527750.0 153600.0 1526550.0 ;
      RECT  152400.0 1527750.0 153600.0 1526550.0 ;
      RECT  150000.0 1527750.0 151200.0 1526550.0 ;
      RECT  150000.0 1537050.0 151200.0 1535850.0 ;
      RECT  152400.0 1537050.0 153600.0 1535850.0 ;
      RECT  152400.0 1537050.0 153600.0 1535850.0 ;
      RECT  150000.0 1537050.0 151200.0 1535850.0 ;
      RECT  154800.0 1527150.0 156000.0 1525950.0 ;
      RECT  154800.0 1537050.0 156000.0 1535850.0 ;
      RECT  150600.0 1532400.0 151800.0 1531200.0 ;
      RECT  150600.0 1532400.0 151800.0 1531200.0 ;
      RECT  153150.0 1532250.0 154050.0 1531350.0 ;
      RECT  148200.0 1525050.0 157800.0 1524150.0 ;
      RECT  148200.0 1538850.0 157800.0 1537950.0 ;
      RECT  120450.0 1531200.0 121650.0 1532400.0 ;
      RECT  122400.0 1533600.0 123600.0 1534800.0 ;
      RECT  139200.0 1532700.0 138000.0 1533900.0 ;
      RECT  130800.0 1550250.0 132000.0 1552200.0 ;
      RECT  130800.0 1538400.0 132000.0 1540350.0 ;
      RECT  126000.0 1539750.0 127200.0 1537950.0 ;
      RECT  126000.0 1549050.0 127200.0 1552650.0 ;
      RECT  128700.0 1539750.0 129600.0 1549050.0 ;
      RECT  126000.0 1549050.0 127200.0 1550250.0 ;
      RECT  128400.0 1549050.0 129600.0 1550250.0 ;
      RECT  128400.0 1549050.0 129600.0 1550250.0 ;
      RECT  126000.0 1549050.0 127200.0 1550250.0 ;
      RECT  126000.0 1539750.0 127200.0 1540950.0 ;
      RECT  128400.0 1539750.0 129600.0 1540950.0 ;
      RECT  128400.0 1539750.0 129600.0 1540950.0 ;
      RECT  126000.0 1539750.0 127200.0 1540950.0 ;
      RECT  130800.0 1549650.0 132000.0 1550850.0 ;
      RECT  130800.0 1539750.0 132000.0 1540950.0 ;
      RECT  126600.0 1544400.0 127800.0 1545600.0 ;
      RECT  126600.0 1544400.0 127800.0 1545600.0 ;
      RECT  129150.0 1544550.0 130050.0 1545450.0 ;
      RECT  124200.0 1551750.0 133800.0 1552650.0 ;
      RECT  124200.0 1537950.0 133800.0 1538850.0 ;
      RECT  135600.0 1540350.0 136800.0 1537950.0 ;
      RECT  135600.0 1549050.0 136800.0 1552650.0 ;
      RECT  140400.0 1549050.0 141600.0 1552650.0 ;
      RECT  142800.0 1550250.0 144000.0 1552200.0 ;
      RECT  142800.0 1538400.0 144000.0 1540350.0 ;
      RECT  135600.0 1549050.0 136800.0 1550250.0 ;
      RECT  138000.0 1549050.0 139200.0 1550250.0 ;
      RECT  138000.0 1549050.0 139200.0 1550250.0 ;
      RECT  135600.0 1549050.0 136800.0 1550250.0 ;
      RECT  138000.0 1549050.0 139200.0 1550250.0 ;
      RECT  140400.0 1549050.0 141600.0 1550250.0 ;
      RECT  140400.0 1549050.0 141600.0 1550250.0 ;
      RECT  138000.0 1549050.0 139200.0 1550250.0 ;
      RECT  135600.0 1540350.0 136800.0 1541550.0 ;
      RECT  138000.0 1540350.0 139200.0 1541550.0 ;
      RECT  138000.0 1540350.0 139200.0 1541550.0 ;
      RECT  135600.0 1540350.0 136800.0 1541550.0 ;
      RECT  138000.0 1540350.0 139200.0 1541550.0 ;
      RECT  140400.0 1540350.0 141600.0 1541550.0 ;
      RECT  140400.0 1540350.0 141600.0 1541550.0 ;
      RECT  138000.0 1540350.0 139200.0 1541550.0 ;
      RECT  142800.0 1549650.0 144000.0 1550850.0 ;
      RECT  142800.0 1539750.0 144000.0 1540950.0 ;
      RECT  140400.0 1542900.0 139200.0 1544100.0 ;
      RECT  137400.0 1545600.0 136200.0 1546800.0 ;
      RECT  138000.0 1549050.0 139200.0 1550250.0 ;
      RECT  140400.0 1540350.0 141600.0 1541550.0 ;
      RECT  141600.0 1545600.0 140400.0 1546800.0 ;
      RECT  136200.0 1545600.0 137400.0 1546800.0 ;
      RECT  139200.0 1542900.0 140400.0 1544100.0 ;
      RECT  140400.0 1545600.0 141600.0 1546800.0 ;
      RECT  133800.0 1551750.0 148200.0 1552650.0 ;
      RECT  133800.0 1537950.0 148200.0 1538850.0 ;
      RECT  154800.0 1550250.0 156000.0 1552200.0 ;
      RECT  154800.0 1538400.0 156000.0 1540350.0 ;
      RECT  150000.0 1539750.0 151200.0 1537950.0 ;
      RECT  150000.0 1549050.0 151200.0 1552650.0 ;
      RECT  152700.0 1539750.0 153600.0 1549050.0 ;
      RECT  150000.0 1549050.0 151200.0 1550250.0 ;
      RECT  152400.0 1549050.0 153600.0 1550250.0 ;
      RECT  152400.0 1549050.0 153600.0 1550250.0 ;
      RECT  150000.0 1549050.0 151200.0 1550250.0 ;
      RECT  150000.0 1539750.0 151200.0 1540950.0 ;
      RECT  152400.0 1539750.0 153600.0 1540950.0 ;
      RECT  152400.0 1539750.0 153600.0 1540950.0 ;
      RECT  150000.0 1539750.0 151200.0 1540950.0 ;
      RECT  154800.0 1549650.0 156000.0 1550850.0 ;
      RECT  154800.0 1539750.0 156000.0 1540950.0 ;
      RECT  150600.0 1544400.0 151800.0 1545600.0 ;
      RECT  150600.0 1544400.0 151800.0 1545600.0 ;
      RECT  153150.0 1544550.0 154050.0 1545450.0 ;
      RECT  148200.0 1551750.0 157800.0 1552650.0 ;
      RECT  148200.0 1537950.0 157800.0 1538850.0 ;
      RECT  120450.0 1544400.0 121650.0 1545600.0 ;
      RECT  122400.0 1542000.0 123600.0 1543200.0 ;
      RECT  139200.0 1542900.0 138000.0 1544100.0 ;
      RECT  130800.0 1554150.0 132000.0 1552200.0 ;
      RECT  130800.0 1566000.0 132000.0 1564050.0 ;
      RECT  126000.0 1564650.0 127200.0 1566450.0 ;
      RECT  126000.0 1555350.0 127200.0 1551750.0 ;
      RECT  128700.0 1564650.0 129600.0 1555350.0 ;
      RECT  126000.0 1555350.0 127200.0 1554150.0 ;
      RECT  128400.0 1555350.0 129600.0 1554150.0 ;
      RECT  128400.0 1555350.0 129600.0 1554150.0 ;
      RECT  126000.0 1555350.0 127200.0 1554150.0 ;
      RECT  126000.0 1564650.0 127200.0 1563450.0 ;
      RECT  128400.0 1564650.0 129600.0 1563450.0 ;
      RECT  128400.0 1564650.0 129600.0 1563450.0 ;
      RECT  126000.0 1564650.0 127200.0 1563450.0 ;
      RECT  130800.0 1554750.0 132000.0 1553550.0 ;
      RECT  130800.0 1564650.0 132000.0 1563450.0 ;
      RECT  126600.0 1560000.0 127800.0 1558800.0 ;
      RECT  126600.0 1560000.0 127800.0 1558800.0 ;
      RECT  129150.0 1559850.0 130050.0 1558950.0 ;
      RECT  124200.0 1552650.0 133800.0 1551750.0 ;
      RECT  124200.0 1566450.0 133800.0 1565550.0 ;
      RECT  135600.0 1564050.0 136800.0 1566450.0 ;
      RECT  135600.0 1555350.0 136800.0 1551750.0 ;
      RECT  140400.0 1555350.0 141600.0 1551750.0 ;
      RECT  142800.0 1554150.0 144000.0 1552200.0 ;
      RECT  142800.0 1566000.0 144000.0 1564050.0 ;
      RECT  135600.0 1555350.0 136800.0 1554150.0 ;
      RECT  138000.0 1555350.0 139200.0 1554150.0 ;
      RECT  138000.0 1555350.0 139200.0 1554150.0 ;
      RECT  135600.0 1555350.0 136800.0 1554150.0 ;
      RECT  138000.0 1555350.0 139200.0 1554150.0 ;
      RECT  140400.0 1555350.0 141600.0 1554150.0 ;
      RECT  140400.0 1555350.0 141600.0 1554150.0 ;
      RECT  138000.0 1555350.0 139200.0 1554150.0 ;
      RECT  135600.0 1564050.0 136800.0 1562850.0 ;
      RECT  138000.0 1564050.0 139200.0 1562850.0 ;
      RECT  138000.0 1564050.0 139200.0 1562850.0 ;
      RECT  135600.0 1564050.0 136800.0 1562850.0 ;
      RECT  138000.0 1564050.0 139200.0 1562850.0 ;
      RECT  140400.0 1564050.0 141600.0 1562850.0 ;
      RECT  140400.0 1564050.0 141600.0 1562850.0 ;
      RECT  138000.0 1564050.0 139200.0 1562850.0 ;
      RECT  142800.0 1554750.0 144000.0 1553550.0 ;
      RECT  142800.0 1564650.0 144000.0 1563450.0 ;
      RECT  140400.0 1561500.0 139200.0 1560300.0 ;
      RECT  137400.0 1558800.0 136200.0 1557600.0 ;
      RECT  138000.0 1555350.0 139200.0 1554150.0 ;
      RECT  140400.0 1564050.0 141600.0 1562850.0 ;
      RECT  141600.0 1558800.0 140400.0 1557600.0 ;
      RECT  136200.0 1558800.0 137400.0 1557600.0 ;
      RECT  139200.0 1561500.0 140400.0 1560300.0 ;
      RECT  140400.0 1558800.0 141600.0 1557600.0 ;
      RECT  133800.0 1552650.0 148200.0 1551750.0 ;
      RECT  133800.0 1566450.0 148200.0 1565550.0 ;
      RECT  154800.0 1554150.0 156000.0 1552200.0 ;
      RECT  154800.0 1566000.0 156000.0 1564050.0 ;
      RECT  150000.0 1564650.0 151200.0 1566450.0 ;
      RECT  150000.0 1555350.0 151200.0 1551750.0 ;
      RECT  152700.0 1564650.0 153600.0 1555350.0 ;
      RECT  150000.0 1555350.0 151200.0 1554150.0 ;
      RECT  152400.0 1555350.0 153600.0 1554150.0 ;
      RECT  152400.0 1555350.0 153600.0 1554150.0 ;
      RECT  150000.0 1555350.0 151200.0 1554150.0 ;
      RECT  150000.0 1564650.0 151200.0 1563450.0 ;
      RECT  152400.0 1564650.0 153600.0 1563450.0 ;
      RECT  152400.0 1564650.0 153600.0 1563450.0 ;
      RECT  150000.0 1564650.0 151200.0 1563450.0 ;
      RECT  154800.0 1554750.0 156000.0 1553550.0 ;
      RECT  154800.0 1564650.0 156000.0 1563450.0 ;
      RECT  150600.0 1560000.0 151800.0 1558800.0 ;
      RECT  150600.0 1560000.0 151800.0 1558800.0 ;
      RECT  153150.0 1559850.0 154050.0 1558950.0 ;
      RECT  148200.0 1552650.0 157800.0 1551750.0 ;
      RECT  148200.0 1566450.0 157800.0 1565550.0 ;
      RECT  120450.0 1558800.0 121650.0 1560000.0 ;
      RECT  122400.0 1561200.0 123600.0 1562400.0 ;
      RECT  139200.0 1560300.0 138000.0 1561500.0 ;
      RECT  130800.0 1577850.0 132000.0 1579800.0 ;
      RECT  130800.0 1566000.0 132000.0 1567950.0 ;
      RECT  126000.0 1567350.0 127200.0 1565550.0 ;
      RECT  126000.0 1576650.0 127200.0 1580250.0 ;
      RECT  128700.0 1567350.0 129600.0 1576650.0 ;
      RECT  126000.0 1576650.0 127200.0 1577850.0 ;
      RECT  128400.0 1576650.0 129600.0 1577850.0 ;
      RECT  128400.0 1576650.0 129600.0 1577850.0 ;
      RECT  126000.0 1576650.0 127200.0 1577850.0 ;
      RECT  126000.0 1567350.0 127200.0 1568550.0 ;
      RECT  128400.0 1567350.0 129600.0 1568550.0 ;
      RECT  128400.0 1567350.0 129600.0 1568550.0 ;
      RECT  126000.0 1567350.0 127200.0 1568550.0 ;
      RECT  130800.0 1577250.0 132000.0 1578450.0 ;
      RECT  130800.0 1567350.0 132000.0 1568550.0 ;
      RECT  126600.0 1572000.0 127800.0 1573200.0 ;
      RECT  126600.0 1572000.0 127800.0 1573200.0 ;
      RECT  129150.0 1572150.0 130050.0 1573050.0 ;
      RECT  124200.0 1579350.0 133800.0 1580250.0 ;
      RECT  124200.0 1565550.0 133800.0 1566450.0 ;
      RECT  135600.0 1567950.0 136800.0 1565550.0 ;
      RECT  135600.0 1576650.0 136800.0 1580250.0 ;
      RECT  140400.0 1576650.0 141600.0 1580250.0 ;
      RECT  142800.0 1577850.0 144000.0 1579800.0 ;
      RECT  142800.0 1566000.0 144000.0 1567950.0 ;
      RECT  135600.0 1576650.0 136800.0 1577850.0 ;
      RECT  138000.0 1576650.0 139200.0 1577850.0 ;
      RECT  138000.0 1576650.0 139200.0 1577850.0 ;
      RECT  135600.0 1576650.0 136800.0 1577850.0 ;
      RECT  138000.0 1576650.0 139200.0 1577850.0 ;
      RECT  140400.0 1576650.0 141600.0 1577850.0 ;
      RECT  140400.0 1576650.0 141600.0 1577850.0 ;
      RECT  138000.0 1576650.0 139200.0 1577850.0 ;
      RECT  135600.0 1567950.0 136800.0 1569150.0 ;
      RECT  138000.0 1567950.0 139200.0 1569150.0 ;
      RECT  138000.0 1567950.0 139200.0 1569150.0 ;
      RECT  135600.0 1567950.0 136800.0 1569150.0 ;
      RECT  138000.0 1567950.0 139200.0 1569150.0 ;
      RECT  140400.0 1567950.0 141600.0 1569150.0 ;
      RECT  140400.0 1567950.0 141600.0 1569150.0 ;
      RECT  138000.0 1567950.0 139200.0 1569150.0 ;
      RECT  142800.0 1577250.0 144000.0 1578450.0 ;
      RECT  142800.0 1567350.0 144000.0 1568550.0 ;
      RECT  140400.0 1570500.0 139200.0 1571700.0 ;
      RECT  137400.0 1573200.0 136200.0 1574400.0 ;
      RECT  138000.0 1576650.0 139200.0 1577850.0 ;
      RECT  140400.0 1567950.0 141600.0 1569150.0 ;
      RECT  141600.0 1573200.0 140400.0 1574400.0 ;
      RECT  136200.0 1573200.0 137400.0 1574400.0 ;
      RECT  139200.0 1570500.0 140400.0 1571700.0 ;
      RECT  140400.0 1573200.0 141600.0 1574400.0 ;
      RECT  133800.0 1579350.0 148200.0 1580250.0 ;
      RECT  133800.0 1565550.0 148200.0 1566450.0 ;
      RECT  154800.0 1577850.0 156000.0 1579800.0 ;
      RECT  154800.0 1566000.0 156000.0 1567950.0 ;
      RECT  150000.0 1567350.0 151200.0 1565550.0 ;
      RECT  150000.0 1576650.0 151200.0 1580250.0 ;
      RECT  152700.0 1567350.0 153600.0 1576650.0 ;
      RECT  150000.0 1576650.0 151200.0 1577850.0 ;
      RECT  152400.0 1576650.0 153600.0 1577850.0 ;
      RECT  152400.0 1576650.0 153600.0 1577850.0 ;
      RECT  150000.0 1576650.0 151200.0 1577850.0 ;
      RECT  150000.0 1567350.0 151200.0 1568550.0 ;
      RECT  152400.0 1567350.0 153600.0 1568550.0 ;
      RECT  152400.0 1567350.0 153600.0 1568550.0 ;
      RECT  150000.0 1567350.0 151200.0 1568550.0 ;
      RECT  154800.0 1577250.0 156000.0 1578450.0 ;
      RECT  154800.0 1567350.0 156000.0 1568550.0 ;
      RECT  150600.0 1572000.0 151800.0 1573200.0 ;
      RECT  150600.0 1572000.0 151800.0 1573200.0 ;
      RECT  153150.0 1572150.0 154050.0 1573050.0 ;
      RECT  148200.0 1579350.0 157800.0 1580250.0 ;
      RECT  148200.0 1565550.0 157800.0 1566450.0 ;
      RECT  120450.0 1572000.0 121650.0 1573200.0 ;
      RECT  122400.0 1569600.0 123600.0 1570800.0 ;
      RECT  139200.0 1570500.0 138000.0 1571700.0 ;
      RECT  130800.0 1581750.0 132000.0 1579800.0 ;
      RECT  130800.0 1593600.0 132000.0 1591650.0 ;
      RECT  126000.0 1592250.0 127200.0 1594050.0 ;
      RECT  126000.0 1582950.0 127200.0 1579350.0 ;
      RECT  128700.0 1592250.0 129600.0 1582950.0 ;
      RECT  126000.0 1582950.0 127200.0 1581750.0 ;
      RECT  128400.0 1582950.0 129600.0 1581750.0 ;
      RECT  128400.0 1582950.0 129600.0 1581750.0 ;
      RECT  126000.0 1582950.0 127200.0 1581750.0 ;
      RECT  126000.0 1592250.0 127200.0 1591050.0 ;
      RECT  128400.0 1592250.0 129600.0 1591050.0 ;
      RECT  128400.0 1592250.0 129600.0 1591050.0 ;
      RECT  126000.0 1592250.0 127200.0 1591050.0 ;
      RECT  130800.0 1582350.0 132000.0 1581150.0 ;
      RECT  130800.0 1592250.0 132000.0 1591050.0 ;
      RECT  126600.0 1587600.0 127800.0 1586400.0 ;
      RECT  126600.0 1587600.0 127800.0 1586400.0 ;
      RECT  129150.0 1587450.0 130050.0 1586550.0 ;
      RECT  124200.0 1580250.0 133800.0 1579350.0 ;
      RECT  124200.0 1594050.0 133800.0 1593150.0 ;
      RECT  135600.0 1591650.0 136800.0 1594050.0 ;
      RECT  135600.0 1582950.0 136800.0 1579350.0 ;
      RECT  140400.0 1582950.0 141600.0 1579350.0 ;
      RECT  142800.0 1581750.0 144000.0 1579800.0 ;
      RECT  142800.0 1593600.0 144000.0 1591650.0 ;
      RECT  135600.0 1582950.0 136800.0 1581750.0 ;
      RECT  138000.0 1582950.0 139200.0 1581750.0 ;
      RECT  138000.0 1582950.0 139200.0 1581750.0 ;
      RECT  135600.0 1582950.0 136800.0 1581750.0 ;
      RECT  138000.0 1582950.0 139200.0 1581750.0 ;
      RECT  140400.0 1582950.0 141600.0 1581750.0 ;
      RECT  140400.0 1582950.0 141600.0 1581750.0 ;
      RECT  138000.0 1582950.0 139200.0 1581750.0 ;
      RECT  135600.0 1591650.0 136800.0 1590450.0 ;
      RECT  138000.0 1591650.0 139200.0 1590450.0 ;
      RECT  138000.0 1591650.0 139200.0 1590450.0 ;
      RECT  135600.0 1591650.0 136800.0 1590450.0 ;
      RECT  138000.0 1591650.0 139200.0 1590450.0 ;
      RECT  140400.0 1591650.0 141600.0 1590450.0 ;
      RECT  140400.0 1591650.0 141600.0 1590450.0 ;
      RECT  138000.0 1591650.0 139200.0 1590450.0 ;
      RECT  142800.0 1582350.0 144000.0 1581150.0 ;
      RECT  142800.0 1592250.0 144000.0 1591050.0 ;
      RECT  140400.0 1589100.0 139200.0 1587900.0 ;
      RECT  137400.0 1586400.0 136200.0 1585200.0 ;
      RECT  138000.0 1582950.0 139200.0 1581750.0 ;
      RECT  140400.0 1591650.0 141600.0 1590450.0 ;
      RECT  141600.0 1586400.0 140400.0 1585200.0 ;
      RECT  136200.0 1586400.0 137400.0 1585200.0 ;
      RECT  139200.0 1589100.0 140400.0 1587900.0 ;
      RECT  140400.0 1586400.0 141600.0 1585200.0 ;
      RECT  133800.0 1580250.0 148200.0 1579350.0 ;
      RECT  133800.0 1594050.0 148200.0 1593150.0 ;
      RECT  154800.0 1581750.0 156000.0 1579800.0 ;
      RECT  154800.0 1593600.0 156000.0 1591650.0 ;
      RECT  150000.0 1592250.0 151200.0 1594050.0 ;
      RECT  150000.0 1582950.0 151200.0 1579350.0 ;
      RECT  152700.0 1592250.0 153600.0 1582950.0 ;
      RECT  150000.0 1582950.0 151200.0 1581750.0 ;
      RECT  152400.0 1582950.0 153600.0 1581750.0 ;
      RECT  152400.0 1582950.0 153600.0 1581750.0 ;
      RECT  150000.0 1582950.0 151200.0 1581750.0 ;
      RECT  150000.0 1592250.0 151200.0 1591050.0 ;
      RECT  152400.0 1592250.0 153600.0 1591050.0 ;
      RECT  152400.0 1592250.0 153600.0 1591050.0 ;
      RECT  150000.0 1592250.0 151200.0 1591050.0 ;
      RECT  154800.0 1582350.0 156000.0 1581150.0 ;
      RECT  154800.0 1592250.0 156000.0 1591050.0 ;
      RECT  150600.0 1587600.0 151800.0 1586400.0 ;
      RECT  150600.0 1587600.0 151800.0 1586400.0 ;
      RECT  153150.0 1587450.0 154050.0 1586550.0 ;
      RECT  148200.0 1580250.0 157800.0 1579350.0 ;
      RECT  148200.0 1594050.0 157800.0 1593150.0 ;
      RECT  120450.0 1586400.0 121650.0 1587600.0 ;
      RECT  122400.0 1588800.0 123600.0 1590000.0 ;
      RECT  139200.0 1587900.0 138000.0 1589100.0 ;
      RECT  130800.0 1605450.0 132000.0 1607400.0 ;
      RECT  130800.0 1593600.0 132000.0 1595550.0 ;
      RECT  126000.0 1594950.0 127200.0 1593150.0 ;
      RECT  126000.0 1604250.0 127200.0 1607850.0 ;
      RECT  128700.0 1594950.0 129600.0 1604250.0 ;
      RECT  126000.0 1604250.0 127200.0 1605450.0 ;
      RECT  128400.0 1604250.0 129600.0 1605450.0 ;
      RECT  128400.0 1604250.0 129600.0 1605450.0 ;
      RECT  126000.0 1604250.0 127200.0 1605450.0 ;
      RECT  126000.0 1594950.0 127200.0 1596150.0 ;
      RECT  128400.0 1594950.0 129600.0 1596150.0 ;
      RECT  128400.0 1594950.0 129600.0 1596150.0 ;
      RECT  126000.0 1594950.0 127200.0 1596150.0 ;
      RECT  130800.0 1604850.0 132000.0 1606050.0 ;
      RECT  130800.0 1594950.0 132000.0 1596150.0 ;
      RECT  126600.0 1599600.0 127800.0 1600800.0 ;
      RECT  126600.0 1599600.0 127800.0 1600800.0 ;
      RECT  129150.0 1599750.0 130050.0 1600650.0 ;
      RECT  124200.0 1606950.0 133800.0 1607850.0 ;
      RECT  124200.0 1593150.0 133800.0 1594050.0 ;
      RECT  135600.0 1595550.0 136800.0 1593150.0 ;
      RECT  135600.0 1604250.0 136800.0 1607850.0 ;
      RECT  140400.0 1604250.0 141600.0 1607850.0 ;
      RECT  142800.0 1605450.0 144000.0 1607400.0 ;
      RECT  142800.0 1593600.0 144000.0 1595550.0 ;
      RECT  135600.0 1604250.0 136800.0 1605450.0 ;
      RECT  138000.0 1604250.0 139200.0 1605450.0 ;
      RECT  138000.0 1604250.0 139200.0 1605450.0 ;
      RECT  135600.0 1604250.0 136800.0 1605450.0 ;
      RECT  138000.0 1604250.0 139200.0 1605450.0 ;
      RECT  140400.0 1604250.0 141600.0 1605450.0 ;
      RECT  140400.0 1604250.0 141600.0 1605450.0 ;
      RECT  138000.0 1604250.0 139200.0 1605450.0 ;
      RECT  135600.0 1595550.0 136800.0 1596750.0 ;
      RECT  138000.0 1595550.0 139200.0 1596750.0 ;
      RECT  138000.0 1595550.0 139200.0 1596750.0 ;
      RECT  135600.0 1595550.0 136800.0 1596750.0 ;
      RECT  138000.0 1595550.0 139200.0 1596750.0 ;
      RECT  140400.0 1595550.0 141600.0 1596750.0 ;
      RECT  140400.0 1595550.0 141600.0 1596750.0 ;
      RECT  138000.0 1595550.0 139200.0 1596750.0 ;
      RECT  142800.0 1604850.0 144000.0 1606050.0 ;
      RECT  142800.0 1594950.0 144000.0 1596150.0 ;
      RECT  140400.0 1598100.0 139200.0 1599300.0 ;
      RECT  137400.0 1600800.0 136200.0 1602000.0 ;
      RECT  138000.0 1604250.0 139200.0 1605450.0 ;
      RECT  140400.0 1595550.0 141600.0 1596750.0 ;
      RECT  141600.0 1600800.0 140400.0 1602000.0 ;
      RECT  136200.0 1600800.0 137400.0 1602000.0 ;
      RECT  139200.0 1598100.0 140400.0 1599300.0 ;
      RECT  140400.0 1600800.0 141600.0 1602000.0 ;
      RECT  133800.0 1606950.0 148200.0 1607850.0 ;
      RECT  133800.0 1593150.0 148200.0 1594050.0 ;
      RECT  154800.0 1605450.0 156000.0 1607400.0 ;
      RECT  154800.0 1593600.0 156000.0 1595550.0 ;
      RECT  150000.0 1594950.0 151200.0 1593150.0 ;
      RECT  150000.0 1604250.0 151200.0 1607850.0 ;
      RECT  152700.0 1594950.0 153600.0 1604250.0 ;
      RECT  150000.0 1604250.0 151200.0 1605450.0 ;
      RECT  152400.0 1604250.0 153600.0 1605450.0 ;
      RECT  152400.0 1604250.0 153600.0 1605450.0 ;
      RECT  150000.0 1604250.0 151200.0 1605450.0 ;
      RECT  150000.0 1594950.0 151200.0 1596150.0 ;
      RECT  152400.0 1594950.0 153600.0 1596150.0 ;
      RECT  152400.0 1594950.0 153600.0 1596150.0 ;
      RECT  150000.0 1594950.0 151200.0 1596150.0 ;
      RECT  154800.0 1604850.0 156000.0 1606050.0 ;
      RECT  154800.0 1594950.0 156000.0 1596150.0 ;
      RECT  150600.0 1599600.0 151800.0 1600800.0 ;
      RECT  150600.0 1599600.0 151800.0 1600800.0 ;
      RECT  153150.0 1599750.0 154050.0 1600650.0 ;
      RECT  148200.0 1606950.0 157800.0 1607850.0 ;
      RECT  148200.0 1593150.0 157800.0 1594050.0 ;
      RECT  120450.0 1599600.0 121650.0 1600800.0 ;
      RECT  122400.0 1597200.0 123600.0 1598400.0 ;
      RECT  139200.0 1598100.0 138000.0 1599300.0 ;
      RECT  130800.0 1609350.0 132000.0 1607400.0 ;
      RECT  130800.0 1621200.0 132000.0 1619250.0 ;
      RECT  126000.0 1619850.0 127200.0 1621650.0 ;
      RECT  126000.0 1610550.0 127200.0 1606950.0 ;
      RECT  128700.0 1619850.0 129600.0 1610550.0 ;
      RECT  126000.0 1610550.0 127200.0 1609350.0 ;
      RECT  128400.0 1610550.0 129600.0 1609350.0 ;
      RECT  128400.0 1610550.0 129600.0 1609350.0 ;
      RECT  126000.0 1610550.0 127200.0 1609350.0 ;
      RECT  126000.0 1619850.0 127200.0 1618650.0 ;
      RECT  128400.0 1619850.0 129600.0 1618650.0 ;
      RECT  128400.0 1619850.0 129600.0 1618650.0 ;
      RECT  126000.0 1619850.0 127200.0 1618650.0 ;
      RECT  130800.0 1609950.0 132000.0 1608750.0 ;
      RECT  130800.0 1619850.0 132000.0 1618650.0 ;
      RECT  126600.0 1615200.0 127800.0 1614000.0 ;
      RECT  126600.0 1615200.0 127800.0 1614000.0 ;
      RECT  129150.0 1615050.0 130050.0 1614150.0 ;
      RECT  124200.0 1607850.0 133800.0 1606950.0 ;
      RECT  124200.0 1621650.0 133800.0 1620750.0 ;
      RECT  135600.0 1619250.0 136800.0 1621650.0 ;
      RECT  135600.0 1610550.0 136800.0 1606950.0 ;
      RECT  140400.0 1610550.0 141600.0 1606950.0 ;
      RECT  142800.0 1609350.0 144000.0 1607400.0 ;
      RECT  142800.0 1621200.0 144000.0 1619250.0 ;
      RECT  135600.0 1610550.0 136800.0 1609350.0 ;
      RECT  138000.0 1610550.0 139200.0 1609350.0 ;
      RECT  138000.0 1610550.0 139200.0 1609350.0 ;
      RECT  135600.0 1610550.0 136800.0 1609350.0 ;
      RECT  138000.0 1610550.0 139200.0 1609350.0 ;
      RECT  140400.0 1610550.0 141600.0 1609350.0 ;
      RECT  140400.0 1610550.0 141600.0 1609350.0 ;
      RECT  138000.0 1610550.0 139200.0 1609350.0 ;
      RECT  135600.0 1619250.0 136800.0 1618050.0 ;
      RECT  138000.0 1619250.0 139200.0 1618050.0 ;
      RECT  138000.0 1619250.0 139200.0 1618050.0 ;
      RECT  135600.0 1619250.0 136800.0 1618050.0 ;
      RECT  138000.0 1619250.0 139200.0 1618050.0 ;
      RECT  140400.0 1619250.0 141600.0 1618050.0 ;
      RECT  140400.0 1619250.0 141600.0 1618050.0 ;
      RECT  138000.0 1619250.0 139200.0 1618050.0 ;
      RECT  142800.0 1609950.0 144000.0 1608750.0 ;
      RECT  142800.0 1619850.0 144000.0 1618650.0 ;
      RECT  140400.0 1616700.0 139200.0 1615500.0 ;
      RECT  137400.0 1614000.0 136200.0 1612800.0 ;
      RECT  138000.0 1610550.0 139200.0 1609350.0 ;
      RECT  140400.0 1619250.0 141600.0 1618050.0 ;
      RECT  141600.0 1614000.0 140400.0 1612800.0 ;
      RECT  136200.0 1614000.0 137400.0 1612800.0 ;
      RECT  139200.0 1616700.0 140400.0 1615500.0 ;
      RECT  140400.0 1614000.0 141600.0 1612800.0 ;
      RECT  133800.0 1607850.0 148200.0 1606950.0 ;
      RECT  133800.0 1621650.0 148200.0 1620750.0 ;
      RECT  154800.0 1609350.0 156000.0 1607400.0 ;
      RECT  154800.0 1621200.0 156000.0 1619250.0 ;
      RECT  150000.0 1619850.0 151200.0 1621650.0 ;
      RECT  150000.0 1610550.0 151200.0 1606950.0 ;
      RECT  152700.0 1619850.0 153600.0 1610550.0 ;
      RECT  150000.0 1610550.0 151200.0 1609350.0 ;
      RECT  152400.0 1610550.0 153600.0 1609350.0 ;
      RECT  152400.0 1610550.0 153600.0 1609350.0 ;
      RECT  150000.0 1610550.0 151200.0 1609350.0 ;
      RECT  150000.0 1619850.0 151200.0 1618650.0 ;
      RECT  152400.0 1619850.0 153600.0 1618650.0 ;
      RECT  152400.0 1619850.0 153600.0 1618650.0 ;
      RECT  150000.0 1619850.0 151200.0 1618650.0 ;
      RECT  154800.0 1609950.0 156000.0 1608750.0 ;
      RECT  154800.0 1619850.0 156000.0 1618650.0 ;
      RECT  150600.0 1615200.0 151800.0 1614000.0 ;
      RECT  150600.0 1615200.0 151800.0 1614000.0 ;
      RECT  153150.0 1615050.0 154050.0 1614150.0 ;
      RECT  148200.0 1607850.0 157800.0 1606950.0 ;
      RECT  148200.0 1621650.0 157800.0 1620750.0 ;
      RECT  120450.0 1614000.0 121650.0 1615200.0 ;
      RECT  122400.0 1616400.0 123600.0 1617600.0 ;
      RECT  139200.0 1615500.0 138000.0 1616700.0 ;
      RECT  130800.0 1633050.0 132000.0 1635000.0 ;
      RECT  130800.0 1621200.0 132000.0 1623150.0 ;
      RECT  126000.0 1622550.0 127200.0 1620750.0 ;
      RECT  126000.0 1631850.0 127200.0 1635450.0 ;
      RECT  128700.0 1622550.0 129600.0 1631850.0 ;
      RECT  126000.0 1631850.0 127200.0 1633050.0 ;
      RECT  128400.0 1631850.0 129600.0 1633050.0 ;
      RECT  128400.0 1631850.0 129600.0 1633050.0 ;
      RECT  126000.0 1631850.0 127200.0 1633050.0 ;
      RECT  126000.0 1622550.0 127200.0 1623750.0 ;
      RECT  128400.0 1622550.0 129600.0 1623750.0 ;
      RECT  128400.0 1622550.0 129600.0 1623750.0 ;
      RECT  126000.0 1622550.0 127200.0 1623750.0 ;
      RECT  130800.0 1632450.0 132000.0 1633650.0 ;
      RECT  130800.0 1622550.0 132000.0 1623750.0 ;
      RECT  126600.0 1627200.0 127800.0 1628400.0 ;
      RECT  126600.0 1627200.0 127800.0 1628400.0 ;
      RECT  129150.0 1627350.0 130050.0 1628250.0 ;
      RECT  124200.0 1634550.0 133800.0 1635450.0 ;
      RECT  124200.0 1620750.0 133800.0 1621650.0 ;
      RECT  135600.0 1623150.0 136800.0 1620750.0 ;
      RECT  135600.0 1631850.0 136800.0 1635450.0 ;
      RECT  140400.0 1631850.0 141600.0 1635450.0 ;
      RECT  142800.0 1633050.0 144000.0 1635000.0 ;
      RECT  142800.0 1621200.0 144000.0 1623150.0 ;
      RECT  135600.0 1631850.0 136800.0 1633050.0 ;
      RECT  138000.0 1631850.0 139200.0 1633050.0 ;
      RECT  138000.0 1631850.0 139200.0 1633050.0 ;
      RECT  135600.0 1631850.0 136800.0 1633050.0 ;
      RECT  138000.0 1631850.0 139200.0 1633050.0 ;
      RECT  140400.0 1631850.0 141600.0 1633050.0 ;
      RECT  140400.0 1631850.0 141600.0 1633050.0 ;
      RECT  138000.0 1631850.0 139200.0 1633050.0 ;
      RECT  135600.0 1623150.0 136800.0 1624350.0 ;
      RECT  138000.0 1623150.0 139200.0 1624350.0 ;
      RECT  138000.0 1623150.0 139200.0 1624350.0 ;
      RECT  135600.0 1623150.0 136800.0 1624350.0 ;
      RECT  138000.0 1623150.0 139200.0 1624350.0 ;
      RECT  140400.0 1623150.0 141600.0 1624350.0 ;
      RECT  140400.0 1623150.0 141600.0 1624350.0 ;
      RECT  138000.0 1623150.0 139200.0 1624350.0 ;
      RECT  142800.0 1632450.0 144000.0 1633650.0 ;
      RECT  142800.0 1622550.0 144000.0 1623750.0 ;
      RECT  140400.0 1625700.0 139200.0 1626900.0 ;
      RECT  137400.0 1628400.0 136200.0 1629600.0 ;
      RECT  138000.0 1631850.0 139200.0 1633050.0 ;
      RECT  140400.0 1623150.0 141600.0 1624350.0 ;
      RECT  141600.0 1628400.0 140400.0 1629600.0 ;
      RECT  136200.0 1628400.0 137400.0 1629600.0 ;
      RECT  139200.0 1625700.0 140400.0 1626900.0 ;
      RECT  140400.0 1628400.0 141600.0 1629600.0 ;
      RECT  133800.0 1634550.0 148200.0 1635450.0 ;
      RECT  133800.0 1620750.0 148200.0 1621650.0 ;
      RECT  154800.0 1633050.0 156000.0 1635000.0 ;
      RECT  154800.0 1621200.0 156000.0 1623150.0 ;
      RECT  150000.0 1622550.0 151200.0 1620750.0 ;
      RECT  150000.0 1631850.0 151200.0 1635450.0 ;
      RECT  152700.0 1622550.0 153600.0 1631850.0 ;
      RECT  150000.0 1631850.0 151200.0 1633050.0 ;
      RECT  152400.0 1631850.0 153600.0 1633050.0 ;
      RECT  152400.0 1631850.0 153600.0 1633050.0 ;
      RECT  150000.0 1631850.0 151200.0 1633050.0 ;
      RECT  150000.0 1622550.0 151200.0 1623750.0 ;
      RECT  152400.0 1622550.0 153600.0 1623750.0 ;
      RECT  152400.0 1622550.0 153600.0 1623750.0 ;
      RECT  150000.0 1622550.0 151200.0 1623750.0 ;
      RECT  154800.0 1632450.0 156000.0 1633650.0 ;
      RECT  154800.0 1622550.0 156000.0 1623750.0 ;
      RECT  150600.0 1627200.0 151800.0 1628400.0 ;
      RECT  150600.0 1627200.0 151800.0 1628400.0 ;
      RECT  153150.0 1627350.0 154050.0 1628250.0 ;
      RECT  148200.0 1634550.0 157800.0 1635450.0 ;
      RECT  148200.0 1620750.0 157800.0 1621650.0 ;
      RECT  120450.0 1627200.0 121650.0 1628400.0 ;
      RECT  122400.0 1624800.0 123600.0 1626000.0 ;
      RECT  139200.0 1625700.0 138000.0 1626900.0 ;
      RECT  130800.0 1636950.0 132000.0 1635000.0 ;
      RECT  130800.0 1648800.0 132000.0 1646850.0 ;
      RECT  126000.0 1647450.0 127200.0 1649250.0 ;
      RECT  126000.0 1638150.0 127200.0 1634550.0 ;
      RECT  128700.0 1647450.0 129600.0 1638150.0 ;
      RECT  126000.0 1638150.0 127200.0 1636950.0 ;
      RECT  128400.0 1638150.0 129600.0 1636950.0 ;
      RECT  128400.0 1638150.0 129600.0 1636950.0 ;
      RECT  126000.0 1638150.0 127200.0 1636950.0 ;
      RECT  126000.0 1647450.0 127200.0 1646250.0 ;
      RECT  128400.0 1647450.0 129600.0 1646250.0 ;
      RECT  128400.0 1647450.0 129600.0 1646250.0 ;
      RECT  126000.0 1647450.0 127200.0 1646250.0 ;
      RECT  130800.0 1637550.0 132000.0 1636350.0 ;
      RECT  130800.0 1647450.0 132000.0 1646250.0 ;
      RECT  126600.0 1642800.0 127800.0 1641600.0 ;
      RECT  126600.0 1642800.0 127800.0 1641600.0 ;
      RECT  129150.0 1642650.0 130050.0 1641750.0 ;
      RECT  124200.0 1635450.0 133800.0 1634550.0 ;
      RECT  124200.0 1649250.0 133800.0 1648350.0 ;
      RECT  135600.0 1646850.0 136800.0 1649250.0 ;
      RECT  135600.0 1638150.0 136800.0 1634550.0 ;
      RECT  140400.0 1638150.0 141600.0 1634550.0 ;
      RECT  142800.0 1636950.0 144000.0 1635000.0 ;
      RECT  142800.0 1648800.0 144000.0 1646850.0 ;
      RECT  135600.0 1638150.0 136800.0 1636950.0 ;
      RECT  138000.0 1638150.0 139200.0 1636950.0 ;
      RECT  138000.0 1638150.0 139200.0 1636950.0 ;
      RECT  135600.0 1638150.0 136800.0 1636950.0 ;
      RECT  138000.0 1638150.0 139200.0 1636950.0 ;
      RECT  140400.0 1638150.0 141600.0 1636950.0 ;
      RECT  140400.0 1638150.0 141600.0 1636950.0 ;
      RECT  138000.0 1638150.0 139200.0 1636950.0 ;
      RECT  135600.0 1646850.0 136800.0 1645650.0 ;
      RECT  138000.0 1646850.0 139200.0 1645650.0 ;
      RECT  138000.0 1646850.0 139200.0 1645650.0 ;
      RECT  135600.0 1646850.0 136800.0 1645650.0 ;
      RECT  138000.0 1646850.0 139200.0 1645650.0 ;
      RECT  140400.0 1646850.0 141600.0 1645650.0 ;
      RECT  140400.0 1646850.0 141600.0 1645650.0 ;
      RECT  138000.0 1646850.0 139200.0 1645650.0 ;
      RECT  142800.0 1637550.0 144000.0 1636350.0 ;
      RECT  142800.0 1647450.0 144000.0 1646250.0 ;
      RECT  140400.0 1644300.0 139200.0 1643100.0 ;
      RECT  137400.0 1641600.0 136200.0 1640400.0 ;
      RECT  138000.0 1638150.0 139200.0 1636950.0 ;
      RECT  140400.0 1646850.0 141600.0 1645650.0 ;
      RECT  141600.0 1641600.0 140400.0 1640400.0 ;
      RECT  136200.0 1641600.0 137400.0 1640400.0 ;
      RECT  139200.0 1644300.0 140400.0 1643100.0 ;
      RECT  140400.0 1641600.0 141600.0 1640400.0 ;
      RECT  133800.0 1635450.0 148200.0 1634550.0 ;
      RECT  133800.0 1649250.0 148200.0 1648350.0 ;
      RECT  154800.0 1636950.0 156000.0 1635000.0 ;
      RECT  154800.0 1648800.0 156000.0 1646850.0 ;
      RECT  150000.0 1647450.0 151200.0 1649250.0 ;
      RECT  150000.0 1638150.0 151200.0 1634550.0 ;
      RECT  152700.0 1647450.0 153600.0 1638150.0 ;
      RECT  150000.0 1638150.0 151200.0 1636950.0 ;
      RECT  152400.0 1638150.0 153600.0 1636950.0 ;
      RECT  152400.0 1638150.0 153600.0 1636950.0 ;
      RECT  150000.0 1638150.0 151200.0 1636950.0 ;
      RECT  150000.0 1647450.0 151200.0 1646250.0 ;
      RECT  152400.0 1647450.0 153600.0 1646250.0 ;
      RECT  152400.0 1647450.0 153600.0 1646250.0 ;
      RECT  150000.0 1647450.0 151200.0 1646250.0 ;
      RECT  154800.0 1637550.0 156000.0 1636350.0 ;
      RECT  154800.0 1647450.0 156000.0 1646250.0 ;
      RECT  150600.0 1642800.0 151800.0 1641600.0 ;
      RECT  150600.0 1642800.0 151800.0 1641600.0 ;
      RECT  153150.0 1642650.0 154050.0 1641750.0 ;
      RECT  148200.0 1635450.0 157800.0 1634550.0 ;
      RECT  148200.0 1649250.0 157800.0 1648350.0 ;
      RECT  120450.0 1641600.0 121650.0 1642800.0 ;
      RECT  122400.0 1644000.0 123600.0 1645200.0 ;
      RECT  139200.0 1643100.0 138000.0 1644300.0 ;
      RECT  130800.0 1660650.0 132000.0 1662600.0 ;
      RECT  130800.0 1648800.0 132000.0 1650750.0 ;
      RECT  126000.0 1650150.0 127200.0 1648350.0 ;
      RECT  126000.0 1659450.0 127200.0 1663050.0 ;
      RECT  128700.0 1650150.0 129600.0 1659450.0 ;
      RECT  126000.0 1659450.0 127200.0 1660650.0 ;
      RECT  128400.0 1659450.0 129600.0 1660650.0 ;
      RECT  128400.0 1659450.0 129600.0 1660650.0 ;
      RECT  126000.0 1659450.0 127200.0 1660650.0 ;
      RECT  126000.0 1650150.0 127200.0 1651350.0 ;
      RECT  128400.0 1650150.0 129600.0 1651350.0 ;
      RECT  128400.0 1650150.0 129600.0 1651350.0 ;
      RECT  126000.0 1650150.0 127200.0 1651350.0 ;
      RECT  130800.0 1660050.0 132000.0 1661250.0 ;
      RECT  130800.0 1650150.0 132000.0 1651350.0 ;
      RECT  126600.0 1654800.0 127800.0 1656000.0 ;
      RECT  126600.0 1654800.0 127800.0 1656000.0 ;
      RECT  129150.0 1654950.0 130050.0 1655850.0 ;
      RECT  124200.0 1662150.0 133800.0 1663050.0 ;
      RECT  124200.0 1648350.0 133800.0 1649250.0 ;
      RECT  135600.0 1650750.0 136800.0 1648350.0 ;
      RECT  135600.0 1659450.0 136800.0 1663050.0 ;
      RECT  140400.0 1659450.0 141600.0 1663050.0 ;
      RECT  142800.0 1660650.0 144000.0 1662600.0 ;
      RECT  142800.0 1648800.0 144000.0 1650750.0 ;
      RECT  135600.0 1659450.0 136800.0 1660650.0 ;
      RECT  138000.0 1659450.0 139200.0 1660650.0 ;
      RECT  138000.0 1659450.0 139200.0 1660650.0 ;
      RECT  135600.0 1659450.0 136800.0 1660650.0 ;
      RECT  138000.0 1659450.0 139200.0 1660650.0 ;
      RECT  140400.0 1659450.0 141600.0 1660650.0 ;
      RECT  140400.0 1659450.0 141600.0 1660650.0 ;
      RECT  138000.0 1659450.0 139200.0 1660650.0 ;
      RECT  135600.0 1650750.0 136800.0 1651950.0 ;
      RECT  138000.0 1650750.0 139200.0 1651950.0 ;
      RECT  138000.0 1650750.0 139200.0 1651950.0 ;
      RECT  135600.0 1650750.0 136800.0 1651950.0 ;
      RECT  138000.0 1650750.0 139200.0 1651950.0 ;
      RECT  140400.0 1650750.0 141600.0 1651950.0 ;
      RECT  140400.0 1650750.0 141600.0 1651950.0 ;
      RECT  138000.0 1650750.0 139200.0 1651950.0 ;
      RECT  142800.0 1660050.0 144000.0 1661250.0 ;
      RECT  142800.0 1650150.0 144000.0 1651350.0 ;
      RECT  140400.0 1653300.0 139200.0 1654500.0 ;
      RECT  137400.0 1656000.0 136200.0 1657200.0 ;
      RECT  138000.0 1659450.0 139200.0 1660650.0 ;
      RECT  140400.0 1650750.0 141600.0 1651950.0 ;
      RECT  141600.0 1656000.0 140400.0 1657200.0 ;
      RECT  136200.0 1656000.0 137400.0 1657200.0 ;
      RECT  139200.0 1653300.0 140400.0 1654500.0 ;
      RECT  140400.0 1656000.0 141600.0 1657200.0 ;
      RECT  133800.0 1662150.0 148200.0 1663050.0 ;
      RECT  133800.0 1648350.0 148200.0 1649250.0 ;
      RECT  154800.0 1660650.0 156000.0 1662600.0 ;
      RECT  154800.0 1648800.0 156000.0 1650750.0 ;
      RECT  150000.0 1650150.0 151200.0 1648350.0 ;
      RECT  150000.0 1659450.0 151200.0 1663050.0 ;
      RECT  152700.0 1650150.0 153600.0 1659450.0 ;
      RECT  150000.0 1659450.0 151200.0 1660650.0 ;
      RECT  152400.0 1659450.0 153600.0 1660650.0 ;
      RECT  152400.0 1659450.0 153600.0 1660650.0 ;
      RECT  150000.0 1659450.0 151200.0 1660650.0 ;
      RECT  150000.0 1650150.0 151200.0 1651350.0 ;
      RECT  152400.0 1650150.0 153600.0 1651350.0 ;
      RECT  152400.0 1650150.0 153600.0 1651350.0 ;
      RECT  150000.0 1650150.0 151200.0 1651350.0 ;
      RECT  154800.0 1660050.0 156000.0 1661250.0 ;
      RECT  154800.0 1650150.0 156000.0 1651350.0 ;
      RECT  150600.0 1654800.0 151800.0 1656000.0 ;
      RECT  150600.0 1654800.0 151800.0 1656000.0 ;
      RECT  153150.0 1654950.0 154050.0 1655850.0 ;
      RECT  148200.0 1662150.0 157800.0 1663050.0 ;
      RECT  148200.0 1648350.0 157800.0 1649250.0 ;
      RECT  120450.0 1654800.0 121650.0 1656000.0 ;
      RECT  122400.0 1652400.0 123600.0 1653600.0 ;
      RECT  139200.0 1653300.0 138000.0 1654500.0 ;
      RECT  130800.0 1664550.0 132000.0 1662600.0 ;
      RECT  130800.0 1676400.0 132000.0 1674450.0 ;
      RECT  126000.0 1675050.0 127200.0 1676850.0 ;
      RECT  126000.0 1665750.0 127200.0 1662150.0 ;
      RECT  128700.0 1675050.0 129600.0 1665750.0 ;
      RECT  126000.0 1665750.0 127200.0 1664550.0 ;
      RECT  128400.0 1665750.0 129600.0 1664550.0 ;
      RECT  128400.0 1665750.0 129600.0 1664550.0 ;
      RECT  126000.0 1665750.0 127200.0 1664550.0 ;
      RECT  126000.0 1675050.0 127200.0 1673850.0 ;
      RECT  128400.0 1675050.0 129600.0 1673850.0 ;
      RECT  128400.0 1675050.0 129600.0 1673850.0 ;
      RECT  126000.0 1675050.0 127200.0 1673850.0 ;
      RECT  130800.0 1665150.0 132000.0 1663950.0 ;
      RECT  130800.0 1675050.0 132000.0 1673850.0 ;
      RECT  126600.0 1670400.0 127800.0 1669200.0 ;
      RECT  126600.0 1670400.0 127800.0 1669200.0 ;
      RECT  129150.0 1670250.0 130050.0 1669350.0 ;
      RECT  124200.0 1663050.0 133800.0 1662150.0 ;
      RECT  124200.0 1676850.0 133800.0 1675950.0 ;
      RECT  135600.0 1674450.0 136800.0 1676850.0 ;
      RECT  135600.0 1665750.0 136800.0 1662150.0 ;
      RECT  140400.0 1665750.0 141600.0 1662150.0 ;
      RECT  142800.0 1664550.0 144000.0 1662600.0 ;
      RECT  142800.0 1676400.0 144000.0 1674450.0 ;
      RECT  135600.0 1665750.0 136800.0 1664550.0 ;
      RECT  138000.0 1665750.0 139200.0 1664550.0 ;
      RECT  138000.0 1665750.0 139200.0 1664550.0 ;
      RECT  135600.0 1665750.0 136800.0 1664550.0 ;
      RECT  138000.0 1665750.0 139200.0 1664550.0 ;
      RECT  140400.0 1665750.0 141600.0 1664550.0 ;
      RECT  140400.0 1665750.0 141600.0 1664550.0 ;
      RECT  138000.0 1665750.0 139200.0 1664550.0 ;
      RECT  135600.0 1674450.0 136800.0 1673250.0 ;
      RECT  138000.0 1674450.0 139200.0 1673250.0 ;
      RECT  138000.0 1674450.0 139200.0 1673250.0 ;
      RECT  135600.0 1674450.0 136800.0 1673250.0 ;
      RECT  138000.0 1674450.0 139200.0 1673250.0 ;
      RECT  140400.0 1674450.0 141600.0 1673250.0 ;
      RECT  140400.0 1674450.0 141600.0 1673250.0 ;
      RECT  138000.0 1674450.0 139200.0 1673250.0 ;
      RECT  142800.0 1665150.0 144000.0 1663950.0 ;
      RECT  142800.0 1675050.0 144000.0 1673850.0 ;
      RECT  140400.0 1671900.0 139200.0 1670700.0 ;
      RECT  137400.0 1669200.0 136200.0 1668000.0 ;
      RECT  138000.0 1665750.0 139200.0 1664550.0 ;
      RECT  140400.0 1674450.0 141600.0 1673250.0 ;
      RECT  141600.0 1669200.0 140400.0 1668000.0 ;
      RECT  136200.0 1669200.0 137400.0 1668000.0 ;
      RECT  139200.0 1671900.0 140400.0 1670700.0 ;
      RECT  140400.0 1669200.0 141600.0 1668000.0 ;
      RECT  133800.0 1663050.0 148200.0 1662150.0 ;
      RECT  133800.0 1676850.0 148200.0 1675950.0 ;
      RECT  154800.0 1664550.0 156000.0 1662600.0 ;
      RECT  154800.0 1676400.0 156000.0 1674450.0 ;
      RECT  150000.0 1675050.0 151200.0 1676850.0 ;
      RECT  150000.0 1665750.0 151200.0 1662150.0 ;
      RECT  152700.0 1675050.0 153600.0 1665750.0 ;
      RECT  150000.0 1665750.0 151200.0 1664550.0 ;
      RECT  152400.0 1665750.0 153600.0 1664550.0 ;
      RECT  152400.0 1665750.0 153600.0 1664550.0 ;
      RECT  150000.0 1665750.0 151200.0 1664550.0 ;
      RECT  150000.0 1675050.0 151200.0 1673850.0 ;
      RECT  152400.0 1675050.0 153600.0 1673850.0 ;
      RECT  152400.0 1675050.0 153600.0 1673850.0 ;
      RECT  150000.0 1675050.0 151200.0 1673850.0 ;
      RECT  154800.0 1665150.0 156000.0 1663950.0 ;
      RECT  154800.0 1675050.0 156000.0 1673850.0 ;
      RECT  150600.0 1670400.0 151800.0 1669200.0 ;
      RECT  150600.0 1670400.0 151800.0 1669200.0 ;
      RECT  153150.0 1670250.0 154050.0 1669350.0 ;
      RECT  148200.0 1663050.0 157800.0 1662150.0 ;
      RECT  148200.0 1676850.0 157800.0 1675950.0 ;
      RECT  120450.0 1669200.0 121650.0 1670400.0 ;
      RECT  122400.0 1671600.0 123600.0 1672800.0 ;
      RECT  139200.0 1670700.0 138000.0 1671900.0 ;
      RECT  130800.0 1688250.0 132000.0 1690200.0 ;
      RECT  130800.0 1676400.0 132000.0 1678350.0 ;
      RECT  126000.0 1677750.0 127200.0 1675950.0 ;
      RECT  126000.0 1687050.0 127200.0 1690650.0 ;
      RECT  128700.0 1677750.0 129600.0 1687050.0 ;
      RECT  126000.0 1687050.0 127200.0 1688250.0 ;
      RECT  128400.0 1687050.0 129600.0 1688250.0 ;
      RECT  128400.0 1687050.0 129600.0 1688250.0 ;
      RECT  126000.0 1687050.0 127200.0 1688250.0 ;
      RECT  126000.0 1677750.0 127200.0 1678950.0 ;
      RECT  128400.0 1677750.0 129600.0 1678950.0 ;
      RECT  128400.0 1677750.0 129600.0 1678950.0 ;
      RECT  126000.0 1677750.0 127200.0 1678950.0 ;
      RECT  130800.0 1687650.0 132000.0 1688850.0 ;
      RECT  130800.0 1677750.0 132000.0 1678950.0 ;
      RECT  126600.0 1682400.0 127800.0 1683600.0 ;
      RECT  126600.0 1682400.0 127800.0 1683600.0 ;
      RECT  129150.0 1682550.0 130050.0 1683450.0 ;
      RECT  124200.0 1689750.0 133800.0 1690650.0 ;
      RECT  124200.0 1675950.0 133800.0 1676850.0 ;
      RECT  135600.0 1678350.0 136800.0 1675950.0 ;
      RECT  135600.0 1687050.0 136800.0 1690650.0 ;
      RECT  140400.0 1687050.0 141600.0 1690650.0 ;
      RECT  142800.0 1688250.0 144000.0 1690200.0 ;
      RECT  142800.0 1676400.0 144000.0 1678350.0 ;
      RECT  135600.0 1687050.0 136800.0 1688250.0 ;
      RECT  138000.0 1687050.0 139200.0 1688250.0 ;
      RECT  138000.0 1687050.0 139200.0 1688250.0 ;
      RECT  135600.0 1687050.0 136800.0 1688250.0 ;
      RECT  138000.0 1687050.0 139200.0 1688250.0 ;
      RECT  140400.0 1687050.0 141600.0 1688250.0 ;
      RECT  140400.0 1687050.0 141600.0 1688250.0 ;
      RECT  138000.0 1687050.0 139200.0 1688250.0 ;
      RECT  135600.0 1678350.0 136800.0 1679550.0 ;
      RECT  138000.0 1678350.0 139200.0 1679550.0 ;
      RECT  138000.0 1678350.0 139200.0 1679550.0 ;
      RECT  135600.0 1678350.0 136800.0 1679550.0 ;
      RECT  138000.0 1678350.0 139200.0 1679550.0 ;
      RECT  140400.0 1678350.0 141600.0 1679550.0 ;
      RECT  140400.0 1678350.0 141600.0 1679550.0 ;
      RECT  138000.0 1678350.0 139200.0 1679550.0 ;
      RECT  142800.0 1687650.0 144000.0 1688850.0 ;
      RECT  142800.0 1677750.0 144000.0 1678950.0 ;
      RECT  140400.0 1680900.0 139200.0 1682100.0 ;
      RECT  137400.0 1683600.0 136200.0 1684800.0 ;
      RECT  138000.0 1687050.0 139200.0 1688250.0 ;
      RECT  140400.0 1678350.0 141600.0 1679550.0 ;
      RECT  141600.0 1683600.0 140400.0 1684800.0 ;
      RECT  136200.0 1683600.0 137400.0 1684800.0 ;
      RECT  139200.0 1680900.0 140400.0 1682100.0 ;
      RECT  140400.0 1683600.0 141600.0 1684800.0 ;
      RECT  133800.0 1689750.0 148200.0 1690650.0 ;
      RECT  133800.0 1675950.0 148200.0 1676850.0 ;
      RECT  154800.0 1688250.0 156000.0 1690200.0 ;
      RECT  154800.0 1676400.0 156000.0 1678350.0 ;
      RECT  150000.0 1677750.0 151200.0 1675950.0 ;
      RECT  150000.0 1687050.0 151200.0 1690650.0 ;
      RECT  152700.0 1677750.0 153600.0 1687050.0 ;
      RECT  150000.0 1687050.0 151200.0 1688250.0 ;
      RECT  152400.0 1687050.0 153600.0 1688250.0 ;
      RECT  152400.0 1687050.0 153600.0 1688250.0 ;
      RECT  150000.0 1687050.0 151200.0 1688250.0 ;
      RECT  150000.0 1677750.0 151200.0 1678950.0 ;
      RECT  152400.0 1677750.0 153600.0 1678950.0 ;
      RECT  152400.0 1677750.0 153600.0 1678950.0 ;
      RECT  150000.0 1677750.0 151200.0 1678950.0 ;
      RECT  154800.0 1687650.0 156000.0 1688850.0 ;
      RECT  154800.0 1677750.0 156000.0 1678950.0 ;
      RECT  150600.0 1682400.0 151800.0 1683600.0 ;
      RECT  150600.0 1682400.0 151800.0 1683600.0 ;
      RECT  153150.0 1682550.0 154050.0 1683450.0 ;
      RECT  148200.0 1689750.0 157800.0 1690650.0 ;
      RECT  148200.0 1675950.0 157800.0 1676850.0 ;
      RECT  120450.0 1682400.0 121650.0 1683600.0 ;
      RECT  122400.0 1680000.0 123600.0 1681200.0 ;
      RECT  139200.0 1680900.0 138000.0 1682100.0 ;
      RECT  130800.0 1692150.0 132000.0 1690200.0 ;
      RECT  130800.0 1704000.0 132000.0 1702050.0 ;
      RECT  126000.0 1702650.0 127200.0 1704450.0 ;
      RECT  126000.0 1693350.0 127200.0 1689750.0 ;
      RECT  128700.0 1702650.0 129600.0 1693350.0 ;
      RECT  126000.0 1693350.0 127200.0 1692150.0 ;
      RECT  128400.0 1693350.0 129600.0 1692150.0 ;
      RECT  128400.0 1693350.0 129600.0 1692150.0 ;
      RECT  126000.0 1693350.0 127200.0 1692150.0 ;
      RECT  126000.0 1702650.0 127200.0 1701450.0 ;
      RECT  128400.0 1702650.0 129600.0 1701450.0 ;
      RECT  128400.0 1702650.0 129600.0 1701450.0 ;
      RECT  126000.0 1702650.0 127200.0 1701450.0 ;
      RECT  130800.0 1692750.0 132000.0 1691550.0 ;
      RECT  130800.0 1702650.0 132000.0 1701450.0 ;
      RECT  126600.0 1698000.0 127800.0 1696800.0 ;
      RECT  126600.0 1698000.0 127800.0 1696800.0 ;
      RECT  129150.0 1697850.0 130050.0 1696950.0 ;
      RECT  124200.0 1690650.0 133800.0 1689750.0 ;
      RECT  124200.0 1704450.0 133800.0 1703550.0 ;
      RECT  135600.0 1702050.0 136800.0 1704450.0 ;
      RECT  135600.0 1693350.0 136800.0 1689750.0 ;
      RECT  140400.0 1693350.0 141600.0 1689750.0 ;
      RECT  142800.0 1692150.0 144000.0 1690200.0 ;
      RECT  142800.0 1704000.0 144000.0 1702050.0 ;
      RECT  135600.0 1693350.0 136800.0 1692150.0 ;
      RECT  138000.0 1693350.0 139200.0 1692150.0 ;
      RECT  138000.0 1693350.0 139200.0 1692150.0 ;
      RECT  135600.0 1693350.0 136800.0 1692150.0 ;
      RECT  138000.0 1693350.0 139200.0 1692150.0 ;
      RECT  140400.0 1693350.0 141600.0 1692150.0 ;
      RECT  140400.0 1693350.0 141600.0 1692150.0 ;
      RECT  138000.0 1693350.0 139200.0 1692150.0 ;
      RECT  135600.0 1702050.0 136800.0 1700850.0 ;
      RECT  138000.0 1702050.0 139200.0 1700850.0 ;
      RECT  138000.0 1702050.0 139200.0 1700850.0 ;
      RECT  135600.0 1702050.0 136800.0 1700850.0 ;
      RECT  138000.0 1702050.0 139200.0 1700850.0 ;
      RECT  140400.0 1702050.0 141600.0 1700850.0 ;
      RECT  140400.0 1702050.0 141600.0 1700850.0 ;
      RECT  138000.0 1702050.0 139200.0 1700850.0 ;
      RECT  142800.0 1692750.0 144000.0 1691550.0 ;
      RECT  142800.0 1702650.0 144000.0 1701450.0 ;
      RECT  140400.0 1699500.0 139200.0 1698300.0 ;
      RECT  137400.0 1696800.0 136200.0 1695600.0 ;
      RECT  138000.0 1693350.0 139200.0 1692150.0 ;
      RECT  140400.0 1702050.0 141600.0 1700850.0 ;
      RECT  141600.0 1696800.0 140400.0 1695600.0 ;
      RECT  136200.0 1696800.0 137400.0 1695600.0 ;
      RECT  139200.0 1699500.0 140400.0 1698300.0 ;
      RECT  140400.0 1696800.0 141600.0 1695600.0 ;
      RECT  133800.0 1690650.0 148200.0 1689750.0 ;
      RECT  133800.0 1704450.0 148200.0 1703550.0 ;
      RECT  154800.0 1692150.0 156000.0 1690200.0 ;
      RECT  154800.0 1704000.0 156000.0 1702050.0 ;
      RECT  150000.0 1702650.0 151200.0 1704450.0 ;
      RECT  150000.0 1693350.0 151200.0 1689750.0 ;
      RECT  152700.0 1702650.0 153600.0 1693350.0 ;
      RECT  150000.0 1693350.0 151200.0 1692150.0 ;
      RECT  152400.0 1693350.0 153600.0 1692150.0 ;
      RECT  152400.0 1693350.0 153600.0 1692150.0 ;
      RECT  150000.0 1693350.0 151200.0 1692150.0 ;
      RECT  150000.0 1702650.0 151200.0 1701450.0 ;
      RECT  152400.0 1702650.0 153600.0 1701450.0 ;
      RECT  152400.0 1702650.0 153600.0 1701450.0 ;
      RECT  150000.0 1702650.0 151200.0 1701450.0 ;
      RECT  154800.0 1692750.0 156000.0 1691550.0 ;
      RECT  154800.0 1702650.0 156000.0 1701450.0 ;
      RECT  150600.0 1698000.0 151800.0 1696800.0 ;
      RECT  150600.0 1698000.0 151800.0 1696800.0 ;
      RECT  153150.0 1697850.0 154050.0 1696950.0 ;
      RECT  148200.0 1690650.0 157800.0 1689750.0 ;
      RECT  148200.0 1704450.0 157800.0 1703550.0 ;
      RECT  120450.0 1696800.0 121650.0 1698000.0 ;
      RECT  122400.0 1699200.0 123600.0 1700400.0 ;
      RECT  139200.0 1698300.0 138000.0 1699500.0 ;
      RECT  130800.0 1715850.0 132000.0 1717800.0 ;
      RECT  130800.0 1704000.0 132000.0 1705950.0 ;
      RECT  126000.0 1705350.0 127200.0 1703550.0 ;
      RECT  126000.0 1714650.0 127200.0 1718250.0 ;
      RECT  128700.0 1705350.0 129600.0 1714650.0 ;
      RECT  126000.0 1714650.0 127200.0 1715850.0 ;
      RECT  128400.0 1714650.0 129600.0 1715850.0 ;
      RECT  128400.0 1714650.0 129600.0 1715850.0 ;
      RECT  126000.0 1714650.0 127200.0 1715850.0 ;
      RECT  126000.0 1705350.0 127200.0 1706550.0 ;
      RECT  128400.0 1705350.0 129600.0 1706550.0 ;
      RECT  128400.0 1705350.0 129600.0 1706550.0 ;
      RECT  126000.0 1705350.0 127200.0 1706550.0 ;
      RECT  130800.0 1715250.0 132000.0 1716450.0 ;
      RECT  130800.0 1705350.0 132000.0 1706550.0 ;
      RECT  126600.0 1710000.0 127800.0 1711200.0 ;
      RECT  126600.0 1710000.0 127800.0 1711200.0 ;
      RECT  129150.0 1710150.0 130050.0 1711050.0 ;
      RECT  124200.0 1717350.0 133800.0 1718250.0 ;
      RECT  124200.0 1703550.0 133800.0 1704450.0 ;
      RECT  135600.0 1705950.0 136800.0 1703550.0 ;
      RECT  135600.0 1714650.0 136800.0 1718250.0 ;
      RECT  140400.0 1714650.0 141600.0 1718250.0 ;
      RECT  142800.0 1715850.0 144000.0 1717800.0 ;
      RECT  142800.0 1704000.0 144000.0 1705950.0 ;
      RECT  135600.0 1714650.0 136800.0 1715850.0 ;
      RECT  138000.0 1714650.0 139200.0 1715850.0 ;
      RECT  138000.0 1714650.0 139200.0 1715850.0 ;
      RECT  135600.0 1714650.0 136800.0 1715850.0 ;
      RECT  138000.0 1714650.0 139200.0 1715850.0 ;
      RECT  140400.0 1714650.0 141600.0 1715850.0 ;
      RECT  140400.0 1714650.0 141600.0 1715850.0 ;
      RECT  138000.0 1714650.0 139200.0 1715850.0 ;
      RECT  135600.0 1705950.0 136800.0 1707150.0 ;
      RECT  138000.0 1705950.0 139200.0 1707150.0 ;
      RECT  138000.0 1705950.0 139200.0 1707150.0 ;
      RECT  135600.0 1705950.0 136800.0 1707150.0 ;
      RECT  138000.0 1705950.0 139200.0 1707150.0 ;
      RECT  140400.0 1705950.0 141600.0 1707150.0 ;
      RECT  140400.0 1705950.0 141600.0 1707150.0 ;
      RECT  138000.0 1705950.0 139200.0 1707150.0 ;
      RECT  142800.0 1715250.0 144000.0 1716450.0 ;
      RECT  142800.0 1705350.0 144000.0 1706550.0 ;
      RECT  140400.0 1708500.0 139200.0 1709700.0 ;
      RECT  137400.0 1711200.0 136200.0 1712400.0 ;
      RECT  138000.0 1714650.0 139200.0 1715850.0 ;
      RECT  140400.0 1705950.0 141600.0 1707150.0 ;
      RECT  141600.0 1711200.0 140400.0 1712400.0 ;
      RECT  136200.0 1711200.0 137400.0 1712400.0 ;
      RECT  139200.0 1708500.0 140400.0 1709700.0 ;
      RECT  140400.0 1711200.0 141600.0 1712400.0 ;
      RECT  133800.0 1717350.0 148200.0 1718250.0 ;
      RECT  133800.0 1703550.0 148200.0 1704450.0 ;
      RECT  154800.0 1715850.0 156000.0 1717800.0 ;
      RECT  154800.0 1704000.0 156000.0 1705950.0 ;
      RECT  150000.0 1705350.0 151200.0 1703550.0 ;
      RECT  150000.0 1714650.0 151200.0 1718250.0 ;
      RECT  152700.0 1705350.0 153600.0 1714650.0 ;
      RECT  150000.0 1714650.0 151200.0 1715850.0 ;
      RECT  152400.0 1714650.0 153600.0 1715850.0 ;
      RECT  152400.0 1714650.0 153600.0 1715850.0 ;
      RECT  150000.0 1714650.0 151200.0 1715850.0 ;
      RECT  150000.0 1705350.0 151200.0 1706550.0 ;
      RECT  152400.0 1705350.0 153600.0 1706550.0 ;
      RECT  152400.0 1705350.0 153600.0 1706550.0 ;
      RECT  150000.0 1705350.0 151200.0 1706550.0 ;
      RECT  154800.0 1715250.0 156000.0 1716450.0 ;
      RECT  154800.0 1705350.0 156000.0 1706550.0 ;
      RECT  150600.0 1710000.0 151800.0 1711200.0 ;
      RECT  150600.0 1710000.0 151800.0 1711200.0 ;
      RECT  153150.0 1710150.0 154050.0 1711050.0 ;
      RECT  148200.0 1717350.0 157800.0 1718250.0 ;
      RECT  148200.0 1703550.0 157800.0 1704450.0 ;
      RECT  120450.0 1710000.0 121650.0 1711200.0 ;
      RECT  122400.0 1707600.0 123600.0 1708800.0 ;
      RECT  139200.0 1708500.0 138000.0 1709700.0 ;
      RECT  130800.0 1719750.0 132000.0 1717800.0 ;
      RECT  130800.0 1731600.0 132000.0 1729650.0 ;
      RECT  126000.0 1730250.0 127200.0 1732050.0 ;
      RECT  126000.0 1720950.0 127200.0 1717350.0 ;
      RECT  128700.0 1730250.0 129600.0 1720950.0 ;
      RECT  126000.0 1720950.0 127200.0 1719750.0 ;
      RECT  128400.0 1720950.0 129600.0 1719750.0 ;
      RECT  128400.0 1720950.0 129600.0 1719750.0 ;
      RECT  126000.0 1720950.0 127200.0 1719750.0 ;
      RECT  126000.0 1730250.0 127200.0 1729050.0 ;
      RECT  128400.0 1730250.0 129600.0 1729050.0 ;
      RECT  128400.0 1730250.0 129600.0 1729050.0 ;
      RECT  126000.0 1730250.0 127200.0 1729050.0 ;
      RECT  130800.0 1720350.0 132000.0 1719150.0 ;
      RECT  130800.0 1730250.0 132000.0 1729050.0 ;
      RECT  126600.0 1725600.0 127800.0 1724400.0 ;
      RECT  126600.0 1725600.0 127800.0 1724400.0 ;
      RECT  129150.0 1725450.0 130050.0 1724550.0 ;
      RECT  124200.0 1718250.0 133800.0 1717350.0 ;
      RECT  124200.0 1732050.0 133800.0 1731150.0 ;
      RECT  135600.0 1729650.0 136800.0 1732050.0 ;
      RECT  135600.0 1720950.0 136800.0 1717350.0 ;
      RECT  140400.0 1720950.0 141600.0 1717350.0 ;
      RECT  142800.0 1719750.0 144000.0 1717800.0 ;
      RECT  142800.0 1731600.0 144000.0 1729650.0 ;
      RECT  135600.0 1720950.0 136800.0 1719750.0 ;
      RECT  138000.0 1720950.0 139200.0 1719750.0 ;
      RECT  138000.0 1720950.0 139200.0 1719750.0 ;
      RECT  135600.0 1720950.0 136800.0 1719750.0 ;
      RECT  138000.0 1720950.0 139200.0 1719750.0 ;
      RECT  140400.0 1720950.0 141600.0 1719750.0 ;
      RECT  140400.0 1720950.0 141600.0 1719750.0 ;
      RECT  138000.0 1720950.0 139200.0 1719750.0 ;
      RECT  135600.0 1729650.0 136800.0 1728450.0 ;
      RECT  138000.0 1729650.0 139200.0 1728450.0 ;
      RECT  138000.0 1729650.0 139200.0 1728450.0 ;
      RECT  135600.0 1729650.0 136800.0 1728450.0 ;
      RECT  138000.0 1729650.0 139200.0 1728450.0 ;
      RECT  140400.0 1729650.0 141600.0 1728450.0 ;
      RECT  140400.0 1729650.0 141600.0 1728450.0 ;
      RECT  138000.0 1729650.0 139200.0 1728450.0 ;
      RECT  142800.0 1720350.0 144000.0 1719150.0 ;
      RECT  142800.0 1730250.0 144000.0 1729050.0 ;
      RECT  140400.0 1727100.0 139200.0 1725900.0 ;
      RECT  137400.0 1724400.0 136200.0 1723200.0 ;
      RECT  138000.0 1720950.0 139200.0 1719750.0 ;
      RECT  140400.0 1729650.0 141600.0 1728450.0 ;
      RECT  141600.0 1724400.0 140400.0 1723200.0 ;
      RECT  136200.0 1724400.0 137400.0 1723200.0 ;
      RECT  139200.0 1727100.0 140400.0 1725900.0 ;
      RECT  140400.0 1724400.0 141600.0 1723200.0 ;
      RECT  133800.0 1718250.0 148200.0 1717350.0 ;
      RECT  133800.0 1732050.0 148200.0 1731150.0 ;
      RECT  154800.0 1719750.0 156000.0 1717800.0 ;
      RECT  154800.0 1731600.0 156000.0 1729650.0 ;
      RECT  150000.0 1730250.0 151200.0 1732050.0 ;
      RECT  150000.0 1720950.0 151200.0 1717350.0 ;
      RECT  152700.0 1730250.0 153600.0 1720950.0 ;
      RECT  150000.0 1720950.0 151200.0 1719750.0 ;
      RECT  152400.0 1720950.0 153600.0 1719750.0 ;
      RECT  152400.0 1720950.0 153600.0 1719750.0 ;
      RECT  150000.0 1720950.0 151200.0 1719750.0 ;
      RECT  150000.0 1730250.0 151200.0 1729050.0 ;
      RECT  152400.0 1730250.0 153600.0 1729050.0 ;
      RECT  152400.0 1730250.0 153600.0 1729050.0 ;
      RECT  150000.0 1730250.0 151200.0 1729050.0 ;
      RECT  154800.0 1720350.0 156000.0 1719150.0 ;
      RECT  154800.0 1730250.0 156000.0 1729050.0 ;
      RECT  150600.0 1725600.0 151800.0 1724400.0 ;
      RECT  150600.0 1725600.0 151800.0 1724400.0 ;
      RECT  153150.0 1725450.0 154050.0 1724550.0 ;
      RECT  148200.0 1718250.0 157800.0 1717350.0 ;
      RECT  148200.0 1732050.0 157800.0 1731150.0 ;
      RECT  120450.0 1724400.0 121650.0 1725600.0 ;
      RECT  122400.0 1726800.0 123600.0 1728000.0 ;
      RECT  139200.0 1725900.0 138000.0 1727100.0 ;
      RECT  130800.0 1743450.0 132000.0 1745400.0 ;
      RECT  130800.0 1731600.0 132000.0 1733550.0 ;
      RECT  126000.0 1732950.0 127200.0 1731150.0 ;
      RECT  126000.0 1742250.0 127200.0 1745850.0 ;
      RECT  128700.0 1732950.0 129600.0 1742250.0 ;
      RECT  126000.0 1742250.0 127200.0 1743450.0 ;
      RECT  128400.0 1742250.0 129600.0 1743450.0 ;
      RECT  128400.0 1742250.0 129600.0 1743450.0 ;
      RECT  126000.0 1742250.0 127200.0 1743450.0 ;
      RECT  126000.0 1732950.0 127200.0 1734150.0 ;
      RECT  128400.0 1732950.0 129600.0 1734150.0 ;
      RECT  128400.0 1732950.0 129600.0 1734150.0 ;
      RECT  126000.0 1732950.0 127200.0 1734150.0 ;
      RECT  130800.0 1742850.0 132000.0 1744050.0 ;
      RECT  130800.0 1732950.0 132000.0 1734150.0 ;
      RECT  126600.0 1737600.0 127800.0 1738800.0 ;
      RECT  126600.0 1737600.0 127800.0 1738800.0 ;
      RECT  129150.0 1737750.0 130050.0 1738650.0 ;
      RECT  124200.0 1744950.0 133800.0 1745850.0 ;
      RECT  124200.0 1731150.0 133800.0 1732050.0 ;
      RECT  135600.0 1733550.0 136800.0 1731150.0 ;
      RECT  135600.0 1742250.0 136800.0 1745850.0 ;
      RECT  140400.0 1742250.0 141600.0 1745850.0 ;
      RECT  142800.0 1743450.0 144000.0 1745400.0 ;
      RECT  142800.0 1731600.0 144000.0 1733550.0 ;
      RECT  135600.0 1742250.0 136800.0 1743450.0 ;
      RECT  138000.0 1742250.0 139200.0 1743450.0 ;
      RECT  138000.0 1742250.0 139200.0 1743450.0 ;
      RECT  135600.0 1742250.0 136800.0 1743450.0 ;
      RECT  138000.0 1742250.0 139200.0 1743450.0 ;
      RECT  140400.0 1742250.0 141600.0 1743450.0 ;
      RECT  140400.0 1742250.0 141600.0 1743450.0 ;
      RECT  138000.0 1742250.0 139200.0 1743450.0 ;
      RECT  135600.0 1733550.0 136800.0 1734750.0 ;
      RECT  138000.0 1733550.0 139200.0 1734750.0 ;
      RECT  138000.0 1733550.0 139200.0 1734750.0 ;
      RECT  135600.0 1733550.0 136800.0 1734750.0 ;
      RECT  138000.0 1733550.0 139200.0 1734750.0 ;
      RECT  140400.0 1733550.0 141600.0 1734750.0 ;
      RECT  140400.0 1733550.0 141600.0 1734750.0 ;
      RECT  138000.0 1733550.0 139200.0 1734750.0 ;
      RECT  142800.0 1742850.0 144000.0 1744050.0 ;
      RECT  142800.0 1732950.0 144000.0 1734150.0 ;
      RECT  140400.0 1736100.0 139200.0 1737300.0 ;
      RECT  137400.0 1738800.0 136200.0 1740000.0 ;
      RECT  138000.0 1742250.0 139200.0 1743450.0 ;
      RECT  140400.0 1733550.0 141600.0 1734750.0 ;
      RECT  141600.0 1738800.0 140400.0 1740000.0 ;
      RECT  136200.0 1738800.0 137400.0 1740000.0 ;
      RECT  139200.0 1736100.0 140400.0 1737300.0 ;
      RECT  140400.0 1738800.0 141600.0 1740000.0 ;
      RECT  133800.0 1744950.0 148200.0 1745850.0 ;
      RECT  133800.0 1731150.0 148200.0 1732050.0 ;
      RECT  154800.0 1743450.0 156000.0 1745400.0 ;
      RECT  154800.0 1731600.0 156000.0 1733550.0 ;
      RECT  150000.0 1732950.0 151200.0 1731150.0 ;
      RECT  150000.0 1742250.0 151200.0 1745850.0 ;
      RECT  152700.0 1732950.0 153600.0 1742250.0 ;
      RECT  150000.0 1742250.0 151200.0 1743450.0 ;
      RECT  152400.0 1742250.0 153600.0 1743450.0 ;
      RECT  152400.0 1742250.0 153600.0 1743450.0 ;
      RECT  150000.0 1742250.0 151200.0 1743450.0 ;
      RECT  150000.0 1732950.0 151200.0 1734150.0 ;
      RECT  152400.0 1732950.0 153600.0 1734150.0 ;
      RECT  152400.0 1732950.0 153600.0 1734150.0 ;
      RECT  150000.0 1732950.0 151200.0 1734150.0 ;
      RECT  154800.0 1742850.0 156000.0 1744050.0 ;
      RECT  154800.0 1732950.0 156000.0 1734150.0 ;
      RECT  150600.0 1737600.0 151800.0 1738800.0 ;
      RECT  150600.0 1737600.0 151800.0 1738800.0 ;
      RECT  153150.0 1737750.0 154050.0 1738650.0 ;
      RECT  148200.0 1744950.0 157800.0 1745850.0 ;
      RECT  148200.0 1731150.0 157800.0 1732050.0 ;
      RECT  120450.0 1737600.0 121650.0 1738800.0 ;
      RECT  122400.0 1735200.0 123600.0 1736400.0 ;
      RECT  139200.0 1736100.0 138000.0 1737300.0 ;
      RECT  130800.0 1747350.0 132000.0 1745400.0 ;
      RECT  130800.0 1759200.0 132000.0 1757250.0 ;
      RECT  126000.0 1757850.0 127200.0 1759650.0 ;
      RECT  126000.0 1748550.0 127200.0 1744950.0 ;
      RECT  128700.0 1757850.0 129600.0 1748550.0 ;
      RECT  126000.0 1748550.0 127200.0 1747350.0 ;
      RECT  128400.0 1748550.0 129600.0 1747350.0 ;
      RECT  128400.0 1748550.0 129600.0 1747350.0 ;
      RECT  126000.0 1748550.0 127200.0 1747350.0 ;
      RECT  126000.0 1757850.0 127200.0 1756650.0 ;
      RECT  128400.0 1757850.0 129600.0 1756650.0 ;
      RECT  128400.0 1757850.0 129600.0 1756650.0 ;
      RECT  126000.0 1757850.0 127200.0 1756650.0 ;
      RECT  130800.0 1747950.0 132000.0 1746750.0 ;
      RECT  130800.0 1757850.0 132000.0 1756650.0 ;
      RECT  126600.0 1753200.0 127800.0 1752000.0 ;
      RECT  126600.0 1753200.0 127800.0 1752000.0 ;
      RECT  129150.0 1753050.0 130050.0 1752150.0 ;
      RECT  124200.0 1745850.0 133800.0 1744950.0 ;
      RECT  124200.0 1759650.0 133800.0 1758750.0 ;
      RECT  135600.0 1757250.0 136800.0 1759650.0 ;
      RECT  135600.0 1748550.0 136800.0 1744950.0 ;
      RECT  140400.0 1748550.0 141600.0 1744950.0 ;
      RECT  142800.0 1747350.0 144000.0 1745400.0 ;
      RECT  142800.0 1759200.0 144000.0 1757250.0 ;
      RECT  135600.0 1748550.0 136800.0 1747350.0 ;
      RECT  138000.0 1748550.0 139200.0 1747350.0 ;
      RECT  138000.0 1748550.0 139200.0 1747350.0 ;
      RECT  135600.0 1748550.0 136800.0 1747350.0 ;
      RECT  138000.0 1748550.0 139200.0 1747350.0 ;
      RECT  140400.0 1748550.0 141600.0 1747350.0 ;
      RECT  140400.0 1748550.0 141600.0 1747350.0 ;
      RECT  138000.0 1748550.0 139200.0 1747350.0 ;
      RECT  135600.0 1757250.0 136800.0 1756050.0 ;
      RECT  138000.0 1757250.0 139200.0 1756050.0 ;
      RECT  138000.0 1757250.0 139200.0 1756050.0 ;
      RECT  135600.0 1757250.0 136800.0 1756050.0 ;
      RECT  138000.0 1757250.0 139200.0 1756050.0 ;
      RECT  140400.0 1757250.0 141600.0 1756050.0 ;
      RECT  140400.0 1757250.0 141600.0 1756050.0 ;
      RECT  138000.0 1757250.0 139200.0 1756050.0 ;
      RECT  142800.0 1747950.0 144000.0 1746750.0 ;
      RECT  142800.0 1757850.0 144000.0 1756650.0 ;
      RECT  140400.0 1754700.0 139200.0 1753500.0 ;
      RECT  137400.0 1752000.0 136200.0 1750800.0 ;
      RECT  138000.0 1748550.0 139200.0 1747350.0 ;
      RECT  140400.0 1757250.0 141600.0 1756050.0 ;
      RECT  141600.0 1752000.0 140400.0 1750800.0 ;
      RECT  136200.0 1752000.0 137400.0 1750800.0 ;
      RECT  139200.0 1754700.0 140400.0 1753500.0 ;
      RECT  140400.0 1752000.0 141600.0 1750800.0 ;
      RECT  133800.0 1745850.0 148200.0 1744950.0 ;
      RECT  133800.0 1759650.0 148200.0 1758750.0 ;
      RECT  154800.0 1747350.0 156000.0 1745400.0 ;
      RECT  154800.0 1759200.0 156000.0 1757250.0 ;
      RECT  150000.0 1757850.0 151200.0 1759650.0 ;
      RECT  150000.0 1748550.0 151200.0 1744950.0 ;
      RECT  152700.0 1757850.0 153600.0 1748550.0 ;
      RECT  150000.0 1748550.0 151200.0 1747350.0 ;
      RECT  152400.0 1748550.0 153600.0 1747350.0 ;
      RECT  152400.0 1748550.0 153600.0 1747350.0 ;
      RECT  150000.0 1748550.0 151200.0 1747350.0 ;
      RECT  150000.0 1757850.0 151200.0 1756650.0 ;
      RECT  152400.0 1757850.0 153600.0 1756650.0 ;
      RECT  152400.0 1757850.0 153600.0 1756650.0 ;
      RECT  150000.0 1757850.0 151200.0 1756650.0 ;
      RECT  154800.0 1747950.0 156000.0 1746750.0 ;
      RECT  154800.0 1757850.0 156000.0 1756650.0 ;
      RECT  150600.0 1753200.0 151800.0 1752000.0 ;
      RECT  150600.0 1753200.0 151800.0 1752000.0 ;
      RECT  153150.0 1753050.0 154050.0 1752150.0 ;
      RECT  148200.0 1745850.0 157800.0 1744950.0 ;
      RECT  148200.0 1759650.0 157800.0 1758750.0 ;
      RECT  120450.0 1752000.0 121650.0 1753200.0 ;
      RECT  122400.0 1754400.0 123600.0 1755600.0 ;
      RECT  139200.0 1753500.0 138000.0 1754700.0 ;
      RECT  130800.0 1771050.0 132000.0 1773000.0 ;
      RECT  130800.0 1759200.0 132000.0 1761150.0 ;
      RECT  126000.0 1760550.0 127200.0 1758750.0 ;
      RECT  126000.0 1769850.0 127200.0 1773450.0 ;
      RECT  128700.0 1760550.0 129600.0 1769850.0 ;
      RECT  126000.0 1769850.0 127200.0 1771050.0 ;
      RECT  128400.0 1769850.0 129600.0 1771050.0 ;
      RECT  128400.0 1769850.0 129600.0 1771050.0 ;
      RECT  126000.0 1769850.0 127200.0 1771050.0 ;
      RECT  126000.0 1760550.0 127200.0 1761750.0 ;
      RECT  128400.0 1760550.0 129600.0 1761750.0 ;
      RECT  128400.0 1760550.0 129600.0 1761750.0 ;
      RECT  126000.0 1760550.0 127200.0 1761750.0 ;
      RECT  130800.0 1770450.0 132000.0 1771650.0 ;
      RECT  130800.0 1760550.0 132000.0 1761750.0 ;
      RECT  126600.0 1765200.0 127800.0 1766400.0 ;
      RECT  126600.0 1765200.0 127800.0 1766400.0 ;
      RECT  129150.0 1765350.0 130050.0 1766250.0 ;
      RECT  124200.0 1772550.0 133800.0 1773450.0 ;
      RECT  124200.0 1758750.0 133800.0 1759650.0 ;
      RECT  135600.0 1761150.0 136800.0 1758750.0 ;
      RECT  135600.0 1769850.0 136800.0 1773450.0 ;
      RECT  140400.0 1769850.0 141600.0 1773450.0 ;
      RECT  142800.0 1771050.0 144000.0 1773000.0 ;
      RECT  142800.0 1759200.0 144000.0 1761150.0 ;
      RECT  135600.0 1769850.0 136800.0 1771050.0 ;
      RECT  138000.0 1769850.0 139200.0 1771050.0 ;
      RECT  138000.0 1769850.0 139200.0 1771050.0 ;
      RECT  135600.0 1769850.0 136800.0 1771050.0 ;
      RECT  138000.0 1769850.0 139200.0 1771050.0 ;
      RECT  140400.0 1769850.0 141600.0 1771050.0 ;
      RECT  140400.0 1769850.0 141600.0 1771050.0 ;
      RECT  138000.0 1769850.0 139200.0 1771050.0 ;
      RECT  135600.0 1761150.0 136800.0 1762350.0 ;
      RECT  138000.0 1761150.0 139200.0 1762350.0 ;
      RECT  138000.0 1761150.0 139200.0 1762350.0 ;
      RECT  135600.0 1761150.0 136800.0 1762350.0 ;
      RECT  138000.0 1761150.0 139200.0 1762350.0 ;
      RECT  140400.0 1761150.0 141600.0 1762350.0 ;
      RECT  140400.0 1761150.0 141600.0 1762350.0 ;
      RECT  138000.0 1761150.0 139200.0 1762350.0 ;
      RECT  142800.0 1770450.0 144000.0 1771650.0 ;
      RECT  142800.0 1760550.0 144000.0 1761750.0 ;
      RECT  140400.0 1763700.0 139200.0 1764900.0 ;
      RECT  137400.0 1766400.0 136200.0 1767600.0 ;
      RECT  138000.0 1769850.0 139200.0 1771050.0 ;
      RECT  140400.0 1761150.0 141600.0 1762350.0 ;
      RECT  141600.0 1766400.0 140400.0 1767600.0 ;
      RECT  136200.0 1766400.0 137400.0 1767600.0 ;
      RECT  139200.0 1763700.0 140400.0 1764900.0 ;
      RECT  140400.0 1766400.0 141600.0 1767600.0 ;
      RECT  133800.0 1772550.0 148200.0 1773450.0 ;
      RECT  133800.0 1758750.0 148200.0 1759650.0 ;
      RECT  154800.0 1771050.0 156000.0 1773000.0 ;
      RECT  154800.0 1759200.0 156000.0 1761150.0 ;
      RECT  150000.0 1760550.0 151200.0 1758750.0 ;
      RECT  150000.0 1769850.0 151200.0 1773450.0 ;
      RECT  152700.0 1760550.0 153600.0 1769850.0 ;
      RECT  150000.0 1769850.0 151200.0 1771050.0 ;
      RECT  152400.0 1769850.0 153600.0 1771050.0 ;
      RECT  152400.0 1769850.0 153600.0 1771050.0 ;
      RECT  150000.0 1769850.0 151200.0 1771050.0 ;
      RECT  150000.0 1760550.0 151200.0 1761750.0 ;
      RECT  152400.0 1760550.0 153600.0 1761750.0 ;
      RECT  152400.0 1760550.0 153600.0 1761750.0 ;
      RECT  150000.0 1760550.0 151200.0 1761750.0 ;
      RECT  154800.0 1770450.0 156000.0 1771650.0 ;
      RECT  154800.0 1760550.0 156000.0 1761750.0 ;
      RECT  150600.0 1765200.0 151800.0 1766400.0 ;
      RECT  150600.0 1765200.0 151800.0 1766400.0 ;
      RECT  153150.0 1765350.0 154050.0 1766250.0 ;
      RECT  148200.0 1772550.0 157800.0 1773450.0 ;
      RECT  148200.0 1758750.0 157800.0 1759650.0 ;
      RECT  120450.0 1765200.0 121650.0 1766400.0 ;
      RECT  122400.0 1762800.0 123600.0 1764000.0 ;
      RECT  139200.0 1763700.0 138000.0 1764900.0 ;
      RECT  130800.0 1774950.0 132000.0 1773000.0 ;
      RECT  130800.0 1786800.0 132000.0 1784850.0 ;
      RECT  126000.0 1785450.0 127200.0 1787250.0 ;
      RECT  126000.0 1776150.0 127200.0 1772550.0 ;
      RECT  128700.0 1785450.0 129600.0 1776150.0 ;
      RECT  126000.0 1776150.0 127200.0 1774950.0 ;
      RECT  128400.0 1776150.0 129600.0 1774950.0 ;
      RECT  128400.0 1776150.0 129600.0 1774950.0 ;
      RECT  126000.0 1776150.0 127200.0 1774950.0 ;
      RECT  126000.0 1785450.0 127200.0 1784250.0 ;
      RECT  128400.0 1785450.0 129600.0 1784250.0 ;
      RECT  128400.0 1785450.0 129600.0 1784250.0 ;
      RECT  126000.0 1785450.0 127200.0 1784250.0 ;
      RECT  130800.0 1775550.0 132000.0 1774350.0 ;
      RECT  130800.0 1785450.0 132000.0 1784250.0 ;
      RECT  126600.0 1780800.0 127800.0 1779600.0 ;
      RECT  126600.0 1780800.0 127800.0 1779600.0 ;
      RECT  129150.0 1780650.0 130050.0 1779750.0 ;
      RECT  124200.0 1773450.0 133800.0 1772550.0 ;
      RECT  124200.0 1787250.0 133800.0 1786350.0 ;
      RECT  135600.0 1784850.0 136800.0 1787250.0 ;
      RECT  135600.0 1776150.0 136800.0 1772550.0 ;
      RECT  140400.0 1776150.0 141600.0 1772550.0 ;
      RECT  142800.0 1774950.0 144000.0 1773000.0 ;
      RECT  142800.0 1786800.0 144000.0 1784850.0 ;
      RECT  135600.0 1776150.0 136800.0 1774950.0 ;
      RECT  138000.0 1776150.0 139200.0 1774950.0 ;
      RECT  138000.0 1776150.0 139200.0 1774950.0 ;
      RECT  135600.0 1776150.0 136800.0 1774950.0 ;
      RECT  138000.0 1776150.0 139200.0 1774950.0 ;
      RECT  140400.0 1776150.0 141600.0 1774950.0 ;
      RECT  140400.0 1776150.0 141600.0 1774950.0 ;
      RECT  138000.0 1776150.0 139200.0 1774950.0 ;
      RECT  135600.0 1784850.0 136800.0 1783650.0 ;
      RECT  138000.0 1784850.0 139200.0 1783650.0 ;
      RECT  138000.0 1784850.0 139200.0 1783650.0 ;
      RECT  135600.0 1784850.0 136800.0 1783650.0 ;
      RECT  138000.0 1784850.0 139200.0 1783650.0 ;
      RECT  140400.0 1784850.0 141600.0 1783650.0 ;
      RECT  140400.0 1784850.0 141600.0 1783650.0 ;
      RECT  138000.0 1784850.0 139200.0 1783650.0 ;
      RECT  142800.0 1775550.0 144000.0 1774350.0 ;
      RECT  142800.0 1785450.0 144000.0 1784250.0 ;
      RECT  140400.0 1782300.0 139200.0 1781100.0 ;
      RECT  137400.0 1779600.0 136200.0 1778400.0 ;
      RECT  138000.0 1776150.0 139200.0 1774950.0 ;
      RECT  140400.0 1784850.0 141600.0 1783650.0 ;
      RECT  141600.0 1779600.0 140400.0 1778400.0 ;
      RECT  136200.0 1779600.0 137400.0 1778400.0 ;
      RECT  139200.0 1782300.0 140400.0 1781100.0 ;
      RECT  140400.0 1779600.0 141600.0 1778400.0 ;
      RECT  133800.0 1773450.0 148200.0 1772550.0 ;
      RECT  133800.0 1787250.0 148200.0 1786350.0 ;
      RECT  154800.0 1774950.0 156000.0 1773000.0 ;
      RECT  154800.0 1786800.0 156000.0 1784850.0 ;
      RECT  150000.0 1785450.0 151200.0 1787250.0 ;
      RECT  150000.0 1776150.0 151200.0 1772550.0 ;
      RECT  152700.0 1785450.0 153600.0 1776150.0 ;
      RECT  150000.0 1776150.0 151200.0 1774950.0 ;
      RECT  152400.0 1776150.0 153600.0 1774950.0 ;
      RECT  152400.0 1776150.0 153600.0 1774950.0 ;
      RECT  150000.0 1776150.0 151200.0 1774950.0 ;
      RECT  150000.0 1785450.0 151200.0 1784250.0 ;
      RECT  152400.0 1785450.0 153600.0 1784250.0 ;
      RECT  152400.0 1785450.0 153600.0 1784250.0 ;
      RECT  150000.0 1785450.0 151200.0 1784250.0 ;
      RECT  154800.0 1775550.0 156000.0 1774350.0 ;
      RECT  154800.0 1785450.0 156000.0 1784250.0 ;
      RECT  150600.0 1780800.0 151800.0 1779600.0 ;
      RECT  150600.0 1780800.0 151800.0 1779600.0 ;
      RECT  153150.0 1780650.0 154050.0 1779750.0 ;
      RECT  148200.0 1773450.0 157800.0 1772550.0 ;
      RECT  148200.0 1787250.0 157800.0 1786350.0 ;
      RECT  120450.0 1779600.0 121650.0 1780800.0 ;
      RECT  122400.0 1782000.0 123600.0 1783200.0 ;
      RECT  139200.0 1781100.0 138000.0 1782300.0 ;
      RECT  130800.0 1798650.0 132000.0 1800600.0 ;
      RECT  130800.0 1786800.0 132000.0 1788750.0 ;
      RECT  126000.0 1788150.0 127200.0 1786350.0 ;
      RECT  126000.0 1797450.0 127200.0 1801050.0 ;
      RECT  128700.0 1788150.0 129600.0 1797450.0 ;
      RECT  126000.0 1797450.0 127200.0 1798650.0 ;
      RECT  128400.0 1797450.0 129600.0 1798650.0 ;
      RECT  128400.0 1797450.0 129600.0 1798650.0 ;
      RECT  126000.0 1797450.0 127200.0 1798650.0 ;
      RECT  126000.0 1788150.0 127200.0 1789350.0 ;
      RECT  128400.0 1788150.0 129600.0 1789350.0 ;
      RECT  128400.0 1788150.0 129600.0 1789350.0 ;
      RECT  126000.0 1788150.0 127200.0 1789350.0 ;
      RECT  130800.0 1798050.0 132000.0 1799250.0 ;
      RECT  130800.0 1788150.0 132000.0 1789350.0 ;
      RECT  126600.0 1792800.0 127800.0 1794000.0 ;
      RECT  126600.0 1792800.0 127800.0 1794000.0 ;
      RECT  129150.0 1792950.0 130050.0 1793850.0 ;
      RECT  124200.0 1800150.0 133800.0 1801050.0 ;
      RECT  124200.0 1786350.0 133800.0 1787250.0 ;
      RECT  135600.0 1788750.0 136800.0 1786350.0 ;
      RECT  135600.0 1797450.0 136800.0 1801050.0 ;
      RECT  140400.0 1797450.0 141600.0 1801050.0 ;
      RECT  142800.0 1798650.0 144000.0 1800600.0 ;
      RECT  142800.0 1786800.0 144000.0 1788750.0 ;
      RECT  135600.0 1797450.0 136800.0 1798650.0 ;
      RECT  138000.0 1797450.0 139200.0 1798650.0 ;
      RECT  138000.0 1797450.0 139200.0 1798650.0 ;
      RECT  135600.0 1797450.0 136800.0 1798650.0 ;
      RECT  138000.0 1797450.0 139200.0 1798650.0 ;
      RECT  140400.0 1797450.0 141600.0 1798650.0 ;
      RECT  140400.0 1797450.0 141600.0 1798650.0 ;
      RECT  138000.0 1797450.0 139200.0 1798650.0 ;
      RECT  135600.0 1788750.0 136800.0 1789950.0 ;
      RECT  138000.0 1788750.0 139200.0 1789950.0 ;
      RECT  138000.0 1788750.0 139200.0 1789950.0 ;
      RECT  135600.0 1788750.0 136800.0 1789950.0 ;
      RECT  138000.0 1788750.0 139200.0 1789950.0 ;
      RECT  140400.0 1788750.0 141600.0 1789950.0 ;
      RECT  140400.0 1788750.0 141600.0 1789950.0 ;
      RECT  138000.0 1788750.0 139200.0 1789950.0 ;
      RECT  142800.0 1798050.0 144000.0 1799250.0 ;
      RECT  142800.0 1788150.0 144000.0 1789350.0 ;
      RECT  140400.0 1791300.0 139200.0 1792500.0 ;
      RECT  137400.0 1794000.0 136200.0 1795200.0 ;
      RECT  138000.0 1797450.0 139200.0 1798650.0 ;
      RECT  140400.0 1788750.0 141600.0 1789950.0 ;
      RECT  141600.0 1794000.0 140400.0 1795200.0 ;
      RECT  136200.0 1794000.0 137400.0 1795200.0 ;
      RECT  139200.0 1791300.0 140400.0 1792500.0 ;
      RECT  140400.0 1794000.0 141600.0 1795200.0 ;
      RECT  133800.0 1800150.0 148200.0 1801050.0 ;
      RECT  133800.0 1786350.0 148200.0 1787250.0 ;
      RECT  154800.0 1798650.0 156000.0 1800600.0 ;
      RECT  154800.0 1786800.0 156000.0 1788750.0 ;
      RECT  150000.0 1788150.0 151200.0 1786350.0 ;
      RECT  150000.0 1797450.0 151200.0 1801050.0 ;
      RECT  152700.0 1788150.0 153600.0 1797450.0 ;
      RECT  150000.0 1797450.0 151200.0 1798650.0 ;
      RECT  152400.0 1797450.0 153600.0 1798650.0 ;
      RECT  152400.0 1797450.0 153600.0 1798650.0 ;
      RECT  150000.0 1797450.0 151200.0 1798650.0 ;
      RECT  150000.0 1788150.0 151200.0 1789350.0 ;
      RECT  152400.0 1788150.0 153600.0 1789350.0 ;
      RECT  152400.0 1788150.0 153600.0 1789350.0 ;
      RECT  150000.0 1788150.0 151200.0 1789350.0 ;
      RECT  154800.0 1798050.0 156000.0 1799250.0 ;
      RECT  154800.0 1788150.0 156000.0 1789350.0 ;
      RECT  150600.0 1792800.0 151800.0 1794000.0 ;
      RECT  150600.0 1792800.0 151800.0 1794000.0 ;
      RECT  153150.0 1792950.0 154050.0 1793850.0 ;
      RECT  148200.0 1800150.0 157800.0 1801050.0 ;
      RECT  148200.0 1786350.0 157800.0 1787250.0 ;
      RECT  120450.0 1792800.0 121650.0 1794000.0 ;
      RECT  122400.0 1790400.0 123600.0 1791600.0 ;
      RECT  139200.0 1791300.0 138000.0 1792500.0 ;
      RECT  130800.0 1802550.0 132000.0 1800600.0 ;
      RECT  130800.0 1814400.0 132000.0 1812450.0 ;
      RECT  126000.0 1813050.0 127200.0 1814850.0 ;
      RECT  126000.0 1803750.0 127200.0 1800150.0 ;
      RECT  128700.0 1813050.0 129600.0 1803750.0 ;
      RECT  126000.0 1803750.0 127200.0 1802550.0 ;
      RECT  128400.0 1803750.0 129600.0 1802550.0 ;
      RECT  128400.0 1803750.0 129600.0 1802550.0 ;
      RECT  126000.0 1803750.0 127200.0 1802550.0 ;
      RECT  126000.0 1813050.0 127200.0 1811850.0 ;
      RECT  128400.0 1813050.0 129600.0 1811850.0 ;
      RECT  128400.0 1813050.0 129600.0 1811850.0 ;
      RECT  126000.0 1813050.0 127200.0 1811850.0 ;
      RECT  130800.0 1803150.0 132000.0 1801950.0 ;
      RECT  130800.0 1813050.0 132000.0 1811850.0 ;
      RECT  126600.0 1808400.0 127800.0 1807200.0 ;
      RECT  126600.0 1808400.0 127800.0 1807200.0 ;
      RECT  129150.0 1808250.0 130050.0 1807350.0 ;
      RECT  124200.0 1801050.0 133800.0 1800150.0 ;
      RECT  124200.0 1814850.0 133800.0 1813950.0 ;
      RECT  135600.0 1812450.0 136800.0 1814850.0 ;
      RECT  135600.0 1803750.0 136800.0 1800150.0 ;
      RECT  140400.0 1803750.0 141600.0 1800150.0 ;
      RECT  142800.0 1802550.0 144000.0 1800600.0 ;
      RECT  142800.0 1814400.0 144000.0 1812450.0 ;
      RECT  135600.0 1803750.0 136800.0 1802550.0 ;
      RECT  138000.0 1803750.0 139200.0 1802550.0 ;
      RECT  138000.0 1803750.0 139200.0 1802550.0 ;
      RECT  135600.0 1803750.0 136800.0 1802550.0 ;
      RECT  138000.0 1803750.0 139200.0 1802550.0 ;
      RECT  140400.0 1803750.0 141600.0 1802550.0 ;
      RECT  140400.0 1803750.0 141600.0 1802550.0 ;
      RECT  138000.0 1803750.0 139200.0 1802550.0 ;
      RECT  135600.0 1812450.0 136800.0 1811250.0 ;
      RECT  138000.0 1812450.0 139200.0 1811250.0 ;
      RECT  138000.0 1812450.0 139200.0 1811250.0 ;
      RECT  135600.0 1812450.0 136800.0 1811250.0 ;
      RECT  138000.0 1812450.0 139200.0 1811250.0 ;
      RECT  140400.0 1812450.0 141600.0 1811250.0 ;
      RECT  140400.0 1812450.0 141600.0 1811250.0 ;
      RECT  138000.0 1812450.0 139200.0 1811250.0 ;
      RECT  142800.0 1803150.0 144000.0 1801950.0 ;
      RECT  142800.0 1813050.0 144000.0 1811850.0 ;
      RECT  140400.0 1809900.0 139200.0 1808700.0 ;
      RECT  137400.0 1807200.0 136200.0 1806000.0 ;
      RECT  138000.0 1803750.0 139200.0 1802550.0 ;
      RECT  140400.0 1812450.0 141600.0 1811250.0 ;
      RECT  141600.0 1807200.0 140400.0 1806000.0 ;
      RECT  136200.0 1807200.0 137400.0 1806000.0 ;
      RECT  139200.0 1809900.0 140400.0 1808700.0 ;
      RECT  140400.0 1807200.0 141600.0 1806000.0 ;
      RECT  133800.0 1801050.0 148200.0 1800150.0 ;
      RECT  133800.0 1814850.0 148200.0 1813950.0 ;
      RECT  154800.0 1802550.0 156000.0 1800600.0 ;
      RECT  154800.0 1814400.0 156000.0 1812450.0 ;
      RECT  150000.0 1813050.0 151200.0 1814850.0 ;
      RECT  150000.0 1803750.0 151200.0 1800150.0 ;
      RECT  152700.0 1813050.0 153600.0 1803750.0 ;
      RECT  150000.0 1803750.0 151200.0 1802550.0 ;
      RECT  152400.0 1803750.0 153600.0 1802550.0 ;
      RECT  152400.0 1803750.0 153600.0 1802550.0 ;
      RECT  150000.0 1803750.0 151200.0 1802550.0 ;
      RECT  150000.0 1813050.0 151200.0 1811850.0 ;
      RECT  152400.0 1813050.0 153600.0 1811850.0 ;
      RECT  152400.0 1813050.0 153600.0 1811850.0 ;
      RECT  150000.0 1813050.0 151200.0 1811850.0 ;
      RECT  154800.0 1803150.0 156000.0 1801950.0 ;
      RECT  154800.0 1813050.0 156000.0 1811850.0 ;
      RECT  150600.0 1808400.0 151800.0 1807200.0 ;
      RECT  150600.0 1808400.0 151800.0 1807200.0 ;
      RECT  153150.0 1808250.0 154050.0 1807350.0 ;
      RECT  148200.0 1801050.0 157800.0 1800150.0 ;
      RECT  148200.0 1814850.0 157800.0 1813950.0 ;
      RECT  120450.0 1807200.0 121650.0 1808400.0 ;
      RECT  122400.0 1809600.0 123600.0 1810800.0 ;
      RECT  139200.0 1808700.0 138000.0 1809900.0 ;
      RECT  130800.0 1826250.0 132000.0 1828200.0 ;
      RECT  130800.0 1814400.0 132000.0 1816350.0 ;
      RECT  126000.0 1815750.0 127200.0 1813950.0 ;
      RECT  126000.0 1825050.0 127200.0 1828650.0 ;
      RECT  128700.0 1815750.0 129600.0 1825050.0 ;
      RECT  126000.0 1825050.0 127200.0 1826250.0 ;
      RECT  128400.0 1825050.0 129600.0 1826250.0 ;
      RECT  128400.0 1825050.0 129600.0 1826250.0 ;
      RECT  126000.0 1825050.0 127200.0 1826250.0 ;
      RECT  126000.0 1815750.0 127200.0 1816950.0 ;
      RECT  128400.0 1815750.0 129600.0 1816950.0 ;
      RECT  128400.0 1815750.0 129600.0 1816950.0 ;
      RECT  126000.0 1815750.0 127200.0 1816950.0 ;
      RECT  130800.0 1825650.0 132000.0 1826850.0 ;
      RECT  130800.0 1815750.0 132000.0 1816950.0 ;
      RECT  126600.0 1820400.0 127800.0 1821600.0 ;
      RECT  126600.0 1820400.0 127800.0 1821600.0 ;
      RECT  129150.0 1820550.0 130050.0 1821450.0 ;
      RECT  124200.0 1827750.0 133800.0 1828650.0 ;
      RECT  124200.0 1813950.0 133800.0 1814850.0 ;
      RECT  135600.0 1816350.0 136800.0 1813950.0 ;
      RECT  135600.0 1825050.0 136800.0 1828650.0 ;
      RECT  140400.0 1825050.0 141600.0 1828650.0 ;
      RECT  142800.0 1826250.0 144000.0 1828200.0 ;
      RECT  142800.0 1814400.0 144000.0 1816350.0 ;
      RECT  135600.0 1825050.0 136800.0 1826250.0 ;
      RECT  138000.0 1825050.0 139200.0 1826250.0 ;
      RECT  138000.0 1825050.0 139200.0 1826250.0 ;
      RECT  135600.0 1825050.0 136800.0 1826250.0 ;
      RECT  138000.0 1825050.0 139200.0 1826250.0 ;
      RECT  140400.0 1825050.0 141600.0 1826250.0 ;
      RECT  140400.0 1825050.0 141600.0 1826250.0 ;
      RECT  138000.0 1825050.0 139200.0 1826250.0 ;
      RECT  135600.0 1816350.0 136800.0 1817550.0 ;
      RECT  138000.0 1816350.0 139200.0 1817550.0 ;
      RECT  138000.0 1816350.0 139200.0 1817550.0 ;
      RECT  135600.0 1816350.0 136800.0 1817550.0 ;
      RECT  138000.0 1816350.0 139200.0 1817550.0 ;
      RECT  140400.0 1816350.0 141600.0 1817550.0 ;
      RECT  140400.0 1816350.0 141600.0 1817550.0 ;
      RECT  138000.0 1816350.0 139200.0 1817550.0 ;
      RECT  142800.0 1825650.0 144000.0 1826850.0 ;
      RECT  142800.0 1815750.0 144000.0 1816950.0 ;
      RECT  140400.0 1818900.0 139200.0 1820100.0 ;
      RECT  137400.0 1821600.0 136200.0 1822800.0 ;
      RECT  138000.0 1825050.0 139200.0 1826250.0 ;
      RECT  140400.0 1816350.0 141600.0 1817550.0 ;
      RECT  141600.0 1821600.0 140400.0 1822800.0 ;
      RECT  136200.0 1821600.0 137400.0 1822800.0 ;
      RECT  139200.0 1818900.0 140400.0 1820100.0 ;
      RECT  140400.0 1821600.0 141600.0 1822800.0 ;
      RECT  133800.0 1827750.0 148200.0 1828650.0 ;
      RECT  133800.0 1813950.0 148200.0 1814850.0 ;
      RECT  154800.0 1826250.0 156000.0 1828200.0 ;
      RECT  154800.0 1814400.0 156000.0 1816350.0 ;
      RECT  150000.0 1815750.0 151200.0 1813950.0 ;
      RECT  150000.0 1825050.0 151200.0 1828650.0 ;
      RECT  152700.0 1815750.0 153600.0 1825050.0 ;
      RECT  150000.0 1825050.0 151200.0 1826250.0 ;
      RECT  152400.0 1825050.0 153600.0 1826250.0 ;
      RECT  152400.0 1825050.0 153600.0 1826250.0 ;
      RECT  150000.0 1825050.0 151200.0 1826250.0 ;
      RECT  150000.0 1815750.0 151200.0 1816950.0 ;
      RECT  152400.0 1815750.0 153600.0 1816950.0 ;
      RECT  152400.0 1815750.0 153600.0 1816950.0 ;
      RECT  150000.0 1815750.0 151200.0 1816950.0 ;
      RECT  154800.0 1825650.0 156000.0 1826850.0 ;
      RECT  154800.0 1815750.0 156000.0 1816950.0 ;
      RECT  150600.0 1820400.0 151800.0 1821600.0 ;
      RECT  150600.0 1820400.0 151800.0 1821600.0 ;
      RECT  153150.0 1820550.0 154050.0 1821450.0 ;
      RECT  148200.0 1827750.0 157800.0 1828650.0 ;
      RECT  148200.0 1813950.0 157800.0 1814850.0 ;
      RECT  120450.0 1820400.0 121650.0 1821600.0 ;
      RECT  122400.0 1818000.0 123600.0 1819200.0 ;
      RECT  139200.0 1818900.0 138000.0 1820100.0 ;
      RECT  130800.0 1830150.0 132000.0 1828200.0 ;
      RECT  130800.0 1842000.0 132000.0 1840050.0 ;
      RECT  126000.0 1840650.0 127200.0 1842450.0 ;
      RECT  126000.0 1831350.0 127200.0 1827750.0 ;
      RECT  128700.0 1840650.0 129600.0 1831350.0 ;
      RECT  126000.0 1831350.0 127200.0 1830150.0 ;
      RECT  128400.0 1831350.0 129600.0 1830150.0 ;
      RECT  128400.0 1831350.0 129600.0 1830150.0 ;
      RECT  126000.0 1831350.0 127200.0 1830150.0 ;
      RECT  126000.0 1840650.0 127200.0 1839450.0 ;
      RECT  128400.0 1840650.0 129600.0 1839450.0 ;
      RECT  128400.0 1840650.0 129600.0 1839450.0 ;
      RECT  126000.0 1840650.0 127200.0 1839450.0 ;
      RECT  130800.0 1830750.0 132000.0 1829550.0 ;
      RECT  130800.0 1840650.0 132000.0 1839450.0 ;
      RECT  126600.0 1836000.0 127800.0 1834800.0 ;
      RECT  126600.0 1836000.0 127800.0 1834800.0 ;
      RECT  129150.0 1835850.0 130050.0 1834950.0 ;
      RECT  124200.0 1828650.0 133800.0 1827750.0 ;
      RECT  124200.0 1842450.0 133800.0 1841550.0 ;
      RECT  135600.0 1840050.0 136800.0 1842450.0 ;
      RECT  135600.0 1831350.0 136800.0 1827750.0 ;
      RECT  140400.0 1831350.0 141600.0 1827750.0 ;
      RECT  142800.0 1830150.0 144000.0 1828200.0 ;
      RECT  142800.0 1842000.0 144000.0 1840050.0 ;
      RECT  135600.0 1831350.0 136800.0 1830150.0 ;
      RECT  138000.0 1831350.0 139200.0 1830150.0 ;
      RECT  138000.0 1831350.0 139200.0 1830150.0 ;
      RECT  135600.0 1831350.0 136800.0 1830150.0 ;
      RECT  138000.0 1831350.0 139200.0 1830150.0 ;
      RECT  140400.0 1831350.0 141600.0 1830150.0 ;
      RECT  140400.0 1831350.0 141600.0 1830150.0 ;
      RECT  138000.0 1831350.0 139200.0 1830150.0 ;
      RECT  135600.0 1840050.0 136800.0 1838850.0 ;
      RECT  138000.0 1840050.0 139200.0 1838850.0 ;
      RECT  138000.0 1840050.0 139200.0 1838850.0 ;
      RECT  135600.0 1840050.0 136800.0 1838850.0 ;
      RECT  138000.0 1840050.0 139200.0 1838850.0 ;
      RECT  140400.0 1840050.0 141600.0 1838850.0 ;
      RECT  140400.0 1840050.0 141600.0 1838850.0 ;
      RECT  138000.0 1840050.0 139200.0 1838850.0 ;
      RECT  142800.0 1830750.0 144000.0 1829550.0 ;
      RECT  142800.0 1840650.0 144000.0 1839450.0 ;
      RECT  140400.0 1837500.0 139200.0 1836300.0 ;
      RECT  137400.0 1834800.0 136200.0 1833600.0 ;
      RECT  138000.0 1831350.0 139200.0 1830150.0 ;
      RECT  140400.0 1840050.0 141600.0 1838850.0 ;
      RECT  141600.0 1834800.0 140400.0 1833600.0 ;
      RECT  136200.0 1834800.0 137400.0 1833600.0 ;
      RECT  139200.0 1837500.0 140400.0 1836300.0 ;
      RECT  140400.0 1834800.0 141600.0 1833600.0 ;
      RECT  133800.0 1828650.0 148200.0 1827750.0 ;
      RECT  133800.0 1842450.0 148200.0 1841550.0 ;
      RECT  154800.0 1830150.0 156000.0 1828200.0 ;
      RECT  154800.0 1842000.0 156000.0 1840050.0 ;
      RECT  150000.0 1840650.0 151200.0 1842450.0 ;
      RECT  150000.0 1831350.0 151200.0 1827750.0 ;
      RECT  152700.0 1840650.0 153600.0 1831350.0 ;
      RECT  150000.0 1831350.0 151200.0 1830150.0 ;
      RECT  152400.0 1831350.0 153600.0 1830150.0 ;
      RECT  152400.0 1831350.0 153600.0 1830150.0 ;
      RECT  150000.0 1831350.0 151200.0 1830150.0 ;
      RECT  150000.0 1840650.0 151200.0 1839450.0 ;
      RECT  152400.0 1840650.0 153600.0 1839450.0 ;
      RECT  152400.0 1840650.0 153600.0 1839450.0 ;
      RECT  150000.0 1840650.0 151200.0 1839450.0 ;
      RECT  154800.0 1830750.0 156000.0 1829550.0 ;
      RECT  154800.0 1840650.0 156000.0 1839450.0 ;
      RECT  150600.0 1836000.0 151800.0 1834800.0 ;
      RECT  150600.0 1836000.0 151800.0 1834800.0 ;
      RECT  153150.0 1835850.0 154050.0 1834950.0 ;
      RECT  148200.0 1828650.0 157800.0 1827750.0 ;
      RECT  148200.0 1842450.0 157800.0 1841550.0 ;
      RECT  120450.0 1834800.0 121650.0 1836000.0 ;
      RECT  122400.0 1837200.0 123600.0 1838400.0 ;
      RECT  139200.0 1836300.0 138000.0 1837500.0 ;
      RECT  130800.0 1853850.0 132000.0 1855800.0 ;
      RECT  130800.0 1842000.0 132000.0 1843950.0 ;
      RECT  126000.0 1843350.0 127200.0 1841550.0 ;
      RECT  126000.0 1852650.0 127200.0 1856250.0 ;
      RECT  128700.0 1843350.0 129600.0 1852650.0 ;
      RECT  126000.0 1852650.0 127200.0 1853850.0 ;
      RECT  128400.0 1852650.0 129600.0 1853850.0 ;
      RECT  128400.0 1852650.0 129600.0 1853850.0 ;
      RECT  126000.0 1852650.0 127200.0 1853850.0 ;
      RECT  126000.0 1843350.0 127200.0 1844550.0 ;
      RECT  128400.0 1843350.0 129600.0 1844550.0 ;
      RECT  128400.0 1843350.0 129600.0 1844550.0 ;
      RECT  126000.0 1843350.0 127200.0 1844550.0 ;
      RECT  130800.0 1853250.0 132000.0 1854450.0 ;
      RECT  130800.0 1843350.0 132000.0 1844550.0 ;
      RECT  126600.0 1848000.0 127800.0 1849200.0 ;
      RECT  126600.0 1848000.0 127800.0 1849200.0 ;
      RECT  129150.0 1848150.0 130050.0 1849050.0 ;
      RECT  124200.0 1855350.0 133800.0 1856250.0 ;
      RECT  124200.0 1841550.0 133800.0 1842450.0 ;
      RECT  135600.0 1843950.0 136800.0 1841550.0 ;
      RECT  135600.0 1852650.0 136800.0 1856250.0 ;
      RECT  140400.0 1852650.0 141600.0 1856250.0 ;
      RECT  142800.0 1853850.0 144000.0 1855800.0 ;
      RECT  142800.0 1842000.0 144000.0 1843950.0 ;
      RECT  135600.0 1852650.0 136800.0 1853850.0 ;
      RECT  138000.0 1852650.0 139200.0 1853850.0 ;
      RECT  138000.0 1852650.0 139200.0 1853850.0 ;
      RECT  135600.0 1852650.0 136800.0 1853850.0 ;
      RECT  138000.0 1852650.0 139200.0 1853850.0 ;
      RECT  140400.0 1852650.0 141600.0 1853850.0 ;
      RECT  140400.0 1852650.0 141600.0 1853850.0 ;
      RECT  138000.0 1852650.0 139200.0 1853850.0 ;
      RECT  135600.0 1843950.0 136800.0 1845150.0 ;
      RECT  138000.0 1843950.0 139200.0 1845150.0 ;
      RECT  138000.0 1843950.0 139200.0 1845150.0 ;
      RECT  135600.0 1843950.0 136800.0 1845150.0 ;
      RECT  138000.0 1843950.0 139200.0 1845150.0 ;
      RECT  140400.0 1843950.0 141600.0 1845150.0 ;
      RECT  140400.0 1843950.0 141600.0 1845150.0 ;
      RECT  138000.0 1843950.0 139200.0 1845150.0 ;
      RECT  142800.0 1853250.0 144000.0 1854450.0 ;
      RECT  142800.0 1843350.0 144000.0 1844550.0 ;
      RECT  140400.0 1846500.0 139200.0 1847700.0 ;
      RECT  137400.0 1849200.0 136200.0 1850400.0 ;
      RECT  138000.0 1852650.0 139200.0 1853850.0 ;
      RECT  140400.0 1843950.0 141600.0 1845150.0 ;
      RECT  141600.0 1849200.0 140400.0 1850400.0 ;
      RECT  136200.0 1849200.0 137400.0 1850400.0 ;
      RECT  139200.0 1846500.0 140400.0 1847700.0 ;
      RECT  140400.0 1849200.0 141600.0 1850400.0 ;
      RECT  133800.0 1855350.0 148200.0 1856250.0 ;
      RECT  133800.0 1841550.0 148200.0 1842450.0 ;
      RECT  154800.0 1853850.0 156000.0 1855800.0 ;
      RECT  154800.0 1842000.0 156000.0 1843950.0 ;
      RECT  150000.0 1843350.0 151200.0 1841550.0 ;
      RECT  150000.0 1852650.0 151200.0 1856250.0 ;
      RECT  152700.0 1843350.0 153600.0 1852650.0 ;
      RECT  150000.0 1852650.0 151200.0 1853850.0 ;
      RECT  152400.0 1852650.0 153600.0 1853850.0 ;
      RECT  152400.0 1852650.0 153600.0 1853850.0 ;
      RECT  150000.0 1852650.0 151200.0 1853850.0 ;
      RECT  150000.0 1843350.0 151200.0 1844550.0 ;
      RECT  152400.0 1843350.0 153600.0 1844550.0 ;
      RECT  152400.0 1843350.0 153600.0 1844550.0 ;
      RECT  150000.0 1843350.0 151200.0 1844550.0 ;
      RECT  154800.0 1853250.0 156000.0 1854450.0 ;
      RECT  154800.0 1843350.0 156000.0 1844550.0 ;
      RECT  150600.0 1848000.0 151800.0 1849200.0 ;
      RECT  150600.0 1848000.0 151800.0 1849200.0 ;
      RECT  153150.0 1848150.0 154050.0 1849050.0 ;
      RECT  148200.0 1855350.0 157800.0 1856250.0 ;
      RECT  148200.0 1841550.0 157800.0 1842450.0 ;
      RECT  120450.0 1848000.0 121650.0 1849200.0 ;
      RECT  122400.0 1845600.0 123600.0 1846800.0 ;
      RECT  139200.0 1846500.0 138000.0 1847700.0 ;
      RECT  130800.0 1857750.0 132000.0 1855800.0 ;
      RECT  130800.0 1869600.0 132000.0 1867650.0 ;
      RECT  126000.0 1868250.0 127200.0 1870050.0 ;
      RECT  126000.0 1858950.0 127200.0 1855350.0 ;
      RECT  128700.0 1868250.0 129600.0 1858950.0 ;
      RECT  126000.0 1858950.0 127200.0 1857750.0 ;
      RECT  128400.0 1858950.0 129600.0 1857750.0 ;
      RECT  128400.0 1858950.0 129600.0 1857750.0 ;
      RECT  126000.0 1858950.0 127200.0 1857750.0 ;
      RECT  126000.0 1868250.0 127200.0 1867050.0 ;
      RECT  128400.0 1868250.0 129600.0 1867050.0 ;
      RECT  128400.0 1868250.0 129600.0 1867050.0 ;
      RECT  126000.0 1868250.0 127200.0 1867050.0 ;
      RECT  130800.0 1858350.0 132000.0 1857150.0 ;
      RECT  130800.0 1868250.0 132000.0 1867050.0 ;
      RECT  126600.0 1863600.0 127800.0 1862400.0 ;
      RECT  126600.0 1863600.0 127800.0 1862400.0 ;
      RECT  129150.0 1863450.0 130050.0 1862550.0 ;
      RECT  124200.0 1856250.0 133800.0 1855350.0 ;
      RECT  124200.0 1870050.0 133800.0 1869150.0 ;
      RECT  135600.0 1867650.0 136800.0 1870050.0 ;
      RECT  135600.0 1858950.0 136800.0 1855350.0 ;
      RECT  140400.0 1858950.0 141600.0 1855350.0 ;
      RECT  142800.0 1857750.0 144000.0 1855800.0 ;
      RECT  142800.0 1869600.0 144000.0 1867650.0 ;
      RECT  135600.0 1858950.0 136800.0 1857750.0 ;
      RECT  138000.0 1858950.0 139200.0 1857750.0 ;
      RECT  138000.0 1858950.0 139200.0 1857750.0 ;
      RECT  135600.0 1858950.0 136800.0 1857750.0 ;
      RECT  138000.0 1858950.0 139200.0 1857750.0 ;
      RECT  140400.0 1858950.0 141600.0 1857750.0 ;
      RECT  140400.0 1858950.0 141600.0 1857750.0 ;
      RECT  138000.0 1858950.0 139200.0 1857750.0 ;
      RECT  135600.0 1867650.0 136800.0 1866450.0 ;
      RECT  138000.0 1867650.0 139200.0 1866450.0 ;
      RECT  138000.0 1867650.0 139200.0 1866450.0 ;
      RECT  135600.0 1867650.0 136800.0 1866450.0 ;
      RECT  138000.0 1867650.0 139200.0 1866450.0 ;
      RECT  140400.0 1867650.0 141600.0 1866450.0 ;
      RECT  140400.0 1867650.0 141600.0 1866450.0 ;
      RECT  138000.0 1867650.0 139200.0 1866450.0 ;
      RECT  142800.0 1858350.0 144000.0 1857150.0 ;
      RECT  142800.0 1868250.0 144000.0 1867050.0 ;
      RECT  140400.0 1865100.0 139200.0 1863900.0 ;
      RECT  137400.0 1862400.0 136200.0 1861200.0 ;
      RECT  138000.0 1858950.0 139200.0 1857750.0 ;
      RECT  140400.0 1867650.0 141600.0 1866450.0 ;
      RECT  141600.0 1862400.0 140400.0 1861200.0 ;
      RECT  136200.0 1862400.0 137400.0 1861200.0 ;
      RECT  139200.0 1865100.0 140400.0 1863900.0 ;
      RECT  140400.0 1862400.0 141600.0 1861200.0 ;
      RECT  133800.0 1856250.0 148200.0 1855350.0 ;
      RECT  133800.0 1870050.0 148200.0 1869150.0 ;
      RECT  154800.0 1857750.0 156000.0 1855800.0 ;
      RECT  154800.0 1869600.0 156000.0 1867650.0 ;
      RECT  150000.0 1868250.0 151200.0 1870050.0 ;
      RECT  150000.0 1858950.0 151200.0 1855350.0 ;
      RECT  152700.0 1868250.0 153600.0 1858950.0 ;
      RECT  150000.0 1858950.0 151200.0 1857750.0 ;
      RECT  152400.0 1858950.0 153600.0 1857750.0 ;
      RECT  152400.0 1858950.0 153600.0 1857750.0 ;
      RECT  150000.0 1858950.0 151200.0 1857750.0 ;
      RECT  150000.0 1868250.0 151200.0 1867050.0 ;
      RECT  152400.0 1868250.0 153600.0 1867050.0 ;
      RECT  152400.0 1868250.0 153600.0 1867050.0 ;
      RECT  150000.0 1868250.0 151200.0 1867050.0 ;
      RECT  154800.0 1858350.0 156000.0 1857150.0 ;
      RECT  154800.0 1868250.0 156000.0 1867050.0 ;
      RECT  150600.0 1863600.0 151800.0 1862400.0 ;
      RECT  150600.0 1863600.0 151800.0 1862400.0 ;
      RECT  153150.0 1863450.0 154050.0 1862550.0 ;
      RECT  148200.0 1856250.0 157800.0 1855350.0 ;
      RECT  148200.0 1870050.0 157800.0 1869150.0 ;
      RECT  120450.0 1862400.0 121650.0 1863600.0 ;
      RECT  122400.0 1864800.0 123600.0 1866000.0 ;
      RECT  139200.0 1863900.0 138000.0 1865100.0 ;
      RECT  130800.0 1881450.0 132000.0 1883400.0 ;
      RECT  130800.0 1869600.0 132000.0 1871550.0 ;
      RECT  126000.0 1870950.0 127200.0 1869150.0 ;
      RECT  126000.0 1880250.0 127200.0 1883850.0 ;
      RECT  128700.0 1870950.0 129600.0 1880250.0 ;
      RECT  126000.0 1880250.0 127200.0 1881450.0 ;
      RECT  128400.0 1880250.0 129600.0 1881450.0 ;
      RECT  128400.0 1880250.0 129600.0 1881450.0 ;
      RECT  126000.0 1880250.0 127200.0 1881450.0 ;
      RECT  126000.0 1870950.0 127200.0 1872150.0 ;
      RECT  128400.0 1870950.0 129600.0 1872150.0 ;
      RECT  128400.0 1870950.0 129600.0 1872150.0 ;
      RECT  126000.0 1870950.0 127200.0 1872150.0 ;
      RECT  130800.0 1880850.0 132000.0 1882050.0 ;
      RECT  130800.0 1870950.0 132000.0 1872150.0 ;
      RECT  126600.0 1875600.0 127800.0 1876800.0 ;
      RECT  126600.0 1875600.0 127800.0 1876800.0 ;
      RECT  129150.0 1875750.0 130050.0 1876650.0 ;
      RECT  124200.0 1882950.0 133800.0 1883850.0 ;
      RECT  124200.0 1869150.0 133800.0 1870050.0 ;
      RECT  135600.0 1871550.0 136800.0 1869150.0 ;
      RECT  135600.0 1880250.0 136800.0 1883850.0 ;
      RECT  140400.0 1880250.0 141600.0 1883850.0 ;
      RECT  142800.0 1881450.0 144000.0 1883400.0 ;
      RECT  142800.0 1869600.0 144000.0 1871550.0 ;
      RECT  135600.0 1880250.0 136800.0 1881450.0 ;
      RECT  138000.0 1880250.0 139200.0 1881450.0 ;
      RECT  138000.0 1880250.0 139200.0 1881450.0 ;
      RECT  135600.0 1880250.0 136800.0 1881450.0 ;
      RECT  138000.0 1880250.0 139200.0 1881450.0 ;
      RECT  140400.0 1880250.0 141600.0 1881450.0 ;
      RECT  140400.0 1880250.0 141600.0 1881450.0 ;
      RECT  138000.0 1880250.0 139200.0 1881450.0 ;
      RECT  135600.0 1871550.0 136800.0 1872750.0 ;
      RECT  138000.0 1871550.0 139200.0 1872750.0 ;
      RECT  138000.0 1871550.0 139200.0 1872750.0 ;
      RECT  135600.0 1871550.0 136800.0 1872750.0 ;
      RECT  138000.0 1871550.0 139200.0 1872750.0 ;
      RECT  140400.0 1871550.0 141600.0 1872750.0 ;
      RECT  140400.0 1871550.0 141600.0 1872750.0 ;
      RECT  138000.0 1871550.0 139200.0 1872750.0 ;
      RECT  142800.0 1880850.0 144000.0 1882050.0 ;
      RECT  142800.0 1870950.0 144000.0 1872150.0 ;
      RECT  140400.0 1874100.0 139200.0 1875300.0 ;
      RECT  137400.0 1876800.0 136200.0 1878000.0 ;
      RECT  138000.0 1880250.0 139200.0 1881450.0 ;
      RECT  140400.0 1871550.0 141600.0 1872750.0 ;
      RECT  141600.0 1876800.0 140400.0 1878000.0 ;
      RECT  136200.0 1876800.0 137400.0 1878000.0 ;
      RECT  139200.0 1874100.0 140400.0 1875300.0 ;
      RECT  140400.0 1876800.0 141600.0 1878000.0 ;
      RECT  133800.0 1882950.0 148200.0 1883850.0 ;
      RECT  133800.0 1869150.0 148200.0 1870050.0 ;
      RECT  154800.0 1881450.0 156000.0 1883400.0 ;
      RECT  154800.0 1869600.0 156000.0 1871550.0 ;
      RECT  150000.0 1870950.0 151200.0 1869150.0 ;
      RECT  150000.0 1880250.0 151200.0 1883850.0 ;
      RECT  152700.0 1870950.0 153600.0 1880250.0 ;
      RECT  150000.0 1880250.0 151200.0 1881450.0 ;
      RECT  152400.0 1880250.0 153600.0 1881450.0 ;
      RECT  152400.0 1880250.0 153600.0 1881450.0 ;
      RECT  150000.0 1880250.0 151200.0 1881450.0 ;
      RECT  150000.0 1870950.0 151200.0 1872150.0 ;
      RECT  152400.0 1870950.0 153600.0 1872150.0 ;
      RECT  152400.0 1870950.0 153600.0 1872150.0 ;
      RECT  150000.0 1870950.0 151200.0 1872150.0 ;
      RECT  154800.0 1880850.0 156000.0 1882050.0 ;
      RECT  154800.0 1870950.0 156000.0 1872150.0 ;
      RECT  150600.0 1875600.0 151800.0 1876800.0 ;
      RECT  150600.0 1875600.0 151800.0 1876800.0 ;
      RECT  153150.0 1875750.0 154050.0 1876650.0 ;
      RECT  148200.0 1882950.0 157800.0 1883850.0 ;
      RECT  148200.0 1869150.0 157800.0 1870050.0 ;
      RECT  120450.0 1875600.0 121650.0 1876800.0 ;
      RECT  122400.0 1873200.0 123600.0 1874400.0 ;
      RECT  139200.0 1874100.0 138000.0 1875300.0 ;
      RECT  130800.0 1885350.0 132000.0 1883400.0 ;
      RECT  130800.0 1897200.0 132000.0 1895250.0 ;
      RECT  126000.0 1895850.0 127200.0 1897650.0 ;
      RECT  126000.0 1886550.0 127200.0 1882950.0 ;
      RECT  128700.0 1895850.0 129600.0 1886550.0 ;
      RECT  126000.0 1886550.0 127200.0 1885350.0 ;
      RECT  128400.0 1886550.0 129600.0 1885350.0 ;
      RECT  128400.0 1886550.0 129600.0 1885350.0 ;
      RECT  126000.0 1886550.0 127200.0 1885350.0 ;
      RECT  126000.0 1895850.0 127200.0 1894650.0 ;
      RECT  128400.0 1895850.0 129600.0 1894650.0 ;
      RECT  128400.0 1895850.0 129600.0 1894650.0 ;
      RECT  126000.0 1895850.0 127200.0 1894650.0 ;
      RECT  130800.0 1885950.0 132000.0 1884750.0 ;
      RECT  130800.0 1895850.0 132000.0 1894650.0 ;
      RECT  126600.0 1891200.0 127800.0 1890000.0 ;
      RECT  126600.0 1891200.0 127800.0 1890000.0 ;
      RECT  129150.0 1891050.0 130050.0 1890150.0 ;
      RECT  124200.0 1883850.0 133800.0 1882950.0 ;
      RECT  124200.0 1897650.0 133800.0 1896750.0 ;
      RECT  135600.0 1895250.0 136800.0 1897650.0 ;
      RECT  135600.0 1886550.0 136800.0 1882950.0 ;
      RECT  140400.0 1886550.0 141600.0 1882950.0 ;
      RECT  142800.0 1885350.0 144000.0 1883400.0 ;
      RECT  142800.0 1897200.0 144000.0 1895250.0 ;
      RECT  135600.0 1886550.0 136800.0 1885350.0 ;
      RECT  138000.0 1886550.0 139200.0 1885350.0 ;
      RECT  138000.0 1886550.0 139200.0 1885350.0 ;
      RECT  135600.0 1886550.0 136800.0 1885350.0 ;
      RECT  138000.0 1886550.0 139200.0 1885350.0 ;
      RECT  140400.0 1886550.0 141600.0 1885350.0 ;
      RECT  140400.0 1886550.0 141600.0 1885350.0 ;
      RECT  138000.0 1886550.0 139200.0 1885350.0 ;
      RECT  135600.0 1895250.0 136800.0 1894050.0 ;
      RECT  138000.0 1895250.0 139200.0 1894050.0 ;
      RECT  138000.0 1895250.0 139200.0 1894050.0 ;
      RECT  135600.0 1895250.0 136800.0 1894050.0 ;
      RECT  138000.0 1895250.0 139200.0 1894050.0 ;
      RECT  140400.0 1895250.0 141600.0 1894050.0 ;
      RECT  140400.0 1895250.0 141600.0 1894050.0 ;
      RECT  138000.0 1895250.0 139200.0 1894050.0 ;
      RECT  142800.0 1885950.0 144000.0 1884750.0 ;
      RECT  142800.0 1895850.0 144000.0 1894650.0 ;
      RECT  140400.0 1892700.0 139200.0 1891500.0 ;
      RECT  137400.0 1890000.0 136200.0 1888800.0 ;
      RECT  138000.0 1886550.0 139200.0 1885350.0 ;
      RECT  140400.0 1895250.0 141600.0 1894050.0 ;
      RECT  141600.0 1890000.0 140400.0 1888800.0 ;
      RECT  136200.0 1890000.0 137400.0 1888800.0 ;
      RECT  139200.0 1892700.0 140400.0 1891500.0 ;
      RECT  140400.0 1890000.0 141600.0 1888800.0 ;
      RECT  133800.0 1883850.0 148200.0 1882950.0 ;
      RECT  133800.0 1897650.0 148200.0 1896750.0 ;
      RECT  154800.0 1885350.0 156000.0 1883400.0 ;
      RECT  154800.0 1897200.0 156000.0 1895250.0 ;
      RECT  150000.0 1895850.0 151200.0 1897650.0 ;
      RECT  150000.0 1886550.0 151200.0 1882950.0 ;
      RECT  152700.0 1895850.0 153600.0 1886550.0 ;
      RECT  150000.0 1886550.0 151200.0 1885350.0 ;
      RECT  152400.0 1886550.0 153600.0 1885350.0 ;
      RECT  152400.0 1886550.0 153600.0 1885350.0 ;
      RECT  150000.0 1886550.0 151200.0 1885350.0 ;
      RECT  150000.0 1895850.0 151200.0 1894650.0 ;
      RECT  152400.0 1895850.0 153600.0 1894650.0 ;
      RECT  152400.0 1895850.0 153600.0 1894650.0 ;
      RECT  150000.0 1895850.0 151200.0 1894650.0 ;
      RECT  154800.0 1885950.0 156000.0 1884750.0 ;
      RECT  154800.0 1895850.0 156000.0 1894650.0 ;
      RECT  150600.0 1891200.0 151800.0 1890000.0 ;
      RECT  150600.0 1891200.0 151800.0 1890000.0 ;
      RECT  153150.0 1891050.0 154050.0 1890150.0 ;
      RECT  148200.0 1883850.0 157800.0 1882950.0 ;
      RECT  148200.0 1897650.0 157800.0 1896750.0 ;
      RECT  120450.0 1890000.0 121650.0 1891200.0 ;
      RECT  122400.0 1892400.0 123600.0 1893600.0 ;
      RECT  139200.0 1891500.0 138000.0 1892700.0 ;
      RECT  130800.0 1909050.0 132000.0 1911000.0 ;
      RECT  130800.0 1897200.0 132000.0 1899150.0 ;
      RECT  126000.0 1898550.0 127200.0 1896750.0 ;
      RECT  126000.0 1907850.0 127200.0 1911450.0 ;
      RECT  128700.0 1898550.0 129600.0 1907850.0 ;
      RECT  126000.0 1907850.0 127200.0 1909050.0 ;
      RECT  128400.0 1907850.0 129600.0 1909050.0 ;
      RECT  128400.0 1907850.0 129600.0 1909050.0 ;
      RECT  126000.0 1907850.0 127200.0 1909050.0 ;
      RECT  126000.0 1898550.0 127200.0 1899750.0 ;
      RECT  128400.0 1898550.0 129600.0 1899750.0 ;
      RECT  128400.0 1898550.0 129600.0 1899750.0 ;
      RECT  126000.0 1898550.0 127200.0 1899750.0 ;
      RECT  130800.0 1908450.0 132000.0 1909650.0 ;
      RECT  130800.0 1898550.0 132000.0 1899750.0 ;
      RECT  126600.0 1903200.0 127800.0 1904400.0 ;
      RECT  126600.0 1903200.0 127800.0 1904400.0 ;
      RECT  129150.0 1903350.0 130050.0 1904250.0 ;
      RECT  124200.0 1910550.0 133800.0 1911450.0 ;
      RECT  124200.0 1896750.0 133800.0 1897650.0 ;
      RECT  135600.0 1899150.0 136800.0 1896750.0 ;
      RECT  135600.0 1907850.0 136800.0 1911450.0 ;
      RECT  140400.0 1907850.0 141600.0 1911450.0 ;
      RECT  142800.0 1909050.0 144000.0 1911000.0 ;
      RECT  142800.0 1897200.0 144000.0 1899150.0 ;
      RECT  135600.0 1907850.0 136800.0 1909050.0 ;
      RECT  138000.0 1907850.0 139200.0 1909050.0 ;
      RECT  138000.0 1907850.0 139200.0 1909050.0 ;
      RECT  135600.0 1907850.0 136800.0 1909050.0 ;
      RECT  138000.0 1907850.0 139200.0 1909050.0 ;
      RECT  140400.0 1907850.0 141600.0 1909050.0 ;
      RECT  140400.0 1907850.0 141600.0 1909050.0 ;
      RECT  138000.0 1907850.0 139200.0 1909050.0 ;
      RECT  135600.0 1899150.0 136800.0 1900350.0 ;
      RECT  138000.0 1899150.0 139200.0 1900350.0 ;
      RECT  138000.0 1899150.0 139200.0 1900350.0 ;
      RECT  135600.0 1899150.0 136800.0 1900350.0 ;
      RECT  138000.0 1899150.0 139200.0 1900350.0 ;
      RECT  140400.0 1899150.0 141600.0 1900350.0 ;
      RECT  140400.0 1899150.0 141600.0 1900350.0 ;
      RECT  138000.0 1899150.0 139200.0 1900350.0 ;
      RECT  142800.0 1908450.0 144000.0 1909650.0 ;
      RECT  142800.0 1898550.0 144000.0 1899750.0 ;
      RECT  140400.0 1901700.0 139200.0 1902900.0 ;
      RECT  137400.0 1904400.0 136200.0 1905600.0 ;
      RECT  138000.0 1907850.0 139200.0 1909050.0 ;
      RECT  140400.0 1899150.0 141600.0 1900350.0 ;
      RECT  141600.0 1904400.0 140400.0 1905600.0 ;
      RECT  136200.0 1904400.0 137400.0 1905600.0 ;
      RECT  139200.0 1901700.0 140400.0 1902900.0 ;
      RECT  140400.0 1904400.0 141600.0 1905600.0 ;
      RECT  133800.0 1910550.0 148200.0 1911450.0 ;
      RECT  133800.0 1896750.0 148200.0 1897650.0 ;
      RECT  154800.0 1909050.0 156000.0 1911000.0 ;
      RECT  154800.0 1897200.0 156000.0 1899150.0 ;
      RECT  150000.0 1898550.0 151200.0 1896750.0 ;
      RECT  150000.0 1907850.0 151200.0 1911450.0 ;
      RECT  152700.0 1898550.0 153600.0 1907850.0 ;
      RECT  150000.0 1907850.0 151200.0 1909050.0 ;
      RECT  152400.0 1907850.0 153600.0 1909050.0 ;
      RECT  152400.0 1907850.0 153600.0 1909050.0 ;
      RECT  150000.0 1907850.0 151200.0 1909050.0 ;
      RECT  150000.0 1898550.0 151200.0 1899750.0 ;
      RECT  152400.0 1898550.0 153600.0 1899750.0 ;
      RECT  152400.0 1898550.0 153600.0 1899750.0 ;
      RECT  150000.0 1898550.0 151200.0 1899750.0 ;
      RECT  154800.0 1908450.0 156000.0 1909650.0 ;
      RECT  154800.0 1898550.0 156000.0 1899750.0 ;
      RECT  150600.0 1903200.0 151800.0 1904400.0 ;
      RECT  150600.0 1903200.0 151800.0 1904400.0 ;
      RECT  153150.0 1903350.0 154050.0 1904250.0 ;
      RECT  148200.0 1910550.0 157800.0 1911450.0 ;
      RECT  148200.0 1896750.0 157800.0 1897650.0 ;
      RECT  120450.0 1903200.0 121650.0 1904400.0 ;
      RECT  122400.0 1900800.0 123600.0 1902000.0 ;
      RECT  139200.0 1901700.0 138000.0 1902900.0 ;
      RECT  130800.0 1912950.0 132000.0 1911000.0 ;
      RECT  130800.0 1924800.0 132000.0 1922850.0 ;
      RECT  126000.0 1923450.0 127200.0 1925250.0 ;
      RECT  126000.0 1914150.0 127200.0 1910550.0 ;
      RECT  128700.0 1923450.0 129600.0 1914150.0 ;
      RECT  126000.0 1914150.0 127200.0 1912950.0 ;
      RECT  128400.0 1914150.0 129600.0 1912950.0 ;
      RECT  128400.0 1914150.0 129600.0 1912950.0 ;
      RECT  126000.0 1914150.0 127200.0 1912950.0 ;
      RECT  126000.0 1923450.0 127200.0 1922250.0 ;
      RECT  128400.0 1923450.0 129600.0 1922250.0 ;
      RECT  128400.0 1923450.0 129600.0 1922250.0 ;
      RECT  126000.0 1923450.0 127200.0 1922250.0 ;
      RECT  130800.0 1913550.0 132000.0 1912350.0 ;
      RECT  130800.0 1923450.0 132000.0 1922250.0 ;
      RECT  126600.0 1918800.0 127800.0 1917600.0 ;
      RECT  126600.0 1918800.0 127800.0 1917600.0 ;
      RECT  129150.0 1918650.0 130050.0 1917750.0 ;
      RECT  124200.0 1911450.0 133800.0 1910550.0 ;
      RECT  124200.0 1925250.0 133800.0 1924350.0 ;
      RECT  135600.0 1922850.0 136800.0 1925250.0 ;
      RECT  135600.0 1914150.0 136800.0 1910550.0 ;
      RECT  140400.0 1914150.0 141600.0 1910550.0 ;
      RECT  142800.0 1912950.0 144000.0 1911000.0 ;
      RECT  142800.0 1924800.0 144000.0 1922850.0 ;
      RECT  135600.0 1914150.0 136800.0 1912950.0 ;
      RECT  138000.0 1914150.0 139200.0 1912950.0 ;
      RECT  138000.0 1914150.0 139200.0 1912950.0 ;
      RECT  135600.0 1914150.0 136800.0 1912950.0 ;
      RECT  138000.0 1914150.0 139200.0 1912950.0 ;
      RECT  140400.0 1914150.0 141600.0 1912950.0 ;
      RECT  140400.0 1914150.0 141600.0 1912950.0 ;
      RECT  138000.0 1914150.0 139200.0 1912950.0 ;
      RECT  135600.0 1922850.0 136800.0 1921650.0 ;
      RECT  138000.0 1922850.0 139200.0 1921650.0 ;
      RECT  138000.0 1922850.0 139200.0 1921650.0 ;
      RECT  135600.0 1922850.0 136800.0 1921650.0 ;
      RECT  138000.0 1922850.0 139200.0 1921650.0 ;
      RECT  140400.0 1922850.0 141600.0 1921650.0 ;
      RECT  140400.0 1922850.0 141600.0 1921650.0 ;
      RECT  138000.0 1922850.0 139200.0 1921650.0 ;
      RECT  142800.0 1913550.0 144000.0 1912350.0 ;
      RECT  142800.0 1923450.0 144000.0 1922250.0 ;
      RECT  140400.0 1920300.0 139200.0 1919100.0 ;
      RECT  137400.0 1917600.0 136200.0 1916400.0 ;
      RECT  138000.0 1914150.0 139200.0 1912950.0 ;
      RECT  140400.0 1922850.0 141600.0 1921650.0 ;
      RECT  141600.0 1917600.0 140400.0 1916400.0 ;
      RECT  136200.0 1917600.0 137400.0 1916400.0 ;
      RECT  139200.0 1920300.0 140400.0 1919100.0 ;
      RECT  140400.0 1917600.0 141600.0 1916400.0 ;
      RECT  133800.0 1911450.0 148200.0 1910550.0 ;
      RECT  133800.0 1925250.0 148200.0 1924350.0 ;
      RECT  154800.0 1912950.0 156000.0 1911000.0 ;
      RECT  154800.0 1924800.0 156000.0 1922850.0 ;
      RECT  150000.0 1923450.0 151200.0 1925250.0 ;
      RECT  150000.0 1914150.0 151200.0 1910550.0 ;
      RECT  152700.0 1923450.0 153600.0 1914150.0 ;
      RECT  150000.0 1914150.0 151200.0 1912950.0 ;
      RECT  152400.0 1914150.0 153600.0 1912950.0 ;
      RECT  152400.0 1914150.0 153600.0 1912950.0 ;
      RECT  150000.0 1914150.0 151200.0 1912950.0 ;
      RECT  150000.0 1923450.0 151200.0 1922250.0 ;
      RECT  152400.0 1923450.0 153600.0 1922250.0 ;
      RECT  152400.0 1923450.0 153600.0 1922250.0 ;
      RECT  150000.0 1923450.0 151200.0 1922250.0 ;
      RECT  154800.0 1913550.0 156000.0 1912350.0 ;
      RECT  154800.0 1923450.0 156000.0 1922250.0 ;
      RECT  150600.0 1918800.0 151800.0 1917600.0 ;
      RECT  150600.0 1918800.0 151800.0 1917600.0 ;
      RECT  153150.0 1918650.0 154050.0 1917750.0 ;
      RECT  148200.0 1911450.0 157800.0 1910550.0 ;
      RECT  148200.0 1925250.0 157800.0 1924350.0 ;
      RECT  120450.0 1917600.0 121650.0 1918800.0 ;
      RECT  122400.0 1920000.0 123600.0 1921200.0 ;
      RECT  139200.0 1919100.0 138000.0 1920300.0 ;
      RECT  130800.0 1936650.0 132000.0 1938600.0 ;
      RECT  130800.0 1924800.0 132000.0 1926750.0 ;
      RECT  126000.0 1926150.0 127200.0 1924350.0 ;
      RECT  126000.0 1935450.0 127200.0 1939050.0 ;
      RECT  128700.0 1926150.0 129600.0 1935450.0 ;
      RECT  126000.0 1935450.0 127200.0 1936650.0 ;
      RECT  128400.0 1935450.0 129600.0 1936650.0 ;
      RECT  128400.0 1935450.0 129600.0 1936650.0 ;
      RECT  126000.0 1935450.0 127200.0 1936650.0 ;
      RECT  126000.0 1926150.0 127200.0 1927350.0 ;
      RECT  128400.0 1926150.0 129600.0 1927350.0 ;
      RECT  128400.0 1926150.0 129600.0 1927350.0 ;
      RECT  126000.0 1926150.0 127200.0 1927350.0 ;
      RECT  130800.0 1936050.0 132000.0 1937250.0 ;
      RECT  130800.0 1926150.0 132000.0 1927350.0 ;
      RECT  126600.0 1930800.0 127800.0 1932000.0 ;
      RECT  126600.0 1930800.0 127800.0 1932000.0 ;
      RECT  129150.0 1930950.0 130050.0 1931850.0 ;
      RECT  124200.0 1938150.0 133800.0 1939050.0 ;
      RECT  124200.0 1924350.0 133800.0 1925250.0 ;
      RECT  135600.0 1926750.0 136800.0 1924350.0 ;
      RECT  135600.0 1935450.0 136800.0 1939050.0 ;
      RECT  140400.0 1935450.0 141600.0 1939050.0 ;
      RECT  142800.0 1936650.0 144000.0 1938600.0 ;
      RECT  142800.0 1924800.0 144000.0 1926750.0 ;
      RECT  135600.0 1935450.0 136800.0 1936650.0 ;
      RECT  138000.0 1935450.0 139200.0 1936650.0 ;
      RECT  138000.0 1935450.0 139200.0 1936650.0 ;
      RECT  135600.0 1935450.0 136800.0 1936650.0 ;
      RECT  138000.0 1935450.0 139200.0 1936650.0 ;
      RECT  140400.0 1935450.0 141600.0 1936650.0 ;
      RECT  140400.0 1935450.0 141600.0 1936650.0 ;
      RECT  138000.0 1935450.0 139200.0 1936650.0 ;
      RECT  135600.0 1926750.0 136800.0 1927950.0 ;
      RECT  138000.0 1926750.0 139200.0 1927950.0 ;
      RECT  138000.0 1926750.0 139200.0 1927950.0 ;
      RECT  135600.0 1926750.0 136800.0 1927950.0 ;
      RECT  138000.0 1926750.0 139200.0 1927950.0 ;
      RECT  140400.0 1926750.0 141600.0 1927950.0 ;
      RECT  140400.0 1926750.0 141600.0 1927950.0 ;
      RECT  138000.0 1926750.0 139200.0 1927950.0 ;
      RECT  142800.0 1936050.0 144000.0 1937250.0 ;
      RECT  142800.0 1926150.0 144000.0 1927350.0 ;
      RECT  140400.0 1929300.0 139200.0 1930500.0 ;
      RECT  137400.0 1932000.0 136200.0 1933200.0 ;
      RECT  138000.0 1935450.0 139200.0 1936650.0 ;
      RECT  140400.0 1926750.0 141600.0 1927950.0 ;
      RECT  141600.0 1932000.0 140400.0 1933200.0 ;
      RECT  136200.0 1932000.0 137400.0 1933200.0 ;
      RECT  139200.0 1929300.0 140400.0 1930500.0 ;
      RECT  140400.0 1932000.0 141600.0 1933200.0 ;
      RECT  133800.0 1938150.0 148200.0 1939050.0 ;
      RECT  133800.0 1924350.0 148200.0 1925250.0 ;
      RECT  154800.0 1936650.0 156000.0 1938600.0 ;
      RECT  154800.0 1924800.0 156000.0 1926750.0 ;
      RECT  150000.0 1926150.0 151200.0 1924350.0 ;
      RECT  150000.0 1935450.0 151200.0 1939050.0 ;
      RECT  152700.0 1926150.0 153600.0 1935450.0 ;
      RECT  150000.0 1935450.0 151200.0 1936650.0 ;
      RECT  152400.0 1935450.0 153600.0 1936650.0 ;
      RECT  152400.0 1935450.0 153600.0 1936650.0 ;
      RECT  150000.0 1935450.0 151200.0 1936650.0 ;
      RECT  150000.0 1926150.0 151200.0 1927350.0 ;
      RECT  152400.0 1926150.0 153600.0 1927350.0 ;
      RECT  152400.0 1926150.0 153600.0 1927350.0 ;
      RECT  150000.0 1926150.0 151200.0 1927350.0 ;
      RECT  154800.0 1936050.0 156000.0 1937250.0 ;
      RECT  154800.0 1926150.0 156000.0 1927350.0 ;
      RECT  150600.0 1930800.0 151800.0 1932000.0 ;
      RECT  150600.0 1930800.0 151800.0 1932000.0 ;
      RECT  153150.0 1930950.0 154050.0 1931850.0 ;
      RECT  148200.0 1938150.0 157800.0 1939050.0 ;
      RECT  148200.0 1924350.0 157800.0 1925250.0 ;
      RECT  120450.0 1930800.0 121650.0 1932000.0 ;
      RECT  122400.0 1928400.0 123600.0 1929600.0 ;
      RECT  139200.0 1929300.0 138000.0 1930500.0 ;
      RECT  130800.0 1940550.0 132000.0 1938600.0 ;
      RECT  130800.0 1952400.0 132000.0 1950450.0 ;
      RECT  126000.0 1951050.0 127200.0 1952850.0 ;
      RECT  126000.0 1941750.0 127200.0 1938150.0 ;
      RECT  128700.0 1951050.0 129600.0 1941750.0 ;
      RECT  126000.0 1941750.0 127200.0 1940550.0 ;
      RECT  128400.0 1941750.0 129600.0 1940550.0 ;
      RECT  128400.0 1941750.0 129600.0 1940550.0 ;
      RECT  126000.0 1941750.0 127200.0 1940550.0 ;
      RECT  126000.0 1951050.0 127200.0 1949850.0 ;
      RECT  128400.0 1951050.0 129600.0 1949850.0 ;
      RECT  128400.0 1951050.0 129600.0 1949850.0 ;
      RECT  126000.0 1951050.0 127200.0 1949850.0 ;
      RECT  130800.0 1941150.0 132000.0 1939950.0 ;
      RECT  130800.0 1951050.0 132000.0 1949850.0 ;
      RECT  126600.0 1946400.0 127800.0 1945200.0 ;
      RECT  126600.0 1946400.0 127800.0 1945200.0 ;
      RECT  129150.0 1946250.0 130050.0 1945350.0 ;
      RECT  124200.0 1939050.0 133800.0 1938150.0 ;
      RECT  124200.0 1952850.0 133800.0 1951950.0 ;
      RECT  135600.0 1950450.0 136800.0 1952850.0 ;
      RECT  135600.0 1941750.0 136800.0 1938150.0 ;
      RECT  140400.0 1941750.0 141600.0 1938150.0 ;
      RECT  142800.0 1940550.0 144000.0 1938600.0 ;
      RECT  142800.0 1952400.0 144000.0 1950450.0 ;
      RECT  135600.0 1941750.0 136800.0 1940550.0 ;
      RECT  138000.0 1941750.0 139200.0 1940550.0 ;
      RECT  138000.0 1941750.0 139200.0 1940550.0 ;
      RECT  135600.0 1941750.0 136800.0 1940550.0 ;
      RECT  138000.0 1941750.0 139200.0 1940550.0 ;
      RECT  140400.0 1941750.0 141600.0 1940550.0 ;
      RECT  140400.0 1941750.0 141600.0 1940550.0 ;
      RECT  138000.0 1941750.0 139200.0 1940550.0 ;
      RECT  135600.0 1950450.0 136800.0 1949250.0 ;
      RECT  138000.0 1950450.0 139200.0 1949250.0 ;
      RECT  138000.0 1950450.0 139200.0 1949250.0 ;
      RECT  135600.0 1950450.0 136800.0 1949250.0 ;
      RECT  138000.0 1950450.0 139200.0 1949250.0 ;
      RECT  140400.0 1950450.0 141600.0 1949250.0 ;
      RECT  140400.0 1950450.0 141600.0 1949250.0 ;
      RECT  138000.0 1950450.0 139200.0 1949250.0 ;
      RECT  142800.0 1941150.0 144000.0 1939950.0 ;
      RECT  142800.0 1951050.0 144000.0 1949850.0 ;
      RECT  140400.0 1947900.0 139200.0 1946700.0 ;
      RECT  137400.0 1945200.0 136200.0 1944000.0 ;
      RECT  138000.0 1941750.0 139200.0 1940550.0 ;
      RECT  140400.0 1950450.0 141600.0 1949250.0 ;
      RECT  141600.0 1945200.0 140400.0 1944000.0 ;
      RECT  136200.0 1945200.0 137400.0 1944000.0 ;
      RECT  139200.0 1947900.0 140400.0 1946700.0 ;
      RECT  140400.0 1945200.0 141600.0 1944000.0 ;
      RECT  133800.0 1939050.0 148200.0 1938150.0 ;
      RECT  133800.0 1952850.0 148200.0 1951950.0 ;
      RECT  154800.0 1940550.0 156000.0 1938600.0 ;
      RECT  154800.0 1952400.0 156000.0 1950450.0 ;
      RECT  150000.0 1951050.0 151200.0 1952850.0 ;
      RECT  150000.0 1941750.0 151200.0 1938150.0 ;
      RECT  152700.0 1951050.0 153600.0 1941750.0 ;
      RECT  150000.0 1941750.0 151200.0 1940550.0 ;
      RECT  152400.0 1941750.0 153600.0 1940550.0 ;
      RECT  152400.0 1941750.0 153600.0 1940550.0 ;
      RECT  150000.0 1941750.0 151200.0 1940550.0 ;
      RECT  150000.0 1951050.0 151200.0 1949850.0 ;
      RECT  152400.0 1951050.0 153600.0 1949850.0 ;
      RECT  152400.0 1951050.0 153600.0 1949850.0 ;
      RECT  150000.0 1951050.0 151200.0 1949850.0 ;
      RECT  154800.0 1941150.0 156000.0 1939950.0 ;
      RECT  154800.0 1951050.0 156000.0 1949850.0 ;
      RECT  150600.0 1946400.0 151800.0 1945200.0 ;
      RECT  150600.0 1946400.0 151800.0 1945200.0 ;
      RECT  153150.0 1946250.0 154050.0 1945350.0 ;
      RECT  148200.0 1939050.0 157800.0 1938150.0 ;
      RECT  148200.0 1952850.0 157800.0 1951950.0 ;
      RECT  120450.0 1945200.0 121650.0 1946400.0 ;
      RECT  122400.0 1947600.0 123600.0 1948800.0 ;
      RECT  139200.0 1946700.0 138000.0 1947900.0 ;
      RECT  130800.0 1964250.0 132000.0 1966200.0 ;
      RECT  130800.0 1952400.0 132000.0 1954350.0 ;
      RECT  126000.0 1953750.0 127200.0 1951950.0 ;
      RECT  126000.0 1963050.0 127200.0 1966650.0 ;
      RECT  128700.0 1953750.0 129600.0 1963050.0 ;
      RECT  126000.0 1963050.0 127200.0 1964250.0 ;
      RECT  128400.0 1963050.0 129600.0 1964250.0 ;
      RECT  128400.0 1963050.0 129600.0 1964250.0 ;
      RECT  126000.0 1963050.0 127200.0 1964250.0 ;
      RECT  126000.0 1953750.0 127200.0 1954950.0 ;
      RECT  128400.0 1953750.0 129600.0 1954950.0 ;
      RECT  128400.0 1953750.0 129600.0 1954950.0 ;
      RECT  126000.0 1953750.0 127200.0 1954950.0 ;
      RECT  130800.0 1963650.0 132000.0 1964850.0 ;
      RECT  130800.0 1953750.0 132000.0 1954950.0 ;
      RECT  126600.0 1958400.0 127800.0 1959600.0 ;
      RECT  126600.0 1958400.0 127800.0 1959600.0 ;
      RECT  129150.0 1958550.0 130050.0 1959450.0 ;
      RECT  124200.0 1965750.0 133800.0 1966650.0 ;
      RECT  124200.0 1951950.0 133800.0 1952850.0 ;
      RECT  135600.0 1954350.0 136800.0 1951950.0 ;
      RECT  135600.0 1963050.0 136800.0 1966650.0 ;
      RECT  140400.0 1963050.0 141600.0 1966650.0 ;
      RECT  142800.0 1964250.0 144000.0 1966200.0 ;
      RECT  142800.0 1952400.0 144000.0 1954350.0 ;
      RECT  135600.0 1963050.0 136800.0 1964250.0 ;
      RECT  138000.0 1963050.0 139200.0 1964250.0 ;
      RECT  138000.0 1963050.0 139200.0 1964250.0 ;
      RECT  135600.0 1963050.0 136800.0 1964250.0 ;
      RECT  138000.0 1963050.0 139200.0 1964250.0 ;
      RECT  140400.0 1963050.0 141600.0 1964250.0 ;
      RECT  140400.0 1963050.0 141600.0 1964250.0 ;
      RECT  138000.0 1963050.0 139200.0 1964250.0 ;
      RECT  135600.0 1954350.0 136800.0 1955550.0 ;
      RECT  138000.0 1954350.0 139200.0 1955550.0 ;
      RECT  138000.0 1954350.0 139200.0 1955550.0 ;
      RECT  135600.0 1954350.0 136800.0 1955550.0 ;
      RECT  138000.0 1954350.0 139200.0 1955550.0 ;
      RECT  140400.0 1954350.0 141600.0 1955550.0 ;
      RECT  140400.0 1954350.0 141600.0 1955550.0 ;
      RECT  138000.0 1954350.0 139200.0 1955550.0 ;
      RECT  142800.0 1963650.0 144000.0 1964850.0 ;
      RECT  142800.0 1953750.0 144000.0 1954950.0 ;
      RECT  140400.0 1956900.0 139200.0 1958100.0 ;
      RECT  137400.0 1959600.0 136200.0 1960800.0 ;
      RECT  138000.0 1963050.0 139200.0 1964250.0 ;
      RECT  140400.0 1954350.0 141600.0 1955550.0 ;
      RECT  141600.0 1959600.0 140400.0 1960800.0 ;
      RECT  136200.0 1959600.0 137400.0 1960800.0 ;
      RECT  139200.0 1956900.0 140400.0 1958100.0 ;
      RECT  140400.0 1959600.0 141600.0 1960800.0 ;
      RECT  133800.0 1965750.0 148200.0 1966650.0 ;
      RECT  133800.0 1951950.0 148200.0 1952850.0 ;
      RECT  154800.0 1964250.0 156000.0 1966200.0 ;
      RECT  154800.0 1952400.0 156000.0 1954350.0 ;
      RECT  150000.0 1953750.0 151200.0 1951950.0 ;
      RECT  150000.0 1963050.0 151200.0 1966650.0 ;
      RECT  152700.0 1953750.0 153600.0 1963050.0 ;
      RECT  150000.0 1963050.0 151200.0 1964250.0 ;
      RECT  152400.0 1963050.0 153600.0 1964250.0 ;
      RECT  152400.0 1963050.0 153600.0 1964250.0 ;
      RECT  150000.0 1963050.0 151200.0 1964250.0 ;
      RECT  150000.0 1953750.0 151200.0 1954950.0 ;
      RECT  152400.0 1953750.0 153600.0 1954950.0 ;
      RECT  152400.0 1953750.0 153600.0 1954950.0 ;
      RECT  150000.0 1953750.0 151200.0 1954950.0 ;
      RECT  154800.0 1963650.0 156000.0 1964850.0 ;
      RECT  154800.0 1953750.0 156000.0 1954950.0 ;
      RECT  150600.0 1958400.0 151800.0 1959600.0 ;
      RECT  150600.0 1958400.0 151800.0 1959600.0 ;
      RECT  153150.0 1958550.0 154050.0 1959450.0 ;
      RECT  148200.0 1965750.0 157800.0 1966650.0 ;
      RECT  148200.0 1951950.0 157800.0 1952850.0 ;
      RECT  120450.0 1958400.0 121650.0 1959600.0 ;
      RECT  122400.0 1956000.0 123600.0 1957200.0 ;
      RECT  139200.0 1956900.0 138000.0 1958100.0 ;
      RECT  130800.0 1968150.0 132000.0 1966200.0 ;
      RECT  130800.0 1980000.0 132000.0 1978050.0 ;
      RECT  126000.0 1978650.0 127200.0 1980450.0 ;
      RECT  126000.0 1969350.0 127200.0 1965750.0 ;
      RECT  128700.0 1978650.0 129600.0 1969350.0 ;
      RECT  126000.0 1969350.0 127200.0 1968150.0 ;
      RECT  128400.0 1969350.0 129600.0 1968150.0 ;
      RECT  128400.0 1969350.0 129600.0 1968150.0 ;
      RECT  126000.0 1969350.0 127200.0 1968150.0 ;
      RECT  126000.0 1978650.0 127200.0 1977450.0 ;
      RECT  128400.0 1978650.0 129600.0 1977450.0 ;
      RECT  128400.0 1978650.0 129600.0 1977450.0 ;
      RECT  126000.0 1978650.0 127200.0 1977450.0 ;
      RECT  130800.0 1968750.0 132000.0 1967550.0 ;
      RECT  130800.0 1978650.0 132000.0 1977450.0 ;
      RECT  126600.0 1974000.0 127800.0 1972800.0 ;
      RECT  126600.0 1974000.0 127800.0 1972800.0 ;
      RECT  129150.0 1973850.0 130050.0 1972950.0 ;
      RECT  124200.0 1966650.0 133800.0 1965750.0 ;
      RECT  124200.0 1980450.0 133800.0 1979550.0 ;
      RECT  135600.0 1978050.0 136800.0 1980450.0 ;
      RECT  135600.0 1969350.0 136800.0 1965750.0 ;
      RECT  140400.0 1969350.0 141600.0 1965750.0 ;
      RECT  142800.0 1968150.0 144000.0 1966200.0 ;
      RECT  142800.0 1980000.0 144000.0 1978050.0 ;
      RECT  135600.0 1969350.0 136800.0 1968150.0 ;
      RECT  138000.0 1969350.0 139200.0 1968150.0 ;
      RECT  138000.0 1969350.0 139200.0 1968150.0 ;
      RECT  135600.0 1969350.0 136800.0 1968150.0 ;
      RECT  138000.0 1969350.0 139200.0 1968150.0 ;
      RECT  140400.0 1969350.0 141600.0 1968150.0 ;
      RECT  140400.0 1969350.0 141600.0 1968150.0 ;
      RECT  138000.0 1969350.0 139200.0 1968150.0 ;
      RECT  135600.0 1978050.0 136800.0 1976850.0 ;
      RECT  138000.0 1978050.0 139200.0 1976850.0 ;
      RECT  138000.0 1978050.0 139200.0 1976850.0 ;
      RECT  135600.0 1978050.0 136800.0 1976850.0 ;
      RECT  138000.0 1978050.0 139200.0 1976850.0 ;
      RECT  140400.0 1978050.0 141600.0 1976850.0 ;
      RECT  140400.0 1978050.0 141600.0 1976850.0 ;
      RECT  138000.0 1978050.0 139200.0 1976850.0 ;
      RECT  142800.0 1968750.0 144000.0 1967550.0 ;
      RECT  142800.0 1978650.0 144000.0 1977450.0 ;
      RECT  140400.0 1975500.0 139200.0 1974300.0 ;
      RECT  137400.0 1972800.0 136200.0 1971600.0 ;
      RECT  138000.0 1969350.0 139200.0 1968150.0 ;
      RECT  140400.0 1978050.0 141600.0 1976850.0 ;
      RECT  141600.0 1972800.0 140400.0 1971600.0 ;
      RECT  136200.0 1972800.0 137400.0 1971600.0 ;
      RECT  139200.0 1975500.0 140400.0 1974300.0 ;
      RECT  140400.0 1972800.0 141600.0 1971600.0 ;
      RECT  133800.0 1966650.0 148200.0 1965750.0 ;
      RECT  133800.0 1980450.0 148200.0 1979550.0 ;
      RECT  154800.0 1968150.0 156000.0 1966200.0 ;
      RECT  154800.0 1980000.0 156000.0 1978050.0 ;
      RECT  150000.0 1978650.0 151200.0 1980450.0 ;
      RECT  150000.0 1969350.0 151200.0 1965750.0 ;
      RECT  152700.0 1978650.0 153600.0 1969350.0 ;
      RECT  150000.0 1969350.0 151200.0 1968150.0 ;
      RECT  152400.0 1969350.0 153600.0 1968150.0 ;
      RECT  152400.0 1969350.0 153600.0 1968150.0 ;
      RECT  150000.0 1969350.0 151200.0 1968150.0 ;
      RECT  150000.0 1978650.0 151200.0 1977450.0 ;
      RECT  152400.0 1978650.0 153600.0 1977450.0 ;
      RECT  152400.0 1978650.0 153600.0 1977450.0 ;
      RECT  150000.0 1978650.0 151200.0 1977450.0 ;
      RECT  154800.0 1968750.0 156000.0 1967550.0 ;
      RECT  154800.0 1978650.0 156000.0 1977450.0 ;
      RECT  150600.0 1974000.0 151800.0 1972800.0 ;
      RECT  150600.0 1974000.0 151800.0 1972800.0 ;
      RECT  153150.0 1973850.0 154050.0 1972950.0 ;
      RECT  148200.0 1966650.0 157800.0 1965750.0 ;
      RECT  148200.0 1980450.0 157800.0 1979550.0 ;
      RECT  120450.0 1972800.0 121650.0 1974000.0 ;
      RECT  122400.0 1975200.0 123600.0 1976400.0 ;
      RECT  139200.0 1974300.0 138000.0 1975500.0 ;
      RECT  130800.0 1991850.0 132000.0 1993800.0 ;
      RECT  130800.0 1980000.0 132000.0 1981950.0 ;
      RECT  126000.0 1981350.0 127200.0 1979550.0 ;
      RECT  126000.0 1990650.0 127200.0 1994250.0 ;
      RECT  128700.0 1981350.0 129600.0 1990650.0 ;
      RECT  126000.0 1990650.0 127200.0 1991850.0 ;
      RECT  128400.0 1990650.0 129600.0 1991850.0 ;
      RECT  128400.0 1990650.0 129600.0 1991850.0 ;
      RECT  126000.0 1990650.0 127200.0 1991850.0 ;
      RECT  126000.0 1981350.0 127200.0 1982550.0 ;
      RECT  128400.0 1981350.0 129600.0 1982550.0 ;
      RECT  128400.0 1981350.0 129600.0 1982550.0 ;
      RECT  126000.0 1981350.0 127200.0 1982550.0 ;
      RECT  130800.0 1991250.0 132000.0 1992450.0 ;
      RECT  130800.0 1981350.0 132000.0 1982550.0 ;
      RECT  126600.0 1986000.0 127800.0 1987200.0 ;
      RECT  126600.0 1986000.0 127800.0 1987200.0 ;
      RECT  129150.0 1986150.0 130050.0 1987050.0 ;
      RECT  124200.0 1993350.0 133800.0 1994250.0 ;
      RECT  124200.0 1979550.0 133800.0 1980450.0 ;
      RECT  135600.0 1981950.0 136800.0 1979550.0 ;
      RECT  135600.0 1990650.0 136800.0 1994250.0 ;
      RECT  140400.0 1990650.0 141600.0 1994250.0 ;
      RECT  142800.0 1991850.0 144000.0 1993800.0 ;
      RECT  142800.0 1980000.0 144000.0 1981950.0 ;
      RECT  135600.0 1990650.0 136800.0 1991850.0 ;
      RECT  138000.0 1990650.0 139200.0 1991850.0 ;
      RECT  138000.0 1990650.0 139200.0 1991850.0 ;
      RECT  135600.0 1990650.0 136800.0 1991850.0 ;
      RECT  138000.0 1990650.0 139200.0 1991850.0 ;
      RECT  140400.0 1990650.0 141600.0 1991850.0 ;
      RECT  140400.0 1990650.0 141600.0 1991850.0 ;
      RECT  138000.0 1990650.0 139200.0 1991850.0 ;
      RECT  135600.0 1981950.0 136800.0 1983150.0 ;
      RECT  138000.0 1981950.0 139200.0 1983150.0 ;
      RECT  138000.0 1981950.0 139200.0 1983150.0 ;
      RECT  135600.0 1981950.0 136800.0 1983150.0 ;
      RECT  138000.0 1981950.0 139200.0 1983150.0 ;
      RECT  140400.0 1981950.0 141600.0 1983150.0 ;
      RECT  140400.0 1981950.0 141600.0 1983150.0 ;
      RECT  138000.0 1981950.0 139200.0 1983150.0 ;
      RECT  142800.0 1991250.0 144000.0 1992450.0 ;
      RECT  142800.0 1981350.0 144000.0 1982550.0 ;
      RECT  140400.0 1984500.0 139200.0 1985700.0 ;
      RECT  137400.0 1987200.0 136200.0 1988400.0 ;
      RECT  138000.0 1990650.0 139200.0 1991850.0 ;
      RECT  140400.0 1981950.0 141600.0 1983150.0 ;
      RECT  141600.0 1987200.0 140400.0 1988400.0 ;
      RECT  136200.0 1987200.0 137400.0 1988400.0 ;
      RECT  139200.0 1984500.0 140400.0 1985700.0 ;
      RECT  140400.0 1987200.0 141600.0 1988400.0 ;
      RECT  133800.0 1993350.0 148200.0 1994250.0 ;
      RECT  133800.0 1979550.0 148200.0 1980450.0 ;
      RECT  154800.0 1991850.0 156000.0 1993800.0 ;
      RECT  154800.0 1980000.0 156000.0 1981950.0 ;
      RECT  150000.0 1981350.0 151200.0 1979550.0 ;
      RECT  150000.0 1990650.0 151200.0 1994250.0 ;
      RECT  152700.0 1981350.0 153600.0 1990650.0 ;
      RECT  150000.0 1990650.0 151200.0 1991850.0 ;
      RECT  152400.0 1990650.0 153600.0 1991850.0 ;
      RECT  152400.0 1990650.0 153600.0 1991850.0 ;
      RECT  150000.0 1990650.0 151200.0 1991850.0 ;
      RECT  150000.0 1981350.0 151200.0 1982550.0 ;
      RECT  152400.0 1981350.0 153600.0 1982550.0 ;
      RECT  152400.0 1981350.0 153600.0 1982550.0 ;
      RECT  150000.0 1981350.0 151200.0 1982550.0 ;
      RECT  154800.0 1991250.0 156000.0 1992450.0 ;
      RECT  154800.0 1981350.0 156000.0 1982550.0 ;
      RECT  150600.0 1986000.0 151800.0 1987200.0 ;
      RECT  150600.0 1986000.0 151800.0 1987200.0 ;
      RECT  153150.0 1986150.0 154050.0 1987050.0 ;
      RECT  148200.0 1993350.0 157800.0 1994250.0 ;
      RECT  148200.0 1979550.0 157800.0 1980450.0 ;
      RECT  120450.0 1986000.0 121650.0 1987200.0 ;
      RECT  122400.0 1983600.0 123600.0 1984800.0 ;
      RECT  139200.0 1984500.0 138000.0 1985700.0 ;
      RECT  130800.0 1995750.0 132000.0 1993800.0 ;
      RECT  130800.0 2007600.0 132000.0 2005650.0 ;
      RECT  126000.0 2006250.0 127200.0 2008050.0 ;
      RECT  126000.0 1996950.0 127200.0 1993350.0 ;
      RECT  128700.0 2006250.0 129600.0 1996950.0 ;
      RECT  126000.0 1996950.0 127200.0 1995750.0 ;
      RECT  128400.0 1996950.0 129600.0 1995750.0 ;
      RECT  128400.0 1996950.0 129600.0 1995750.0 ;
      RECT  126000.0 1996950.0 127200.0 1995750.0 ;
      RECT  126000.0 2006250.0 127200.0 2005050.0 ;
      RECT  128400.0 2006250.0 129600.0 2005050.0 ;
      RECT  128400.0 2006250.0 129600.0 2005050.0 ;
      RECT  126000.0 2006250.0 127200.0 2005050.0 ;
      RECT  130800.0 1996350.0 132000.0 1995150.0 ;
      RECT  130800.0 2006250.0 132000.0 2005050.0 ;
      RECT  126600.0 2001600.0 127800.0 2000400.0 ;
      RECT  126600.0 2001600.0 127800.0 2000400.0 ;
      RECT  129150.0 2001450.0 130050.0 2000550.0 ;
      RECT  124200.0 1994250.0 133800.0 1993350.0 ;
      RECT  124200.0 2008050.0 133800.0 2007150.0 ;
      RECT  135600.0 2005650.0 136800.0 2008050.0 ;
      RECT  135600.0 1996950.0 136800.0 1993350.0 ;
      RECT  140400.0 1996950.0 141600.0 1993350.0 ;
      RECT  142800.0 1995750.0 144000.0 1993800.0 ;
      RECT  142800.0 2007600.0 144000.0 2005650.0 ;
      RECT  135600.0 1996950.0 136800.0 1995750.0 ;
      RECT  138000.0 1996950.0 139200.0 1995750.0 ;
      RECT  138000.0 1996950.0 139200.0 1995750.0 ;
      RECT  135600.0 1996950.0 136800.0 1995750.0 ;
      RECT  138000.0 1996950.0 139200.0 1995750.0 ;
      RECT  140400.0 1996950.0 141600.0 1995750.0 ;
      RECT  140400.0 1996950.0 141600.0 1995750.0 ;
      RECT  138000.0 1996950.0 139200.0 1995750.0 ;
      RECT  135600.0 2005650.0 136800.0 2004450.0 ;
      RECT  138000.0 2005650.0 139200.0 2004450.0 ;
      RECT  138000.0 2005650.0 139200.0 2004450.0 ;
      RECT  135600.0 2005650.0 136800.0 2004450.0 ;
      RECT  138000.0 2005650.0 139200.0 2004450.0 ;
      RECT  140400.0 2005650.0 141600.0 2004450.0 ;
      RECT  140400.0 2005650.0 141600.0 2004450.0 ;
      RECT  138000.0 2005650.0 139200.0 2004450.0 ;
      RECT  142800.0 1996350.0 144000.0 1995150.0 ;
      RECT  142800.0 2006250.0 144000.0 2005050.0 ;
      RECT  140400.0 2003100.0 139200.0 2001900.0 ;
      RECT  137400.0 2000400.0 136200.0 1999200.0 ;
      RECT  138000.0 1996950.0 139200.0 1995750.0 ;
      RECT  140400.0 2005650.0 141600.0 2004450.0 ;
      RECT  141600.0 2000400.0 140400.0 1999200.0 ;
      RECT  136200.0 2000400.0 137400.0 1999200.0 ;
      RECT  139200.0 2003100.0 140400.0 2001900.0 ;
      RECT  140400.0 2000400.0 141600.0 1999200.0 ;
      RECT  133800.0 1994250.0 148200.0 1993350.0 ;
      RECT  133800.0 2008050.0 148200.0 2007150.0 ;
      RECT  154800.0 1995750.0 156000.0 1993800.0 ;
      RECT  154800.0 2007600.0 156000.0 2005650.0 ;
      RECT  150000.0 2006250.0 151200.0 2008050.0 ;
      RECT  150000.0 1996950.0 151200.0 1993350.0 ;
      RECT  152700.0 2006250.0 153600.0 1996950.0 ;
      RECT  150000.0 1996950.0 151200.0 1995750.0 ;
      RECT  152400.0 1996950.0 153600.0 1995750.0 ;
      RECT  152400.0 1996950.0 153600.0 1995750.0 ;
      RECT  150000.0 1996950.0 151200.0 1995750.0 ;
      RECT  150000.0 2006250.0 151200.0 2005050.0 ;
      RECT  152400.0 2006250.0 153600.0 2005050.0 ;
      RECT  152400.0 2006250.0 153600.0 2005050.0 ;
      RECT  150000.0 2006250.0 151200.0 2005050.0 ;
      RECT  154800.0 1996350.0 156000.0 1995150.0 ;
      RECT  154800.0 2006250.0 156000.0 2005050.0 ;
      RECT  150600.0 2001600.0 151800.0 2000400.0 ;
      RECT  150600.0 2001600.0 151800.0 2000400.0 ;
      RECT  153150.0 2001450.0 154050.0 2000550.0 ;
      RECT  148200.0 1994250.0 157800.0 1993350.0 ;
      RECT  148200.0 2008050.0 157800.0 2007150.0 ;
      RECT  120450.0 2000400.0 121650.0 2001600.0 ;
      RECT  122400.0 2002800.0 123600.0 2004000.0 ;
      RECT  139200.0 2001900.0 138000.0 2003100.0 ;
      RECT  130800.0 2019450.0 132000.0 2021400.0 ;
      RECT  130800.0 2007600.0 132000.0 2009550.0 ;
      RECT  126000.0 2008950.0 127200.0 2007150.0 ;
      RECT  126000.0 2018250.0 127200.0 2021850.0 ;
      RECT  128700.0 2008950.0 129600.0 2018250.0 ;
      RECT  126000.0 2018250.0 127200.0 2019450.0 ;
      RECT  128400.0 2018250.0 129600.0 2019450.0 ;
      RECT  128400.0 2018250.0 129600.0 2019450.0 ;
      RECT  126000.0 2018250.0 127200.0 2019450.0 ;
      RECT  126000.0 2008950.0 127200.0 2010150.0 ;
      RECT  128400.0 2008950.0 129600.0 2010150.0 ;
      RECT  128400.0 2008950.0 129600.0 2010150.0 ;
      RECT  126000.0 2008950.0 127200.0 2010150.0 ;
      RECT  130800.0 2018850.0 132000.0 2020050.0 ;
      RECT  130800.0 2008950.0 132000.0 2010150.0 ;
      RECT  126600.0 2013600.0 127800.0 2014800.0 ;
      RECT  126600.0 2013600.0 127800.0 2014800.0 ;
      RECT  129150.0 2013750.0 130050.0 2014650.0 ;
      RECT  124200.0 2020950.0 133800.0 2021850.0 ;
      RECT  124200.0 2007150.0 133800.0 2008050.0 ;
      RECT  135600.0 2009550.0 136800.0 2007150.0 ;
      RECT  135600.0 2018250.0 136800.0 2021850.0 ;
      RECT  140400.0 2018250.0 141600.0 2021850.0 ;
      RECT  142800.0 2019450.0 144000.0 2021400.0 ;
      RECT  142800.0 2007600.0 144000.0 2009550.0 ;
      RECT  135600.0 2018250.0 136800.0 2019450.0 ;
      RECT  138000.0 2018250.0 139200.0 2019450.0 ;
      RECT  138000.0 2018250.0 139200.0 2019450.0 ;
      RECT  135600.0 2018250.0 136800.0 2019450.0 ;
      RECT  138000.0 2018250.0 139200.0 2019450.0 ;
      RECT  140400.0 2018250.0 141600.0 2019450.0 ;
      RECT  140400.0 2018250.0 141600.0 2019450.0 ;
      RECT  138000.0 2018250.0 139200.0 2019450.0 ;
      RECT  135600.0 2009550.0 136800.0 2010750.0 ;
      RECT  138000.0 2009550.0 139200.0 2010750.0 ;
      RECT  138000.0 2009550.0 139200.0 2010750.0 ;
      RECT  135600.0 2009550.0 136800.0 2010750.0 ;
      RECT  138000.0 2009550.0 139200.0 2010750.0 ;
      RECT  140400.0 2009550.0 141600.0 2010750.0 ;
      RECT  140400.0 2009550.0 141600.0 2010750.0 ;
      RECT  138000.0 2009550.0 139200.0 2010750.0 ;
      RECT  142800.0 2018850.0 144000.0 2020050.0 ;
      RECT  142800.0 2008950.0 144000.0 2010150.0 ;
      RECT  140400.0 2012100.0 139200.0 2013300.0 ;
      RECT  137400.0 2014800.0 136200.0 2016000.0 ;
      RECT  138000.0 2018250.0 139200.0 2019450.0 ;
      RECT  140400.0 2009550.0 141600.0 2010750.0 ;
      RECT  141600.0 2014800.0 140400.0 2016000.0 ;
      RECT  136200.0 2014800.0 137400.0 2016000.0 ;
      RECT  139200.0 2012100.0 140400.0 2013300.0 ;
      RECT  140400.0 2014800.0 141600.0 2016000.0 ;
      RECT  133800.0 2020950.0 148200.0 2021850.0 ;
      RECT  133800.0 2007150.0 148200.0 2008050.0 ;
      RECT  154800.0 2019450.0 156000.0 2021400.0 ;
      RECT  154800.0 2007600.0 156000.0 2009550.0 ;
      RECT  150000.0 2008950.0 151200.0 2007150.0 ;
      RECT  150000.0 2018250.0 151200.0 2021850.0 ;
      RECT  152700.0 2008950.0 153600.0 2018250.0 ;
      RECT  150000.0 2018250.0 151200.0 2019450.0 ;
      RECT  152400.0 2018250.0 153600.0 2019450.0 ;
      RECT  152400.0 2018250.0 153600.0 2019450.0 ;
      RECT  150000.0 2018250.0 151200.0 2019450.0 ;
      RECT  150000.0 2008950.0 151200.0 2010150.0 ;
      RECT  152400.0 2008950.0 153600.0 2010150.0 ;
      RECT  152400.0 2008950.0 153600.0 2010150.0 ;
      RECT  150000.0 2008950.0 151200.0 2010150.0 ;
      RECT  154800.0 2018850.0 156000.0 2020050.0 ;
      RECT  154800.0 2008950.0 156000.0 2010150.0 ;
      RECT  150600.0 2013600.0 151800.0 2014800.0 ;
      RECT  150600.0 2013600.0 151800.0 2014800.0 ;
      RECT  153150.0 2013750.0 154050.0 2014650.0 ;
      RECT  148200.0 2020950.0 157800.0 2021850.0 ;
      RECT  148200.0 2007150.0 157800.0 2008050.0 ;
      RECT  120450.0 2013600.0 121650.0 2014800.0 ;
      RECT  122400.0 2011200.0 123600.0 2012400.0 ;
      RECT  139200.0 2012100.0 138000.0 2013300.0 ;
      RECT  130800.0 2023350.0 132000.0 2021400.0 ;
      RECT  130800.0 2035200.0 132000.0 2033250.0 ;
      RECT  126000.0 2033850.0 127200.0 2035650.0 ;
      RECT  126000.0 2024550.0 127200.0 2020950.0 ;
      RECT  128700.0 2033850.0 129600.0 2024550.0 ;
      RECT  126000.0 2024550.0 127200.0 2023350.0 ;
      RECT  128400.0 2024550.0 129600.0 2023350.0 ;
      RECT  128400.0 2024550.0 129600.0 2023350.0 ;
      RECT  126000.0 2024550.0 127200.0 2023350.0 ;
      RECT  126000.0 2033850.0 127200.0 2032650.0 ;
      RECT  128400.0 2033850.0 129600.0 2032650.0 ;
      RECT  128400.0 2033850.0 129600.0 2032650.0 ;
      RECT  126000.0 2033850.0 127200.0 2032650.0 ;
      RECT  130800.0 2023950.0 132000.0 2022750.0 ;
      RECT  130800.0 2033850.0 132000.0 2032650.0 ;
      RECT  126600.0 2029200.0 127800.0 2028000.0 ;
      RECT  126600.0 2029200.0 127800.0 2028000.0 ;
      RECT  129150.0 2029050.0 130050.0 2028150.0 ;
      RECT  124200.0 2021850.0 133800.0 2020950.0 ;
      RECT  124200.0 2035650.0 133800.0 2034750.0 ;
      RECT  135600.0 2033250.0 136800.0 2035650.0 ;
      RECT  135600.0 2024550.0 136800.0 2020950.0 ;
      RECT  140400.0 2024550.0 141600.0 2020950.0 ;
      RECT  142800.0 2023350.0 144000.0 2021400.0 ;
      RECT  142800.0 2035200.0 144000.0 2033250.0 ;
      RECT  135600.0 2024550.0 136800.0 2023350.0 ;
      RECT  138000.0 2024550.0 139200.0 2023350.0 ;
      RECT  138000.0 2024550.0 139200.0 2023350.0 ;
      RECT  135600.0 2024550.0 136800.0 2023350.0 ;
      RECT  138000.0 2024550.0 139200.0 2023350.0 ;
      RECT  140400.0 2024550.0 141600.0 2023350.0 ;
      RECT  140400.0 2024550.0 141600.0 2023350.0 ;
      RECT  138000.0 2024550.0 139200.0 2023350.0 ;
      RECT  135600.0 2033250.0 136800.0 2032050.0 ;
      RECT  138000.0 2033250.0 139200.0 2032050.0 ;
      RECT  138000.0 2033250.0 139200.0 2032050.0 ;
      RECT  135600.0 2033250.0 136800.0 2032050.0 ;
      RECT  138000.0 2033250.0 139200.0 2032050.0 ;
      RECT  140400.0 2033250.0 141600.0 2032050.0 ;
      RECT  140400.0 2033250.0 141600.0 2032050.0 ;
      RECT  138000.0 2033250.0 139200.0 2032050.0 ;
      RECT  142800.0 2023950.0 144000.0 2022750.0 ;
      RECT  142800.0 2033850.0 144000.0 2032650.0 ;
      RECT  140400.0 2030700.0 139200.0 2029500.0 ;
      RECT  137400.0 2028000.0 136200.0 2026800.0 ;
      RECT  138000.0 2024550.0 139200.0 2023350.0 ;
      RECT  140400.0 2033250.0 141600.0 2032050.0 ;
      RECT  141600.0 2028000.0 140400.0 2026800.0 ;
      RECT  136200.0 2028000.0 137400.0 2026800.0 ;
      RECT  139200.0 2030700.0 140400.0 2029500.0 ;
      RECT  140400.0 2028000.0 141600.0 2026800.0 ;
      RECT  133800.0 2021850.0 148200.0 2020950.0 ;
      RECT  133800.0 2035650.0 148200.0 2034750.0 ;
      RECT  154800.0 2023350.0 156000.0 2021400.0 ;
      RECT  154800.0 2035200.0 156000.0 2033250.0 ;
      RECT  150000.0 2033850.0 151200.0 2035650.0 ;
      RECT  150000.0 2024550.0 151200.0 2020950.0 ;
      RECT  152700.0 2033850.0 153600.0 2024550.0 ;
      RECT  150000.0 2024550.0 151200.0 2023350.0 ;
      RECT  152400.0 2024550.0 153600.0 2023350.0 ;
      RECT  152400.0 2024550.0 153600.0 2023350.0 ;
      RECT  150000.0 2024550.0 151200.0 2023350.0 ;
      RECT  150000.0 2033850.0 151200.0 2032650.0 ;
      RECT  152400.0 2033850.0 153600.0 2032650.0 ;
      RECT  152400.0 2033850.0 153600.0 2032650.0 ;
      RECT  150000.0 2033850.0 151200.0 2032650.0 ;
      RECT  154800.0 2023950.0 156000.0 2022750.0 ;
      RECT  154800.0 2033850.0 156000.0 2032650.0 ;
      RECT  150600.0 2029200.0 151800.0 2028000.0 ;
      RECT  150600.0 2029200.0 151800.0 2028000.0 ;
      RECT  153150.0 2029050.0 154050.0 2028150.0 ;
      RECT  148200.0 2021850.0 157800.0 2020950.0 ;
      RECT  148200.0 2035650.0 157800.0 2034750.0 ;
      RECT  120450.0 2028000.0 121650.0 2029200.0 ;
      RECT  122400.0 2030400.0 123600.0 2031600.0 ;
      RECT  139200.0 2029500.0 138000.0 2030700.0 ;
      RECT  130800.0 2047050.0 132000.0 2049000.0 ;
      RECT  130800.0 2035200.0 132000.0 2037150.0 ;
      RECT  126000.0 2036550.0 127200.0 2034750.0 ;
      RECT  126000.0 2045850.0 127200.0 2049450.0 ;
      RECT  128700.0 2036550.0 129600.0 2045850.0 ;
      RECT  126000.0 2045850.0 127200.0 2047050.0 ;
      RECT  128400.0 2045850.0 129600.0 2047050.0 ;
      RECT  128400.0 2045850.0 129600.0 2047050.0 ;
      RECT  126000.0 2045850.0 127200.0 2047050.0 ;
      RECT  126000.0 2036550.0 127200.0 2037750.0 ;
      RECT  128400.0 2036550.0 129600.0 2037750.0 ;
      RECT  128400.0 2036550.0 129600.0 2037750.0 ;
      RECT  126000.0 2036550.0 127200.0 2037750.0 ;
      RECT  130800.0 2046450.0 132000.0 2047650.0 ;
      RECT  130800.0 2036550.0 132000.0 2037750.0 ;
      RECT  126600.0 2041200.0 127800.0 2042400.0 ;
      RECT  126600.0 2041200.0 127800.0 2042400.0 ;
      RECT  129150.0 2041350.0 130050.0 2042250.0 ;
      RECT  124200.0 2048550.0 133800.0 2049450.0 ;
      RECT  124200.0 2034750.0 133800.0 2035650.0 ;
      RECT  135600.0 2037150.0 136800.0 2034750.0 ;
      RECT  135600.0 2045850.0 136800.0 2049450.0 ;
      RECT  140400.0 2045850.0 141600.0 2049450.0 ;
      RECT  142800.0 2047050.0 144000.0 2049000.0 ;
      RECT  142800.0 2035200.0 144000.0 2037150.0 ;
      RECT  135600.0 2045850.0 136800.0 2047050.0 ;
      RECT  138000.0 2045850.0 139200.0 2047050.0 ;
      RECT  138000.0 2045850.0 139200.0 2047050.0 ;
      RECT  135600.0 2045850.0 136800.0 2047050.0 ;
      RECT  138000.0 2045850.0 139200.0 2047050.0 ;
      RECT  140400.0 2045850.0 141600.0 2047050.0 ;
      RECT  140400.0 2045850.0 141600.0 2047050.0 ;
      RECT  138000.0 2045850.0 139200.0 2047050.0 ;
      RECT  135600.0 2037150.0 136800.0 2038350.0 ;
      RECT  138000.0 2037150.0 139200.0 2038350.0 ;
      RECT  138000.0 2037150.0 139200.0 2038350.0 ;
      RECT  135600.0 2037150.0 136800.0 2038350.0 ;
      RECT  138000.0 2037150.0 139200.0 2038350.0 ;
      RECT  140400.0 2037150.0 141600.0 2038350.0 ;
      RECT  140400.0 2037150.0 141600.0 2038350.0 ;
      RECT  138000.0 2037150.0 139200.0 2038350.0 ;
      RECT  142800.0 2046450.0 144000.0 2047650.0 ;
      RECT  142800.0 2036550.0 144000.0 2037750.0 ;
      RECT  140400.0 2039700.0 139200.0 2040900.0 ;
      RECT  137400.0 2042400.0 136200.0 2043600.0 ;
      RECT  138000.0 2045850.0 139200.0 2047050.0 ;
      RECT  140400.0 2037150.0 141600.0 2038350.0 ;
      RECT  141600.0 2042400.0 140400.0 2043600.0 ;
      RECT  136200.0 2042400.0 137400.0 2043600.0 ;
      RECT  139200.0 2039700.0 140400.0 2040900.0 ;
      RECT  140400.0 2042400.0 141600.0 2043600.0 ;
      RECT  133800.0 2048550.0 148200.0 2049450.0 ;
      RECT  133800.0 2034750.0 148200.0 2035650.0 ;
      RECT  154800.0 2047050.0 156000.0 2049000.0 ;
      RECT  154800.0 2035200.0 156000.0 2037150.0 ;
      RECT  150000.0 2036550.0 151200.0 2034750.0 ;
      RECT  150000.0 2045850.0 151200.0 2049450.0 ;
      RECT  152700.0 2036550.0 153600.0 2045850.0 ;
      RECT  150000.0 2045850.0 151200.0 2047050.0 ;
      RECT  152400.0 2045850.0 153600.0 2047050.0 ;
      RECT  152400.0 2045850.0 153600.0 2047050.0 ;
      RECT  150000.0 2045850.0 151200.0 2047050.0 ;
      RECT  150000.0 2036550.0 151200.0 2037750.0 ;
      RECT  152400.0 2036550.0 153600.0 2037750.0 ;
      RECT  152400.0 2036550.0 153600.0 2037750.0 ;
      RECT  150000.0 2036550.0 151200.0 2037750.0 ;
      RECT  154800.0 2046450.0 156000.0 2047650.0 ;
      RECT  154800.0 2036550.0 156000.0 2037750.0 ;
      RECT  150600.0 2041200.0 151800.0 2042400.0 ;
      RECT  150600.0 2041200.0 151800.0 2042400.0 ;
      RECT  153150.0 2041350.0 154050.0 2042250.0 ;
      RECT  148200.0 2048550.0 157800.0 2049450.0 ;
      RECT  148200.0 2034750.0 157800.0 2035650.0 ;
      RECT  120450.0 2041200.0 121650.0 2042400.0 ;
      RECT  122400.0 2038800.0 123600.0 2040000.0 ;
      RECT  139200.0 2039700.0 138000.0 2040900.0 ;
      RECT  130800.0 2050950.0 132000.0 2049000.0 ;
      RECT  130800.0 2062800.0 132000.0 2060850.0 ;
      RECT  126000.0 2061450.0 127200.0 2063250.0 ;
      RECT  126000.0 2052150.0 127200.0 2048550.0 ;
      RECT  128700.0 2061450.0 129600.0 2052150.0 ;
      RECT  126000.0 2052150.0 127200.0 2050950.0 ;
      RECT  128400.0 2052150.0 129600.0 2050950.0 ;
      RECT  128400.0 2052150.0 129600.0 2050950.0 ;
      RECT  126000.0 2052150.0 127200.0 2050950.0 ;
      RECT  126000.0 2061450.0 127200.0 2060250.0 ;
      RECT  128400.0 2061450.0 129600.0 2060250.0 ;
      RECT  128400.0 2061450.0 129600.0 2060250.0 ;
      RECT  126000.0 2061450.0 127200.0 2060250.0 ;
      RECT  130800.0 2051550.0 132000.0 2050350.0 ;
      RECT  130800.0 2061450.0 132000.0 2060250.0 ;
      RECT  126600.0 2056800.0 127800.0 2055600.0 ;
      RECT  126600.0 2056800.0 127800.0 2055600.0 ;
      RECT  129150.0 2056650.0 130050.0 2055750.0 ;
      RECT  124200.0 2049450.0 133800.0 2048550.0 ;
      RECT  124200.0 2063250.0 133800.0 2062350.0 ;
      RECT  135600.0 2060850.0 136800.0 2063250.0 ;
      RECT  135600.0 2052150.0 136800.0 2048550.0 ;
      RECT  140400.0 2052150.0 141600.0 2048550.0 ;
      RECT  142800.0 2050950.0 144000.0 2049000.0 ;
      RECT  142800.0 2062800.0 144000.0 2060850.0 ;
      RECT  135600.0 2052150.0 136800.0 2050950.0 ;
      RECT  138000.0 2052150.0 139200.0 2050950.0 ;
      RECT  138000.0 2052150.0 139200.0 2050950.0 ;
      RECT  135600.0 2052150.0 136800.0 2050950.0 ;
      RECT  138000.0 2052150.0 139200.0 2050950.0 ;
      RECT  140400.0 2052150.0 141600.0 2050950.0 ;
      RECT  140400.0 2052150.0 141600.0 2050950.0 ;
      RECT  138000.0 2052150.0 139200.0 2050950.0 ;
      RECT  135600.0 2060850.0 136800.0 2059650.0 ;
      RECT  138000.0 2060850.0 139200.0 2059650.0 ;
      RECT  138000.0 2060850.0 139200.0 2059650.0 ;
      RECT  135600.0 2060850.0 136800.0 2059650.0 ;
      RECT  138000.0 2060850.0 139200.0 2059650.0 ;
      RECT  140400.0 2060850.0 141600.0 2059650.0 ;
      RECT  140400.0 2060850.0 141600.0 2059650.0 ;
      RECT  138000.0 2060850.0 139200.0 2059650.0 ;
      RECT  142800.0 2051550.0 144000.0 2050350.0 ;
      RECT  142800.0 2061450.0 144000.0 2060250.0 ;
      RECT  140400.0 2058300.0 139200.0 2057100.0 ;
      RECT  137400.0 2055600.0 136200.0 2054400.0 ;
      RECT  138000.0 2052150.0 139200.0 2050950.0 ;
      RECT  140400.0 2060850.0 141600.0 2059650.0 ;
      RECT  141600.0 2055600.0 140400.0 2054400.0 ;
      RECT  136200.0 2055600.0 137400.0 2054400.0 ;
      RECT  139200.0 2058300.0 140400.0 2057100.0 ;
      RECT  140400.0 2055600.0 141600.0 2054400.0 ;
      RECT  133800.0 2049450.0 148200.0 2048550.0 ;
      RECT  133800.0 2063250.0 148200.0 2062350.0 ;
      RECT  154800.0 2050950.0 156000.0 2049000.0 ;
      RECT  154800.0 2062800.0 156000.0 2060850.0 ;
      RECT  150000.0 2061450.0 151200.0 2063250.0 ;
      RECT  150000.0 2052150.0 151200.0 2048550.0 ;
      RECT  152700.0 2061450.0 153600.0 2052150.0 ;
      RECT  150000.0 2052150.0 151200.0 2050950.0 ;
      RECT  152400.0 2052150.0 153600.0 2050950.0 ;
      RECT  152400.0 2052150.0 153600.0 2050950.0 ;
      RECT  150000.0 2052150.0 151200.0 2050950.0 ;
      RECT  150000.0 2061450.0 151200.0 2060250.0 ;
      RECT  152400.0 2061450.0 153600.0 2060250.0 ;
      RECT  152400.0 2061450.0 153600.0 2060250.0 ;
      RECT  150000.0 2061450.0 151200.0 2060250.0 ;
      RECT  154800.0 2051550.0 156000.0 2050350.0 ;
      RECT  154800.0 2061450.0 156000.0 2060250.0 ;
      RECT  150600.0 2056800.0 151800.0 2055600.0 ;
      RECT  150600.0 2056800.0 151800.0 2055600.0 ;
      RECT  153150.0 2056650.0 154050.0 2055750.0 ;
      RECT  148200.0 2049450.0 157800.0 2048550.0 ;
      RECT  148200.0 2063250.0 157800.0 2062350.0 ;
      RECT  120450.0 2055600.0 121650.0 2056800.0 ;
      RECT  122400.0 2058000.0 123600.0 2059200.0 ;
      RECT  139200.0 2057100.0 138000.0 2058300.0 ;
      RECT  130800.0 2074650.0 132000.0 2076600.0 ;
      RECT  130800.0 2062800.0 132000.0 2064750.0 ;
      RECT  126000.0 2064150.0 127200.0 2062350.0 ;
      RECT  126000.0 2073450.0 127200.0 2077050.0 ;
      RECT  128700.0 2064150.0 129600.0 2073450.0 ;
      RECT  126000.0 2073450.0 127200.0 2074650.0 ;
      RECT  128400.0 2073450.0 129600.0 2074650.0 ;
      RECT  128400.0 2073450.0 129600.0 2074650.0 ;
      RECT  126000.0 2073450.0 127200.0 2074650.0 ;
      RECT  126000.0 2064150.0 127200.0 2065350.0 ;
      RECT  128400.0 2064150.0 129600.0 2065350.0 ;
      RECT  128400.0 2064150.0 129600.0 2065350.0 ;
      RECT  126000.0 2064150.0 127200.0 2065350.0 ;
      RECT  130800.0 2074050.0 132000.0 2075250.0 ;
      RECT  130800.0 2064150.0 132000.0 2065350.0 ;
      RECT  126600.0 2068800.0 127800.0 2070000.0 ;
      RECT  126600.0 2068800.0 127800.0 2070000.0 ;
      RECT  129150.0 2068950.0 130050.0 2069850.0 ;
      RECT  124200.0 2076150.0 133800.0 2077050.0 ;
      RECT  124200.0 2062350.0 133800.0 2063250.0 ;
      RECT  135600.0 2064750.0 136800.0 2062350.0 ;
      RECT  135600.0 2073450.0 136800.0 2077050.0 ;
      RECT  140400.0 2073450.0 141600.0 2077050.0 ;
      RECT  142800.0 2074650.0 144000.0 2076600.0 ;
      RECT  142800.0 2062800.0 144000.0 2064750.0 ;
      RECT  135600.0 2073450.0 136800.0 2074650.0 ;
      RECT  138000.0 2073450.0 139200.0 2074650.0 ;
      RECT  138000.0 2073450.0 139200.0 2074650.0 ;
      RECT  135600.0 2073450.0 136800.0 2074650.0 ;
      RECT  138000.0 2073450.0 139200.0 2074650.0 ;
      RECT  140400.0 2073450.0 141600.0 2074650.0 ;
      RECT  140400.0 2073450.0 141600.0 2074650.0 ;
      RECT  138000.0 2073450.0 139200.0 2074650.0 ;
      RECT  135600.0 2064750.0 136800.0 2065950.0 ;
      RECT  138000.0 2064750.0 139200.0 2065950.0 ;
      RECT  138000.0 2064750.0 139200.0 2065950.0 ;
      RECT  135600.0 2064750.0 136800.0 2065950.0 ;
      RECT  138000.0 2064750.0 139200.0 2065950.0 ;
      RECT  140400.0 2064750.0 141600.0 2065950.0 ;
      RECT  140400.0 2064750.0 141600.0 2065950.0 ;
      RECT  138000.0 2064750.0 139200.0 2065950.0 ;
      RECT  142800.0 2074050.0 144000.0 2075250.0 ;
      RECT  142800.0 2064150.0 144000.0 2065350.0 ;
      RECT  140400.0 2067300.0 139200.0 2068500.0 ;
      RECT  137400.0 2070000.0 136200.0 2071200.0 ;
      RECT  138000.0 2073450.0 139200.0 2074650.0 ;
      RECT  140400.0 2064750.0 141600.0 2065950.0 ;
      RECT  141600.0 2070000.0 140400.0 2071200.0 ;
      RECT  136200.0 2070000.0 137400.0 2071200.0 ;
      RECT  139200.0 2067300.0 140400.0 2068500.0 ;
      RECT  140400.0 2070000.0 141600.0 2071200.0 ;
      RECT  133800.0 2076150.0 148200.0 2077050.0 ;
      RECT  133800.0 2062350.0 148200.0 2063250.0 ;
      RECT  154800.0 2074650.0 156000.0 2076600.0 ;
      RECT  154800.0 2062800.0 156000.0 2064750.0 ;
      RECT  150000.0 2064150.0 151200.0 2062350.0 ;
      RECT  150000.0 2073450.0 151200.0 2077050.0 ;
      RECT  152700.0 2064150.0 153600.0 2073450.0 ;
      RECT  150000.0 2073450.0 151200.0 2074650.0 ;
      RECT  152400.0 2073450.0 153600.0 2074650.0 ;
      RECT  152400.0 2073450.0 153600.0 2074650.0 ;
      RECT  150000.0 2073450.0 151200.0 2074650.0 ;
      RECT  150000.0 2064150.0 151200.0 2065350.0 ;
      RECT  152400.0 2064150.0 153600.0 2065350.0 ;
      RECT  152400.0 2064150.0 153600.0 2065350.0 ;
      RECT  150000.0 2064150.0 151200.0 2065350.0 ;
      RECT  154800.0 2074050.0 156000.0 2075250.0 ;
      RECT  154800.0 2064150.0 156000.0 2065350.0 ;
      RECT  150600.0 2068800.0 151800.0 2070000.0 ;
      RECT  150600.0 2068800.0 151800.0 2070000.0 ;
      RECT  153150.0 2068950.0 154050.0 2069850.0 ;
      RECT  148200.0 2076150.0 157800.0 2077050.0 ;
      RECT  148200.0 2062350.0 157800.0 2063250.0 ;
      RECT  120450.0 2068800.0 121650.0 2070000.0 ;
      RECT  122400.0 2066400.0 123600.0 2067600.0 ;
      RECT  139200.0 2067300.0 138000.0 2068500.0 ;
      RECT  130800.0 2078550.0 132000.0 2076600.0 ;
      RECT  130800.0 2090400.0 132000.0 2088450.0 ;
      RECT  126000.0 2089050.0 127200.0 2090850.0 ;
      RECT  126000.0 2079750.0 127200.0 2076150.0 ;
      RECT  128700.0 2089050.0 129600.0 2079750.0 ;
      RECT  126000.0 2079750.0 127200.0 2078550.0 ;
      RECT  128400.0 2079750.0 129600.0 2078550.0 ;
      RECT  128400.0 2079750.0 129600.0 2078550.0 ;
      RECT  126000.0 2079750.0 127200.0 2078550.0 ;
      RECT  126000.0 2089050.0 127200.0 2087850.0 ;
      RECT  128400.0 2089050.0 129600.0 2087850.0 ;
      RECT  128400.0 2089050.0 129600.0 2087850.0 ;
      RECT  126000.0 2089050.0 127200.0 2087850.0 ;
      RECT  130800.0 2079150.0 132000.0 2077950.0 ;
      RECT  130800.0 2089050.0 132000.0 2087850.0 ;
      RECT  126600.0 2084400.0 127800.0 2083200.0 ;
      RECT  126600.0 2084400.0 127800.0 2083200.0 ;
      RECT  129150.0 2084250.0 130050.0 2083350.0 ;
      RECT  124200.0 2077050.0 133800.0 2076150.0 ;
      RECT  124200.0 2090850.0 133800.0 2089950.0 ;
      RECT  135600.0 2088450.0 136800.0 2090850.0 ;
      RECT  135600.0 2079750.0 136800.0 2076150.0 ;
      RECT  140400.0 2079750.0 141600.0 2076150.0 ;
      RECT  142800.0 2078550.0 144000.0 2076600.0 ;
      RECT  142800.0 2090400.0 144000.0 2088450.0 ;
      RECT  135600.0 2079750.0 136800.0 2078550.0 ;
      RECT  138000.0 2079750.0 139200.0 2078550.0 ;
      RECT  138000.0 2079750.0 139200.0 2078550.0 ;
      RECT  135600.0 2079750.0 136800.0 2078550.0 ;
      RECT  138000.0 2079750.0 139200.0 2078550.0 ;
      RECT  140400.0 2079750.0 141600.0 2078550.0 ;
      RECT  140400.0 2079750.0 141600.0 2078550.0 ;
      RECT  138000.0 2079750.0 139200.0 2078550.0 ;
      RECT  135600.0 2088450.0 136800.0 2087250.0 ;
      RECT  138000.0 2088450.0 139200.0 2087250.0 ;
      RECT  138000.0 2088450.0 139200.0 2087250.0 ;
      RECT  135600.0 2088450.0 136800.0 2087250.0 ;
      RECT  138000.0 2088450.0 139200.0 2087250.0 ;
      RECT  140400.0 2088450.0 141600.0 2087250.0 ;
      RECT  140400.0 2088450.0 141600.0 2087250.0 ;
      RECT  138000.0 2088450.0 139200.0 2087250.0 ;
      RECT  142800.0 2079150.0 144000.0 2077950.0 ;
      RECT  142800.0 2089050.0 144000.0 2087850.0 ;
      RECT  140400.0 2085900.0 139200.0 2084700.0 ;
      RECT  137400.0 2083200.0 136200.0 2082000.0 ;
      RECT  138000.0 2079750.0 139200.0 2078550.0 ;
      RECT  140400.0 2088450.0 141600.0 2087250.0 ;
      RECT  141600.0 2083200.0 140400.0 2082000.0 ;
      RECT  136200.0 2083200.0 137400.0 2082000.0 ;
      RECT  139200.0 2085900.0 140400.0 2084700.0 ;
      RECT  140400.0 2083200.0 141600.0 2082000.0 ;
      RECT  133800.0 2077050.0 148200.0 2076150.0 ;
      RECT  133800.0 2090850.0 148200.0 2089950.0 ;
      RECT  154800.0 2078550.0 156000.0 2076600.0 ;
      RECT  154800.0 2090400.0 156000.0 2088450.0 ;
      RECT  150000.0 2089050.0 151200.0 2090850.0 ;
      RECT  150000.0 2079750.0 151200.0 2076150.0 ;
      RECT  152700.0 2089050.0 153600.0 2079750.0 ;
      RECT  150000.0 2079750.0 151200.0 2078550.0 ;
      RECT  152400.0 2079750.0 153600.0 2078550.0 ;
      RECT  152400.0 2079750.0 153600.0 2078550.0 ;
      RECT  150000.0 2079750.0 151200.0 2078550.0 ;
      RECT  150000.0 2089050.0 151200.0 2087850.0 ;
      RECT  152400.0 2089050.0 153600.0 2087850.0 ;
      RECT  152400.0 2089050.0 153600.0 2087850.0 ;
      RECT  150000.0 2089050.0 151200.0 2087850.0 ;
      RECT  154800.0 2079150.0 156000.0 2077950.0 ;
      RECT  154800.0 2089050.0 156000.0 2087850.0 ;
      RECT  150600.0 2084400.0 151800.0 2083200.0 ;
      RECT  150600.0 2084400.0 151800.0 2083200.0 ;
      RECT  153150.0 2084250.0 154050.0 2083350.0 ;
      RECT  148200.0 2077050.0 157800.0 2076150.0 ;
      RECT  148200.0 2090850.0 157800.0 2089950.0 ;
      RECT  120450.0 2083200.0 121650.0 2084400.0 ;
      RECT  122400.0 2085600.0 123600.0 2086800.0 ;
      RECT  139200.0 2084700.0 138000.0 2085900.0 ;
      RECT  130800.0 2102250.0 132000.0 2104200.0 ;
      RECT  130800.0 2090400.0 132000.0 2092350.0 ;
      RECT  126000.0 2091750.0 127200.0 2089950.0 ;
      RECT  126000.0 2101050.0 127200.0 2104650.0 ;
      RECT  128700.0 2091750.0 129600.0 2101050.0 ;
      RECT  126000.0 2101050.0 127200.0 2102250.0 ;
      RECT  128400.0 2101050.0 129600.0 2102250.0 ;
      RECT  128400.0 2101050.0 129600.0 2102250.0 ;
      RECT  126000.0 2101050.0 127200.0 2102250.0 ;
      RECT  126000.0 2091750.0 127200.0 2092950.0 ;
      RECT  128400.0 2091750.0 129600.0 2092950.0 ;
      RECT  128400.0 2091750.0 129600.0 2092950.0 ;
      RECT  126000.0 2091750.0 127200.0 2092950.0 ;
      RECT  130800.0 2101650.0 132000.0 2102850.0 ;
      RECT  130800.0 2091750.0 132000.0 2092950.0 ;
      RECT  126600.0 2096400.0 127800.0 2097600.0 ;
      RECT  126600.0 2096400.0 127800.0 2097600.0 ;
      RECT  129150.0 2096550.0 130050.0 2097450.0 ;
      RECT  124200.0 2103750.0 133800.0 2104650.0 ;
      RECT  124200.0 2089950.0 133800.0 2090850.0 ;
      RECT  135600.0 2092350.0 136800.0 2089950.0 ;
      RECT  135600.0 2101050.0 136800.0 2104650.0 ;
      RECT  140400.0 2101050.0 141600.0 2104650.0 ;
      RECT  142800.0 2102250.0 144000.0 2104200.0 ;
      RECT  142800.0 2090400.0 144000.0 2092350.0 ;
      RECT  135600.0 2101050.0 136800.0 2102250.0 ;
      RECT  138000.0 2101050.0 139200.0 2102250.0 ;
      RECT  138000.0 2101050.0 139200.0 2102250.0 ;
      RECT  135600.0 2101050.0 136800.0 2102250.0 ;
      RECT  138000.0 2101050.0 139200.0 2102250.0 ;
      RECT  140400.0 2101050.0 141600.0 2102250.0 ;
      RECT  140400.0 2101050.0 141600.0 2102250.0 ;
      RECT  138000.0 2101050.0 139200.0 2102250.0 ;
      RECT  135600.0 2092350.0 136800.0 2093550.0 ;
      RECT  138000.0 2092350.0 139200.0 2093550.0 ;
      RECT  138000.0 2092350.0 139200.0 2093550.0 ;
      RECT  135600.0 2092350.0 136800.0 2093550.0 ;
      RECT  138000.0 2092350.0 139200.0 2093550.0 ;
      RECT  140400.0 2092350.0 141600.0 2093550.0 ;
      RECT  140400.0 2092350.0 141600.0 2093550.0 ;
      RECT  138000.0 2092350.0 139200.0 2093550.0 ;
      RECT  142800.0 2101650.0 144000.0 2102850.0 ;
      RECT  142800.0 2091750.0 144000.0 2092950.0 ;
      RECT  140400.0 2094900.0 139200.0 2096100.0 ;
      RECT  137400.0 2097600.0 136200.0 2098800.0 ;
      RECT  138000.0 2101050.0 139200.0 2102250.0 ;
      RECT  140400.0 2092350.0 141600.0 2093550.0 ;
      RECT  141600.0 2097600.0 140400.0 2098800.0 ;
      RECT  136200.0 2097600.0 137400.0 2098800.0 ;
      RECT  139200.0 2094900.0 140400.0 2096100.0 ;
      RECT  140400.0 2097600.0 141600.0 2098800.0 ;
      RECT  133800.0 2103750.0 148200.0 2104650.0 ;
      RECT  133800.0 2089950.0 148200.0 2090850.0 ;
      RECT  154800.0 2102250.0 156000.0 2104200.0 ;
      RECT  154800.0 2090400.0 156000.0 2092350.0 ;
      RECT  150000.0 2091750.0 151200.0 2089950.0 ;
      RECT  150000.0 2101050.0 151200.0 2104650.0 ;
      RECT  152700.0 2091750.0 153600.0 2101050.0 ;
      RECT  150000.0 2101050.0 151200.0 2102250.0 ;
      RECT  152400.0 2101050.0 153600.0 2102250.0 ;
      RECT  152400.0 2101050.0 153600.0 2102250.0 ;
      RECT  150000.0 2101050.0 151200.0 2102250.0 ;
      RECT  150000.0 2091750.0 151200.0 2092950.0 ;
      RECT  152400.0 2091750.0 153600.0 2092950.0 ;
      RECT  152400.0 2091750.0 153600.0 2092950.0 ;
      RECT  150000.0 2091750.0 151200.0 2092950.0 ;
      RECT  154800.0 2101650.0 156000.0 2102850.0 ;
      RECT  154800.0 2091750.0 156000.0 2092950.0 ;
      RECT  150600.0 2096400.0 151800.0 2097600.0 ;
      RECT  150600.0 2096400.0 151800.0 2097600.0 ;
      RECT  153150.0 2096550.0 154050.0 2097450.0 ;
      RECT  148200.0 2103750.0 157800.0 2104650.0 ;
      RECT  148200.0 2089950.0 157800.0 2090850.0 ;
      RECT  120450.0 2096400.0 121650.0 2097600.0 ;
      RECT  122400.0 2094000.0 123600.0 2095200.0 ;
      RECT  139200.0 2094900.0 138000.0 2096100.0 ;
      RECT  130800.0 2106150.0 132000.0 2104200.0 ;
      RECT  130800.0 2118000.0 132000.0 2116050.0 ;
      RECT  126000.0 2116650.0 127200.0 2118450.0 ;
      RECT  126000.0 2107350.0 127200.0 2103750.0 ;
      RECT  128700.0 2116650.0 129600.0 2107350.0 ;
      RECT  126000.0 2107350.0 127200.0 2106150.0 ;
      RECT  128400.0 2107350.0 129600.0 2106150.0 ;
      RECT  128400.0 2107350.0 129600.0 2106150.0 ;
      RECT  126000.0 2107350.0 127200.0 2106150.0 ;
      RECT  126000.0 2116650.0 127200.0 2115450.0 ;
      RECT  128400.0 2116650.0 129600.0 2115450.0 ;
      RECT  128400.0 2116650.0 129600.0 2115450.0 ;
      RECT  126000.0 2116650.0 127200.0 2115450.0 ;
      RECT  130800.0 2106750.0 132000.0 2105550.0 ;
      RECT  130800.0 2116650.0 132000.0 2115450.0 ;
      RECT  126600.0 2112000.0 127800.0 2110800.0 ;
      RECT  126600.0 2112000.0 127800.0 2110800.0 ;
      RECT  129150.0 2111850.0 130050.0 2110950.0 ;
      RECT  124200.0 2104650.0 133800.0 2103750.0 ;
      RECT  124200.0 2118450.0 133800.0 2117550.0 ;
      RECT  135600.0 2116050.0 136800.0 2118450.0 ;
      RECT  135600.0 2107350.0 136800.0 2103750.0 ;
      RECT  140400.0 2107350.0 141600.0 2103750.0 ;
      RECT  142800.0 2106150.0 144000.0 2104200.0 ;
      RECT  142800.0 2118000.0 144000.0 2116050.0 ;
      RECT  135600.0 2107350.0 136800.0 2106150.0 ;
      RECT  138000.0 2107350.0 139200.0 2106150.0 ;
      RECT  138000.0 2107350.0 139200.0 2106150.0 ;
      RECT  135600.0 2107350.0 136800.0 2106150.0 ;
      RECT  138000.0 2107350.0 139200.0 2106150.0 ;
      RECT  140400.0 2107350.0 141600.0 2106150.0 ;
      RECT  140400.0 2107350.0 141600.0 2106150.0 ;
      RECT  138000.0 2107350.0 139200.0 2106150.0 ;
      RECT  135600.0 2116050.0 136800.0 2114850.0 ;
      RECT  138000.0 2116050.0 139200.0 2114850.0 ;
      RECT  138000.0 2116050.0 139200.0 2114850.0 ;
      RECT  135600.0 2116050.0 136800.0 2114850.0 ;
      RECT  138000.0 2116050.0 139200.0 2114850.0 ;
      RECT  140400.0 2116050.0 141600.0 2114850.0 ;
      RECT  140400.0 2116050.0 141600.0 2114850.0 ;
      RECT  138000.0 2116050.0 139200.0 2114850.0 ;
      RECT  142800.0 2106750.0 144000.0 2105550.0 ;
      RECT  142800.0 2116650.0 144000.0 2115450.0 ;
      RECT  140400.0 2113500.0 139200.0 2112300.0 ;
      RECT  137400.0 2110800.0 136200.0 2109600.0 ;
      RECT  138000.0 2107350.0 139200.0 2106150.0 ;
      RECT  140400.0 2116050.0 141600.0 2114850.0 ;
      RECT  141600.0 2110800.0 140400.0 2109600.0 ;
      RECT  136200.0 2110800.0 137400.0 2109600.0 ;
      RECT  139200.0 2113500.0 140400.0 2112300.0 ;
      RECT  140400.0 2110800.0 141600.0 2109600.0 ;
      RECT  133800.0 2104650.0 148200.0 2103750.0 ;
      RECT  133800.0 2118450.0 148200.0 2117550.0 ;
      RECT  154800.0 2106150.0 156000.0 2104200.0 ;
      RECT  154800.0 2118000.0 156000.0 2116050.0 ;
      RECT  150000.0 2116650.0 151200.0 2118450.0 ;
      RECT  150000.0 2107350.0 151200.0 2103750.0 ;
      RECT  152700.0 2116650.0 153600.0 2107350.0 ;
      RECT  150000.0 2107350.0 151200.0 2106150.0 ;
      RECT  152400.0 2107350.0 153600.0 2106150.0 ;
      RECT  152400.0 2107350.0 153600.0 2106150.0 ;
      RECT  150000.0 2107350.0 151200.0 2106150.0 ;
      RECT  150000.0 2116650.0 151200.0 2115450.0 ;
      RECT  152400.0 2116650.0 153600.0 2115450.0 ;
      RECT  152400.0 2116650.0 153600.0 2115450.0 ;
      RECT  150000.0 2116650.0 151200.0 2115450.0 ;
      RECT  154800.0 2106750.0 156000.0 2105550.0 ;
      RECT  154800.0 2116650.0 156000.0 2115450.0 ;
      RECT  150600.0 2112000.0 151800.0 2110800.0 ;
      RECT  150600.0 2112000.0 151800.0 2110800.0 ;
      RECT  153150.0 2111850.0 154050.0 2110950.0 ;
      RECT  148200.0 2104650.0 157800.0 2103750.0 ;
      RECT  148200.0 2118450.0 157800.0 2117550.0 ;
      RECT  120450.0 2110800.0 121650.0 2112000.0 ;
      RECT  122400.0 2113200.0 123600.0 2114400.0 ;
      RECT  139200.0 2112300.0 138000.0 2113500.0 ;
      RECT  130800.0 2129850.0 132000.0 2131800.0 ;
      RECT  130800.0 2118000.0 132000.0 2119950.0 ;
      RECT  126000.0 2119350.0 127200.0 2117550.0 ;
      RECT  126000.0 2128650.0 127200.0 2132250.0 ;
      RECT  128700.0 2119350.0 129600.0 2128650.0 ;
      RECT  126000.0 2128650.0 127200.0 2129850.0 ;
      RECT  128400.0 2128650.0 129600.0 2129850.0 ;
      RECT  128400.0 2128650.0 129600.0 2129850.0 ;
      RECT  126000.0 2128650.0 127200.0 2129850.0 ;
      RECT  126000.0 2119350.0 127200.0 2120550.0 ;
      RECT  128400.0 2119350.0 129600.0 2120550.0 ;
      RECT  128400.0 2119350.0 129600.0 2120550.0 ;
      RECT  126000.0 2119350.0 127200.0 2120550.0 ;
      RECT  130800.0 2129250.0 132000.0 2130450.0 ;
      RECT  130800.0 2119350.0 132000.0 2120550.0 ;
      RECT  126600.0 2124000.0 127800.0 2125200.0 ;
      RECT  126600.0 2124000.0 127800.0 2125200.0 ;
      RECT  129150.0 2124150.0 130050.0 2125050.0 ;
      RECT  124200.0 2131350.0 133800.0 2132250.0 ;
      RECT  124200.0 2117550.0 133800.0 2118450.0 ;
      RECT  135600.0 2119950.0 136800.0 2117550.0 ;
      RECT  135600.0 2128650.0 136800.0 2132250.0 ;
      RECT  140400.0 2128650.0 141600.0 2132250.0 ;
      RECT  142800.0 2129850.0 144000.0 2131800.0 ;
      RECT  142800.0 2118000.0 144000.0 2119950.0 ;
      RECT  135600.0 2128650.0 136800.0 2129850.0 ;
      RECT  138000.0 2128650.0 139200.0 2129850.0 ;
      RECT  138000.0 2128650.0 139200.0 2129850.0 ;
      RECT  135600.0 2128650.0 136800.0 2129850.0 ;
      RECT  138000.0 2128650.0 139200.0 2129850.0 ;
      RECT  140400.0 2128650.0 141600.0 2129850.0 ;
      RECT  140400.0 2128650.0 141600.0 2129850.0 ;
      RECT  138000.0 2128650.0 139200.0 2129850.0 ;
      RECT  135600.0 2119950.0 136800.0 2121150.0 ;
      RECT  138000.0 2119950.0 139200.0 2121150.0 ;
      RECT  138000.0 2119950.0 139200.0 2121150.0 ;
      RECT  135600.0 2119950.0 136800.0 2121150.0 ;
      RECT  138000.0 2119950.0 139200.0 2121150.0 ;
      RECT  140400.0 2119950.0 141600.0 2121150.0 ;
      RECT  140400.0 2119950.0 141600.0 2121150.0 ;
      RECT  138000.0 2119950.0 139200.0 2121150.0 ;
      RECT  142800.0 2129250.0 144000.0 2130450.0 ;
      RECT  142800.0 2119350.0 144000.0 2120550.0 ;
      RECT  140400.0 2122500.0 139200.0 2123700.0 ;
      RECT  137400.0 2125200.0 136200.0 2126400.0 ;
      RECT  138000.0 2128650.0 139200.0 2129850.0 ;
      RECT  140400.0 2119950.0 141600.0 2121150.0 ;
      RECT  141600.0 2125200.0 140400.0 2126400.0 ;
      RECT  136200.0 2125200.0 137400.0 2126400.0 ;
      RECT  139200.0 2122500.0 140400.0 2123700.0 ;
      RECT  140400.0 2125200.0 141600.0 2126400.0 ;
      RECT  133800.0 2131350.0 148200.0 2132250.0 ;
      RECT  133800.0 2117550.0 148200.0 2118450.0 ;
      RECT  154800.0 2129850.0 156000.0 2131800.0 ;
      RECT  154800.0 2118000.0 156000.0 2119950.0 ;
      RECT  150000.0 2119350.0 151200.0 2117550.0 ;
      RECT  150000.0 2128650.0 151200.0 2132250.0 ;
      RECT  152700.0 2119350.0 153600.0 2128650.0 ;
      RECT  150000.0 2128650.0 151200.0 2129850.0 ;
      RECT  152400.0 2128650.0 153600.0 2129850.0 ;
      RECT  152400.0 2128650.0 153600.0 2129850.0 ;
      RECT  150000.0 2128650.0 151200.0 2129850.0 ;
      RECT  150000.0 2119350.0 151200.0 2120550.0 ;
      RECT  152400.0 2119350.0 153600.0 2120550.0 ;
      RECT  152400.0 2119350.0 153600.0 2120550.0 ;
      RECT  150000.0 2119350.0 151200.0 2120550.0 ;
      RECT  154800.0 2129250.0 156000.0 2130450.0 ;
      RECT  154800.0 2119350.0 156000.0 2120550.0 ;
      RECT  150600.0 2124000.0 151800.0 2125200.0 ;
      RECT  150600.0 2124000.0 151800.0 2125200.0 ;
      RECT  153150.0 2124150.0 154050.0 2125050.0 ;
      RECT  148200.0 2131350.0 157800.0 2132250.0 ;
      RECT  148200.0 2117550.0 157800.0 2118450.0 ;
      RECT  120450.0 2124000.0 121650.0 2125200.0 ;
      RECT  122400.0 2121600.0 123600.0 2122800.0 ;
      RECT  139200.0 2122500.0 138000.0 2123700.0 ;
      RECT  130800.0 2133750.0 132000.0 2131800.0 ;
      RECT  130800.0 2145600.0 132000.0 2143650.0 ;
      RECT  126000.0 2144250.0 127200.0 2146050.0 ;
      RECT  126000.0 2134950.0 127200.0 2131350.0 ;
      RECT  128700.0 2144250.0 129600.0 2134950.0 ;
      RECT  126000.0 2134950.0 127200.0 2133750.0 ;
      RECT  128400.0 2134950.0 129600.0 2133750.0 ;
      RECT  128400.0 2134950.0 129600.0 2133750.0 ;
      RECT  126000.0 2134950.0 127200.0 2133750.0 ;
      RECT  126000.0 2144250.0 127200.0 2143050.0 ;
      RECT  128400.0 2144250.0 129600.0 2143050.0 ;
      RECT  128400.0 2144250.0 129600.0 2143050.0 ;
      RECT  126000.0 2144250.0 127200.0 2143050.0 ;
      RECT  130800.0 2134350.0 132000.0 2133150.0 ;
      RECT  130800.0 2144250.0 132000.0 2143050.0 ;
      RECT  126600.0 2139600.0 127800.0 2138400.0 ;
      RECT  126600.0 2139600.0 127800.0 2138400.0 ;
      RECT  129150.0 2139450.0 130050.0 2138550.0 ;
      RECT  124200.0 2132250.0 133800.0 2131350.0 ;
      RECT  124200.0 2146050.0 133800.0 2145150.0 ;
      RECT  135600.0 2143650.0 136800.0 2146050.0 ;
      RECT  135600.0 2134950.0 136800.0 2131350.0 ;
      RECT  140400.0 2134950.0 141600.0 2131350.0 ;
      RECT  142800.0 2133750.0 144000.0 2131800.0 ;
      RECT  142800.0 2145600.0 144000.0 2143650.0 ;
      RECT  135600.0 2134950.0 136800.0 2133750.0 ;
      RECT  138000.0 2134950.0 139200.0 2133750.0 ;
      RECT  138000.0 2134950.0 139200.0 2133750.0 ;
      RECT  135600.0 2134950.0 136800.0 2133750.0 ;
      RECT  138000.0 2134950.0 139200.0 2133750.0 ;
      RECT  140400.0 2134950.0 141600.0 2133750.0 ;
      RECT  140400.0 2134950.0 141600.0 2133750.0 ;
      RECT  138000.0 2134950.0 139200.0 2133750.0 ;
      RECT  135600.0 2143650.0 136800.0 2142450.0 ;
      RECT  138000.0 2143650.0 139200.0 2142450.0 ;
      RECT  138000.0 2143650.0 139200.0 2142450.0 ;
      RECT  135600.0 2143650.0 136800.0 2142450.0 ;
      RECT  138000.0 2143650.0 139200.0 2142450.0 ;
      RECT  140400.0 2143650.0 141600.0 2142450.0 ;
      RECT  140400.0 2143650.0 141600.0 2142450.0 ;
      RECT  138000.0 2143650.0 139200.0 2142450.0 ;
      RECT  142800.0 2134350.0 144000.0 2133150.0 ;
      RECT  142800.0 2144250.0 144000.0 2143050.0 ;
      RECT  140400.0 2141100.0 139200.0 2139900.0 ;
      RECT  137400.0 2138400.0 136200.0 2137200.0 ;
      RECT  138000.0 2134950.0 139200.0 2133750.0 ;
      RECT  140400.0 2143650.0 141600.0 2142450.0 ;
      RECT  141600.0 2138400.0 140400.0 2137200.0 ;
      RECT  136200.0 2138400.0 137400.0 2137200.0 ;
      RECT  139200.0 2141100.0 140400.0 2139900.0 ;
      RECT  140400.0 2138400.0 141600.0 2137200.0 ;
      RECT  133800.0 2132250.0 148200.0 2131350.0 ;
      RECT  133800.0 2146050.0 148200.0 2145150.0 ;
      RECT  154800.0 2133750.0 156000.0 2131800.0 ;
      RECT  154800.0 2145600.0 156000.0 2143650.0 ;
      RECT  150000.0 2144250.0 151200.0 2146050.0 ;
      RECT  150000.0 2134950.0 151200.0 2131350.0 ;
      RECT  152700.0 2144250.0 153600.0 2134950.0 ;
      RECT  150000.0 2134950.0 151200.0 2133750.0 ;
      RECT  152400.0 2134950.0 153600.0 2133750.0 ;
      RECT  152400.0 2134950.0 153600.0 2133750.0 ;
      RECT  150000.0 2134950.0 151200.0 2133750.0 ;
      RECT  150000.0 2144250.0 151200.0 2143050.0 ;
      RECT  152400.0 2144250.0 153600.0 2143050.0 ;
      RECT  152400.0 2144250.0 153600.0 2143050.0 ;
      RECT  150000.0 2144250.0 151200.0 2143050.0 ;
      RECT  154800.0 2134350.0 156000.0 2133150.0 ;
      RECT  154800.0 2144250.0 156000.0 2143050.0 ;
      RECT  150600.0 2139600.0 151800.0 2138400.0 ;
      RECT  150600.0 2139600.0 151800.0 2138400.0 ;
      RECT  153150.0 2139450.0 154050.0 2138550.0 ;
      RECT  148200.0 2132250.0 157800.0 2131350.0 ;
      RECT  148200.0 2146050.0 157800.0 2145150.0 ;
      RECT  120450.0 2138400.0 121650.0 2139600.0 ;
      RECT  122400.0 2140800.0 123600.0 2142000.0 ;
      RECT  139200.0 2139900.0 138000.0 2141100.0 ;
      RECT  117900.0 382950.0 123000.0 383850.0 ;
      RECT  117900.0 402150.0 123000.0 403050.0 ;
      RECT  117900.0 410550.0 123000.0 411450.0 ;
      RECT  117900.0 429750.0 123000.0 430650.0 ;
      RECT  117900.0 438150.0 123000.0 439050.0 ;
      RECT  117900.0 457350.0 123000.0 458250.0 ;
      RECT  117900.0 465750.0 123000.0 466650.0 ;
      RECT  117900.0 484950.0 123000.0 485850.0 ;
      RECT  117900.0 493350.0 123000.0 494250.0 ;
      RECT  117900.0 512550.0 123000.0 513450.0 ;
      RECT  117900.0 520950.0 123000.0 521850.0 ;
      RECT  117900.0 540150.0 123000.0 541050.0 ;
      RECT  117900.0 548550.0 123000.0 549450.0 ;
      RECT  117900.0 567750.0 123000.0 568650.0 ;
      RECT  117900.0 576150.0 123000.0 577050.0 ;
      RECT  117900.0 595350.0 123000.0 596250.0 ;
      RECT  117900.0 603750.0 123000.0 604650.0 ;
      RECT  117900.0 622950.0 123000.0 623850.0 ;
      RECT  117900.0 631350.0 123000.0 632250.0 ;
      RECT  117900.0 650550.0 123000.0 651450.0 ;
      RECT  117900.0 658950.0 123000.0 659850.0 ;
      RECT  117900.0 678150.0 123000.0 679050.0 ;
      RECT  117900.0 686550.0 123000.0 687450.0 ;
      RECT  117900.0 705750.0 123000.0 706650.0 ;
      RECT  117900.0 714150.0 123000.0 715050.0 ;
      RECT  117900.0 733350.0 123000.0 734250.0 ;
      RECT  117900.0 741750.0 123000.0 742650.0 ;
      RECT  117900.0 760950.0 123000.0 761850.0 ;
      RECT  117900.0 769350.0 123000.0 770250.0 ;
      RECT  117900.0 788550.0 123000.0 789450.0 ;
      RECT  117900.0 796950.0 123000.0 797850.0 ;
      RECT  117900.0 816150.0 123000.0 817050.0 ;
      RECT  117900.0 824550.0 123000.0 825450.0 ;
      RECT  117900.0 843750.0 123000.0 844650.0 ;
      RECT  117900.0 852150.0 123000.0 853050.0 ;
      RECT  117900.0 871350.0 123000.0 872250.0 ;
      RECT  117900.0 879750.0 123000.0 880650.0 ;
      RECT  117900.0 898950.0 123000.0 899850.0 ;
      RECT  117900.0 907350.0 123000.0 908250.0 ;
      RECT  117900.0 926550.0 123000.0 927450.0 ;
      RECT  117900.0 934950.0 123000.0 935850.0 ;
      RECT  117900.0 954150.0 123000.0 955050.0 ;
      RECT  117900.0 962550.0 123000.0 963450.0 ;
      RECT  117900.0 981750.0 123000.0 982650.0 ;
      RECT  117900.0 990150.0 123000.0 991050.0 ;
      RECT  117900.0 1009350.0 123000.0 1010250.0 ;
      RECT  117900.0 1017750.0 123000.0 1018650.0 ;
      RECT  117900.0 1036950.0 123000.0 1037850.0 ;
      RECT  117900.0 1045350.0 123000.0 1046250.0 ;
      RECT  117900.0 1064550.0 123000.0 1065450.0 ;
      RECT  117900.0 1072950.0 123000.0 1073850.0 ;
      RECT  117900.0 1092150.0 123000.0 1093050.0 ;
      RECT  117900.0 1100550.0 123000.0 1101450.0 ;
      RECT  117900.0 1119750.0 123000.0 1120650.0 ;
      RECT  117900.0 1128150.0 123000.0 1129050.0 ;
      RECT  117900.0 1147350.0 123000.0 1148250.0 ;
      RECT  117900.0 1155750.0 123000.0 1156650.0 ;
      RECT  117900.0 1174950.0 123000.0 1175850.0 ;
      RECT  117900.0 1183350.0 123000.0 1184250.0 ;
      RECT  117900.0 1202550.0 123000.0 1203450.0 ;
      RECT  117900.0 1210950.0 123000.0 1211850.0 ;
      RECT  117900.0 1230150.0 123000.0 1231050.0 ;
      RECT  117900.0 1238550.0 123000.0 1239450.0 ;
      RECT  117900.0 1257750.0 123000.0 1258650.0 ;
      RECT  117900.0 1266150.0 123000.0 1267050.0 ;
      RECT  117900.0 1285350.0 123000.0 1286250.0 ;
      RECT  117900.0 1293750.0 123000.0 1294650.0 ;
      RECT  117900.0 1312950.0 123000.0 1313850.0 ;
      RECT  117900.0 1321350.0 123000.0 1322250.0 ;
      RECT  117900.0 1340550.0 123000.0 1341450.0 ;
      RECT  117900.0 1348950.0 123000.0 1349850.0 ;
      RECT  117900.0 1368150.0 123000.0 1369050.0 ;
      RECT  117900.0 1376550.0 123000.0 1377450.0 ;
      RECT  117900.0 1395750.0 123000.0 1396650.0 ;
      RECT  117900.0 1404150.0 123000.0 1405050.0 ;
      RECT  117900.0 1423350.0 123000.0 1424250.0 ;
      RECT  117900.0 1431750.0 123000.0 1432650.0 ;
      RECT  117900.0 1450950.0 123000.0 1451850.0 ;
      RECT  117900.0 1459350.0 123000.0 1460250.0 ;
      RECT  117900.0 1478550.0 123000.0 1479450.0 ;
      RECT  117900.0 1486950.0 123000.0 1487850.0 ;
      RECT  117900.0 1506150.0 123000.0 1507050.0 ;
      RECT  117900.0 1514550.0 123000.0 1515450.0 ;
      RECT  117900.0 1533750.0 123000.0 1534650.0 ;
      RECT  117900.0 1542150.0 123000.0 1543050.0 ;
      RECT  117900.0 1561350.0 123000.0 1562250.0 ;
      RECT  117900.0 1569750.0 123000.0 1570650.0 ;
      RECT  117900.0 1588950.0 123000.0 1589850.0 ;
      RECT  117900.0 1597350.0 123000.0 1598250.0 ;
      RECT  117900.0 1616550.0 123000.0 1617450.0 ;
      RECT  117900.0 1624950.0 123000.0 1625850.0 ;
      RECT  117900.0 1644150.0 123000.0 1645050.0 ;
      RECT  117900.0 1652550.0 123000.0 1653450.0 ;
      RECT  117900.0 1671750.0 123000.0 1672650.0 ;
      RECT  117900.0 1680150.0 123000.0 1681050.0 ;
      RECT  117900.0 1699350.0 123000.0 1700250.0 ;
      RECT  117900.0 1707750.0 123000.0 1708650.0 ;
      RECT  117900.0 1726950.0 123000.0 1727850.0 ;
      RECT  117900.0 1735350.0 123000.0 1736250.0 ;
      RECT  117900.0 1754550.0 123000.0 1755450.0 ;
      RECT  117900.0 1762950.0 123000.0 1763850.0 ;
      RECT  117900.0 1782150.0 123000.0 1783050.0 ;
      RECT  117900.0 1790550.0 123000.0 1791450.0 ;
      RECT  117900.0 1809750.0 123000.0 1810650.0 ;
      RECT  117900.0 1818150.0 123000.0 1819050.0 ;
      RECT  117900.0 1837350.0 123000.0 1838250.0 ;
      RECT  117900.0 1845750.0 123000.0 1846650.0 ;
      RECT  117900.0 1864950.0 123000.0 1865850.0 ;
      RECT  117900.0 1873350.0 123000.0 1874250.0 ;
      RECT  117900.0 1892550.0 123000.0 1893450.0 ;
      RECT  117900.0 1900950.0 123000.0 1901850.0 ;
      RECT  117900.0 1920150.0 123000.0 1921050.0 ;
      RECT  117900.0 1928550.0 123000.0 1929450.0 ;
      RECT  117900.0 1947750.0 123000.0 1948650.0 ;
      RECT  117900.0 1956150.0 123000.0 1957050.0 ;
      RECT  117900.0 1975350.0 123000.0 1976250.0 ;
      RECT  117900.0 1983750.0 123000.0 1984650.0 ;
      RECT  117900.0 2002950.0 123000.0 2003850.0 ;
      RECT  117900.0 2011350.0 123000.0 2012250.0 ;
      RECT  117900.0 2030550.0 123000.0 2031450.0 ;
      RECT  117900.0 2038950.0 123000.0 2039850.0 ;
      RECT  117900.0 2058150.0 123000.0 2059050.0 ;
      RECT  117900.0 2066550.0 123000.0 2067450.0 ;
      RECT  117900.0 2085750.0 123000.0 2086650.0 ;
      RECT  117900.0 2094150.0 123000.0 2095050.0 ;
      RECT  117900.0 2113350.0 123000.0 2114250.0 ;
      RECT  117900.0 2121750.0 123000.0 2122650.0 ;
      RECT  117900.0 2140950.0 123000.0 2141850.0 ;
      RECT  153150.0 385350.0 154050.0 386250.0 ;
      RECT  153150.0 399750.0 154050.0 400650.0 ;
      RECT  153150.0 412950.0 154050.0 413850.0 ;
      RECT  153150.0 427350.0 154050.0 428250.0 ;
      RECT  153150.0 440550.0 154050.0 441450.0 ;
      RECT  153150.0 454950.0 154050.0 455850.0 ;
      RECT  153150.0 468150.0 154050.0 469050.0 ;
      RECT  153150.0 482550.0 154050.0 483450.0 ;
      RECT  153150.0 495750.0 154050.0 496650.0 ;
      RECT  153150.0 510150.0 154050.0 511050.0 ;
      RECT  153150.0 523350.0 154050.0 524250.0 ;
      RECT  153150.0 537750.0 154050.0 538650.0 ;
      RECT  153150.0 550950.0 154050.0 551850.0 ;
      RECT  153150.0 565350.0 154050.0 566250.0 ;
      RECT  153150.0 578550.0 154050.0 579450.0 ;
      RECT  153150.0 592950.0 154050.0 593850.0 ;
      RECT  153150.0 606150.0 154050.0 607050.0 ;
      RECT  153150.0 620550.0 154050.0 621450.0 ;
      RECT  153150.0 633750.0 154050.0 634650.0 ;
      RECT  153150.0 648150.0 154050.0 649050.0 ;
      RECT  153150.0 661350.0 154050.0 662250.0 ;
      RECT  153150.0 675750.0 154050.0 676650.0 ;
      RECT  153150.0 688950.0 154050.0 689850.0 ;
      RECT  153150.0 703350.0 154050.0 704250.0 ;
      RECT  153150.0 716550.0 154050.0 717450.0 ;
      RECT  153150.0 730950.0 154050.0 731850.0 ;
      RECT  153150.0 744150.0 154050.0 745050.0 ;
      RECT  153150.0 758550.0 154050.0 759450.0 ;
      RECT  153150.0 771750.0 154050.0 772650.0 ;
      RECT  153150.0 786150.0 154050.0 787050.0 ;
      RECT  153150.0 799350.0 154050.0 800250.0 ;
      RECT  153150.0 813750.0 154050.0 814650.0 ;
      RECT  153150.0 826950.0 154050.0 827850.0 ;
      RECT  153150.0 841350.0 154050.0 842250.0 ;
      RECT  153150.0 854550.0 154050.0 855450.0 ;
      RECT  153150.0 868950.0 154050.0 869850.0 ;
      RECT  153150.0 882150.0 154050.0 883050.0 ;
      RECT  153150.0 896550.0 154050.0 897450.0 ;
      RECT  153150.0 909750.0 154050.0 910650.0 ;
      RECT  153150.0 924150.0 154050.0 925050.0 ;
      RECT  153150.0 937350.0 154050.0 938250.0 ;
      RECT  153150.0 951750.0 154050.0 952650.0 ;
      RECT  153150.0 964950.0 154050.0 965850.0 ;
      RECT  153150.0 979350.0 154050.0 980250.0 ;
      RECT  153150.0 992550.0 154050.0 993450.0 ;
      RECT  153150.0 1006950.0 154050.0 1007850.0 ;
      RECT  153150.0 1020150.0 154050.0 1021050.0 ;
      RECT  153150.0 1034550.0 154050.0 1035450.0 ;
      RECT  153150.0 1047750.0 154050.0 1048650.0 ;
      RECT  153150.0 1062150.0 154050.0 1063050.0 ;
      RECT  153150.0 1075350.0 154050.0 1076250.0 ;
      RECT  153150.0 1089750.0 154050.0 1090650.0 ;
      RECT  153150.0 1102950.0 154050.0 1103850.0 ;
      RECT  153150.0 1117350.0 154050.0 1118250.0 ;
      RECT  153150.0 1130550.0 154050.0 1131450.0 ;
      RECT  153150.0 1144950.0 154050.0 1145850.0 ;
      RECT  153150.0 1158150.0 154050.0 1159050.0 ;
      RECT  153150.0 1172550.0 154050.0 1173450.0 ;
      RECT  153150.0 1185750.0 154050.0 1186650.0 ;
      RECT  153150.0 1200150.0 154050.0 1201050.0 ;
      RECT  153150.0 1213350.0 154050.0 1214250.0 ;
      RECT  153150.0 1227750.0 154050.0 1228650.0 ;
      RECT  153150.0 1240950.0 154050.0 1241850.0 ;
      RECT  153150.0 1255350.0 154050.0 1256250.0 ;
      RECT  153150.0 1268550.0 154050.0 1269450.0 ;
      RECT  153150.0 1282950.0 154050.0 1283850.0 ;
      RECT  153150.0 1296150.0 154050.0 1297050.0 ;
      RECT  153150.0 1310550.0 154050.0 1311450.0 ;
      RECT  153150.0 1323750.0 154050.0 1324650.0 ;
      RECT  153150.0 1338150.0 154050.0 1339050.0 ;
      RECT  153150.0 1351350.0 154050.0 1352250.0 ;
      RECT  153150.0 1365750.0 154050.0 1366650.0 ;
      RECT  153150.0 1378950.0 154050.0 1379850.0 ;
      RECT  153150.0 1393350.0 154050.0 1394250.0 ;
      RECT  153150.0 1406550.0 154050.0 1407450.0 ;
      RECT  153150.0 1420950.0 154050.0 1421850.0 ;
      RECT  153150.0 1434150.0 154050.0 1435050.0 ;
      RECT  153150.0 1448550.0 154050.0 1449450.0 ;
      RECT  153150.0 1461750.0 154050.0 1462650.0 ;
      RECT  153150.0 1476150.0 154050.0 1477050.0 ;
      RECT  153150.0 1489350.0 154050.0 1490250.0 ;
      RECT  153150.0 1503750.0 154050.0 1504650.0 ;
      RECT  153150.0 1516950.0 154050.0 1517850.0 ;
      RECT  153150.0 1531350.0 154050.0 1532250.0 ;
      RECT  153150.0 1544550.0 154050.0 1545450.0 ;
      RECT  153150.0 1558950.0 154050.0 1559850.0 ;
      RECT  153150.0 1572150.0 154050.0 1573050.0 ;
      RECT  153150.0 1586550.0 154050.0 1587450.0 ;
      RECT  153150.0 1599750.0 154050.0 1600650.0 ;
      RECT  153150.0 1614150.0 154050.0 1615050.0 ;
      RECT  153150.0 1627350.0 154050.0 1628250.0 ;
      RECT  153150.0 1641750.0 154050.0 1642650.0 ;
      RECT  153150.0 1654950.0 154050.0 1655850.0 ;
      RECT  153150.0 1669350.0 154050.0 1670250.0 ;
      RECT  153150.0 1682550.0 154050.0 1683450.0 ;
      RECT  153150.0 1696950.0 154050.0 1697850.0 ;
      RECT  153150.0 1710150.0 154050.0 1711050.0 ;
      RECT  153150.0 1724550.0 154050.0 1725450.0 ;
      RECT  153150.0 1737750.0 154050.0 1738650.0 ;
      RECT  153150.0 1752150.0 154050.0 1753050.0 ;
      RECT  153150.0 1765350.0 154050.0 1766250.0 ;
      RECT  153150.0 1779750.0 154050.0 1780650.0 ;
      RECT  153150.0 1792950.0 154050.0 1793850.0 ;
      RECT  153150.0 1807350.0 154050.0 1808250.0 ;
      RECT  153150.0 1820550.0 154050.0 1821450.0 ;
      RECT  153150.0 1834950.0 154050.0 1835850.0 ;
      RECT  153150.0 1848150.0 154050.0 1849050.0 ;
      RECT  153150.0 1862550.0 154050.0 1863450.0 ;
      RECT  153150.0 1875750.0 154050.0 1876650.0 ;
      RECT  153150.0 1890150.0 154050.0 1891050.0 ;
      RECT  153150.0 1903350.0 154050.0 1904250.0 ;
      RECT  153150.0 1917750.0 154050.0 1918650.0 ;
      RECT  153150.0 1930950.0 154050.0 1931850.0 ;
      RECT  153150.0 1945350.0 154050.0 1946250.0 ;
      RECT  153150.0 1958550.0 154050.0 1959450.0 ;
      RECT  153150.0 1972950.0 154050.0 1973850.0 ;
      RECT  153150.0 1986150.0 154050.0 1987050.0 ;
      RECT  153150.0 2000550.0 154050.0 2001450.0 ;
      RECT  153150.0 2013750.0 154050.0 2014650.0 ;
      RECT  153150.0 2028150.0 154050.0 2029050.0 ;
      RECT  153150.0 2041350.0 154050.0 2042250.0 ;
      RECT  153150.0 2055750.0 154050.0 2056650.0 ;
      RECT  153150.0 2068950.0 154050.0 2069850.0 ;
      RECT  153150.0 2083350.0 154050.0 2084250.0 ;
      RECT  153150.0 2096550.0 154050.0 2097450.0 ;
      RECT  153150.0 2110950.0 154050.0 2111850.0 ;
      RECT  153150.0 2124150.0 154050.0 2125050.0 ;
      RECT  153150.0 2138550.0 154050.0 2139450.0 ;
      RECT  117900.0 392550.0 124200.0 393450.0 ;
      RECT  117900.0 420150.0 124200.0 421050.0 ;
      RECT  117900.0 447750.0 124200.0 448650.0 ;
      RECT  117900.0 475350.0 124200.0 476250.0 ;
      RECT  117900.0 502950.0 124200.0 503850.0 ;
      RECT  117900.0 530550.0 124200.0 531450.0 ;
      RECT  117900.0 558150.0 124200.0 559050.0 ;
      RECT  117900.0 585750.0 124200.0 586650.0 ;
      RECT  117900.0 613350.0 124200.0 614250.0 ;
      RECT  117900.0 640950.0 124200.0 641850.0 ;
      RECT  117900.0 668550.0 124200.0 669450.0 ;
      RECT  117900.0 696150.0 124200.0 697050.0 ;
      RECT  117900.0 723750.0 124200.0 724650.0 ;
      RECT  117900.0 751350.0 124200.0 752250.0 ;
      RECT  117900.0 778950.0 124200.0 779850.0 ;
      RECT  117900.0 806550.0 124200.0 807450.0 ;
      RECT  117900.0 834150.0 124200.0 835050.0 ;
      RECT  117900.0 861750.0 124200.0 862650.0 ;
      RECT  117900.0 889350.0 124200.0 890250.0 ;
      RECT  117900.0 916950.0 124200.0 917850.0 ;
      RECT  117900.0 944550.0 124200.0 945450.0 ;
      RECT  117900.0 972150.0 124200.0 973050.0 ;
      RECT  117900.0 999750.0 124200.0 1000650.0 ;
      RECT  117900.0 1027350.0 124200.0 1028250.0 ;
      RECT  117900.0 1054950.0 124200.0 1055850.0 ;
      RECT  117900.0 1082550.0 124200.0 1083450.0 ;
      RECT  117900.0 1110150.0 124200.0 1111050.0 ;
      RECT  117900.0 1137750.0 124200.0 1138650.0 ;
      RECT  117900.0 1165350.0 124200.0 1166250.0 ;
      RECT  117900.0 1192950.0 124200.0 1193850.0 ;
      RECT  117900.0 1220550.0 124200.0 1221450.0 ;
      RECT  117900.0 1248150.0 124200.0 1249050.0 ;
      RECT  117900.0 1275750.0 124200.0 1276650.0 ;
      RECT  117900.0 1303350.0 124200.0 1304250.0 ;
      RECT  117900.0 1330950.0 124200.0 1331850.0 ;
      RECT  117900.0 1358550.0 124200.0 1359450.0 ;
      RECT  117900.0 1386150.0 124200.0 1387050.0 ;
      RECT  117900.0 1413750.0 124200.0 1414650.0 ;
      RECT  117900.0 1441350.0 124200.0 1442250.0 ;
      RECT  117900.0 1468950.0 124200.0 1469850.0 ;
      RECT  117900.0 1496550.0 124200.0 1497450.0 ;
      RECT  117900.0 1524150.0 124200.0 1525050.0 ;
      RECT  117900.0 1551750.0 124200.0 1552650.0 ;
      RECT  117900.0 1579350.0 124200.0 1580250.0 ;
      RECT  117900.0 1606950.0 124200.0 1607850.0 ;
      RECT  117900.0 1634550.0 124200.0 1635450.0 ;
      RECT  117900.0 1662150.0 124200.0 1663050.0 ;
      RECT  117900.0 1689750.0 124200.0 1690650.0 ;
      RECT  117900.0 1717350.0 124200.0 1718250.0 ;
      RECT  117900.0 1744950.0 124200.0 1745850.0 ;
      RECT  117900.0 1772550.0 124200.0 1773450.0 ;
      RECT  117900.0 1800150.0 124200.0 1801050.0 ;
      RECT  117900.0 1827750.0 124200.0 1828650.0 ;
      RECT  117900.0 1855350.0 124200.0 1856250.0 ;
      RECT  117900.0 1882950.0 124200.0 1883850.0 ;
      RECT  117900.0 1910550.0 124200.0 1911450.0 ;
      RECT  117900.0 1938150.0 124200.0 1939050.0 ;
      RECT  117900.0 1965750.0 124200.0 1966650.0 ;
      RECT  117900.0 1993350.0 124200.0 1994250.0 ;
      RECT  117900.0 2020950.0 124200.0 2021850.0 ;
      RECT  117900.0 2048550.0 124200.0 2049450.0 ;
      RECT  117900.0 2076150.0 124200.0 2077050.0 ;
      RECT  117900.0 2103750.0 124200.0 2104650.0 ;
      RECT  117900.0 2131350.0 124200.0 2132250.0 ;
      RECT  117900.0 378750.0 124200.0 379650.0 ;
      RECT  117900.0 406350.0 124200.0 407250.0 ;
      RECT  117900.0 433950.0 124200.0 434850.0 ;
      RECT  117900.0 461550.0 124200.0 462450.0 ;
      RECT  117900.0 489150.0 124200.0 490050.0 ;
      RECT  117900.0 516750.0 124200.0 517650.0 ;
      RECT  117900.0 544350.0 124200.0 545250.0 ;
      RECT  117900.0 571950.0 124200.0 572850.0 ;
      RECT  117900.0 599550.0 124200.0 600450.0 ;
      RECT  117900.0 627150.0 124200.0 628050.0 ;
      RECT  117900.0 654750.0 124200.0 655650.0 ;
      RECT  117900.0 682350.0 124200.0 683250.0 ;
      RECT  117900.0 709950.0 124200.0 710850.0 ;
      RECT  117900.0 737550.0 124200.0 738450.0 ;
      RECT  117900.0 765150.0 124200.0 766050.0 ;
      RECT  117900.0 792750.0 124200.0 793650.0 ;
      RECT  117900.0 820350.0 124200.0 821250.0 ;
      RECT  117900.0 847950.0 124200.0 848850.0 ;
      RECT  117900.0 875550.0 124200.0 876450.0 ;
      RECT  117900.0 903150.0 124200.0 904050.0 ;
      RECT  117900.0 930750.0 124200.0 931650.0 ;
      RECT  117900.0 958350.0 124200.0 959250.0 ;
      RECT  117900.0 985950.0 124200.0 986850.0 ;
      RECT  117900.0 1013550.0 124200.0 1014450.0 ;
      RECT  117900.0 1041150.0 124200.0 1042050.0 ;
      RECT  117900.0 1068750.0 124200.0 1069650.0 ;
      RECT  117900.0 1096350.0 124200.0 1097250.0 ;
      RECT  117900.0 1123950.0 124200.0 1124850.0 ;
      RECT  117900.0 1151550.0 124200.0 1152450.0 ;
      RECT  117900.0 1179150.0 124200.0 1180050.0 ;
      RECT  117900.0 1206750.0 124200.0 1207650.0 ;
      RECT  117900.0 1234350.0 124200.0 1235250.0 ;
      RECT  117900.0 1261950.0 124200.0 1262850.0 ;
      RECT  117900.0 1289550.0 124200.0 1290450.0 ;
      RECT  117900.0 1317150.0 124200.0 1318050.0 ;
      RECT  117900.0 1344750.0 124200.0 1345650.0 ;
      RECT  117900.0 1372350.0 124200.0 1373250.0 ;
      RECT  117900.0 1399950.0 124200.0 1400850.0 ;
      RECT  117900.0 1427550.0 124200.0 1428450.0 ;
      RECT  117900.0 1455150.0 124200.0 1456050.0 ;
      RECT  117900.0 1482750.0 124200.0 1483650.0 ;
      RECT  117900.0 1510350.0 124200.0 1511250.0 ;
      RECT  117900.0 1537950.0 124200.0 1538850.0 ;
      RECT  117900.0 1565550.0 124200.0 1566450.0 ;
      RECT  117900.0 1593150.0 124200.0 1594050.0 ;
      RECT  117900.0 1620750.0 124200.0 1621650.0 ;
      RECT  117900.0 1648350.0 124200.0 1649250.0 ;
      RECT  117900.0 1675950.0 124200.0 1676850.0 ;
      RECT  117900.0 1703550.0 124200.0 1704450.0 ;
      RECT  117900.0 1731150.0 124200.0 1732050.0 ;
      RECT  117900.0 1758750.0 124200.0 1759650.0 ;
      RECT  117900.0 1786350.0 124200.0 1787250.0 ;
      RECT  117900.0 1813950.0 124200.0 1814850.0 ;
      RECT  117900.0 1841550.0 124200.0 1842450.0 ;
      RECT  117900.0 1869150.0 124200.0 1870050.0 ;
      RECT  117900.0 1896750.0 124200.0 1897650.0 ;
      RECT  117900.0 1924350.0 124200.0 1925250.0 ;
      RECT  117900.0 1951950.0 124200.0 1952850.0 ;
      RECT  117900.0 1979550.0 124200.0 1980450.0 ;
      RECT  117900.0 2007150.0 124200.0 2008050.0 ;
      RECT  117900.0 2034750.0 124200.0 2035650.0 ;
      RECT  117900.0 2062350.0 124200.0 2063250.0 ;
      RECT  117900.0 2089950.0 124200.0 2090850.0 ;
      RECT  117900.0 2117550.0 124200.0 2118450.0 ;
      RECT  117900.0 2145150.0 124200.0 2146050.0 ;
      RECT  59100.0 153000.0 119100.0 142800.0 ;
      RECT  59100.0 132600.0 119100.0 142800.0 ;
      RECT  59100.0 132600.0 119100.0 122400.0 ;
      RECT  59100.0 112200.0 119100.0 122400.0 ;
      RECT  59100.0 112200.0 119100.0 102000.0 ;
      RECT  59100.0 91800.0 119100.0 102000.0 ;
      RECT  59100.0 91800.0 119100.0 81600.0 ;
      RECT  59100.0 71400.0 119100.0 81600.0 ;
      RECT  59100.0 71400.0 119100.0 61200.0 ;
      RECT  61500.0 153000.0 62400.0 61200.0 ;
      RECT  115500.0 153000.0 116400.0 61200.0 ;
      RECT  193950.0 379800.0 195150.0 378600.0 ;
      RECT  193950.0 407400.0 195150.0 406200.0 ;
      RECT  193950.0 435000.0 195150.0 433800.0 ;
      RECT  193950.0 462600.0 195150.0 461400.0 ;
      RECT  193950.0 490200.0 195150.0 489000.0 ;
      RECT  193950.0 517800.0 195150.0 516600.0 ;
      RECT  193950.0 545400.0 195150.0 544200.0 ;
      RECT  193950.0 573000.0 195150.0 571800.0 ;
      RECT  193950.0 600600.0 195150.0 599400.0 ;
      RECT  193950.0 628200.0 195150.0 627000.0 ;
      RECT  193950.0 655800.0 195150.0 654600.0 ;
      RECT  193950.0 683400.0 195150.0 682200.0 ;
      RECT  193950.0 711000.0 195150.0 709800.0 ;
      RECT  193950.0 738600.0 195150.0 737400.0 ;
      RECT  193950.0 766200.0 195150.0 765000.0 ;
      RECT  193950.0 793800.0 195150.0 792600.0 ;
      RECT  193950.0 821400.0 195150.0 820200.0 ;
      RECT  193950.0 849000.0 195150.0 847800.0 ;
      RECT  193950.0 876600.0 195150.0 875400.0 ;
      RECT  193950.0 904200.0 195150.0 903000.0 ;
      RECT  193950.0 931800.0 195150.0 930600.0 ;
      RECT  193950.0 959400.0 195150.0 958200.0 ;
      RECT  193950.0 987000.0 195150.0 985800.0 ;
      RECT  193950.0 1014600.0 195150.0 1013400.0 ;
      RECT  193950.0 1042200.0 195150.0 1041000.0 ;
      RECT  193950.0 1069800.0 195150.0 1068600.0 ;
      RECT  193950.0 1097400.0 195150.0 1096200.0 ;
      RECT  193950.0 1125000.0 195150.0 1123800.0 ;
      RECT  193950.0 1152600.0 195150.0 1151400.0 ;
      RECT  193950.0 1180200.0 195150.0 1179000.0 ;
      RECT  193950.0 1207800.0 195150.0 1206600.0 ;
      RECT  193950.0 1235400.0 195150.0 1234200.0 ;
      RECT  193950.0 1263000.0 195150.0 1261800.0 ;
      RECT  193950.0 1290600.0 195150.0 1289400.0 ;
      RECT  193950.0 1318200.0 195150.0 1317000.0 ;
      RECT  193950.0 1345800.0 195150.0 1344600.0 ;
      RECT  193950.0 1373400.0 195150.0 1372200.0 ;
      RECT  193950.0 1401000.0 195150.0 1399800.0 ;
      RECT  193950.0 1428600.0 195150.0 1427400.0 ;
      RECT  193950.0 1456200.0 195150.0 1455000.0 ;
      RECT  193950.0 1483800.0 195150.0 1482600.0 ;
      RECT  193950.0 1511400.0 195150.0 1510200.0 ;
      RECT  193950.0 1539000.0 195150.0 1537800.0 ;
      RECT  193950.0 1566600.0 195150.0 1565400.0 ;
      RECT  193950.0 1594200.0 195150.0 1593000.0 ;
      RECT  193950.0 1621800.0 195150.0 1620600.0 ;
      RECT  193950.0 1649400.0 195150.0 1648200.0 ;
      RECT  193950.0 1677000.0 195150.0 1675800.0 ;
      RECT  193950.0 1704600.0 195150.0 1703400.0 ;
      RECT  193950.0 1732200.0 195150.0 1731000.0 ;
      RECT  193950.0 1759800.0 195150.0 1758600.0 ;
      RECT  193950.0 1787400.0 195150.0 1786200.0 ;
      RECT  193950.0 1815000.0 195150.0 1813800.0 ;
      RECT  193950.0 1842600.0 195150.0 1841400.0 ;
      RECT  193950.0 1870200.0 195150.0 1869000.0 ;
      RECT  193950.0 1897800.0 195150.0 1896600.0 ;
      RECT  193950.0 1925400.0 195150.0 1924200.0 ;
      RECT  193950.0 1953000.0 195150.0 1951800.0 ;
      RECT  193950.0 1980600.0 195150.0 1979400.0 ;
      RECT  193950.0 2008200.0 195150.0 2007000.0 ;
      RECT  193950.0 2035800.0 195150.0 2034600.0 ;
      RECT  193950.0 2063400.0 195150.0 2062200.0 ;
      RECT  193950.0 2091000.0 195150.0 2089800.0 ;
      RECT  193950.0 2118600.0 195150.0 2117400.0 ;
      RECT  193950.0 2146200.0 195150.0 2145000.0 ;
      RECT  147300.0 160650.0 146100.0 161850.0 ;
      RECT  162600.0 160500.0 161400.0 161700.0 ;
      RECT  144300.0 174450.0 143100.0 175650.0 ;
      RECT  165300.0 174300.0 164100.0 175500.0 ;
      RECT  147300.0 215850.0 146100.0 217050.0 ;
      RECT  168000.0 215700.0 166800.0 216900.0 ;
      RECT  144300.0 229650.0 143100.0 230850.0 ;
      RECT  170700.0 229500.0 169500.0 230700.0 ;
      RECT  157500.0 271050.0 156300.0 272250.0 ;
      RECT  173400.0 270900.0 172200.0 272100.0 ;
      RECT  154500.0 284850.0 153300.0 286050.0 ;
      RECT  176100.0 284700.0 174900.0 285900.0 ;
      RECT  151500.0 298650.0 150300.0 299850.0 ;
      RECT  178800.0 298500.0 177600.0 299700.0 ;
      RECT  159600.0 157800.0 158400.0 159000.0 ;
      RECT  159600.0 185400.0 158400.0 186600.0 ;
      RECT  159600.0 213000.0 158400.0 214200.0 ;
      RECT  159600.0 240600.0 158400.0 241800.0 ;
      RECT  159600.0 268200.0 158400.0 269400.0 ;
      RECT  159600.0 295800.0 158400.0 297000.0 ;
      RECT  159600.0 323400.0 158400.0 324600.0 ;
      RECT  159600.0 351000.0 158400.0 352200.0 ;
      RECT  181500.0 351150.0 180300.0 352350.0 ;
      RECT  184200.0 349050.0 183000.0 350250.0 ;
      RECT  186900.0 346950.0 185700.0 348150.0 ;
      RECT  189600.0 344850.0 188400.0 346050.0 ;
      RECT  181500.0 6600.0 180300.0 7800.0 ;
      RECT  184200.0 21000.0 183000.0 22200.0 ;
      RECT  186900.0 34200.0 185700.0 35400.0 ;
      RECT  189600.0 48600.0 188400.0 49800.0 ;
      RECT  193950.0 1200.0 195150.0 -6.83897383169e-11 ;
      RECT  193950.0 28800.0 195150.0 27600.0 ;
      RECT  193950.0 56400.0 195150.0 55200.0 ;
      RECT  118500.0 146550.0 117300.0 147750.0 ;
      RECT  162600.0 146550.0 161400.0 147750.0 ;
      RECT  118500.0 137850.0 117300.0 139050.0 ;
      RECT  165300.0 137850.0 164100.0 139050.0 ;
      RECT  118500.0 126150.0 117300.0 127350.0 ;
      RECT  168000.0 126150.0 166800.0 127350.0 ;
      RECT  118500.0 117450.0 117300.0 118650.0 ;
      RECT  170700.0 117450.0 169500.0 118650.0 ;
      RECT  118500.0 105750.0 117300.0 106950.0 ;
      RECT  173400.0 105750.0 172200.0 106950.0 ;
      RECT  118500.0 97050.0 117300.0 98250.0 ;
      RECT  176100.0 97050.0 174900.0 98250.0 ;
      RECT  118500.0 85350.0 117300.0 86550.0 ;
      RECT  178800.0 85350.0 177600.0 86550.0 ;
      RECT  120300.0 142200.0 119100.0 143400.0 ;
      RECT  195150.0 142350.0 193950.0 143550.0 ;
      RECT  120300.0 121800.0 119100.0 123000.0 ;
      RECT  195150.0 121950.0 193950.0 123150.0 ;
      RECT  120300.0 101400.0 119100.0 102600.0 ;
      RECT  195150.0 101550.0 193950.0 102750.0 ;
      RECT  120300.0 81000.0 119100.0 82200.0 ;
      RECT  195150.0 81150.0 193950.0 82350.0 ;
      RECT  120300.0 60600.0 119100.0 61800.0 ;
      RECT  195150.0 60750.0 193950.0 61950.0 ;
      RECT  210300.0 171300.0 209100.0 172500.0 ;
      RECT  204900.0 166800.0 203700.0 168000.0 ;
      RECT  207600.0 164400.0 206400.0 165600.0 ;
      RECT  210300.0 2153850.0 209100.0 2155050.0 ;
      RECT  213000.0 236100.0 211800.0 237300.0 ;
      RECT  215700.0 334200.0 214500.0 335400.0 ;
      RECT  202200.0 154500.0 201000.0 155700.0 ;
      RECT  121650.0 2147100.0 120450.0 2148300.0 ;
      RECT  202200.0 2147100.0 201000.0 2148300.0 ;
      RECT  198450.0 162450.0 197250.0 163650.0 ;
      RECT  198450.0 332250.0 197250.0 333450.0 ;
      RECT  198450.0 234150.0 197250.0 235350.0 ;
      RECT  1529700.0 600.0 1534200.0 2166000.0 ;
      RECT  52800.0 600.0 57300.0 2166000.0 ;
      RECT  43650.0 387600.0 42750.0 397200.0 ;
      RECT  43800.0 403800.0 42900.0 404700.0 ;
      RECT  43350.0 403800.0 43200.0 404700.0 ;
      RECT  43800.0 404250.0 42900.0 411600.0 ;
      RECT  43800.0 423450.0 42900.0 430800.0 ;
      RECT  35550.0 438600.0 30600.0 439500.0 ;
      RECT  43650.0 387150.0 42750.0 388050.0 ;
      RECT  43650.0 403800.0 42750.0 404700.0 ;
      RECT  29250.0 542100.0 28350.0 555450.0 ;
      RECT  43800.0 452700.0 42900.0 464850.0 ;
      RECT  33300.0 384600.0 30600.0 385500.0 ;
      RECT  29700.0 464850.0 28800.0 491700.0 ;
      RECT  27000.0 470250.0 26100.0 494700.0 ;
      RECT  41700.0 483750.0 40800.0 492300.0 ;
      RECT  43650.0 481050.0 42750.0 494700.0 ;
      RECT  45600.0 472950.0 44700.0 497100.0 ;
      RECT  41700.0 506850.0 40800.0 507750.0 ;
      RECT  41700.0 498300.0 40800.0 507300.0 ;
      RECT  43200.0 506850.0 41250.0 507750.0 ;
      RECT  43800.0 509250.0 42900.0 510150.0 ;
      RECT  43350.0 509250.0 43200.0 510150.0 ;
      RECT  43800.0 509700.0 42900.0 567300.0 ;
      RECT  14100.0 483750.0 13200.0 501900.0 ;
      RECT  16050.0 472950.0 15150.0 504300.0 ;
      RECT  18000.0 475650.0 17100.0 506700.0 ;
      RECT  14100.0 516450.0 13200.0 517350.0 ;
      RECT  14100.0 507900.0 13200.0 516900.0 ;
      RECT  15600.0 516450.0 13650.0 517350.0 ;
      RECT  16050.0 519300.0 15150.0 526500.0 ;
      RECT  16050.0 528900.0 15150.0 536100.0 ;
      RECT  29250.0 541650.0 28350.0 542550.0 ;
      RECT  28800.0 541650.0 28350.0 542550.0 ;
      RECT  29250.0 539700.0 28350.0 542100.0 ;
      RECT  29250.0 529500.0 28350.0 536700.0 ;
      RECT  29700.0 496800.0 28800.0 503100.0 ;
      RECT  30450.0 513000.0 29550.0 520200.0 ;
      RECT  16050.0 538500.0 15150.0 542700.0 ;
      RECT  29250.0 522900.0 28350.0 527100.0 ;
      RECT  50250.0 382200.0 49350.0 542100.0 ;
      RECT  50250.0 467550.0 49350.0 488700.0 ;
      RECT  36450.0 382200.0 35550.0 542100.0 ;
      RECT  36450.0 478350.0 35550.0 488700.0 ;
      RECT  22650.0 488700.0 21750.0 542100.0 ;
      RECT  22650.0 467550.0 21750.0 488700.0 ;
      RECT  8850.0 488700.0 7950.0 542100.0 ;
      RECT  8850.0 478350.0 7950.0 488700.0 ;
      RECT  8850.0 541650.0 7950.0 542550.0 ;
      RECT  8850.0 540000.0 7950.0 542100.0 ;
      RECT  8400.0 541650.0 3600.0 542550.0 ;
      RECT  7.1054273576e-12 382200.0 10200.0 442200.0 ;
      RECT  20400.0 382200.0 10200.0 442200.0 ;
      RECT  20400.0 382200.0 30600.0 442200.0 ;
      RECT  7.1054273576e-12 384600.0 30600.0 385500.0 ;
      RECT  1.42108547152e-11 438600.0 30600.0 439500.0 ;
      RECT  37950.0 391200.0 36000.0 392400.0 ;
      RECT  49800.0 391200.0 47850.0 392400.0 ;
      RECT  48450.0 386700.0 39150.0 387600.0 ;
      RECT  38550.0 384150.0 36600.0 385050.0 ;
      RECT  38550.0 388950.0 36600.0 389850.0 ;
      RECT  39150.0 384000.0 37950.0 385200.0 ;
      RECT  39150.0 388800.0 37950.0 390000.0 ;
      RECT  39150.0 386400.0 37950.0 387600.0 ;
      RECT  39150.0 386400.0 37950.0 387600.0 ;
      RECT  37050.0 384150.0 36150.0 389850.0 ;
      RECT  49800.0 384150.0 47850.0 385050.0 ;
      RECT  49800.0 388950.0 47850.0 389850.0 ;
      RECT  48450.0 384000.0 47250.0 385200.0 ;
      RECT  48450.0 388800.0 47250.0 390000.0 ;
      RECT  48450.0 386400.0 47250.0 387600.0 ;
      RECT  48450.0 386400.0 47250.0 387600.0 ;
      RECT  50250.0 384150.0 49350.0 389850.0 ;
      RECT  38550.0 391200.0 37350.0 392400.0 ;
      RECT  48450.0 391200.0 47250.0 392400.0 ;
      RECT  43800.0 384600.0 42600.0 385800.0 ;
      RECT  43800.0 384600.0 42600.0 385800.0 ;
      RECT  43650.0 387150.0 42750.0 388050.0 ;
      RECT  36450.0 382200.0 35550.0 394200.0 ;
      RECT  50250.0 382200.0 49350.0 394200.0 ;
      RECT  37950.0 405600.0 36000.0 406800.0 ;
      RECT  49800.0 405600.0 47850.0 406800.0 ;
      RECT  37350.0 396150.0 35550.0 401850.0 ;
      RECT  46050.0 403350.0 41250.0 404250.0 ;
      RECT  38850.0 396150.0 36900.0 397050.0 ;
      RECT  38850.0 400950.0 36900.0 401850.0 ;
      RECT  40800.0 398550.0 38850.0 399450.0 ;
      RECT  40800.0 403350.0 38850.0 404250.0 ;
      RECT  39450.0 396000.0 38250.0 397200.0 ;
      RECT  39450.0 400800.0 38250.0 402000.0 ;
      RECT  39450.0 398400.0 38250.0 399600.0 ;
      RECT  39450.0 403200.0 38250.0 404400.0 ;
      RECT  41250.0 398550.0 40350.0 404250.0 ;
      RECT  37350.0 396150.0 36450.0 401850.0 ;
      RECT  49500.0 396150.0 47550.0 397050.0 ;
      RECT  49500.0 400950.0 47550.0 401850.0 ;
      RECT  47550.0 398550.0 45600.0 399450.0 ;
      RECT  47550.0 403350.0 45600.0 404250.0 ;
      RECT  48150.0 396000.0 46950.0 397200.0 ;
      RECT  48150.0 400800.0 46950.0 402000.0 ;
      RECT  48150.0 398400.0 46950.0 399600.0 ;
      RECT  48150.0 403200.0 46950.0 404400.0 ;
      RECT  46050.0 398550.0 45150.0 404250.0 ;
      RECT  49950.0 396150.0 49050.0 401850.0 ;
      RECT  38550.0 405600.0 37350.0 406800.0 ;
      RECT  48450.0 405600.0 47250.0 406800.0 ;
      RECT  43800.0 396600.0 42600.0 397800.0 ;
      RECT  43800.0 396600.0 42600.0 397800.0 ;
      RECT  43650.0 403800.0 42750.0 404700.0 ;
      RECT  36450.0 394200.0 35550.0 408600.0 ;
      RECT  50250.0 394200.0 49350.0 408600.0 ;
      RECT  37950.0 424800.0 36000.0 426000.0 ;
      RECT  49800.0 424800.0 47850.0 426000.0 ;
      RECT  37800.0 410550.0 35550.0 421050.0 ;
      RECT  45900.0 422550.0 41700.0 423450.0 ;
      RECT  39300.0 410550.0 37350.0 411450.0 ;
      RECT  39300.0 415350.0 37350.0 416250.0 ;
      RECT  39300.0 420150.0 37350.0 421050.0 ;
      RECT  41250.0 412950.0 39300.0 413850.0 ;
      RECT  41250.0 417750.0 39300.0 418650.0 ;
      RECT  41250.0 422550.0 39300.0 423450.0 ;
      RECT  39900.0 410400.0 38700.0 411600.0 ;
      RECT  39900.0 415200.0 38700.0 416400.0 ;
      RECT  39900.0 420000.0 38700.0 421200.0 ;
      RECT  39900.0 412800.0 38700.0 414000.0 ;
      RECT  39900.0 417600.0 38700.0 418800.0 ;
      RECT  39900.0 422400.0 38700.0 423600.0 ;
      RECT  41700.0 412950.0 40800.0 423450.0 ;
      RECT  37800.0 410550.0 36900.0 421050.0 ;
      RECT  49350.0 410550.0 47400.0 411450.0 ;
      RECT  49350.0 415350.0 47400.0 416250.0 ;
      RECT  49350.0 420150.0 47400.0 421050.0 ;
      RECT  47400.0 412950.0 45450.0 413850.0 ;
      RECT  47400.0 417750.0 45450.0 418650.0 ;
      RECT  47400.0 422550.0 45450.0 423450.0 ;
      RECT  48000.0 410400.0 46800.0 411600.0 ;
      RECT  48000.0 415200.0 46800.0 416400.0 ;
      RECT  48000.0 420000.0 46800.0 421200.0 ;
      RECT  48000.0 412800.0 46800.0 414000.0 ;
      RECT  48000.0 417600.0 46800.0 418800.0 ;
      RECT  48000.0 422400.0 46800.0 423600.0 ;
      RECT  45900.0 412950.0 45000.0 423450.0 ;
      RECT  49800.0 410550.0 48900.0 421050.0 ;
      RECT  38550.0 424800.0 37350.0 426000.0 ;
      RECT  48450.0 424800.0 47250.0 426000.0 ;
      RECT  43950.0 411000.0 42750.0 412200.0 ;
      RECT  43950.0 411000.0 42750.0 412200.0 ;
      RECT  43800.0 423000.0 42900.0 423900.0 ;
      RECT  36450.0 408600.0 35550.0 427800.0 ;
      RECT  50250.0 408600.0 49350.0 427800.0 ;
      RECT  37950.0 456000.0 36000.0 457200.0 ;
      RECT  49800.0 456000.0 47850.0 457200.0 ;
      RECT  37800.0 429750.0 35550.0 454650.0 ;
      RECT  45900.0 451350.0 41700.0 452250.0 ;
      RECT  39300.0 429750.0 37350.0 430650.0 ;
      RECT  39300.0 434550.0 37350.0 435450.0 ;
      RECT  39300.0 439350.0 37350.0 440250.0 ;
      RECT  39300.0 444150.0 37350.0 445050.0 ;
      RECT  39300.0 448950.0 37350.0 449850.0 ;
      RECT  39300.0 453750.0 37350.0 454650.0 ;
      RECT  41250.0 432150.0 39300.0 433050.0 ;
      RECT  41250.0 436950.0 39300.0 437850.0 ;
      RECT  41250.0 441750.0 39300.0 442650.0 ;
      RECT  41250.0 446550.0 39300.0 447450.0 ;
      RECT  41250.0 451350.0 39300.0 452250.0 ;
      RECT  39900.0 429600.0 38700.0 430800.0 ;
      RECT  39900.0 434400.0 38700.0 435600.0 ;
      RECT  39900.0 439200.0 38700.0 440400.0 ;
      RECT  39900.0 444000.0 38700.0 445200.0 ;
      RECT  39900.0 448800.0 38700.0 450000.0 ;
      RECT  39900.0 453600.0 38700.0 454800.0 ;
      RECT  39900.0 432000.0 38700.0 433200.0 ;
      RECT  39900.0 436800.0 38700.0 438000.0 ;
      RECT  39900.0 441600.0 38700.0 442800.0 ;
      RECT  39900.0 446400.0 38700.0 447600.0 ;
      RECT  39900.0 451200.0 38700.0 452400.0 ;
      RECT  41700.0 432150.0 40800.0 452250.0 ;
      RECT  37800.0 429750.0 36900.0 454650.0 ;
      RECT  49350.0 429750.0 47400.0 430650.0 ;
      RECT  49350.0 434550.0 47400.0 435450.0 ;
      RECT  49350.0 439350.0 47400.0 440250.0 ;
      RECT  49350.0 444150.0 47400.0 445050.0 ;
      RECT  49350.0 448950.0 47400.0 449850.0 ;
      RECT  49350.0 453750.0 47400.0 454650.0 ;
      RECT  47400.0 432150.0 45450.0 433050.0 ;
      RECT  47400.0 436950.0 45450.0 437850.0 ;
      RECT  47400.0 441750.0 45450.0 442650.0 ;
      RECT  47400.0 446550.0 45450.0 447450.0 ;
      RECT  47400.0 451350.0 45450.0 452250.0 ;
      RECT  48000.0 429600.0 46800.0 430800.0 ;
      RECT  48000.0 434400.0 46800.0 435600.0 ;
      RECT  48000.0 439200.0 46800.0 440400.0 ;
      RECT  48000.0 444000.0 46800.0 445200.0 ;
      RECT  48000.0 448800.0 46800.0 450000.0 ;
      RECT  48000.0 453600.0 46800.0 454800.0 ;
      RECT  48000.0 432000.0 46800.0 433200.0 ;
      RECT  48000.0 436800.0 46800.0 438000.0 ;
      RECT  48000.0 441600.0 46800.0 442800.0 ;
      RECT  48000.0 446400.0 46800.0 447600.0 ;
      RECT  48000.0 451200.0 46800.0 452400.0 ;
      RECT  45900.0 432150.0 45000.0 452250.0 ;
      RECT  49800.0 429750.0 48900.0 454650.0 ;
      RECT  38550.0 456000.0 37350.0 457200.0 ;
      RECT  48450.0 456000.0 47250.0 457200.0 ;
      RECT  43950.0 430200.0 42750.0 431400.0 ;
      RECT  43950.0 430200.0 42750.0 431400.0 ;
      RECT  43800.0 451800.0 42900.0 452700.0 ;
      RECT  36450.0 427800.0 35550.0 459000.0 ;
      RECT  50250.0 427800.0 49350.0 459000.0 ;
      RECT  47850.0 490500.0 50250.0 491700.0 ;
      RECT  39150.0 490500.0 35550.0 491700.0 ;
      RECT  39150.0 495300.0 35550.0 496500.0 ;
      RECT  37950.0 500100.0 36000.0 501300.0 ;
      RECT  49800.0 500100.0 47850.0 501300.0 ;
      RECT  39150.0 490500.0 37950.0 491700.0 ;
      RECT  39150.0 492900.0 37950.0 494100.0 ;
      RECT  39150.0 492900.0 37950.0 494100.0 ;
      RECT  39150.0 490500.0 37950.0 491700.0 ;
      RECT  39150.0 492900.0 37950.0 494100.0 ;
      RECT  39150.0 495300.0 37950.0 496500.0 ;
      RECT  39150.0 495300.0 37950.0 496500.0 ;
      RECT  39150.0 492900.0 37950.0 494100.0 ;
      RECT  39150.0 495300.0 37950.0 496500.0 ;
      RECT  39150.0 497700.0 37950.0 498900.0 ;
      RECT  39150.0 497700.0 37950.0 498900.0 ;
      RECT  39150.0 495300.0 37950.0 496500.0 ;
      RECT  47850.0 490500.0 46650.0 491700.0 ;
      RECT  47850.0 492900.0 46650.0 494100.0 ;
      RECT  47850.0 492900.0 46650.0 494100.0 ;
      RECT  47850.0 490500.0 46650.0 491700.0 ;
      RECT  47850.0 492900.0 46650.0 494100.0 ;
      RECT  47850.0 495300.0 46650.0 496500.0 ;
      RECT  47850.0 495300.0 46650.0 496500.0 ;
      RECT  47850.0 492900.0 46650.0 494100.0 ;
      RECT  47850.0 495300.0 46650.0 496500.0 ;
      RECT  47850.0 497700.0 46650.0 498900.0 ;
      RECT  47850.0 497700.0 46650.0 498900.0 ;
      RECT  47850.0 495300.0 46650.0 496500.0 ;
      RECT  38550.0 500100.0 37350.0 501300.0 ;
      RECT  48450.0 500100.0 47250.0 501300.0 ;
      RECT  45750.0 497700.0 44550.0 496500.0 ;
      RECT  43800.0 495300.0 42600.0 494100.0 ;
      RECT  41850.0 492900.0 40650.0 491700.0 ;
      RECT  39150.0 492900.0 37950.0 494100.0 ;
      RECT  39150.0 497700.0 37950.0 498900.0 ;
      RECT  47850.0 497700.0 46650.0 498900.0 ;
      RECT  41850.0 497700.0 40650.0 498900.0 ;
      RECT  41850.0 491700.0 40650.0 492900.0 ;
      RECT  43800.0 494100.0 42600.0 495300.0 ;
      RECT  45750.0 496500.0 44550.0 497700.0 ;
      RECT  41850.0 497700.0 40650.0 498900.0 ;
      RECT  36450.0 488700.0 35550.0 504300.0 ;
      RECT  50250.0 488700.0 49350.0 504300.0 ;
      RECT  37950.0 510900.0 36000.0 512100.0 ;
      RECT  49800.0 510900.0 47850.0 512100.0 ;
      RECT  48450.0 506100.0 50250.0 507300.0 ;
      RECT  39150.0 506100.0 35550.0 507300.0 ;
      RECT  48450.0 508800.0 39150.0 509700.0 ;
      RECT  39150.0 506100.0 37950.0 507300.0 ;
      RECT  39150.0 508500.0 37950.0 509700.0 ;
      RECT  39150.0 508500.0 37950.0 509700.0 ;
      RECT  39150.0 506100.0 37950.0 507300.0 ;
      RECT  48450.0 506100.0 47250.0 507300.0 ;
      RECT  48450.0 508500.0 47250.0 509700.0 ;
      RECT  48450.0 508500.0 47250.0 509700.0 ;
      RECT  48450.0 506100.0 47250.0 507300.0 ;
      RECT  38550.0 510900.0 37350.0 512100.0 ;
      RECT  48450.0 510900.0 47250.0 512100.0 ;
      RECT  43800.0 506700.0 42600.0 507900.0 ;
      RECT  43800.0 506700.0 42600.0 507900.0 ;
      RECT  43650.0 509250.0 42750.0 510150.0 ;
      RECT  36450.0 504300.0 35550.0 513900.0 ;
      RECT  50250.0 504300.0 49350.0 513900.0 ;
      RECT  23550.0 490500.0 21750.0 491700.0 ;
      RECT  23550.0 495300.0 21750.0 496500.0 ;
      RECT  32250.0 490500.0 36450.0 491700.0 ;
      RECT  34050.0 497700.0 36000.0 498900.0 ;
      RECT  22200.0 497700.0 24150.0 498900.0 ;
      RECT  32250.0 490500.0 33450.0 491700.0 ;
      RECT  32250.0 492900.0 33450.0 494100.0 ;
      RECT  32250.0 492900.0 33450.0 494100.0 ;
      RECT  32250.0 490500.0 33450.0 491700.0 ;
      RECT  32250.0 492900.0 33450.0 494100.0 ;
      RECT  32250.0 495300.0 33450.0 496500.0 ;
      RECT  32250.0 495300.0 33450.0 496500.0 ;
      RECT  32250.0 492900.0 33450.0 494100.0 ;
      RECT  23550.0 490500.0 24750.0 491700.0 ;
      RECT  23550.0 492900.0 24750.0 494100.0 ;
      RECT  23550.0 492900.0 24750.0 494100.0 ;
      RECT  23550.0 490500.0 24750.0 491700.0 ;
      RECT  23550.0 492900.0 24750.0 494100.0 ;
      RECT  23550.0 495300.0 24750.0 496500.0 ;
      RECT  23550.0 495300.0 24750.0 496500.0 ;
      RECT  23550.0 492900.0 24750.0 494100.0 ;
      RECT  33450.0 497700.0 34650.0 498900.0 ;
      RECT  23550.0 497700.0 24750.0 498900.0 ;
      RECT  25950.0 495300.0 27150.0 494100.0 ;
      RECT  28650.0 492300.0 29850.0 491100.0 ;
      RECT  32250.0 495300.0 33450.0 496500.0 ;
      RECT  23550.0 494100.0 24750.0 492900.0 ;
      RECT  28650.0 497400.0 29850.0 496200.0 ;
      RECT  28650.0 491100.0 29850.0 492300.0 ;
      RECT  25950.0 494100.0 27150.0 495300.0 ;
      RECT  28650.0 496200.0 29850.0 497400.0 ;
      RECT  35550.0 488700.0 36450.0 503100.0 ;
      RECT  21750.0 488700.0 22650.0 503100.0 ;
      RECT  24150.0 507600.0 21750.0 508800.0 ;
      RECT  32850.0 507600.0 36450.0 508800.0 ;
      RECT  32850.0 512400.0 36450.0 513600.0 ;
      RECT  34050.0 514800.0 36000.0 516000.0 ;
      RECT  22200.0 514800.0 24150.0 516000.0 ;
      RECT  32850.0 507600.0 34050.0 508800.0 ;
      RECT  32850.0 510000.0 34050.0 511200.0 ;
      RECT  32850.0 510000.0 34050.0 511200.0 ;
      RECT  32850.0 507600.0 34050.0 508800.0 ;
      RECT  32850.0 510000.0 34050.0 511200.0 ;
      RECT  32850.0 512400.0 34050.0 513600.0 ;
      RECT  32850.0 512400.0 34050.0 513600.0 ;
      RECT  32850.0 510000.0 34050.0 511200.0 ;
      RECT  24150.0 507600.0 25350.0 508800.0 ;
      RECT  24150.0 510000.0 25350.0 511200.0 ;
      RECT  24150.0 510000.0 25350.0 511200.0 ;
      RECT  24150.0 507600.0 25350.0 508800.0 ;
      RECT  24150.0 510000.0 25350.0 511200.0 ;
      RECT  24150.0 512400.0 25350.0 513600.0 ;
      RECT  24150.0 512400.0 25350.0 513600.0 ;
      RECT  24150.0 510000.0 25350.0 511200.0 ;
      RECT  33450.0 514800.0 34650.0 516000.0 ;
      RECT  23550.0 514800.0 24750.0 516000.0 ;
      RECT  26700.0 512400.0 27900.0 511200.0 ;
      RECT  29400.0 509400.0 30600.0 508200.0 ;
      RECT  32850.0 510000.0 34050.0 511200.0 ;
      RECT  24150.0 512400.0 25350.0 513600.0 ;
      RECT  29400.0 513600.0 30600.0 512400.0 ;
      RECT  29400.0 508200.0 30600.0 509400.0 ;
      RECT  26700.0 511200.0 27900.0 512400.0 ;
      RECT  29400.0 512400.0 30600.0 513600.0 ;
      RECT  35550.0 505800.0 36450.0 520200.0 ;
      RECT  21750.0 505800.0 22650.0 520200.0 ;
      RECT  34050.0 525900.0 36000.0 524700.0 ;
      RECT  22200.0 525900.0 24150.0 524700.0 ;
      RECT  23550.0 530700.0 21750.0 529500.0 ;
      RECT  32850.0 530700.0 36450.0 529500.0 ;
      RECT  23550.0 528000.0 32850.0 527100.0 ;
      RECT  32850.0 530700.0 34050.0 529500.0 ;
      RECT  32850.0 528300.0 34050.0 527100.0 ;
      RECT  32850.0 528300.0 34050.0 527100.0 ;
      RECT  32850.0 530700.0 34050.0 529500.0 ;
      RECT  23550.0 530700.0 24750.0 529500.0 ;
      RECT  23550.0 528300.0 24750.0 527100.0 ;
      RECT  23550.0 528300.0 24750.0 527100.0 ;
      RECT  23550.0 530700.0 24750.0 529500.0 ;
      RECT  33450.0 525900.0 34650.0 524700.0 ;
      RECT  23550.0 525900.0 24750.0 524700.0 ;
      RECT  28200.0 530100.0 29400.0 528900.0 ;
      RECT  28200.0 530100.0 29400.0 528900.0 ;
      RECT  28350.0 527550.0 29250.0 526650.0 ;
      RECT  35550.0 532500.0 36450.0 522900.0 ;
      RECT  21750.0 532500.0 22650.0 522900.0 ;
      RECT  34050.0 535500.0 36000.0 534300.0 ;
      RECT  22200.0 535500.0 24150.0 534300.0 ;
      RECT  23550.0 540300.0 21750.0 539100.0 ;
      RECT  32850.0 540300.0 36450.0 539100.0 ;
      RECT  23550.0 537600.0 32850.0 536700.0 ;
      RECT  32850.0 540300.0 34050.0 539100.0 ;
      RECT  32850.0 537900.0 34050.0 536700.0 ;
      RECT  32850.0 537900.0 34050.0 536700.0 ;
      RECT  32850.0 540300.0 34050.0 539100.0 ;
      RECT  23550.0 540300.0 24750.0 539100.0 ;
      RECT  23550.0 537900.0 24750.0 536700.0 ;
      RECT  23550.0 537900.0 24750.0 536700.0 ;
      RECT  23550.0 540300.0 24750.0 539100.0 ;
      RECT  33450.0 535500.0 34650.0 534300.0 ;
      RECT  23550.0 535500.0 24750.0 534300.0 ;
      RECT  28200.0 539700.0 29400.0 538500.0 ;
      RECT  28200.0 539700.0 29400.0 538500.0 ;
      RECT  28350.0 537150.0 29250.0 536250.0 ;
      RECT  35550.0 542100.0 36450.0 532500.0 ;
      RECT  21750.0 542100.0 22650.0 532500.0 ;
      RECT  20250.0 500100.0 22650.0 501300.0 ;
      RECT  11550.0 500100.0 7950.0 501300.0 ;
      RECT  11550.0 504900.0 7950.0 506100.0 ;
      RECT  10350.0 509700.0 8400.0 510900.0 ;
      RECT  22200.0 509700.0 20250.0 510900.0 ;
      RECT  11550.0 500100.0 10350.0 501300.0 ;
      RECT  11550.0 502500.0 10350.0 503700.0 ;
      RECT  11550.0 502500.0 10350.0 503700.0 ;
      RECT  11550.0 500100.0 10350.0 501300.0 ;
      RECT  11550.0 502500.0 10350.0 503700.0 ;
      RECT  11550.0 504900.0 10350.0 506100.0 ;
      RECT  11550.0 504900.0 10350.0 506100.0 ;
      RECT  11550.0 502500.0 10350.0 503700.0 ;
      RECT  11550.0 504900.0 10350.0 506100.0 ;
      RECT  11550.0 507300.0 10350.0 508500.0 ;
      RECT  11550.0 507300.0 10350.0 508500.0 ;
      RECT  11550.0 504900.0 10350.0 506100.0 ;
      RECT  20250.0 500100.0 19050.0 501300.0 ;
      RECT  20250.0 502500.0 19050.0 503700.0 ;
      RECT  20250.0 502500.0 19050.0 503700.0 ;
      RECT  20250.0 500100.0 19050.0 501300.0 ;
      RECT  20250.0 502500.0 19050.0 503700.0 ;
      RECT  20250.0 504900.0 19050.0 506100.0 ;
      RECT  20250.0 504900.0 19050.0 506100.0 ;
      RECT  20250.0 502500.0 19050.0 503700.0 ;
      RECT  20250.0 504900.0 19050.0 506100.0 ;
      RECT  20250.0 507300.0 19050.0 508500.0 ;
      RECT  20250.0 507300.0 19050.0 508500.0 ;
      RECT  20250.0 504900.0 19050.0 506100.0 ;
      RECT  10950.0 509700.0 9750.0 510900.0 ;
      RECT  20850.0 509700.0 19650.0 510900.0 ;
      RECT  18150.0 507300.0 16950.0 506100.0 ;
      RECT  16200.0 504900.0 15000.0 503700.0 ;
      RECT  14250.0 502500.0 13050.0 501300.0 ;
      RECT  11550.0 502500.0 10350.0 503700.0 ;
      RECT  11550.0 507300.0 10350.0 508500.0 ;
      RECT  20250.0 507300.0 19050.0 508500.0 ;
      RECT  14250.0 507300.0 13050.0 508500.0 ;
      RECT  14250.0 501300.0 13050.0 502500.0 ;
      RECT  16200.0 503700.0 15000.0 504900.0 ;
      RECT  18150.0 506100.0 16950.0 507300.0 ;
      RECT  14250.0 507300.0 13050.0 508500.0 ;
      RECT  8850.0 498300.0 7950.0 513900.0 ;
      RECT  22650.0 498300.0 21750.0 513900.0 ;
      RECT  10350.0 520500.0 8400.0 521700.0 ;
      RECT  22200.0 520500.0 20250.0 521700.0 ;
      RECT  20850.0 515700.0 22650.0 516900.0 ;
      RECT  11550.0 515700.0 7950.0 516900.0 ;
      RECT  20850.0 518400.0 11550.0 519300.0 ;
      RECT  11550.0 515700.0 10350.0 516900.0 ;
      RECT  11550.0 518100.0 10350.0 519300.0 ;
      RECT  11550.0 518100.0 10350.0 519300.0 ;
      RECT  11550.0 515700.0 10350.0 516900.0 ;
      RECT  20850.0 515700.0 19650.0 516900.0 ;
      RECT  20850.0 518100.0 19650.0 519300.0 ;
      RECT  20850.0 518100.0 19650.0 519300.0 ;
      RECT  20850.0 515700.0 19650.0 516900.0 ;
      RECT  10950.0 520500.0 9750.0 521700.0 ;
      RECT  20850.0 520500.0 19650.0 521700.0 ;
      RECT  16200.0 516300.0 15000.0 517500.0 ;
      RECT  16200.0 516300.0 15000.0 517500.0 ;
      RECT  16050.0 518850.0 15150.0 519750.0 ;
      RECT  8850.0 513900.0 7950.0 523500.0 ;
      RECT  22650.0 513900.0 21750.0 523500.0 ;
      RECT  10350.0 530100.0 8400.0 531300.0 ;
      RECT  22200.0 530100.0 20250.0 531300.0 ;
      RECT  20850.0 525300.0 22650.0 526500.0 ;
      RECT  11550.0 525300.0 7950.0 526500.0 ;
      RECT  20850.0 528000.0 11550.0 528900.0 ;
      RECT  11550.0 525300.0 10350.0 526500.0 ;
      RECT  11550.0 527700.0 10350.0 528900.0 ;
      RECT  11550.0 527700.0 10350.0 528900.0 ;
      RECT  11550.0 525300.0 10350.0 526500.0 ;
      RECT  20850.0 525300.0 19650.0 526500.0 ;
      RECT  20850.0 527700.0 19650.0 528900.0 ;
      RECT  20850.0 527700.0 19650.0 528900.0 ;
      RECT  20850.0 525300.0 19650.0 526500.0 ;
      RECT  10950.0 530100.0 9750.0 531300.0 ;
      RECT  20850.0 530100.0 19650.0 531300.0 ;
      RECT  16200.0 525900.0 15000.0 527100.0 ;
      RECT  16200.0 525900.0 15000.0 527100.0 ;
      RECT  16050.0 528450.0 15150.0 529350.0 ;
      RECT  8850.0 523500.0 7950.0 533100.0 ;
      RECT  22650.0 523500.0 21750.0 533100.0 ;
      RECT  10350.0 539700.0 8400.0 540900.0 ;
      RECT  22200.0 539700.0 20250.0 540900.0 ;
      RECT  20850.0 534900.0 22650.0 536100.0 ;
      RECT  11550.0 534900.0 7950.0 536100.0 ;
      RECT  20850.0 537600.0 11550.0 538500.0 ;
      RECT  11550.0 534900.0 10350.0 536100.0 ;
      RECT  11550.0 537300.0 10350.0 538500.0 ;
      RECT  11550.0 537300.0 10350.0 538500.0 ;
      RECT  11550.0 534900.0 10350.0 536100.0 ;
      RECT  20850.0 534900.0 19650.0 536100.0 ;
      RECT  20850.0 537300.0 19650.0 538500.0 ;
      RECT  20850.0 537300.0 19650.0 538500.0 ;
      RECT  20850.0 534900.0 19650.0 536100.0 ;
      RECT  10950.0 539700.0 9750.0 540900.0 ;
      RECT  20850.0 539700.0 19650.0 540900.0 ;
      RECT  16200.0 535500.0 15000.0 536700.0 ;
      RECT  16200.0 535500.0 15000.0 536700.0 ;
      RECT  16050.0 538050.0 15150.0 538950.0 ;
      RECT  8850.0 533100.0 7950.0 542700.0 ;
      RECT  22650.0 533100.0 21750.0 542700.0 ;
      RECT  22650.0 659550.0 21750.0 941100.0 ;
      RECT  21750.0 576750.0 17400.0 577650.0 ;
      RECT  21750.0 600150.0 17400.0 601050.0 ;
      RECT  21750.0 604350.0 17400.0 605250.0 ;
      RECT  21750.0 627750.0 17400.0 628650.0 ;
      RECT  21750.0 631950.0 17400.0 632850.0 ;
      RECT  21750.0 655350.0 17400.0 656250.0 ;
      RECT  21750.0 659550.0 17400.0 660450.0 ;
      RECT  21750.0 682950.0 17400.0 683850.0 ;
      RECT  21750.0 687150.0 17400.0 688050.0 ;
      RECT  21750.0 710550.0 17400.0 711450.0 ;
      RECT  21750.0 714750.0 17400.0 715650.0 ;
      RECT  21750.0 738150.0 17400.0 739050.0 ;
      RECT  21750.0 742350.0 17400.0 743250.0 ;
      RECT  21750.0 765750.0 17400.0 766650.0 ;
      RECT  21750.0 769950.0 17400.0 770850.0 ;
      RECT  21750.0 793350.0 17400.0 794250.0 ;
      RECT  21750.0 797550.0 17400.0 798450.0 ;
      RECT  21750.0 820950.0 17400.0 821850.0 ;
      RECT  21750.0 825150.0 17400.0 826050.0 ;
      RECT  21750.0 848550.0 17400.0 849450.0 ;
      RECT  21750.0 852750.0 17400.0 853650.0 ;
      RECT  21750.0 876150.0 17400.0 877050.0 ;
      RECT  21750.0 880350.0 17400.0 881250.0 ;
      RECT  21750.0 903750.0 17400.0 904650.0 ;
      RECT  21750.0 907950.0 17400.0 908850.0 ;
      RECT  21750.0 931350.0 17400.0 932250.0 ;
      RECT  22650.0 551250.0 16800.0 552150.0 ;
      RECT  16800.0 551250.0 6600.0 552150.0 ;
      RECT  4500.0 588300.0 16800.0 589200.0 ;
      RECT  4500.0 615900.0 16800.0 616800.0 ;
      RECT  4500.0 643500.0 16800.0 644400.0 ;
      RECT  4500.0 671100.0 16800.0 672000.0 ;
      RECT  4500.0 698700.0 16800.0 699600.0 ;
      RECT  4500.0 726300.0 16800.0 727200.0 ;
      RECT  4500.0 753900.0 16800.0 754800.0 ;
      RECT  4500.0 781500.0 16800.0 782400.0 ;
      RECT  4500.0 809100.0 16800.0 810000.0 ;
      RECT  4500.0 836700.0 16800.0 837600.0 ;
      RECT  4500.0 864300.0 16800.0 865200.0 ;
      RECT  4500.0 891900.0 16800.0 892800.0 ;
      RECT  4500.0 919500.0 16800.0 920400.0 ;
      RECT  4500.0 560700.0 16800.0 561600.0 ;
      RECT  29250.0 577500.0 28350.0 590100.0 ;
      RECT  29250.0 572550.0 28350.0 573450.0 ;
      RECT  29250.0 573000.0 28350.0 577500.0 ;
      RECT  28800.0 572550.0 17400.0 573450.0 ;
      RECT  36000.0 578250.0 33750.0 579150.0 ;
      RECT  33600.0 563550.0 32700.0 564450.0 ;
      RECT  29250.0 563550.0 28350.0 564450.0 ;
      RECT  33600.0 564000.0 32700.0 575700.0 ;
      RECT  33150.0 563550.0 28800.0 564450.0 ;
      RECT  29250.0 558900.0 28350.0 564000.0 ;
      RECT  28800.0 563550.0 19950.0 564450.0 ;
      RECT  19950.0 555450.0 13200.0 556350.0 ;
      RECT  29400.0 557700.0 28200.0 558900.0 ;
      RECT  29250.0 590100.0 28350.0 593850.0 ;
      RECT  34050.0 554700.0 36000.0 553500.0 ;
      RECT  22200.0 554700.0 24150.0 553500.0 ;
      RECT  23550.0 559500.0 21750.0 558300.0 ;
      RECT  32850.0 559500.0 36450.0 558300.0 ;
      RECT  23550.0 556800.0 32850.0 555900.0 ;
      RECT  32850.0 559500.0 34050.0 558300.0 ;
      RECT  32850.0 557100.0 34050.0 555900.0 ;
      RECT  32850.0 557100.0 34050.0 555900.0 ;
      RECT  32850.0 559500.0 34050.0 558300.0 ;
      RECT  23550.0 559500.0 24750.0 558300.0 ;
      RECT  23550.0 557100.0 24750.0 555900.0 ;
      RECT  23550.0 557100.0 24750.0 555900.0 ;
      RECT  23550.0 559500.0 24750.0 558300.0 ;
      RECT  33450.0 554700.0 34650.0 553500.0 ;
      RECT  23550.0 554700.0 24750.0 553500.0 ;
      RECT  28200.0 558900.0 29400.0 557700.0 ;
      RECT  28200.0 558900.0 29400.0 557700.0 ;
      RECT  28350.0 556350.0 29250.0 555450.0 ;
      RECT  35550.0 561300.0 36450.0 551700.0 ;
      RECT  21750.0 561300.0 22650.0 551700.0 ;
      RECT  32550.0 575700.0 33750.0 576900.0 ;
      RECT  32550.0 578100.0 33750.0 579300.0 ;
      RECT  32550.0 578100.0 33750.0 579300.0 ;
      RECT  32550.0 575700.0 33750.0 576900.0 ;
      RECT  21750.0 658650.0 22650.0 659550.0 ;
      RECT  49350.0 658650.0 50250.0 659550.0 ;
      RECT  21750.0 657300.0 22650.0 659100.0 ;
      RECT  22200.0 658650.0 49800.0 659550.0 ;
      RECT  49350.0 657300.0 50250.0 659100.0 ;
      RECT  37950.0 596700.0 36000.0 597900.0 ;
      RECT  49800.0 596700.0 47850.0 597900.0 ;
      RECT  48450.0 591900.0 50250.0 593100.0 ;
      RECT  39150.0 591900.0 35550.0 593100.0 ;
      RECT  48450.0 594600.0 39150.0 595500.0 ;
      RECT  39150.0 591900.0 37950.0 593100.0 ;
      RECT  39150.0 594300.0 37950.0 595500.0 ;
      RECT  39150.0 594300.0 37950.0 595500.0 ;
      RECT  39150.0 591900.0 37950.0 593100.0 ;
      RECT  48450.0 591900.0 47250.0 593100.0 ;
      RECT  48450.0 594300.0 47250.0 595500.0 ;
      RECT  48450.0 594300.0 47250.0 595500.0 ;
      RECT  48450.0 591900.0 47250.0 593100.0 ;
      RECT  38550.0 596700.0 37350.0 597900.0 ;
      RECT  48450.0 596700.0 47250.0 597900.0 ;
      RECT  43800.0 592500.0 42600.0 593700.0 ;
      RECT  43800.0 592500.0 42600.0 593700.0 ;
      RECT  43650.0 595050.0 42750.0 595950.0 ;
      RECT  36450.0 590100.0 35550.0 599700.0 ;
      RECT  50250.0 590100.0 49350.0 599700.0 ;
      RECT  37950.0 606300.0 36000.0 607500.0 ;
      RECT  49800.0 606300.0 47850.0 607500.0 ;
      RECT  48450.0 601500.0 50250.0 602700.0 ;
      RECT  39150.0 601500.0 35550.0 602700.0 ;
      RECT  48450.0 604200.0 39150.0 605100.0 ;
      RECT  39150.0 601500.0 37950.0 602700.0 ;
      RECT  39150.0 603900.0 37950.0 605100.0 ;
      RECT  39150.0 603900.0 37950.0 605100.0 ;
      RECT  39150.0 601500.0 37950.0 602700.0 ;
      RECT  48450.0 601500.0 47250.0 602700.0 ;
      RECT  48450.0 603900.0 47250.0 605100.0 ;
      RECT  48450.0 603900.0 47250.0 605100.0 ;
      RECT  48450.0 601500.0 47250.0 602700.0 ;
      RECT  38550.0 606300.0 37350.0 607500.0 ;
      RECT  48450.0 606300.0 47250.0 607500.0 ;
      RECT  43800.0 602100.0 42600.0 603300.0 ;
      RECT  43800.0 602100.0 42600.0 603300.0 ;
      RECT  43650.0 604650.0 42750.0 605550.0 ;
      RECT  36450.0 599700.0 35550.0 609300.0 ;
      RECT  50250.0 599700.0 49350.0 609300.0 ;
      RECT  42600.0 602100.0 43800.0 603300.0 ;
      RECT  37950.0 615900.0 36000.0 617100.0 ;
      RECT  49800.0 615900.0 47850.0 617100.0 ;
      RECT  48450.0 611100.0 50250.0 612300.0 ;
      RECT  39150.0 611100.0 35550.0 612300.0 ;
      RECT  48450.0 613800.0 39150.0 614700.0 ;
      RECT  39150.0 611100.0 37950.0 612300.0 ;
      RECT  39150.0 613500.0 37950.0 614700.0 ;
      RECT  39150.0 613500.0 37950.0 614700.0 ;
      RECT  39150.0 611100.0 37950.0 612300.0 ;
      RECT  48450.0 611100.0 47250.0 612300.0 ;
      RECT  48450.0 613500.0 47250.0 614700.0 ;
      RECT  48450.0 613500.0 47250.0 614700.0 ;
      RECT  48450.0 611100.0 47250.0 612300.0 ;
      RECT  38550.0 615900.0 37350.0 617100.0 ;
      RECT  48450.0 615900.0 47250.0 617100.0 ;
      RECT  43800.0 611700.0 42600.0 612900.0 ;
      RECT  43800.0 611700.0 42600.0 612900.0 ;
      RECT  43650.0 614250.0 42750.0 615150.0 ;
      RECT  36450.0 609300.0 35550.0 618900.0 ;
      RECT  50250.0 609300.0 49350.0 618900.0 ;
      RECT  42600.0 611700.0 43800.0 612900.0 ;
      RECT  37950.0 625500.0 36000.0 626700.0 ;
      RECT  49800.0 625500.0 47850.0 626700.0 ;
      RECT  48450.0 620700.0 50250.0 621900.0 ;
      RECT  39150.0 620700.0 35550.0 621900.0 ;
      RECT  48450.0 623400.0 39150.0 624300.0 ;
      RECT  39150.0 620700.0 37950.0 621900.0 ;
      RECT  39150.0 623100.0 37950.0 624300.0 ;
      RECT  39150.0 623100.0 37950.0 624300.0 ;
      RECT  39150.0 620700.0 37950.0 621900.0 ;
      RECT  48450.0 620700.0 47250.0 621900.0 ;
      RECT  48450.0 623100.0 47250.0 624300.0 ;
      RECT  48450.0 623100.0 47250.0 624300.0 ;
      RECT  48450.0 620700.0 47250.0 621900.0 ;
      RECT  38550.0 625500.0 37350.0 626700.0 ;
      RECT  48450.0 625500.0 47250.0 626700.0 ;
      RECT  43800.0 621300.0 42600.0 622500.0 ;
      RECT  43800.0 621300.0 42600.0 622500.0 ;
      RECT  43650.0 623850.0 42750.0 624750.0 ;
      RECT  36450.0 618900.0 35550.0 628500.0 ;
      RECT  50250.0 618900.0 49350.0 628500.0 ;
      RECT  42600.0 621300.0 43800.0 622500.0 ;
      RECT  37950.0 635100.0 36000.0 636300.0 ;
      RECT  49800.0 635100.0 47850.0 636300.0 ;
      RECT  48450.0 630300.0 50250.0 631500.0 ;
      RECT  39150.0 630300.0 35550.0 631500.0 ;
      RECT  48450.0 633000.0 39150.0 633900.0 ;
      RECT  39150.0 630300.0 37950.0 631500.0 ;
      RECT  39150.0 632700.0 37950.0 633900.0 ;
      RECT  39150.0 632700.0 37950.0 633900.0 ;
      RECT  39150.0 630300.0 37950.0 631500.0 ;
      RECT  48450.0 630300.0 47250.0 631500.0 ;
      RECT  48450.0 632700.0 47250.0 633900.0 ;
      RECT  48450.0 632700.0 47250.0 633900.0 ;
      RECT  48450.0 630300.0 47250.0 631500.0 ;
      RECT  38550.0 635100.0 37350.0 636300.0 ;
      RECT  48450.0 635100.0 47250.0 636300.0 ;
      RECT  43800.0 630900.0 42600.0 632100.0 ;
      RECT  43800.0 630900.0 42600.0 632100.0 ;
      RECT  43650.0 633450.0 42750.0 634350.0 ;
      RECT  36450.0 628500.0 35550.0 638100.0 ;
      RECT  50250.0 628500.0 49350.0 638100.0 ;
      RECT  42600.0 630900.0 43800.0 632100.0 ;
      RECT  37950.0 644700.0 36000.0 645900.0 ;
      RECT  49800.0 644700.0 47850.0 645900.0 ;
      RECT  48450.0 639900.0 50250.0 641100.0 ;
      RECT  39150.0 639900.0 35550.0 641100.0 ;
      RECT  48450.0 642600.0 39150.0 643500.0 ;
      RECT  39150.0 639900.0 37950.0 641100.0 ;
      RECT  39150.0 642300.0 37950.0 643500.0 ;
      RECT  39150.0 642300.0 37950.0 643500.0 ;
      RECT  39150.0 639900.0 37950.0 641100.0 ;
      RECT  48450.0 639900.0 47250.0 641100.0 ;
      RECT  48450.0 642300.0 47250.0 643500.0 ;
      RECT  48450.0 642300.0 47250.0 643500.0 ;
      RECT  48450.0 639900.0 47250.0 641100.0 ;
      RECT  38550.0 644700.0 37350.0 645900.0 ;
      RECT  48450.0 644700.0 47250.0 645900.0 ;
      RECT  43800.0 640500.0 42600.0 641700.0 ;
      RECT  43800.0 640500.0 42600.0 641700.0 ;
      RECT  43650.0 643050.0 42750.0 643950.0 ;
      RECT  36450.0 638100.0 35550.0 647700.0 ;
      RECT  50250.0 638100.0 49350.0 647700.0 ;
      RECT  42600.0 640500.0 43800.0 641700.0 ;
      RECT  37950.0 654300.0 36000.0 655500.0 ;
      RECT  49800.0 654300.0 47850.0 655500.0 ;
      RECT  48450.0 649500.0 50250.0 650700.0 ;
      RECT  39150.0 649500.0 35550.0 650700.0 ;
      RECT  48450.0 652200.0 39150.0 653100.0 ;
      RECT  39150.0 649500.0 37950.0 650700.0 ;
      RECT  39150.0 651900.0 37950.0 653100.0 ;
      RECT  39150.0 651900.0 37950.0 653100.0 ;
      RECT  39150.0 649500.0 37950.0 650700.0 ;
      RECT  48450.0 649500.0 47250.0 650700.0 ;
      RECT  48450.0 651900.0 47250.0 653100.0 ;
      RECT  48450.0 651900.0 47250.0 653100.0 ;
      RECT  48450.0 649500.0 47250.0 650700.0 ;
      RECT  38550.0 654300.0 37350.0 655500.0 ;
      RECT  48450.0 654300.0 47250.0 655500.0 ;
      RECT  43800.0 650100.0 42600.0 651300.0 ;
      RECT  43800.0 650100.0 42600.0 651300.0 ;
      RECT  43650.0 652650.0 42750.0 653550.0 ;
      RECT  36450.0 647700.0 35550.0 657300.0 ;
      RECT  50250.0 647700.0 49350.0 657300.0 ;
      RECT  42600.0 650100.0 43800.0 651300.0 ;
      RECT  34050.0 641100.0 36000.0 639900.0 ;
      RECT  22200.0 641100.0 24150.0 639900.0 ;
      RECT  23550.0 645900.0 21750.0 644700.0 ;
      RECT  32850.0 645900.0 36450.0 644700.0 ;
      RECT  23550.0 643200.0 32850.0 642300.0 ;
      RECT  32850.0 645900.0 34050.0 644700.0 ;
      RECT  32850.0 643500.0 34050.0 642300.0 ;
      RECT  32850.0 643500.0 34050.0 642300.0 ;
      RECT  32850.0 645900.0 34050.0 644700.0 ;
      RECT  23550.0 645900.0 24750.0 644700.0 ;
      RECT  23550.0 643500.0 24750.0 642300.0 ;
      RECT  23550.0 643500.0 24750.0 642300.0 ;
      RECT  23550.0 645900.0 24750.0 644700.0 ;
      RECT  33450.0 641100.0 34650.0 639900.0 ;
      RECT  23550.0 641100.0 24750.0 639900.0 ;
      RECT  28200.0 645300.0 29400.0 644100.0 ;
      RECT  28200.0 645300.0 29400.0 644100.0 ;
      RECT  28350.0 642750.0 29250.0 641850.0 ;
      RECT  35550.0 647700.0 36450.0 638100.0 ;
      RECT  21750.0 647700.0 22650.0 638100.0 ;
      RECT  28200.0 644100.0 29400.0 645300.0 ;
      RECT  34050.0 631500.0 36000.0 630300.0 ;
      RECT  22200.0 631500.0 24150.0 630300.0 ;
      RECT  23550.0 636300.0 21750.0 635100.0 ;
      RECT  32850.0 636300.0 36450.0 635100.0 ;
      RECT  23550.0 633600.0 32850.0 632700.0 ;
      RECT  32850.0 636300.0 34050.0 635100.0 ;
      RECT  32850.0 633900.0 34050.0 632700.0 ;
      RECT  32850.0 633900.0 34050.0 632700.0 ;
      RECT  32850.0 636300.0 34050.0 635100.0 ;
      RECT  23550.0 636300.0 24750.0 635100.0 ;
      RECT  23550.0 633900.0 24750.0 632700.0 ;
      RECT  23550.0 633900.0 24750.0 632700.0 ;
      RECT  23550.0 636300.0 24750.0 635100.0 ;
      RECT  33450.0 631500.0 34650.0 630300.0 ;
      RECT  23550.0 631500.0 24750.0 630300.0 ;
      RECT  28200.0 635700.0 29400.0 634500.0 ;
      RECT  28200.0 635700.0 29400.0 634500.0 ;
      RECT  28350.0 633150.0 29250.0 632250.0 ;
      RECT  35550.0 638100.0 36450.0 628500.0 ;
      RECT  21750.0 638100.0 22650.0 628500.0 ;
      RECT  28200.0 634500.0 29400.0 635700.0 ;
      RECT  34050.0 621900.0 36000.0 620700.0 ;
      RECT  22200.0 621900.0 24150.0 620700.0 ;
      RECT  23550.0 626700.0 21750.0 625500.0 ;
      RECT  32850.0 626700.0 36450.0 625500.0 ;
      RECT  23550.0 624000.0 32850.0 623100.0 ;
      RECT  32850.0 626700.0 34050.0 625500.0 ;
      RECT  32850.0 624300.0 34050.0 623100.0 ;
      RECT  32850.0 624300.0 34050.0 623100.0 ;
      RECT  32850.0 626700.0 34050.0 625500.0 ;
      RECT  23550.0 626700.0 24750.0 625500.0 ;
      RECT  23550.0 624300.0 24750.0 623100.0 ;
      RECT  23550.0 624300.0 24750.0 623100.0 ;
      RECT  23550.0 626700.0 24750.0 625500.0 ;
      RECT  33450.0 621900.0 34650.0 620700.0 ;
      RECT  23550.0 621900.0 24750.0 620700.0 ;
      RECT  28200.0 626100.0 29400.0 624900.0 ;
      RECT  28200.0 626100.0 29400.0 624900.0 ;
      RECT  28350.0 623550.0 29250.0 622650.0 ;
      RECT  35550.0 628500.0 36450.0 618900.0 ;
      RECT  21750.0 628500.0 22650.0 618900.0 ;
      RECT  28200.0 624900.0 29400.0 626100.0 ;
      RECT  34050.0 612300.0 36000.0 611100.0 ;
      RECT  22200.0 612300.0 24150.0 611100.0 ;
      RECT  23550.0 617100.0 21750.0 615900.0 ;
      RECT  32850.0 617100.0 36450.0 615900.0 ;
      RECT  23550.0 614400.0 32850.0 613500.0 ;
      RECT  32850.0 617100.0 34050.0 615900.0 ;
      RECT  32850.0 614700.0 34050.0 613500.0 ;
      RECT  32850.0 614700.0 34050.0 613500.0 ;
      RECT  32850.0 617100.0 34050.0 615900.0 ;
      RECT  23550.0 617100.0 24750.0 615900.0 ;
      RECT  23550.0 614700.0 24750.0 613500.0 ;
      RECT  23550.0 614700.0 24750.0 613500.0 ;
      RECT  23550.0 617100.0 24750.0 615900.0 ;
      RECT  33450.0 612300.0 34650.0 611100.0 ;
      RECT  23550.0 612300.0 24750.0 611100.0 ;
      RECT  28200.0 616500.0 29400.0 615300.0 ;
      RECT  28200.0 616500.0 29400.0 615300.0 ;
      RECT  28350.0 613950.0 29250.0 613050.0 ;
      RECT  35550.0 618900.0 36450.0 609300.0 ;
      RECT  21750.0 618900.0 22650.0 609300.0 ;
      RECT  28200.0 615300.0 29400.0 616500.0 ;
      RECT  34050.0 602700.0 36000.0 601500.0 ;
      RECT  22200.0 602700.0 24150.0 601500.0 ;
      RECT  23550.0 607500.0 21750.0 606300.0 ;
      RECT  32850.0 607500.0 36450.0 606300.0 ;
      RECT  23550.0 604800.0 32850.0 603900.0 ;
      RECT  32850.0 607500.0 34050.0 606300.0 ;
      RECT  32850.0 605100.0 34050.0 603900.0 ;
      RECT  32850.0 605100.0 34050.0 603900.0 ;
      RECT  32850.0 607500.0 34050.0 606300.0 ;
      RECT  23550.0 607500.0 24750.0 606300.0 ;
      RECT  23550.0 605100.0 24750.0 603900.0 ;
      RECT  23550.0 605100.0 24750.0 603900.0 ;
      RECT  23550.0 607500.0 24750.0 606300.0 ;
      RECT  33450.0 602700.0 34650.0 601500.0 ;
      RECT  23550.0 602700.0 24750.0 601500.0 ;
      RECT  28200.0 606900.0 29400.0 605700.0 ;
      RECT  28200.0 606900.0 29400.0 605700.0 ;
      RECT  28350.0 604350.0 29250.0 603450.0 ;
      RECT  35550.0 609300.0 36450.0 599700.0 ;
      RECT  21750.0 609300.0 22650.0 599700.0 ;
      RECT  28200.0 605700.0 29400.0 606900.0 ;
      RECT  34050.0 593100.0 36000.0 591900.0 ;
      RECT  22200.0 593100.0 24150.0 591900.0 ;
      RECT  23550.0 597900.0 21750.0 596700.0 ;
      RECT  32850.0 597900.0 36450.0 596700.0 ;
      RECT  23550.0 595200.0 32850.0 594300.0 ;
      RECT  32850.0 597900.0 34050.0 596700.0 ;
      RECT  32850.0 595500.0 34050.0 594300.0 ;
      RECT  32850.0 595500.0 34050.0 594300.0 ;
      RECT  32850.0 597900.0 34050.0 596700.0 ;
      RECT  23550.0 597900.0 24750.0 596700.0 ;
      RECT  23550.0 595500.0 24750.0 594300.0 ;
      RECT  23550.0 595500.0 24750.0 594300.0 ;
      RECT  23550.0 597900.0 24750.0 596700.0 ;
      RECT  33450.0 593100.0 34650.0 591900.0 ;
      RECT  23550.0 593100.0 24750.0 591900.0 ;
      RECT  28200.0 597300.0 29400.0 596100.0 ;
      RECT  28200.0 597300.0 29400.0 596100.0 ;
      RECT  28350.0 594750.0 29250.0 593850.0 ;
      RECT  35550.0 599700.0 36450.0 590100.0 ;
      RECT  21750.0 599700.0 22650.0 590100.0 ;
      RECT  28200.0 596100.0 29400.0 597300.0 ;
      RECT  42600.0 594900.0 43800.0 596100.0 ;
      RECT  42600.0 623700.0 43800.0 624900.0 ;
      RECT  42600.0 652500.0 43800.0 653700.0 ;
      RECT  28200.0 622500.0 29400.0 623700.0 ;
      RECT  42600.0 592500.0 43800.0 593700.0 ;
      RECT  28350.0 590100.0 29250.0 593850.0 ;
      RECT  35550.0 590100.0 36450.0 657300.0 ;
      RECT  21750.0 590100.0 22650.0 657300.0 ;
      RECT  49350.0 590100.0 50250.0 657300.0 ;
      RECT  16800.0 575100.0 6600.0 561300.0 ;
      RECT  16800.0 575100.0 6600.0 588900.0 ;
      RECT  16800.0 602700.0 6600.0 588900.0 ;
      RECT  16800.0 602700.0 6600.0 616500.0 ;
      RECT  16800.0 630300.0 6600.0 616500.0 ;
      RECT  16800.0 630300.0 6600.0 644100.0 ;
      RECT  16800.0 657900.0 6600.0 644100.0 ;
      RECT  16800.0 657900.0 6600.0 671700.0 ;
      RECT  16800.0 685500.0 6600.0 671700.0 ;
      RECT  16800.0 685500.0 6600.0 699300.0 ;
      RECT  16800.0 713100.0 6600.0 699300.0 ;
      RECT  16800.0 713100.0 6600.0 726900.0 ;
      RECT  16800.0 740700.0 6600.0 726900.0 ;
      RECT  16800.0 740700.0 6600.0 754500.0 ;
      RECT  16800.0 768300.0 6600.0 754500.0 ;
      RECT  16800.0 768300.0 6600.0 782100.0 ;
      RECT  16800.0 795900.0 6600.0 782100.0 ;
      RECT  16800.0 795900.0 6600.0 809700.0 ;
      RECT  16800.0 823500.0 6600.0 809700.0 ;
      RECT  16800.0 823500.0 6600.0 837300.0 ;
      RECT  16800.0 851100.0 6600.0 837300.0 ;
      RECT  16800.0 851100.0 6600.0 864900.0 ;
      RECT  16800.0 878700.0 6600.0 864900.0 ;
      RECT  16800.0 878700.0 6600.0 892500.0 ;
      RECT  16800.0 906300.0 6600.0 892500.0 ;
      RECT  16800.0 906300.0 6600.0 920100.0 ;
      RECT  16800.0 933900.0 6600.0 920100.0 ;
      RECT  17400.0 576600.0 6000.0 577800.0 ;
      RECT  17400.0 600000.0 6000.0 601200.0 ;
      RECT  17400.0 604200.0 6000.0 605400.0 ;
      RECT  17400.0 627600.0 6000.0 628800.0 ;
      RECT  17400.0 631800.0 6000.0 633000.0 ;
      RECT  17400.0 655200.0 6000.0 656400.0 ;
      RECT  17400.0 659400.0 6000.0 660600.0 ;
      RECT  17400.0 682800.0 6000.0 684000.0 ;
      RECT  17400.0 687000.0 6000.0 688200.0 ;
      RECT  17400.0 710400.0 6000.0 711600.0 ;
      RECT  17400.0 714600.0 6000.0 715800.0 ;
      RECT  17400.0 738000.0 6000.0 739200.0 ;
      RECT  17400.0 742200.0 6000.0 743400.0 ;
      RECT  17400.0 765600.0 6000.0 766800.0 ;
      RECT  17400.0 769800.0 6000.0 771000.0 ;
      RECT  17400.0 793200.0 6000.0 794400.0 ;
      RECT  17400.0 797400.0 6000.0 798600.0 ;
      RECT  17400.0 820800.0 6000.0 822000.0 ;
      RECT  17400.0 825000.0 6000.0 826200.0 ;
      RECT  17400.0 848400.0 6000.0 849600.0 ;
      RECT  17400.0 852600.0 6000.0 853800.0 ;
      RECT  17400.0 876000.0 6000.0 877200.0 ;
      RECT  17400.0 880200.0 6000.0 881400.0 ;
      RECT  17400.0 903600.0 6000.0 904800.0 ;
      RECT  17400.0 907800.0 6000.0 909000.0 ;
      RECT  17400.0 931200.0 6000.0 932400.0 ;
      RECT  17400.0 588300.0 6000.0 589200.0 ;
      RECT  17400.0 615900.0 6000.0 616800.0 ;
      RECT  17400.0 643500.0 6000.0 644400.0 ;
      RECT  17400.0 671100.0 6000.0 672000.0 ;
      RECT  17400.0 698700.0 6000.0 699600.0 ;
      RECT  17400.0 726300.0 6000.0 727200.0 ;
      RECT  17400.0 753900.0 6000.0 754800.0 ;
      RECT  17400.0 781500.0 6000.0 782400.0 ;
      RECT  17400.0 809100.0 6000.0 810000.0 ;
      RECT  17400.0 836700.0 6000.0 837600.0 ;
      RECT  17400.0 864300.0 6000.0 865200.0 ;
      RECT  17400.0 891900.0 6000.0 892800.0 ;
      RECT  17400.0 919500.0 6000.0 920400.0 ;
      RECT  22350.0 576600.0 21150.0 577800.0 ;
      RECT  22350.0 600000.0 21150.0 601200.0 ;
      RECT  22350.0 604200.0 21150.0 605400.0 ;
      RECT  22350.0 627600.0 21150.0 628800.0 ;
      RECT  22350.0 631800.0 21150.0 633000.0 ;
      RECT  22350.0 655200.0 21150.0 656400.0 ;
      RECT  22350.0 659400.0 21150.0 660600.0 ;
      RECT  22350.0 682800.0 21150.0 684000.0 ;
      RECT  22350.0 687000.0 21150.0 688200.0 ;
      RECT  22350.0 710400.0 21150.0 711600.0 ;
      RECT  22350.0 714600.0 21150.0 715800.0 ;
      RECT  22350.0 738000.0 21150.0 739200.0 ;
      RECT  22350.0 742200.0 21150.0 743400.0 ;
      RECT  22350.0 765600.0 21150.0 766800.0 ;
      RECT  22350.0 769800.0 21150.0 771000.0 ;
      RECT  22350.0 793200.0 21150.0 794400.0 ;
      RECT  22350.0 797400.0 21150.0 798600.0 ;
      RECT  22350.0 820800.0 21150.0 822000.0 ;
      RECT  22350.0 825000.0 21150.0 826200.0 ;
      RECT  22350.0 848400.0 21150.0 849600.0 ;
      RECT  22350.0 852600.0 21150.0 853800.0 ;
      RECT  22350.0 876000.0 21150.0 877200.0 ;
      RECT  22350.0 880200.0 21150.0 881400.0 ;
      RECT  22350.0 903600.0 21150.0 904800.0 ;
      RECT  22350.0 907800.0 21150.0 909000.0 ;
      RECT  22350.0 931200.0 21150.0 932400.0 ;
      RECT  22200.0 590100.0 21000.0 591300.0 ;
      RECT  22800.0 550500.0 21600.0 551700.0 ;
      RECT  16200.0 551100.0 17400.0 552300.0 ;
      RECT  6000.0 551100.0 7200.0 552300.0 ;
      RECT  29400.0 576900.0 28200.0 578100.0 ;
      RECT  19350.0 563400.0 20550.0 564600.0 ;
      RECT  19350.0 555300.0 20550.0 556500.0 ;
      RECT  12600.0 555300.0 13800.0 556500.0 ;
      RECT  43800.0 542100.0 42900.0 592500.0 ;
      RECT  29250.0 542100.0 28350.0 555450.0 ;
      RECT  4500.0 542100.0 3600.0 936150.0 ;
      RECT  36450.0 542100.0 35550.0 590100.0 ;
      RECT  22650.0 542100.0 21750.0 551700.0 ;
      RECT  50250.0 542100.0 49350.0 590100.0 ;
      RECT  43950.0 465450.0 42750.0 464250.0 ;
      RECT  43950.0 424500.0 42750.0 423300.0 ;
      RECT  33900.0 385650.0 32700.0 384450.0 ;
      RECT  29850.0 465450.0 28650.0 464250.0 ;
      RECT  27150.0 470850.0 25950.0 469650.0 ;
      RECT  30600.0 508200.0 29400.0 507000.0 ;
      RECT  27900.0 511200.0 26700.0 510000.0 ;
      RECT  41850.0 484350.0 40650.0 483150.0 ;
      RECT  43800.0 481650.0 42600.0 480450.0 ;
      RECT  45750.0 473550.0 44550.0 472350.0 ;
      RECT  14250.0 484350.0 13050.0 483150.0 ;
      RECT  16200.0 473550.0 15000.0 472350.0 ;
      RECT  18150.0 476250.0 16950.0 475050.0 ;
      RECT  29850.0 502500.0 28650.0 503700.0 ;
      RECT  30600.0 519600.0 29400.0 520800.0 ;
      RECT  16200.0 542100.0 15000.0 543300.0 ;
      RECT  29400.0 522300.0 28200.0 523500.0 ;
      RECT  50400.0 468150.0 49200.0 466950.0 ;
      RECT  36600.0 478950.0 35400.0 477750.0 ;
      RECT  22800.0 468150.0 21600.0 466950.0 ;
      RECT  9000.0 478950.0 7800.0 477750.0 ;
      RECT  43800.0 382200.0 42600.0 385800.0 ;
      RECT  36450.0 382200.0 35550.0 383100.0 ;
      RECT  50250.0 382200.0 49350.0 383100.0 ;
      RECT  55650.0 477750.0 54450.0 478950.0 ;
   LAYER  metal2 ;
      RECT  214650.0 520200.0 215550.0 522900.0 ;
      RECT  211950.0 540000.0 212850.0 542700.0 ;
      RECT  206550.0 500400.0 207450.0 503100.0 ;
      RECT  203850.0 517500.0 204750.0 520200.0 ;
      RECT  209250.0 481050.0 210150.0 483750.0 ;
      RECT  201150.0 462150.0 202050.0 464850.0 ;
      RECT  49800.0 477900.0 55050.0 478800.0 ;
      RECT  195750.0 464850.0 196650.0 467550.0 ;
      RECT  201150.0 600.0 202050.0 2166000.0 ;
      RECT  203850.0 600.0 204750.0 2166000.0 ;
      RECT  206550.0 600.0 207450.0 2166000.0 ;
      RECT  209250.0 600.0 210150.0 2166000.0 ;
      RECT  211950.0 600.0 212850.0 2166000.0 ;
      RECT  214650.0 600.0 215550.0 2166000.0 ;
      RECT  161550.0 600.0 162450.0 379200.0 ;
      RECT  164250.0 600.0 165150.0 379200.0 ;
      RECT  166950.0 600.0 167850.0 379200.0 ;
      RECT  169650.0 600.0 170550.0 379200.0 ;
      RECT  172350.0 600.0 173250.0 379200.0 ;
      RECT  175050.0 600.0 175950.0 379200.0 ;
      RECT  177750.0 600.0 178650.0 379200.0 ;
      RECT  180450.0 600.0 181350.0 379200.0 ;
      RECT  183150.0 600.0 184050.0 379200.0 ;
      RECT  185850.0 600.0 186750.0 379200.0 ;
      RECT  188550.0 600.0 189450.0 379200.0 ;
      RECT  227550.0 2148000.0 228450.0 2149200.0 ;
      RECT  237750.0 2148000.0 238650.0 2149200.0 ;
      RECT  247950.0 2148000.0 248850.0 2149200.0 ;
      RECT  258150.0 2148000.0 259050.0 2149200.0 ;
      RECT  268350.0 2148000.0 269250.0 2149200.0 ;
      RECT  278550.0 2148000.0 279450.0 2149200.0 ;
      RECT  288750.0 2148000.0 289650.0 2149200.0 ;
      RECT  298950.0 2148000.0 299850.0 2149200.0 ;
      RECT  309150.0 2148000.0 310050.0 2149200.0 ;
      RECT  319350.0 2148000.0 320250.0 2149200.0 ;
      RECT  329550.0 2148000.0 330450.0 2149200.0 ;
      RECT  339750.0 2148000.0 340650.0 2149200.0 ;
      RECT  349950.0 2148000.0 350850.0 2149200.0 ;
      RECT  360150.0 2148000.0 361050.0 2149200.0 ;
      RECT  370350.0 2148000.0 371250.0 2149200.0 ;
      RECT  380550.0 2148000.0 381450.0 2149200.0 ;
      RECT  390750.0 2148000.0 391650.0 2149200.0 ;
      RECT  400950.0 2148000.0 401850.0 2149200.0 ;
      RECT  411150.0 2148000.0 412050.0 2149200.0 ;
      RECT  421350.0 2148000.0 422250.0 2149200.0 ;
      RECT  431550.0 2148000.0 432450.0 2149200.0 ;
      RECT  441750.0 2148000.0 442650.0 2149200.0 ;
      RECT  451950.0 2148000.0 452850.0 2149200.0 ;
      RECT  462150.0 2148000.0 463050.0 2149200.0 ;
      RECT  472350.0 2148000.0 473250.0 2149200.0 ;
      RECT  482550.0 2148000.0 483450.0 2149200.0 ;
      RECT  492750.0 2148000.0 493650.0 2149200.0 ;
      RECT  502950.0 2148000.0 503850.0 2149200.0 ;
      RECT  513150.0 2148000.0 514050.0 2149200.0 ;
      RECT  523350.0 2148000.0 524250.0 2149200.0 ;
      RECT  533550.0 2148000.0 534450.0 2149200.0 ;
      RECT  543750.0 2148000.0 544650.0 2149200.0 ;
      RECT  553950.0 2148000.0 554850.0 2149200.0 ;
      RECT  564150.0 2148000.0 565050.0 2149200.0 ;
      RECT  574350.0 2148000.0 575250.0 2149200.0 ;
      RECT  584550.0 2148000.0 585450.0 2149200.0 ;
      RECT  594750.0 2148000.0 595650.0 2149200.0 ;
      RECT  604950.0 2148000.0 605850.0 2149200.0 ;
      RECT  615150.0 2148000.0 616050.0 2149200.0 ;
      RECT  625350.0 2148000.0 626250.0 2149200.0 ;
      RECT  635550.0 2148000.0 636450.0 2149200.0 ;
      RECT  645750.0 2148000.0 646650.0 2149200.0 ;
      RECT  655950.0 2148000.0 656850.0 2149200.0 ;
      RECT  666150.0 2148000.0 667050.0 2149200.0 ;
      RECT  676350.0 2148000.0 677250.0 2149200.0 ;
      RECT  686550.0 2148000.0 687450.0 2149200.0 ;
      RECT  696750.0 2148000.0 697650.0 2149200.0 ;
      RECT  706950.0 2148000.0 707850.0 2149200.0 ;
      RECT  717150.0 2148000.0 718050.0 2149200.0 ;
      RECT  727350.0 2148000.0 728250.0 2149200.0 ;
      RECT  737550.0 2148000.0 738450.0 2149200.0 ;
      RECT  747750.0 2148000.0 748650.0 2149200.0 ;
      RECT  757950.0 2148000.0 758850.0 2149200.0 ;
      RECT  768150.0 2148000.0 769050.0 2149200.0 ;
      RECT  778350.0 2148000.0 779250.0 2149200.0 ;
      RECT  788550.0 2148000.0 789450.0 2149200.0 ;
      RECT  798750.0 2148000.0 799650.0 2149200.0 ;
      RECT  808950.0 2148000.0 809850.0 2149200.0 ;
      RECT  819150.0 2148000.0 820050.0 2149200.0 ;
      RECT  829350.0 2148000.0 830250.0 2149200.0 ;
      RECT  839550.0 2148000.0 840450.0 2149200.0 ;
      RECT  849750.0 2148000.0 850650.0 2149200.0 ;
      RECT  859950.0 2148000.0 860850.0 2149200.0 ;
      RECT  870150.0 2148000.0 871050.0 2149200.0 ;
      RECT  880350.0 2148000.0 881250.0 2149200.0 ;
      RECT  890550.0 2148000.0 891450.0 2149200.0 ;
      RECT  900750.0 2148000.0 901650.0 2149200.0 ;
      RECT  910950.0 2148000.0 911850.0 2149200.0 ;
      RECT  921150.0 2148000.0 922050.0 2149200.0 ;
      RECT  931350.0 2148000.0 932250.0 2149200.0 ;
      RECT  941550.0 2148000.0 942450.0 2149200.0 ;
      RECT  951750.0 2148000.0 952650.0 2149200.0 ;
      RECT  961950.0 2148000.0 962850.0 2149200.0 ;
      RECT  972150.0 2148000.0 973050.0 2149200.0 ;
      RECT  982350.0 2148000.0 983250.0 2149200.0 ;
      RECT  992550.0 2148000.0 993450.0 2149200.0 ;
      RECT  1002750.0 2148000.0 1003650.0 2149200.0 ;
      RECT  1012950.0 2148000.0 1013850.0 2149200.0 ;
      RECT  1023150.0 2148000.0 1024050.0 2149200.0 ;
      RECT  1033350.0 2148000.0 1034250.0 2149200.0 ;
      RECT  1043550.0 2148000.0 1044450.0 2149200.0 ;
      RECT  1053750.0 2148000.0 1054650.0 2149200.0 ;
      RECT  1063950.0 2148000.0 1064850.0 2149200.0 ;
      RECT  1074150.0 2148000.0 1075050.0 2149200.0 ;
      RECT  1084350.0 2148000.0 1085250.0 2149200.0 ;
      RECT  1094550.0 2148000.0 1095450.0 2149200.0 ;
      RECT  1104750.0 2148000.0 1105650.0 2149200.0 ;
      RECT  1114950.0 2148000.0 1115850.0 2149200.0 ;
      RECT  1125150.0 2148000.0 1126050.0 2149200.0 ;
      RECT  1135350.0 2148000.0 1136250.0 2149200.0 ;
      RECT  1145550.0 2148000.0 1146450.0 2149200.0 ;
      RECT  1155750.0 2148000.0 1156650.0 2149200.0 ;
      RECT  1165950.0 2148000.0 1166850.0 2149200.0 ;
      RECT  1176150.0 2148000.0 1177050.0 2149200.0 ;
      RECT  1186350.0 2148000.0 1187250.0 2149200.0 ;
      RECT  1196550.0 2148000.0 1197450.0 2149200.0 ;
      RECT  1206750.0 2148000.0 1207650.0 2149200.0 ;
      RECT  1216950.0 2148000.0 1217850.0 2149200.0 ;
      RECT  1227150.0 2148000.0 1228050.0 2149200.0 ;
      RECT  1237350.0 2148000.0 1238250.0 2149200.0 ;
      RECT  1247550.0 2148000.0 1248450.0 2149200.0 ;
      RECT  1257750.0 2148000.0 1258650.0 2149200.0 ;
      RECT  1267950.0 2148000.0 1268850.0 2149200.0 ;
      RECT  1278150.0 2148000.0 1279050.0 2149200.0 ;
      RECT  1288350.0 2148000.0 1289250.0 2149200.0 ;
      RECT  1298550.0 2148000.0 1299450.0 2149200.0 ;
      RECT  1308750.0 2148000.0 1309650.0 2149200.0 ;
      RECT  1318950.0 2148000.0 1319850.0 2149200.0 ;
      RECT  1329150.0 2148000.0 1330050.0 2149200.0 ;
      RECT  1339350.0 2148000.0 1340250.0 2149200.0 ;
      RECT  1349550.0 2148000.0 1350450.0 2149200.0 ;
      RECT  1359750.0 2148000.0 1360650.0 2149200.0 ;
      RECT  1369950.0 2148000.0 1370850.0 2149200.0 ;
      RECT  1380150.0 2148000.0 1381050.0 2149200.0 ;
      RECT  1390350.0 2148000.0 1391250.0 2149200.0 ;
      RECT  1400550.0 2148000.0 1401450.0 2149200.0 ;
      RECT  1410750.0 2148000.0 1411650.0 2149200.0 ;
      RECT  1420950.0 2148000.0 1421850.0 2149200.0 ;
      RECT  1431150.0 2148000.0 1432050.0 2149200.0 ;
      RECT  1441350.0 2148000.0 1442250.0 2149200.0 ;
      RECT  1451550.0 2148000.0 1452450.0 2149200.0 ;
      RECT  1461750.0 2148000.0 1462650.0 2149200.0 ;
      RECT  1471950.0 2148000.0 1472850.0 2149200.0 ;
      RECT  1482150.0 2148000.0 1483050.0 2149200.0 ;
      RECT  1492350.0 2148000.0 1493250.0 2149200.0 ;
      RECT  1502550.0 2148000.0 1503450.0 2149200.0 ;
      RECT  1512750.0 2148000.0 1513650.0 2149200.0 ;
      RECT  1522950.0 2148000.0 1523850.0 2149200.0 ;
      RECT  226050.0 144900.0 226950.0 145800.0 ;
      RECT  222900.0 144900.0 226500.0 145800.0 ;
      RECT  226050.0 145350.0 226950.0 147150.0 ;
      RECT  266850.0 144900.0 267750.0 145800.0 ;
      RECT  263700.0 144900.0 267300.0 145800.0 ;
      RECT  266850.0 145350.0 267750.0 147150.0 ;
      RECT  307650.0 144900.0 308550.0 145800.0 ;
      RECT  304500.0 144900.0 308100.0 145800.0 ;
      RECT  307650.0 145350.0 308550.0 147150.0 ;
      RECT  348450.0 144900.0 349350.0 145800.0 ;
      RECT  345300.0 144900.0 348900.0 145800.0 ;
      RECT  348450.0 145350.0 349350.0 147150.0 ;
      RECT  389250.0 144900.0 390150.0 145800.0 ;
      RECT  386100.0 144900.0 389700.0 145800.0 ;
      RECT  389250.0 145350.0 390150.0 147150.0 ;
      RECT  430050.0 144900.0 430950.0 145800.0 ;
      RECT  426900.0 144900.0 430500.0 145800.0 ;
      RECT  430050.0 145350.0 430950.0 147150.0 ;
      RECT  470850.0 144900.0 471750.0 145800.0 ;
      RECT  467700.0 144900.0 471300.0 145800.0 ;
      RECT  470850.0 145350.0 471750.0 147150.0 ;
      RECT  511650.0 144900.0 512550.0 145800.0 ;
      RECT  508500.0 144900.0 512100.0 145800.0 ;
      RECT  511650.0 145350.0 512550.0 147150.0 ;
      RECT  552450.0 144900.0 553350.0 145800.0 ;
      RECT  549300.0 144900.0 552900.0 145800.0 ;
      RECT  552450.0 145350.0 553350.0 147150.0 ;
      RECT  593250.0 144900.0 594150.0 145800.0 ;
      RECT  590100.0 144900.0 593700.0 145800.0 ;
      RECT  593250.0 145350.0 594150.0 147150.0 ;
      RECT  634050.0 144900.0 634950.0 145800.0 ;
      RECT  630900.0 144900.0 634500.0 145800.0 ;
      RECT  634050.0 145350.0 634950.0 147150.0 ;
      RECT  674850.0 144900.0 675750.0 145800.0 ;
      RECT  671700.0 144900.0 675300.0 145800.0 ;
      RECT  674850.0 145350.0 675750.0 147150.0 ;
      RECT  715650.0 144900.0 716550.0 145800.0 ;
      RECT  712500.0 144900.0 716100.0 145800.0 ;
      RECT  715650.0 145350.0 716550.0 147150.0 ;
      RECT  756450.0 144900.0 757350.0 145800.0 ;
      RECT  753300.0 144900.0 756900.0 145800.0 ;
      RECT  756450.0 145350.0 757350.0 147150.0 ;
      RECT  797250.0 144900.0 798150.0 145800.0 ;
      RECT  794100.0 144900.0 797700.0 145800.0 ;
      RECT  797250.0 145350.0 798150.0 147150.0 ;
      RECT  838050.0 144900.0 838950.0 145800.0 ;
      RECT  834900.0 144900.0 838500.0 145800.0 ;
      RECT  838050.0 145350.0 838950.0 147150.0 ;
      RECT  878850.0 144900.0 879750.0 145800.0 ;
      RECT  875700.0 144900.0 879300.0 145800.0 ;
      RECT  878850.0 145350.0 879750.0 147150.0 ;
      RECT  919650.0 144900.0 920550.0 145800.0 ;
      RECT  916500.0 144900.0 920100.0 145800.0 ;
      RECT  919650.0 145350.0 920550.0 147150.0 ;
      RECT  960450.0 144900.0 961350.0 145800.0 ;
      RECT  957300.0 144900.0 960900.0 145800.0 ;
      RECT  960450.0 145350.0 961350.0 147150.0 ;
      RECT  1001250.0 144900.0 1002150.0 145800.0 ;
      RECT  998100.0 144900.0 1001700.0 145800.0 ;
      RECT  1001250.0 145350.0 1002150.0 147150.0 ;
      RECT  1042050.0 144900.0 1042950.0 145800.0 ;
      RECT  1038900.0 144900.0 1042500.0 145800.0 ;
      RECT  1042050.0 145350.0 1042950.0 147150.0 ;
      RECT  1082850.0 144900.0 1083750.0 145800.0 ;
      RECT  1079700.0 144900.0 1083300.0 145800.0 ;
      RECT  1082850.0 145350.0 1083750.0 147150.0 ;
      RECT  1123650.0 144900.0 1124550.0 145800.0 ;
      RECT  1120500.0 144900.0 1124100.0 145800.0 ;
      RECT  1123650.0 145350.0 1124550.0 147150.0 ;
      RECT  1164450.0 144900.0 1165350.0 145800.0 ;
      RECT  1161300.0 144900.0 1164900.0 145800.0 ;
      RECT  1164450.0 145350.0 1165350.0 147150.0 ;
      RECT  1205250.0 144900.0 1206150.0 145800.0 ;
      RECT  1202100.0 144900.0 1205700.0 145800.0 ;
      RECT  1205250.0 145350.0 1206150.0 147150.0 ;
      RECT  1246050.0 144900.0 1246950.0 145800.0 ;
      RECT  1242900.0 144900.0 1246500.0 145800.0 ;
      RECT  1246050.0 145350.0 1246950.0 147150.0 ;
      RECT  1286850.0 144900.0 1287750.0 145800.0 ;
      RECT  1283700.0 144900.0 1287300.0 145800.0 ;
      RECT  1286850.0 145350.0 1287750.0 147150.0 ;
      RECT  1327650.0 144900.0 1328550.0 145800.0 ;
      RECT  1324500.0 144900.0 1328100.0 145800.0 ;
      RECT  1327650.0 145350.0 1328550.0 147150.0 ;
      RECT  1368450.0 144900.0 1369350.0 145800.0 ;
      RECT  1365300.0 144900.0 1368900.0 145800.0 ;
      RECT  1368450.0 145350.0 1369350.0 147150.0 ;
      RECT  1409250.0 144900.0 1410150.0 145800.0 ;
      RECT  1406100.0 144900.0 1409700.0 145800.0 ;
      RECT  1409250.0 145350.0 1410150.0 147150.0 ;
      RECT  1450050.0 144900.0 1450950.0 145800.0 ;
      RECT  1446900.0 144900.0 1450500.0 145800.0 ;
      RECT  1450050.0 145350.0 1450950.0 147150.0 ;
      RECT  1490850.0 144900.0 1491750.0 145800.0 ;
      RECT  1487700.0 144900.0 1491300.0 145800.0 ;
      RECT  1490850.0 145350.0 1491750.0 147150.0 ;
      RECT  120600.0 2145600.0 121500.0 2147700.0 ;
      RECT  221400.0 379200.0 231600.0 393000.0 ;
      RECT  221400.0 406800.0 231600.0 393000.0 ;
      RECT  221400.0 406800.0 231600.0 420600.0 ;
      RECT  221400.0 434400.0 231600.0 420600.0 ;
      RECT  221400.0 434400.0 231600.0 448200.0 ;
      RECT  221400.0 462000.0 231600.0 448200.0 ;
      RECT  221400.0 462000.0 231600.0 475800.0 ;
      RECT  221400.0 489600.0 231600.0 475800.0 ;
      RECT  221400.0 489600.0 231600.0 503400.0 ;
      RECT  221400.0 517200.0 231600.0 503400.0 ;
      RECT  221400.0 517200.0 231600.0 531000.0 ;
      RECT  221400.0 544800.0 231600.0 531000.0 ;
      RECT  221400.0 544800.0 231600.0 558600.0 ;
      RECT  221400.0 572400.0 231600.0 558600.0 ;
      RECT  221400.0 572400.0 231600.0 586200.0 ;
      RECT  221400.0 600000.0 231600.0 586200.0 ;
      RECT  221400.0 600000.0 231600.0 613800.0 ;
      RECT  221400.0 627600.0 231600.0 613800.0 ;
      RECT  221400.0 627600.0 231600.0 641400.0 ;
      RECT  221400.0 655200.0 231600.0 641400.0 ;
      RECT  221400.0 655200.0 231600.0 669000.0 ;
      RECT  221400.0 682800.0 231600.0 669000.0 ;
      RECT  221400.0 682800.0 231600.0 696600.0 ;
      RECT  221400.0 710400.0 231600.0 696600.0 ;
      RECT  221400.0 710400.0 231600.0 724200.0 ;
      RECT  221400.0 738000.0 231600.0 724200.0 ;
      RECT  221400.0 738000.0 231600.0 751800.0 ;
      RECT  221400.0 765600.0 231600.0 751800.0 ;
      RECT  221400.0 765600.0 231600.0 779400.0 ;
      RECT  221400.0 793200.0 231600.0 779400.0 ;
      RECT  221400.0 793200.0 231600.0 807000.0 ;
      RECT  221400.0 820800.0 231600.0 807000.0 ;
      RECT  221400.0 820800.0 231600.0 834600.0 ;
      RECT  221400.0 848400.0 231600.0 834600.0 ;
      RECT  221400.0 848400.0 231600.0 862200.0 ;
      RECT  221400.0 876000.0 231600.0 862200.0 ;
      RECT  221400.0 876000.0 231600.0 889800.0 ;
      RECT  221400.0 903600.0 231600.0 889800.0 ;
      RECT  221400.0 903600.0 231600.0 917400.0 ;
      RECT  221400.0 931200.0 231600.0 917400.0 ;
      RECT  221400.0 931200.0 231600.0 945000.0 ;
      RECT  221400.0 958800.0 231600.0 945000.0 ;
      RECT  221400.0 958800.0 231600.0 972600.0 ;
      RECT  221400.0 986400.0 231600.0 972600.0 ;
      RECT  221400.0 986400.0 231600.0 1000200.0 ;
      RECT  221400.0 1014000.0 231600.0 1000200.0 ;
      RECT  221400.0 1014000.0 231600.0 1027800.0 ;
      RECT  221400.0 1041600.0 231600.0 1027800.0 ;
      RECT  221400.0 1041600.0 231600.0 1055400.0 ;
      RECT  221400.0 1069200.0 231600.0 1055400.0 ;
      RECT  221400.0 1069200.0 231600.0 1083000.0 ;
      RECT  221400.0 1096800.0 231600.0 1083000.0 ;
      RECT  221400.0 1096800.0 231600.0 1110600.0 ;
      RECT  221400.0 1124400.0 231600.0 1110600.0 ;
      RECT  221400.0 1124400.0 231600.0 1138200.0 ;
      RECT  221400.0 1152000.0 231600.0 1138200.0 ;
      RECT  221400.0 1152000.0 231600.0 1165800.0 ;
      RECT  221400.0 1179600.0 231600.0 1165800.0 ;
      RECT  221400.0 1179600.0 231600.0 1193400.0 ;
      RECT  221400.0 1207200.0 231600.0 1193400.0 ;
      RECT  221400.0 1207200.0 231600.0 1221000.0 ;
      RECT  221400.0 1234800.0 231600.0 1221000.0 ;
      RECT  221400.0 1234800.0 231600.0 1248600.0 ;
      RECT  221400.0 1262400.0 231600.0 1248600.0 ;
      RECT  221400.0 1262400.0 231600.0 1276200.0 ;
      RECT  221400.0 1290000.0 231600.0 1276200.0 ;
      RECT  221400.0 1290000.0 231600.0 1303800.0 ;
      RECT  221400.0 1317600.0 231600.0 1303800.0 ;
      RECT  221400.0 1317600.0 231600.0 1331400.0 ;
      RECT  221400.0 1345200.0 231600.0 1331400.0 ;
      RECT  221400.0 1345200.0 231600.0 1359000.0 ;
      RECT  221400.0 1372800.0 231600.0 1359000.0 ;
      RECT  221400.0 1372800.0 231600.0 1386600.0 ;
      RECT  221400.0 1400400.0 231600.0 1386600.0 ;
      RECT  221400.0 1400400.0 231600.0 1414200.0 ;
      RECT  221400.0 1428000.0 231600.0 1414200.0 ;
      RECT  221400.0 1428000.0 231600.0 1441800.0 ;
      RECT  221400.0 1455600.0 231600.0 1441800.0 ;
      RECT  221400.0 1455600.0 231600.0 1469400.0 ;
      RECT  221400.0 1483200.0 231600.0 1469400.0 ;
      RECT  221400.0 1483200.0 231600.0 1497000.0 ;
      RECT  221400.0 1510800.0 231600.0 1497000.0 ;
      RECT  221400.0 1510800.0 231600.0 1524600.0 ;
      RECT  221400.0 1538400.0 231600.0 1524600.0 ;
      RECT  221400.0 1538400.0 231600.0 1552200.0 ;
      RECT  221400.0 1566000.0 231600.0 1552200.0 ;
      RECT  221400.0 1566000.0 231600.0 1579800.0 ;
      RECT  221400.0 1593600.0 231600.0 1579800.0 ;
      RECT  221400.0 1593600.0 231600.0 1607400.0 ;
      RECT  221400.0 1621200.0 231600.0 1607400.0 ;
      RECT  221400.0 1621200.0 231600.0 1635000.0 ;
      RECT  221400.0 1648800.0 231600.0 1635000.0 ;
      RECT  221400.0 1648800.0 231600.0 1662600.0 ;
      RECT  221400.0 1676400.0 231600.0 1662600.0 ;
      RECT  221400.0 1676400.0 231600.0 1690200.0 ;
      RECT  221400.0 1704000.0 231600.0 1690200.0 ;
      RECT  221400.0 1704000.0 231600.0 1717800.0 ;
      RECT  221400.0 1731600.0 231600.0 1717800.0 ;
      RECT  221400.0 1731600.0 231600.0 1745400.0 ;
      RECT  221400.0 1759200.0 231600.0 1745400.0 ;
      RECT  221400.0 1759200.0 231600.0 1773000.0 ;
      RECT  221400.0 1786800.0 231600.0 1773000.0 ;
      RECT  221400.0 1786800.0 231600.0 1800600.0 ;
      RECT  221400.0 1814400.0 231600.0 1800600.0 ;
      RECT  221400.0 1814400.0 231600.0 1828200.0 ;
      RECT  221400.0 1842000.0 231600.0 1828200.0 ;
      RECT  221400.0 1842000.0 231600.0 1855800.0 ;
      RECT  221400.0 1869600.0 231600.0 1855800.0 ;
      RECT  221400.0 1869600.0 231600.0 1883400.0 ;
      RECT  221400.0 1897200.0 231600.0 1883400.0 ;
      RECT  221400.0 1897200.0 231600.0 1911000.0 ;
      RECT  221400.0 1924800.0 231600.0 1911000.0 ;
      RECT  221400.0 1924800.0 231600.0 1938600.0 ;
      RECT  221400.0 1952400.0 231600.0 1938600.0 ;
      RECT  221400.0 1952400.0 231600.0 1966200.0 ;
      RECT  221400.0 1980000.0 231600.0 1966200.0 ;
      RECT  221400.0 1980000.0 231600.0 1993800.0 ;
      RECT  221400.0 2007600.0 231600.0 1993800.0 ;
      RECT  221400.0 2007600.0 231600.0 2021400.0 ;
      RECT  221400.0 2035200.0 231600.0 2021400.0 ;
      RECT  221400.0 2035200.0 231600.0 2049000.0 ;
      RECT  221400.0 2062800.0 231600.0 2049000.0 ;
      RECT  221400.0 2062800.0 231600.0 2076600.0 ;
      RECT  221400.0 2090400.0 231600.0 2076600.0 ;
      RECT  221400.0 2090400.0 231600.0 2104200.0 ;
      RECT  221400.0 2118000.0 231600.0 2104200.0 ;
      RECT  221400.0 2118000.0 231600.0 2131800.0 ;
      RECT  221400.0 2145600.0 231600.0 2131800.0 ;
      RECT  231600.0 379200.0 241800.0 393000.0 ;
      RECT  231600.0 406800.0 241800.0 393000.0 ;
      RECT  231600.0 406800.0 241800.0 420600.0 ;
      RECT  231600.0 434400.0 241800.0 420600.0 ;
      RECT  231600.0 434400.0 241800.0 448200.0 ;
      RECT  231600.0 462000.0 241800.0 448200.0 ;
      RECT  231600.0 462000.0 241800.0 475800.0 ;
      RECT  231600.0 489600.0 241800.0 475800.0 ;
      RECT  231600.0 489600.0 241800.0 503400.0 ;
      RECT  231600.0 517200.0 241800.0 503400.0 ;
      RECT  231600.0 517200.0 241800.0 531000.0 ;
      RECT  231600.0 544800.0 241800.0 531000.0 ;
      RECT  231600.0 544800.0 241800.0 558600.0 ;
      RECT  231600.0 572400.0 241800.0 558600.0 ;
      RECT  231600.0 572400.0 241800.0 586200.0 ;
      RECT  231600.0 600000.0 241800.0 586200.0 ;
      RECT  231600.0 600000.0 241800.0 613800.0 ;
      RECT  231600.0 627600.0 241800.0 613800.0 ;
      RECT  231600.0 627600.0 241800.0 641400.0 ;
      RECT  231600.0 655200.0 241800.0 641400.0 ;
      RECT  231600.0 655200.0 241800.0 669000.0 ;
      RECT  231600.0 682800.0 241800.0 669000.0 ;
      RECT  231600.0 682800.0 241800.0 696600.0 ;
      RECT  231600.0 710400.0 241800.0 696600.0 ;
      RECT  231600.0 710400.0 241800.0 724200.0 ;
      RECT  231600.0 738000.0 241800.0 724200.0 ;
      RECT  231600.0 738000.0 241800.0 751800.0 ;
      RECT  231600.0 765600.0 241800.0 751800.0 ;
      RECT  231600.0 765600.0 241800.0 779400.0 ;
      RECT  231600.0 793200.0 241800.0 779400.0 ;
      RECT  231600.0 793200.0 241800.0 807000.0 ;
      RECT  231600.0 820800.0 241800.0 807000.0 ;
      RECT  231600.0 820800.0 241800.0 834600.0 ;
      RECT  231600.0 848400.0 241800.0 834600.0 ;
      RECT  231600.0 848400.0 241800.0 862200.0 ;
      RECT  231600.0 876000.0 241800.0 862200.0 ;
      RECT  231600.0 876000.0 241800.0 889800.0 ;
      RECT  231600.0 903600.0 241800.0 889800.0 ;
      RECT  231600.0 903600.0 241800.0 917400.0 ;
      RECT  231600.0 931200.0 241800.0 917400.0 ;
      RECT  231600.0 931200.0 241800.0 945000.0 ;
      RECT  231600.0 958800.0 241800.0 945000.0 ;
      RECT  231600.0 958800.0 241800.0 972600.0 ;
      RECT  231600.0 986400.0 241800.0 972600.0 ;
      RECT  231600.0 986400.0 241800.0 1000200.0 ;
      RECT  231600.0 1014000.0 241800.0 1000200.0 ;
      RECT  231600.0 1014000.0 241800.0 1027800.0 ;
      RECT  231600.0 1041600.0 241800.0 1027800.0 ;
      RECT  231600.0 1041600.0 241800.0 1055400.0 ;
      RECT  231600.0 1069200.0 241800.0 1055400.0 ;
      RECT  231600.0 1069200.0 241800.0 1083000.0 ;
      RECT  231600.0 1096800.0 241800.0 1083000.0 ;
      RECT  231600.0 1096800.0 241800.0 1110600.0 ;
      RECT  231600.0 1124400.0 241800.0 1110600.0 ;
      RECT  231600.0 1124400.0 241800.0 1138200.0 ;
      RECT  231600.0 1152000.0 241800.0 1138200.0 ;
      RECT  231600.0 1152000.0 241800.0 1165800.0 ;
      RECT  231600.0 1179600.0 241800.0 1165800.0 ;
      RECT  231600.0 1179600.0 241800.0 1193400.0 ;
      RECT  231600.0 1207200.0 241800.0 1193400.0 ;
      RECT  231600.0 1207200.0 241800.0 1221000.0 ;
      RECT  231600.0 1234800.0 241800.0 1221000.0 ;
      RECT  231600.0 1234800.0 241800.0 1248600.0 ;
      RECT  231600.0 1262400.0 241800.0 1248600.0 ;
      RECT  231600.0 1262400.0 241800.0 1276200.0 ;
      RECT  231600.0 1290000.0 241800.0 1276200.0 ;
      RECT  231600.0 1290000.0 241800.0 1303800.0 ;
      RECT  231600.0 1317600.0 241800.0 1303800.0 ;
      RECT  231600.0 1317600.0 241800.0 1331400.0 ;
      RECT  231600.0 1345200.0 241800.0 1331400.0 ;
      RECT  231600.0 1345200.0 241800.0 1359000.0 ;
      RECT  231600.0 1372800.0 241800.0 1359000.0 ;
      RECT  231600.0 1372800.0 241800.0 1386600.0 ;
      RECT  231600.0 1400400.0 241800.0 1386600.0 ;
      RECT  231600.0 1400400.0 241800.0 1414200.0 ;
      RECT  231600.0 1428000.0 241800.0 1414200.0 ;
      RECT  231600.0 1428000.0 241800.0 1441800.0 ;
      RECT  231600.0 1455600.0 241800.0 1441800.0 ;
      RECT  231600.0 1455600.0 241800.0 1469400.0 ;
      RECT  231600.0 1483200.0 241800.0 1469400.0 ;
      RECT  231600.0 1483200.0 241800.0 1497000.0 ;
      RECT  231600.0 1510800.0 241800.0 1497000.0 ;
      RECT  231600.0 1510800.0 241800.0 1524600.0 ;
      RECT  231600.0 1538400.0 241800.0 1524600.0 ;
      RECT  231600.0 1538400.0 241800.0 1552200.0 ;
      RECT  231600.0 1566000.0 241800.0 1552200.0 ;
      RECT  231600.0 1566000.0 241800.0 1579800.0 ;
      RECT  231600.0 1593600.0 241800.0 1579800.0 ;
      RECT  231600.0 1593600.0 241800.0 1607400.0 ;
      RECT  231600.0 1621200.0 241800.0 1607400.0 ;
      RECT  231600.0 1621200.0 241800.0 1635000.0 ;
      RECT  231600.0 1648800.0 241800.0 1635000.0 ;
      RECT  231600.0 1648800.0 241800.0 1662600.0 ;
      RECT  231600.0 1676400.0 241800.0 1662600.0 ;
      RECT  231600.0 1676400.0 241800.0 1690200.0 ;
      RECT  231600.0 1704000.0 241800.0 1690200.0 ;
      RECT  231600.0 1704000.0 241800.0 1717800.0 ;
      RECT  231600.0 1731600.0 241800.0 1717800.0 ;
      RECT  231600.0 1731600.0 241800.0 1745400.0 ;
      RECT  231600.0 1759200.0 241800.0 1745400.0 ;
      RECT  231600.0 1759200.0 241800.0 1773000.0 ;
      RECT  231600.0 1786800.0 241800.0 1773000.0 ;
      RECT  231600.0 1786800.0 241800.0 1800600.0 ;
      RECT  231600.0 1814400.0 241800.0 1800600.0 ;
      RECT  231600.0 1814400.0 241800.0 1828200.0 ;
      RECT  231600.0 1842000.0 241800.0 1828200.0 ;
      RECT  231600.0 1842000.0 241800.0 1855800.0 ;
      RECT  231600.0 1869600.0 241800.0 1855800.0 ;
      RECT  231600.0 1869600.0 241800.0 1883400.0 ;
      RECT  231600.0 1897200.0 241800.0 1883400.0 ;
      RECT  231600.0 1897200.0 241800.0 1911000.0 ;
      RECT  231600.0 1924800.0 241800.0 1911000.0 ;
      RECT  231600.0 1924800.0 241800.0 1938600.0 ;
      RECT  231600.0 1952400.0 241800.0 1938600.0 ;
      RECT  231600.0 1952400.0 241800.0 1966200.0 ;
      RECT  231600.0 1980000.0 241800.0 1966200.0 ;
      RECT  231600.0 1980000.0 241800.0 1993800.0 ;
      RECT  231600.0 2007600.0 241800.0 1993800.0 ;
      RECT  231600.0 2007600.0 241800.0 2021400.0 ;
      RECT  231600.0 2035200.0 241800.0 2021400.0 ;
      RECT  231600.0 2035200.0 241800.0 2049000.0 ;
      RECT  231600.0 2062800.0 241800.0 2049000.0 ;
      RECT  231600.0 2062800.0 241800.0 2076600.0 ;
      RECT  231600.0 2090400.0 241800.0 2076600.0 ;
      RECT  231600.0 2090400.0 241800.0 2104200.0 ;
      RECT  231600.0 2118000.0 241800.0 2104200.0 ;
      RECT  231600.0 2118000.0 241800.0 2131800.0 ;
      RECT  231600.0 2145600.0 241800.0 2131800.0 ;
      RECT  241800.0 379200.0 252000.0 393000.0 ;
      RECT  241800.0 406800.0 252000.0 393000.0 ;
      RECT  241800.0 406800.0 252000.0 420600.0 ;
      RECT  241800.0 434400.0 252000.0 420600.0 ;
      RECT  241800.0 434400.0 252000.0 448200.0 ;
      RECT  241800.0 462000.0 252000.0 448200.0 ;
      RECT  241800.0 462000.0 252000.0 475800.0 ;
      RECT  241800.0 489600.0 252000.0 475800.0 ;
      RECT  241800.0 489600.0 252000.0 503400.0 ;
      RECT  241800.0 517200.0 252000.0 503400.0 ;
      RECT  241800.0 517200.0 252000.0 531000.0 ;
      RECT  241800.0 544800.0 252000.0 531000.0 ;
      RECT  241800.0 544800.0 252000.0 558600.0 ;
      RECT  241800.0 572400.0 252000.0 558600.0 ;
      RECT  241800.0 572400.0 252000.0 586200.0 ;
      RECT  241800.0 600000.0 252000.0 586200.0 ;
      RECT  241800.0 600000.0 252000.0 613800.0 ;
      RECT  241800.0 627600.0 252000.0 613800.0 ;
      RECT  241800.0 627600.0 252000.0 641400.0 ;
      RECT  241800.0 655200.0 252000.0 641400.0 ;
      RECT  241800.0 655200.0 252000.0 669000.0 ;
      RECT  241800.0 682800.0 252000.0 669000.0 ;
      RECT  241800.0 682800.0 252000.0 696600.0 ;
      RECT  241800.0 710400.0 252000.0 696600.0 ;
      RECT  241800.0 710400.0 252000.0 724200.0 ;
      RECT  241800.0 738000.0 252000.0 724200.0 ;
      RECT  241800.0 738000.0 252000.0 751800.0 ;
      RECT  241800.0 765600.0 252000.0 751800.0 ;
      RECT  241800.0 765600.0 252000.0 779400.0 ;
      RECT  241800.0 793200.0 252000.0 779400.0 ;
      RECT  241800.0 793200.0 252000.0 807000.0 ;
      RECT  241800.0 820800.0 252000.0 807000.0 ;
      RECT  241800.0 820800.0 252000.0 834600.0 ;
      RECT  241800.0 848400.0 252000.0 834600.0 ;
      RECT  241800.0 848400.0 252000.0 862200.0 ;
      RECT  241800.0 876000.0 252000.0 862200.0 ;
      RECT  241800.0 876000.0 252000.0 889800.0 ;
      RECT  241800.0 903600.0 252000.0 889800.0 ;
      RECT  241800.0 903600.0 252000.0 917400.0 ;
      RECT  241800.0 931200.0 252000.0 917400.0 ;
      RECT  241800.0 931200.0 252000.0 945000.0 ;
      RECT  241800.0 958800.0 252000.0 945000.0 ;
      RECT  241800.0 958800.0 252000.0 972600.0 ;
      RECT  241800.0 986400.0 252000.0 972600.0 ;
      RECT  241800.0 986400.0 252000.0 1000200.0 ;
      RECT  241800.0 1014000.0 252000.0 1000200.0 ;
      RECT  241800.0 1014000.0 252000.0 1027800.0 ;
      RECT  241800.0 1041600.0 252000.0 1027800.0 ;
      RECT  241800.0 1041600.0 252000.0 1055400.0 ;
      RECT  241800.0 1069200.0 252000.0 1055400.0 ;
      RECT  241800.0 1069200.0 252000.0 1083000.0 ;
      RECT  241800.0 1096800.0 252000.0 1083000.0 ;
      RECT  241800.0 1096800.0 252000.0 1110600.0 ;
      RECT  241800.0 1124400.0 252000.0 1110600.0 ;
      RECT  241800.0 1124400.0 252000.0 1138200.0 ;
      RECT  241800.0 1152000.0 252000.0 1138200.0 ;
      RECT  241800.0 1152000.0 252000.0 1165800.0 ;
      RECT  241800.0 1179600.0 252000.0 1165800.0 ;
      RECT  241800.0 1179600.0 252000.0 1193400.0 ;
      RECT  241800.0 1207200.0 252000.0 1193400.0 ;
      RECT  241800.0 1207200.0 252000.0 1221000.0 ;
      RECT  241800.0 1234800.0 252000.0 1221000.0 ;
      RECT  241800.0 1234800.0 252000.0 1248600.0 ;
      RECT  241800.0 1262400.0 252000.0 1248600.0 ;
      RECT  241800.0 1262400.0 252000.0 1276200.0 ;
      RECT  241800.0 1290000.0 252000.0 1276200.0 ;
      RECT  241800.0 1290000.0 252000.0 1303800.0 ;
      RECT  241800.0 1317600.0 252000.0 1303800.0 ;
      RECT  241800.0 1317600.0 252000.0 1331400.0 ;
      RECT  241800.0 1345200.0 252000.0 1331400.0 ;
      RECT  241800.0 1345200.0 252000.0 1359000.0 ;
      RECT  241800.0 1372800.0 252000.0 1359000.0 ;
      RECT  241800.0 1372800.0 252000.0 1386600.0 ;
      RECT  241800.0 1400400.0 252000.0 1386600.0 ;
      RECT  241800.0 1400400.0 252000.0 1414200.0 ;
      RECT  241800.0 1428000.0 252000.0 1414200.0 ;
      RECT  241800.0 1428000.0 252000.0 1441800.0 ;
      RECT  241800.0 1455600.0 252000.0 1441800.0 ;
      RECT  241800.0 1455600.0 252000.0 1469400.0 ;
      RECT  241800.0 1483200.0 252000.0 1469400.0 ;
      RECT  241800.0 1483200.0 252000.0 1497000.0 ;
      RECT  241800.0 1510800.0 252000.0 1497000.0 ;
      RECT  241800.0 1510800.0 252000.0 1524600.0 ;
      RECT  241800.0 1538400.0 252000.0 1524600.0 ;
      RECT  241800.0 1538400.0 252000.0 1552200.0 ;
      RECT  241800.0 1566000.0 252000.0 1552200.0 ;
      RECT  241800.0 1566000.0 252000.0 1579800.0 ;
      RECT  241800.0 1593600.0 252000.0 1579800.0 ;
      RECT  241800.0 1593600.0 252000.0 1607400.0 ;
      RECT  241800.0 1621200.0 252000.0 1607400.0 ;
      RECT  241800.0 1621200.0 252000.0 1635000.0 ;
      RECT  241800.0 1648800.0 252000.0 1635000.0 ;
      RECT  241800.0 1648800.0 252000.0 1662600.0 ;
      RECT  241800.0 1676400.0 252000.0 1662600.0 ;
      RECT  241800.0 1676400.0 252000.0 1690200.0 ;
      RECT  241800.0 1704000.0 252000.0 1690200.0 ;
      RECT  241800.0 1704000.0 252000.0 1717800.0 ;
      RECT  241800.0 1731600.0 252000.0 1717800.0 ;
      RECT  241800.0 1731600.0 252000.0 1745400.0 ;
      RECT  241800.0 1759200.0 252000.0 1745400.0 ;
      RECT  241800.0 1759200.0 252000.0 1773000.0 ;
      RECT  241800.0 1786800.0 252000.0 1773000.0 ;
      RECT  241800.0 1786800.0 252000.0 1800600.0 ;
      RECT  241800.0 1814400.0 252000.0 1800600.0 ;
      RECT  241800.0 1814400.0 252000.0 1828200.0 ;
      RECT  241800.0 1842000.0 252000.0 1828200.0 ;
      RECT  241800.0 1842000.0 252000.0 1855800.0 ;
      RECT  241800.0 1869600.0 252000.0 1855800.0 ;
      RECT  241800.0 1869600.0 252000.0 1883400.0 ;
      RECT  241800.0 1897200.0 252000.0 1883400.0 ;
      RECT  241800.0 1897200.0 252000.0 1911000.0 ;
      RECT  241800.0 1924800.0 252000.0 1911000.0 ;
      RECT  241800.0 1924800.0 252000.0 1938600.0 ;
      RECT  241800.0 1952400.0 252000.0 1938600.0 ;
      RECT  241800.0 1952400.0 252000.0 1966200.0 ;
      RECT  241800.0 1980000.0 252000.0 1966200.0 ;
      RECT  241800.0 1980000.0 252000.0 1993800.0 ;
      RECT  241800.0 2007600.0 252000.0 1993800.0 ;
      RECT  241800.0 2007600.0 252000.0 2021400.0 ;
      RECT  241800.0 2035200.0 252000.0 2021400.0 ;
      RECT  241800.0 2035200.0 252000.0 2049000.0 ;
      RECT  241800.0 2062800.0 252000.0 2049000.0 ;
      RECT  241800.0 2062800.0 252000.0 2076600.0 ;
      RECT  241800.0 2090400.0 252000.0 2076600.0 ;
      RECT  241800.0 2090400.0 252000.0 2104200.0 ;
      RECT  241800.0 2118000.0 252000.0 2104200.0 ;
      RECT  241800.0 2118000.0 252000.0 2131800.0 ;
      RECT  241800.0 2145600.0 252000.0 2131800.0 ;
      RECT  252000.0 379200.0 262200.0 393000.0 ;
      RECT  252000.0 406800.0 262200.0 393000.0 ;
      RECT  252000.0 406800.0 262200.0 420600.0 ;
      RECT  252000.0 434400.0 262200.0 420600.0 ;
      RECT  252000.0 434400.0 262200.0 448200.0 ;
      RECT  252000.0 462000.0 262200.0 448200.0 ;
      RECT  252000.0 462000.0 262200.0 475800.0 ;
      RECT  252000.0 489600.0 262200.0 475800.0 ;
      RECT  252000.0 489600.0 262200.0 503400.0 ;
      RECT  252000.0 517200.0 262200.0 503400.0 ;
      RECT  252000.0 517200.0 262200.0 531000.0 ;
      RECT  252000.0 544800.0 262200.0 531000.0 ;
      RECT  252000.0 544800.0 262200.0 558600.0 ;
      RECT  252000.0 572400.0 262200.0 558600.0 ;
      RECT  252000.0 572400.0 262200.0 586200.0 ;
      RECT  252000.0 600000.0 262200.0 586200.0 ;
      RECT  252000.0 600000.0 262200.0 613800.0 ;
      RECT  252000.0 627600.0 262200.0 613800.0 ;
      RECT  252000.0 627600.0 262200.0 641400.0 ;
      RECT  252000.0 655200.0 262200.0 641400.0 ;
      RECT  252000.0 655200.0 262200.0 669000.0 ;
      RECT  252000.0 682800.0 262200.0 669000.0 ;
      RECT  252000.0 682800.0 262200.0 696600.0 ;
      RECT  252000.0 710400.0 262200.0 696600.0 ;
      RECT  252000.0 710400.0 262200.0 724200.0 ;
      RECT  252000.0 738000.0 262200.0 724200.0 ;
      RECT  252000.0 738000.0 262200.0 751800.0 ;
      RECT  252000.0 765600.0 262200.0 751800.0 ;
      RECT  252000.0 765600.0 262200.0 779400.0 ;
      RECT  252000.0 793200.0 262200.0 779400.0 ;
      RECT  252000.0 793200.0 262200.0 807000.0 ;
      RECT  252000.0 820800.0 262200.0 807000.0 ;
      RECT  252000.0 820800.0 262200.0 834600.0 ;
      RECT  252000.0 848400.0 262200.0 834600.0 ;
      RECT  252000.0 848400.0 262200.0 862200.0 ;
      RECT  252000.0 876000.0 262200.0 862200.0 ;
      RECT  252000.0 876000.0 262200.0 889800.0 ;
      RECT  252000.0 903600.0 262200.0 889800.0 ;
      RECT  252000.0 903600.0 262200.0 917400.0 ;
      RECT  252000.0 931200.0 262200.0 917400.0 ;
      RECT  252000.0 931200.0 262200.0 945000.0 ;
      RECT  252000.0 958800.0 262200.0 945000.0 ;
      RECT  252000.0 958800.0 262200.0 972600.0 ;
      RECT  252000.0 986400.0 262200.0 972600.0 ;
      RECT  252000.0 986400.0 262200.0 1000200.0 ;
      RECT  252000.0 1014000.0 262200.0 1000200.0 ;
      RECT  252000.0 1014000.0 262200.0 1027800.0 ;
      RECT  252000.0 1041600.0 262200.0 1027800.0 ;
      RECT  252000.0 1041600.0 262200.0 1055400.0 ;
      RECT  252000.0 1069200.0 262200.0 1055400.0 ;
      RECT  252000.0 1069200.0 262200.0 1083000.0 ;
      RECT  252000.0 1096800.0 262200.0 1083000.0 ;
      RECT  252000.0 1096800.0 262200.0 1110600.0 ;
      RECT  252000.0 1124400.0 262200.0 1110600.0 ;
      RECT  252000.0 1124400.0 262200.0 1138200.0 ;
      RECT  252000.0 1152000.0 262200.0 1138200.0 ;
      RECT  252000.0 1152000.0 262200.0 1165800.0 ;
      RECT  252000.0 1179600.0 262200.0 1165800.0 ;
      RECT  252000.0 1179600.0 262200.0 1193400.0 ;
      RECT  252000.0 1207200.0 262200.0 1193400.0 ;
      RECT  252000.0 1207200.0 262200.0 1221000.0 ;
      RECT  252000.0 1234800.0 262200.0 1221000.0 ;
      RECT  252000.0 1234800.0 262200.0 1248600.0 ;
      RECT  252000.0 1262400.0 262200.0 1248600.0 ;
      RECT  252000.0 1262400.0 262200.0 1276200.0 ;
      RECT  252000.0 1290000.0 262200.0 1276200.0 ;
      RECT  252000.0 1290000.0 262200.0 1303800.0 ;
      RECT  252000.0 1317600.0 262200.0 1303800.0 ;
      RECT  252000.0 1317600.0 262200.0 1331400.0 ;
      RECT  252000.0 1345200.0 262200.0 1331400.0 ;
      RECT  252000.0 1345200.0 262200.0 1359000.0 ;
      RECT  252000.0 1372800.0 262200.0 1359000.0 ;
      RECT  252000.0 1372800.0 262200.0 1386600.0 ;
      RECT  252000.0 1400400.0 262200.0 1386600.0 ;
      RECT  252000.0 1400400.0 262200.0 1414200.0 ;
      RECT  252000.0 1428000.0 262200.0 1414200.0 ;
      RECT  252000.0 1428000.0 262200.0 1441800.0 ;
      RECT  252000.0 1455600.0 262200.0 1441800.0 ;
      RECT  252000.0 1455600.0 262200.0 1469400.0 ;
      RECT  252000.0 1483200.0 262200.0 1469400.0 ;
      RECT  252000.0 1483200.0 262200.0 1497000.0 ;
      RECT  252000.0 1510800.0 262200.0 1497000.0 ;
      RECT  252000.0 1510800.0 262200.0 1524600.0 ;
      RECT  252000.0 1538400.0 262200.0 1524600.0 ;
      RECT  252000.0 1538400.0 262200.0 1552200.0 ;
      RECT  252000.0 1566000.0 262200.0 1552200.0 ;
      RECT  252000.0 1566000.0 262200.0 1579800.0 ;
      RECT  252000.0 1593600.0 262200.0 1579800.0 ;
      RECT  252000.0 1593600.0 262200.0 1607400.0 ;
      RECT  252000.0 1621200.0 262200.0 1607400.0 ;
      RECT  252000.0 1621200.0 262200.0 1635000.0 ;
      RECT  252000.0 1648800.0 262200.0 1635000.0 ;
      RECT  252000.0 1648800.0 262200.0 1662600.0 ;
      RECT  252000.0 1676400.0 262200.0 1662600.0 ;
      RECT  252000.0 1676400.0 262200.0 1690200.0 ;
      RECT  252000.0 1704000.0 262200.0 1690200.0 ;
      RECT  252000.0 1704000.0 262200.0 1717800.0 ;
      RECT  252000.0 1731600.0 262200.0 1717800.0 ;
      RECT  252000.0 1731600.0 262200.0 1745400.0 ;
      RECT  252000.0 1759200.0 262200.0 1745400.0 ;
      RECT  252000.0 1759200.0 262200.0 1773000.0 ;
      RECT  252000.0 1786800.0 262200.0 1773000.0 ;
      RECT  252000.0 1786800.0 262200.0 1800600.0 ;
      RECT  252000.0 1814400.0 262200.0 1800600.0 ;
      RECT  252000.0 1814400.0 262200.0 1828200.0 ;
      RECT  252000.0 1842000.0 262200.0 1828200.0 ;
      RECT  252000.0 1842000.0 262200.0 1855800.0 ;
      RECT  252000.0 1869600.0 262200.0 1855800.0 ;
      RECT  252000.0 1869600.0 262200.0 1883400.0 ;
      RECT  252000.0 1897200.0 262200.0 1883400.0 ;
      RECT  252000.0 1897200.0 262200.0 1911000.0 ;
      RECT  252000.0 1924800.0 262200.0 1911000.0 ;
      RECT  252000.0 1924800.0 262200.0 1938600.0 ;
      RECT  252000.0 1952400.0 262200.0 1938600.0 ;
      RECT  252000.0 1952400.0 262200.0 1966200.0 ;
      RECT  252000.0 1980000.0 262200.0 1966200.0 ;
      RECT  252000.0 1980000.0 262200.0 1993800.0 ;
      RECT  252000.0 2007600.0 262200.0 1993800.0 ;
      RECT  252000.0 2007600.0 262200.0 2021400.0 ;
      RECT  252000.0 2035200.0 262200.0 2021400.0 ;
      RECT  252000.0 2035200.0 262200.0 2049000.0 ;
      RECT  252000.0 2062800.0 262200.0 2049000.0 ;
      RECT  252000.0 2062800.0 262200.0 2076600.0 ;
      RECT  252000.0 2090400.0 262200.0 2076600.0 ;
      RECT  252000.0 2090400.0 262200.0 2104200.0 ;
      RECT  252000.0 2118000.0 262200.0 2104200.0 ;
      RECT  252000.0 2118000.0 262200.0 2131800.0 ;
      RECT  252000.0 2145600.0 262200.0 2131800.0 ;
      RECT  262200.0 379200.0 272400.0 393000.0 ;
      RECT  262200.0 406800.0 272400.0 393000.0 ;
      RECT  262200.0 406800.0 272400.0 420600.0 ;
      RECT  262200.0 434400.0 272400.0 420600.0 ;
      RECT  262200.0 434400.0 272400.0 448200.0 ;
      RECT  262200.0 462000.0 272400.0 448200.0 ;
      RECT  262200.0 462000.0 272400.0 475800.0 ;
      RECT  262200.0 489600.0 272400.0 475800.0 ;
      RECT  262200.0 489600.0 272400.0 503400.0 ;
      RECT  262200.0 517200.0 272400.0 503400.0 ;
      RECT  262200.0 517200.0 272400.0 531000.0 ;
      RECT  262200.0 544800.0 272400.0 531000.0 ;
      RECT  262200.0 544800.0 272400.0 558600.0 ;
      RECT  262200.0 572400.0 272400.0 558600.0 ;
      RECT  262200.0 572400.0 272400.0 586200.0 ;
      RECT  262200.0 600000.0 272400.0 586200.0 ;
      RECT  262200.0 600000.0 272400.0 613800.0 ;
      RECT  262200.0 627600.0 272400.0 613800.0 ;
      RECT  262200.0 627600.0 272400.0 641400.0 ;
      RECT  262200.0 655200.0 272400.0 641400.0 ;
      RECT  262200.0 655200.0 272400.0 669000.0 ;
      RECT  262200.0 682800.0 272400.0 669000.0 ;
      RECT  262200.0 682800.0 272400.0 696600.0 ;
      RECT  262200.0 710400.0 272400.0 696600.0 ;
      RECT  262200.0 710400.0 272400.0 724200.0 ;
      RECT  262200.0 738000.0 272400.0 724200.0 ;
      RECT  262200.0 738000.0 272400.0 751800.0 ;
      RECT  262200.0 765600.0 272400.0 751800.0 ;
      RECT  262200.0 765600.0 272400.0 779400.0 ;
      RECT  262200.0 793200.0 272400.0 779400.0 ;
      RECT  262200.0 793200.0 272400.0 807000.0 ;
      RECT  262200.0 820800.0 272400.0 807000.0 ;
      RECT  262200.0 820800.0 272400.0 834600.0 ;
      RECT  262200.0 848400.0 272400.0 834600.0 ;
      RECT  262200.0 848400.0 272400.0 862200.0 ;
      RECT  262200.0 876000.0 272400.0 862200.0 ;
      RECT  262200.0 876000.0 272400.0 889800.0 ;
      RECT  262200.0 903600.0 272400.0 889800.0 ;
      RECT  262200.0 903600.0 272400.0 917400.0 ;
      RECT  262200.0 931200.0 272400.0 917400.0 ;
      RECT  262200.0 931200.0 272400.0 945000.0 ;
      RECT  262200.0 958800.0 272400.0 945000.0 ;
      RECT  262200.0 958800.0 272400.0 972600.0 ;
      RECT  262200.0 986400.0 272400.0 972600.0 ;
      RECT  262200.0 986400.0 272400.0 1000200.0 ;
      RECT  262200.0 1014000.0 272400.0 1000200.0 ;
      RECT  262200.0 1014000.0 272400.0 1027800.0 ;
      RECT  262200.0 1041600.0 272400.0 1027800.0 ;
      RECT  262200.0 1041600.0 272400.0 1055400.0 ;
      RECT  262200.0 1069200.0 272400.0 1055400.0 ;
      RECT  262200.0 1069200.0 272400.0 1083000.0 ;
      RECT  262200.0 1096800.0 272400.0 1083000.0 ;
      RECT  262200.0 1096800.0 272400.0 1110600.0 ;
      RECT  262200.0 1124400.0 272400.0 1110600.0 ;
      RECT  262200.0 1124400.0 272400.0 1138200.0 ;
      RECT  262200.0 1152000.0 272400.0 1138200.0 ;
      RECT  262200.0 1152000.0 272400.0 1165800.0 ;
      RECT  262200.0 1179600.0 272400.0 1165800.0 ;
      RECT  262200.0 1179600.0 272400.0 1193400.0 ;
      RECT  262200.0 1207200.0 272400.0 1193400.0 ;
      RECT  262200.0 1207200.0 272400.0 1221000.0 ;
      RECT  262200.0 1234800.0 272400.0 1221000.0 ;
      RECT  262200.0 1234800.0 272400.0 1248600.0 ;
      RECT  262200.0 1262400.0 272400.0 1248600.0 ;
      RECT  262200.0 1262400.0 272400.0 1276200.0 ;
      RECT  262200.0 1290000.0 272400.0 1276200.0 ;
      RECT  262200.0 1290000.0 272400.0 1303800.0 ;
      RECT  262200.0 1317600.0 272400.0 1303800.0 ;
      RECT  262200.0 1317600.0 272400.0 1331400.0 ;
      RECT  262200.0 1345200.0 272400.0 1331400.0 ;
      RECT  262200.0 1345200.0 272400.0 1359000.0 ;
      RECT  262200.0 1372800.0 272400.0 1359000.0 ;
      RECT  262200.0 1372800.0 272400.0 1386600.0 ;
      RECT  262200.0 1400400.0 272400.0 1386600.0 ;
      RECT  262200.0 1400400.0 272400.0 1414200.0 ;
      RECT  262200.0 1428000.0 272400.0 1414200.0 ;
      RECT  262200.0 1428000.0 272400.0 1441800.0 ;
      RECT  262200.0 1455600.0 272400.0 1441800.0 ;
      RECT  262200.0 1455600.0 272400.0 1469400.0 ;
      RECT  262200.0 1483200.0 272400.0 1469400.0 ;
      RECT  262200.0 1483200.0 272400.0 1497000.0 ;
      RECT  262200.0 1510800.0 272400.0 1497000.0 ;
      RECT  262200.0 1510800.0 272400.0 1524600.0 ;
      RECT  262200.0 1538400.0 272400.0 1524600.0 ;
      RECT  262200.0 1538400.0 272400.0 1552200.0 ;
      RECT  262200.0 1566000.0 272400.0 1552200.0 ;
      RECT  262200.0 1566000.0 272400.0 1579800.0 ;
      RECT  262200.0 1593600.0 272400.0 1579800.0 ;
      RECT  262200.0 1593600.0 272400.0 1607400.0 ;
      RECT  262200.0 1621200.0 272400.0 1607400.0 ;
      RECT  262200.0 1621200.0 272400.0 1635000.0 ;
      RECT  262200.0 1648800.0 272400.0 1635000.0 ;
      RECT  262200.0 1648800.0 272400.0 1662600.0 ;
      RECT  262200.0 1676400.0 272400.0 1662600.0 ;
      RECT  262200.0 1676400.0 272400.0 1690200.0 ;
      RECT  262200.0 1704000.0 272400.0 1690200.0 ;
      RECT  262200.0 1704000.0 272400.0 1717800.0 ;
      RECT  262200.0 1731600.0 272400.0 1717800.0 ;
      RECT  262200.0 1731600.0 272400.0 1745400.0 ;
      RECT  262200.0 1759200.0 272400.0 1745400.0 ;
      RECT  262200.0 1759200.0 272400.0 1773000.0 ;
      RECT  262200.0 1786800.0 272400.0 1773000.0 ;
      RECT  262200.0 1786800.0 272400.0 1800600.0 ;
      RECT  262200.0 1814400.0 272400.0 1800600.0 ;
      RECT  262200.0 1814400.0 272400.0 1828200.0 ;
      RECT  262200.0 1842000.0 272400.0 1828200.0 ;
      RECT  262200.0 1842000.0 272400.0 1855800.0 ;
      RECT  262200.0 1869600.0 272400.0 1855800.0 ;
      RECT  262200.0 1869600.0 272400.0 1883400.0 ;
      RECT  262200.0 1897200.0 272400.0 1883400.0 ;
      RECT  262200.0 1897200.0 272400.0 1911000.0 ;
      RECT  262200.0 1924800.0 272400.0 1911000.0 ;
      RECT  262200.0 1924800.0 272400.0 1938600.0 ;
      RECT  262200.0 1952400.0 272400.0 1938600.0 ;
      RECT  262200.0 1952400.0 272400.0 1966200.0 ;
      RECT  262200.0 1980000.0 272400.0 1966200.0 ;
      RECT  262200.0 1980000.0 272400.0 1993800.0 ;
      RECT  262200.0 2007600.0 272400.0 1993800.0 ;
      RECT  262200.0 2007600.0 272400.0 2021400.0 ;
      RECT  262200.0 2035200.0 272400.0 2021400.0 ;
      RECT  262200.0 2035200.0 272400.0 2049000.0 ;
      RECT  262200.0 2062800.0 272400.0 2049000.0 ;
      RECT  262200.0 2062800.0 272400.0 2076600.0 ;
      RECT  262200.0 2090400.0 272400.0 2076600.0 ;
      RECT  262200.0 2090400.0 272400.0 2104200.0 ;
      RECT  262200.0 2118000.0 272400.0 2104200.0 ;
      RECT  262200.0 2118000.0 272400.0 2131800.0 ;
      RECT  262200.0 2145600.0 272400.0 2131800.0 ;
      RECT  272400.0 379200.0 282600.0 393000.0 ;
      RECT  272400.0 406800.0 282600.0 393000.0 ;
      RECT  272400.0 406800.0 282600.0 420600.0 ;
      RECT  272400.0 434400.0 282600.0 420600.0 ;
      RECT  272400.0 434400.0 282600.0 448200.0 ;
      RECT  272400.0 462000.0 282600.0 448200.0 ;
      RECT  272400.0 462000.0 282600.0 475800.0 ;
      RECT  272400.0 489600.0 282600.0 475800.0 ;
      RECT  272400.0 489600.0 282600.0 503400.0 ;
      RECT  272400.0 517200.0 282600.0 503400.0 ;
      RECT  272400.0 517200.0 282600.0 531000.0 ;
      RECT  272400.0 544800.0 282600.0 531000.0 ;
      RECT  272400.0 544800.0 282600.0 558600.0 ;
      RECT  272400.0 572400.0 282600.0 558600.0 ;
      RECT  272400.0 572400.0 282600.0 586200.0 ;
      RECT  272400.0 600000.0 282600.0 586200.0 ;
      RECT  272400.0 600000.0 282600.0 613800.0 ;
      RECT  272400.0 627600.0 282600.0 613800.0 ;
      RECT  272400.0 627600.0 282600.0 641400.0 ;
      RECT  272400.0 655200.0 282600.0 641400.0 ;
      RECT  272400.0 655200.0 282600.0 669000.0 ;
      RECT  272400.0 682800.0 282600.0 669000.0 ;
      RECT  272400.0 682800.0 282600.0 696600.0 ;
      RECT  272400.0 710400.0 282600.0 696600.0 ;
      RECT  272400.0 710400.0 282600.0 724200.0 ;
      RECT  272400.0 738000.0 282600.0 724200.0 ;
      RECT  272400.0 738000.0 282600.0 751800.0 ;
      RECT  272400.0 765600.0 282600.0 751800.0 ;
      RECT  272400.0 765600.0 282600.0 779400.0 ;
      RECT  272400.0 793200.0 282600.0 779400.0 ;
      RECT  272400.0 793200.0 282600.0 807000.0 ;
      RECT  272400.0 820800.0 282600.0 807000.0 ;
      RECT  272400.0 820800.0 282600.0 834600.0 ;
      RECT  272400.0 848400.0 282600.0 834600.0 ;
      RECT  272400.0 848400.0 282600.0 862200.0 ;
      RECT  272400.0 876000.0 282600.0 862200.0 ;
      RECT  272400.0 876000.0 282600.0 889800.0 ;
      RECT  272400.0 903600.0 282600.0 889800.0 ;
      RECT  272400.0 903600.0 282600.0 917400.0 ;
      RECT  272400.0 931200.0 282600.0 917400.0 ;
      RECT  272400.0 931200.0 282600.0 945000.0 ;
      RECT  272400.0 958800.0 282600.0 945000.0 ;
      RECT  272400.0 958800.0 282600.0 972600.0 ;
      RECT  272400.0 986400.0 282600.0 972600.0 ;
      RECT  272400.0 986400.0 282600.0 1000200.0 ;
      RECT  272400.0 1014000.0 282600.0 1000200.0 ;
      RECT  272400.0 1014000.0 282600.0 1027800.0 ;
      RECT  272400.0 1041600.0 282600.0 1027800.0 ;
      RECT  272400.0 1041600.0 282600.0 1055400.0 ;
      RECT  272400.0 1069200.0 282600.0 1055400.0 ;
      RECT  272400.0 1069200.0 282600.0 1083000.0 ;
      RECT  272400.0 1096800.0 282600.0 1083000.0 ;
      RECT  272400.0 1096800.0 282600.0 1110600.0 ;
      RECT  272400.0 1124400.0 282600.0 1110600.0 ;
      RECT  272400.0 1124400.0 282600.0 1138200.0 ;
      RECT  272400.0 1152000.0 282600.0 1138200.0 ;
      RECT  272400.0 1152000.0 282600.0 1165800.0 ;
      RECT  272400.0 1179600.0 282600.0 1165800.0 ;
      RECT  272400.0 1179600.0 282600.0 1193400.0 ;
      RECT  272400.0 1207200.0 282600.0 1193400.0 ;
      RECT  272400.0 1207200.0 282600.0 1221000.0 ;
      RECT  272400.0 1234800.0 282600.0 1221000.0 ;
      RECT  272400.0 1234800.0 282600.0 1248600.0 ;
      RECT  272400.0 1262400.0 282600.0 1248600.0 ;
      RECT  272400.0 1262400.0 282600.0 1276200.0 ;
      RECT  272400.0 1290000.0 282600.0 1276200.0 ;
      RECT  272400.0 1290000.0 282600.0 1303800.0 ;
      RECT  272400.0 1317600.0 282600.0 1303800.0 ;
      RECT  272400.0 1317600.0 282600.0 1331400.0 ;
      RECT  272400.0 1345200.0 282600.0 1331400.0 ;
      RECT  272400.0 1345200.0 282600.0 1359000.0 ;
      RECT  272400.0 1372800.0 282600.0 1359000.0 ;
      RECT  272400.0 1372800.0 282600.0 1386600.0 ;
      RECT  272400.0 1400400.0 282600.0 1386600.0 ;
      RECT  272400.0 1400400.0 282600.0 1414200.0 ;
      RECT  272400.0 1428000.0 282600.0 1414200.0 ;
      RECT  272400.0 1428000.0 282600.0 1441800.0 ;
      RECT  272400.0 1455600.0 282600.0 1441800.0 ;
      RECT  272400.0 1455600.0 282600.0 1469400.0 ;
      RECT  272400.0 1483200.0 282600.0 1469400.0 ;
      RECT  272400.0 1483200.0 282600.0 1497000.0 ;
      RECT  272400.0 1510800.0 282600.0 1497000.0 ;
      RECT  272400.0 1510800.0 282600.0 1524600.0 ;
      RECT  272400.0 1538400.0 282600.0 1524600.0 ;
      RECT  272400.0 1538400.0 282600.0 1552200.0 ;
      RECT  272400.0 1566000.0 282600.0 1552200.0 ;
      RECT  272400.0 1566000.0 282600.0 1579800.0 ;
      RECT  272400.0 1593600.0 282600.0 1579800.0 ;
      RECT  272400.0 1593600.0 282600.0 1607400.0 ;
      RECT  272400.0 1621200.0 282600.0 1607400.0 ;
      RECT  272400.0 1621200.0 282600.0 1635000.0 ;
      RECT  272400.0 1648800.0 282600.0 1635000.0 ;
      RECT  272400.0 1648800.0 282600.0 1662600.0 ;
      RECT  272400.0 1676400.0 282600.0 1662600.0 ;
      RECT  272400.0 1676400.0 282600.0 1690200.0 ;
      RECT  272400.0 1704000.0 282600.0 1690200.0 ;
      RECT  272400.0 1704000.0 282600.0 1717800.0 ;
      RECT  272400.0 1731600.0 282600.0 1717800.0 ;
      RECT  272400.0 1731600.0 282600.0 1745400.0 ;
      RECT  272400.0 1759200.0 282600.0 1745400.0 ;
      RECT  272400.0 1759200.0 282600.0 1773000.0 ;
      RECT  272400.0 1786800.0 282600.0 1773000.0 ;
      RECT  272400.0 1786800.0 282600.0 1800600.0 ;
      RECT  272400.0 1814400.0 282600.0 1800600.0 ;
      RECT  272400.0 1814400.0 282600.0 1828200.0 ;
      RECT  272400.0 1842000.0 282600.0 1828200.0 ;
      RECT  272400.0 1842000.0 282600.0 1855800.0 ;
      RECT  272400.0 1869600.0 282600.0 1855800.0 ;
      RECT  272400.0 1869600.0 282600.0 1883400.0 ;
      RECT  272400.0 1897200.0 282600.0 1883400.0 ;
      RECT  272400.0 1897200.0 282600.0 1911000.0 ;
      RECT  272400.0 1924800.0 282600.0 1911000.0 ;
      RECT  272400.0 1924800.0 282600.0 1938600.0 ;
      RECT  272400.0 1952400.0 282600.0 1938600.0 ;
      RECT  272400.0 1952400.0 282600.0 1966200.0 ;
      RECT  272400.0 1980000.0 282600.0 1966200.0 ;
      RECT  272400.0 1980000.0 282600.0 1993800.0 ;
      RECT  272400.0 2007600.0 282600.0 1993800.0 ;
      RECT  272400.0 2007600.0 282600.0 2021400.0 ;
      RECT  272400.0 2035200.0 282600.0 2021400.0 ;
      RECT  272400.0 2035200.0 282600.0 2049000.0 ;
      RECT  272400.0 2062800.0 282600.0 2049000.0 ;
      RECT  272400.0 2062800.0 282600.0 2076600.0 ;
      RECT  272400.0 2090400.0 282600.0 2076600.0 ;
      RECT  272400.0 2090400.0 282600.0 2104200.0 ;
      RECT  272400.0 2118000.0 282600.0 2104200.0 ;
      RECT  272400.0 2118000.0 282600.0 2131800.0 ;
      RECT  272400.0 2145600.0 282600.0 2131800.0 ;
      RECT  282600.0 379200.0 292800.0 393000.0 ;
      RECT  282600.0 406800.0 292800.0 393000.0 ;
      RECT  282600.0 406800.0 292800.0 420600.0 ;
      RECT  282600.0 434400.0 292800.0 420600.0 ;
      RECT  282600.0 434400.0 292800.0 448200.0 ;
      RECT  282600.0 462000.0 292800.0 448200.0 ;
      RECT  282600.0 462000.0 292800.0 475800.0 ;
      RECT  282600.0 489600.0 292800.0 475800.0 ;
      RECT  282600.0 489600.0 292800.0 503400.0 ;
      RECT  282600.0 517200.0 292800.0 503400.0 ;
      RECT  282600.0 517200.0 292800.0 531000.0 ;
      RECT  282600.0 544800.0 292800.0 531000.0 ;
      RECT  282600.0 544800.0 292800.0 558600.0 ;
      RECT  282600.0 572400.0 292800.0 558600.0 ;
      RECT  282600.0 572400.0 292800.0 586200.0 ;
      RECT  282600.0 600000.0 292800.0 586200.0 ;
      RECT  282600.0 600000.0 292800.0 613800.0 ;
      RECT  282600.0 627600.0 292800.0 613800.0 ;
      RECT  282600.0 627600.0 292800.0 641400.0 ;
      RECT  282600.0 655200.0 292800.0 641400.0 ;
      RECT  282600.0 655200.0 292800.0 669000.0 ;
      RECT  282600.0 682800.0 292800.0 669000.0 ;
      RECT  282600.0 682800.0 292800.0 696600.0 ;
      RECT  282600.0 710400.0 292800.0 696600.0 ;
      RECT  282600.0 710400.0 292800.0 724200.0 ;
      RECT  282600.0 738000.0 292800.0 724200.0 ;
      RECT  282600.0 738000.0 292800.0 751800.0 ;
      RECT  282600.0 765600.0 292800.0 751800.0 ;
      RECT  282600.0 765600.0 292800.0 779400.0 ;
      RECT  282600.0 793200.0 292800.0 779400.0 ;
      RECT  282600.0 793200.0 292800.0 807000.0 ;
      RECT  282600.0 820800.0 292800.0 807000.0 ;
      RECT  282600.0 820800.0 292800.0 834600.0 ;
      RECT  282600.0 848400.0 292800.0 834600.0 ;
      RECT  282600.0 848400.0 292800.0 862200.0 ;
      RECT  282600.0 876000.0 292800.0 862200.0 ;
      RECT  282600.0 876000.0 292800.0 889800.0 ;
      RECT  282600.0 903600.0 292800.0 889800.0 ;
      RECT  282600.0 903600.0 292800.0 917400.0 ;
      RECT  282600.0 931200.0 292800.0 917400.0 ;
      RECT  282600.0 931200.0 292800.0 945000.0 ;
      RECT  282600.0 958800.0 292800.0 945000.0 ;
      RECT  282600.0 958800.0 292800.0 972600.0 ;
      RECT  282600.0 986400.0 292800.0 972600.0 ;
      RECT  282600.0 986400.0 292800.0 1000200.0 ;
      RECT  282600.0 1014000.0 292800.0 1000200.0 ;
      RECT  282600.0 1014000.0 292800.0 1027800.0 ;
      RECT  282600.0 1041600.0 292800.0 1027800.0 ;
      RECT  282600.0 1041600.0 292800.0 1055400.0 ;
      RECT  282600.0 1069200.0 292800.0 1055400.0 ;
      RECT  282600.0 1069200.0 292800.0 1083000.0 ;
      RECT  282600.0 1096800.0 292800.0 1083000.0 ;
      RECT  282600.0 1096800.0 292800.0 1110600.0 ;
      RECT  282600.0 1124400.0 292800.0 1110600.0 ;
      RECT  282600.0 1124400.0 292800.0 1138200.0 ;
      RECT  282600.0 1152000.0 292800.0 1138200.0 ;
      RECT  282600.0 1152000.0 292800.0 1165800.0 ;
      RECT  282600.0 1179600.0 292800.0 1165800.0 ;
      RECT  282600.0 1179600.0 292800.0 1193400.0 ;
      RECT  282600.0 1207200.0 292800.0 1193400.0 ;
      RECT  282600.0 1207200.0 292800.0 1221000.0 ;
      RECT  282600.0 1234800.0 292800.0 1221000.0 ;
      RECT  282600.0 1234800.0 292800.0 1248600.0 ;
      RECT  282600.0 1262400.0 292800.0 1248600.0 ;
      RECT  282600.0 1262400.0 292800.0 1276200.0 ;
      RECT  282600.0 1290000.0 292800.0 1276200.0 ;
      RECT  282600.0 1290000.0 292800.0 1303800.0 ;
      RECT  282600.0 1317600.0 292800.0 1303800.0 ;
      RECT  282600.0 1317600.0 292800.0 1331400.0 ;
      RECT  282600.0 1345200.0 292800.0 1331400.0 ;
      RECT  282600.0 1345200.0 292800.0 1359000.0 ;
      RECT  282600.0 1372800.0 292800.0 1359000.0 ;
      RECT  282600.0 1372800.0 292800.0 1386600.0 ;
      RECT  282600.0 1400400.0 292800.0 1386600.0 ;
      RECT  282600.0 1400400.0 292800.0 1414200.0 ;
      RECT  282600.0 1428000.0 292800.0 1414200.0 ;
      RECT  282600.0 1428000.0 292800.0 1441800.0 ;
      RECT  282600.0 1455600.0 292800.0 1441800.0 ;
      RECT  282600.0 1455600.0 292800.0 1469400.0 ;
      RECT  282600.0 1483200.0 292800.0 1469400.0 ;
      RECT  282600.0 1483200.0 292800.0 1497000.0 ;
      RECT  282600.0 1510800.0 292800.0 1497000.0 ;
      RECT  282600.0 1510800.0 292800.0 1524600.0 ;
      RECT  282600.0 1538400.0 292800.0 1524600.0 ;
      RECT  282600.0 1538400.0 292800.0 1552200.0 ;
      RECT  282600.0 1566000.0 292800.0 1552200.0 ;
      RECT  282600.0 1566000.0 292800.0 1579800.0 ;
      RECT  282600.0 1593600.0 292800.0 1579800.0 ;
      RECT  282600.0 1593600.0 292800.0 1607400.0 ;
      RECT  282600.0 1621200.0 292800.0 1607400.0 ;
      RECT  282600.0 1621200.0 292800.0 1635000.0 ;
      RECT  282600.0 1648800.0 292800.0 1635000.0 ;
      RECT  282600.0 1648800.0 292800.0 1662600.0 ;
      RECT  282600.0 1676400.0 292800.0 1662600.0 ;
      RECT  282600.0 1676400.0 292800.0 1690200.0 ;
      RECT  282600.0 1704000.0 292800.0 1690200.0 ;
      RECT  282600.0 1704000.0 292800.0 1717800.0 ;
      RECT  282600.0 1731600.0 292800.0 1717800.0 ;
      RECT  282600.0 1731600.0 292800.0 1745400.0 ;
      RECT  282600.0 1759200.0 292800.0 1745400.0 ;
      RECT  282600.0 1759200.0 292800.0 1773000.0 ;
      RECT  282600.0 1786800.0 292800.0 1773000.0 ;
      RECT  282600.0 1786800.0 292800.0 1800600.0 ;
      RECT  282600.0 1814400.0 292800.0 1800600.0 ;
      RECT  282600.0 1814400.0 292800.0 1828200.0 ;
      RECT  282600.0 1842000.0 292800.0 1828200.0 ;
      RECT  282600.0 1842000.0 292800.0 1855800.0 ;
      RECT  282600.0 1869600.0 292800.0 1855800.0 ;
      RECT  282600.0 1869600.0 292800.0 1883400.0 ;
      RECT  282600.0 1897200.0 292800.0 1883400.0 ;
      RECT  282600.0 1897200.0 292800.0 1911000.0 ;
      RECT  282600.0 1924800.0 292800.0 1911000.0 ;
      RECT  282600.0 1924800.0 292800.0 1938600.0 ;
      RECT  282600.0 1952400.0 292800.0 1938600.0 ;
      RECT  282600.0 1952400.0 292800.0 1966200.0 ;
      RECT  282600.0 1980000.0 292800.0 1966200.0 ;
      RECT  282600.0 1980000.0 292800.0 1993800.0 ;
      RECT  282600.0 2007600.0 292800.0 1993800.0 ;
      RECT  282600.0 2007600.0 292800.0 2021400.0 ;
      RECT  282600.0 2035200.0 292800.0 2021400.0 ;
      RECT  282600.0 2035200.0 292800.0 2049000.0 ;
      RECT  282600.0 2062800.0 292800.0 2049000.0 ;
      RECT  282600.0 2062800.0 292800.0 2076600.0 ;
      RECT  282600.0 2090400.0 292800.0 2076600.0 ;
      RECT  282600.0 2090400.0 292800.0 2104200.0 ;
      RECT  282600.0 2118000.0 292800.0 2104200.0 ;
      RECT  282600.0 2118000.0 292800.0 2131800.0 ;
      RECT  282600.0 2145600.0 292800.0 2131800.0 ;
      RECT  292800.0 379200.0 303000.0 393000.0 ;
      RECT  292800.0 406800.0 303000.0 393000.0 ;
      RECT  292800.0 406800.0 303000.0 420600.0 ;
      RECT  292800.0 434400.0 303000.0 420600.0 ;
      RECT  292800.0 434400.0 303000.0 448200.0 ;
      RECT  292800.0 462000.0 303000.0 448200.0 ;
      RECT  292800.0 462000.0 303000.0 475800.0 ;
      RECT  292800.0 489600.0 303000.0 475800.0 ;
      RECT  292800.0 489600.0 303000.0 503400.0 ;
      RECT  292800.0 517200.0 303000.0 503400.0 ;
      RECT  292800.0 517200.0 303000.0 531000.0 ;
      RECT  292800.0 544800.0 303000.0 531000.0 ;
      RECT  292800.0 544800.0 303000.0 558600.0 ;
      RECT  292800.0 572400.0 303000.0 558600.0 ;
      RECT  292800.0 572400.0 303000.0 586200.0 ;
      RECT  292800.0 600000.0 303000.0 586200.0 ;
      RECT  292800.0 600000.0 303000.0 613800.0 ;
      RECT  292800.0 627600.0 303000.0 613800.0 ;
      RECT  292800.0 627600.0 303000.0 641400.0 ;
      RECT  292800.0 655200.0 303000.0 641400.0 ;
      RECT  292800.0 655200.0 303000.0 669000.0 ;
      RECT  292800.0 682800.0 303000.0 669000.0 ;
      RECT  292800.0 682800.0 303000.0 696600.0 ;
      RECT  292800.0 710400.0 303000.0 696600.0 ;
      RECT  292800.0 710400.0 303000.0 724200.0 ;
      RECT  292800.0 738000.0 303000.0 724200.0 ;
      RECT  292800.0 738000.0 303000.0 751800.0 ;
      RECT  292800.0 765600.0 303000.0 751800.0 ;
      RECT  292800.0 765600.0 303000.0 779400.0 ;
      RECT  292800.0 793200.0 303000.0 779400.0 ;
      RECT  292800.0 793200.0 303000.0 807000.0 ;
      RECT  292800.0 820800.0 303000.0 807000.0 ;
      RECT  292800.0 820800.0 303000.0 834600.0 ;
      RECT  292800.0 848400.0 303000.0 834600.0 ;
      RECT  292800.0 848400.0 303000.0 862200.0 ;
      RECT  292800.0 876000.0 303000.0 862200.0 ;
      RECT  292800.0 876000.0 303000.0 889800.0 ;
      RECT  292800.0 903600.0 303000.0 889800.0 ;
      RECT  292800.0 903600.0 303000.0 917400.0 ;
      RECT  292800.0 931200.0 303000.0 917400.0 ;
      RECT  292800.0 931200.0 303000.0 945000.0 ;
      RECT  292800.0 958800.0 303000.0 945000.0 ;
      RECT  292800.0 958800.0 303000.0 972600.0 ;
      RECT  292800.0 986400.0 303000.0 972600.0 ;
      RECT  292800.0 986400.0 303000.0 1000200.0 ;
      RECT  292800.0 1014000.0 303000.0 1000200.0 ;
      RECT  292800.0 1014000.0 303000.0 1027800.0 ;
      RECT  292800.0 1041600.0 303000.0 1027800.0 ;
      RECT  292800.0 1041600.0 303000.0 1055400.0 ;
      RECT  292800.0 1069200.0 303000.0 1055400.0 ;
      RECT  292800.0 1069200.0 303000.0 1083000.0 ;
      RECT  292800.0 1096800.0 303000.0 1083000.0 ;
      RECT  292800.0 1096800.0 303000.0 1110600.0 ;
      RECT  292800.0 1124400.0 303000.0 1110600.0 ;
      RECT  292800.0 1124400.0 303000.0 1138200.0 ;
      RECT  292800.0 1152000.0 303000.0 1138200.0 ;
      RECT  292800.0 1152000.0 303000.0 1165800.0 ;
      RECT  292800.0 1179600.0 303000.0 1165800.0 ;
      RECT  292800.0 1179600.0 303000.0 1193400.0 ;
      RECT  292800.0 1207200.0 303000.0 1193400.0 ;
      RECT  292800.0 1207200.0 303000.0 1221000.0 ;
      RECT  292800.0 1234800.0 303000.0 1221000.0 ;
      RECT  292800.0 1234800.0 303000.0 1248600.0 ;
      RECT  292800.0 1262400.0 303000.0 1248600.0 ;
      RECT  292800.0 1262400.0 303000.0 1276200.0 ;
      RECT  292800.0 1290000.0 303000.0 1276200.0 ;
      RECT  292800.0 1290000.0 303000.0 1303800.0 ;
      RECT  292800.0 1317600.0 303000.0 1303800.0 ;
      RECT  292800.0 1317600.0 303000.0 1331400.0 ;
      RECT  292800.0 1345200.0 303000.0 1331400.0 ;
      RECT  292800.0 1345200.0 303000.0 1359000.0 ;
      RECT  292800.0 1372800.0 303000.0 1359000.0 ;
      RECT  292800.0 1372800.0 303000.0 1386600.0 ;
      RECT  292800.0 1400400.0 303000.0 1386600.0 ;
      RECT  292800.0 1400400.0 303000.0 1414200.0 ;
      RECT  292800.0 1428000.0 303000.0 1414200.0 ;
      RECT  292800.0 1428000.0 303000.0 1441800.0 ;
      RECT  292800.0 1455600.0 303000.0 1441800.0 ;
      RECT  292800.0 1455600.0 303000.0 1469400.0 ;
      RECT  292800.0 1483200.0 303000.0 1469400.0 ;
      RECT  292800.0 1483200.0 303000.0 1497000.0 ;
      RECT  292800.0 1510800.0 303000.0 1497000.0 ;
      RECT  292800.0 1510800.0 303000.0 1524600.0 ;
      RECT  292800.0 1538400.0 303000.0 1524600.0 ;
      RECT  292800.0 1538400.0 303000.0 1552200.0 ;
      RECT  292800.0 1566000.0 303000.0 1552200.0 ;
      RECT  292800.0 1566000.0 303000.0 1579800.0 ;
      RECT  292800.0 1593600.0 303000.0 1579800.0 ;
      RECT  292800.0 1593600.0 303000.0 1607400.0 ;
      RECT  292800.0 1621200.0 303000.0 1607400.0 ;
      RECT  292800.0 1621200.0 303000.0 1635000.0 ;
      RECT  292800.0 1648800.0 303000.0 1635000.0 ;
      RECT  292800.0 1648800.0 303000.0 1662600.0 ;
      RECT  292800.0 1676400.0 303000.0 1662600.0 ;
      RECT  292800.0 1676400.0 303000.0 1690200.0 ;
      RECT  292800.0 1704000.0 303000.0 1690200.0 ;
      RECT  292800.0 1704000.0 303000.0 1717800.0 ;
      RECT  292800.0 1731600.0 303000.0 1717800.0 ;
      RECT  292800.0 1731600.0 303000.0 1745400.0 ;
      RECT  292800.0 1759200.0 303000.0 1745400.0 ;
      RECT  292800.0 1759200.0 303000.0 1773000.0 ;
      RECT  292800.0 1786800.0 303000.0 1773000.0 ;
      RECT  292800.0 1786800.0 303000.0 1800600.0 ;
      RECT  292800.0 1814400.0 303000.0 1800600.0 ;
      RECT  292800.0 1814400.0 303000.0 1828200.0 ;
      RECT  292800.0 1842000.0 303000.0 1828200.0 ;
      RECT  292800.0 1842000.0 303000.0 1855800.0 ;
      RECT  292800.0 1869600.0 303000.0 1855800.0 ;
      RECT  292800.0 1869600.0 303000.0 1883400.0 ;
      RECT  292800.0 1897200.0 303000.0 1883400.0 ;
      RECT  292800.0 1897200.0 303000.0 1911000.0 ;
      RECT  292800.0 1924800.0 303000.0 1911000.0 ;
      RECT  292800.0 1924800.0 303000.0 1938600.0 ;
      RECT  292800.0 1952400.0 303000.0 1938600.0 ;
      RECT  292800.0 1952400.0 303000.0 1966200.0 ;
      RECT  292800.0 1980000.0 303000.0 1966200.0 ;
      RECT  292800.0 1980000.0 303000.0 1993800.0 ;
      RECT  292800.0 2007600.0 303000.0 1993800.0 ;
      RECT  292800.0 2007600.0 303000.0 2021400.0 ;
      RECT  292800.0 2035200.0 303000.0 2021400.0 ;
      RECT  292800.0 2035200.0 303000.0 2049000.0 ;
      RECT  292800.0 2062800.0 303000.0 2049000.0 ;
      RECT  292800.0 2062800.0 303000.0 2076600.0 ;
      RECT  292800.0 2090400.0 303000.0 2076600.0 ;
      RECT  292800.0 2090400.0 303000.0 2104200.0 ;
      RECT  292800.0 2118000.0 303000.0 2104200.0 ;
      RECT  292800.0 2118000.0 303000.0 2131800.0 ;
      RECT  292800.0 2145600.0 303000.0 2131800.0 ;
      RECT  303000.0 379200.0 313200.0 393000.0 ;
      RECT  303000.0 406800.0 313200.0 393000.0 ;
      RECT  303000.0 406800.0 313200.0 420600.0 ;
      RECT  303000.0 434400.0 313200.0 420600.0 ;
      RECT  303000.0 434400.0 313200.0 448200.0 ;
      RECT  303000.0 462000.0 313200.0 448200.0 ;
      RECT  303000.0 462000.0 313200.0 475800.0 ;
      RECT  303000.0 489600.0 313200.0 475800.0 ;
      RECT  303000.0 489600.0 313200.0 503400.0 ;
      RECT  303000.0 517200.0 313200.0 503400.0 ;
      RECT  303000.0 517200.0 313200.0 531000.0 ;
      RECT  303000.0 544800.0 313200.0 531000.0 ;
      RECT  303000.0 544800.0 313200.0 558600.0 ;
      RECT  303000.0 572400.0 313200.0 558600.0 ;
      RECT  303000.0 572400.0 313200.0 586200.0 ;
      RECT  303000.0 600000.0 313200.0 586200.0 ;
      RECT  303000.0 600000.0 313200.0 613800.0 ;
      RECT  303000.0 627600.0 313200.0 613800.0 ;
      RECT  303000.0 627600.0 313200.0 641400.0 ;
      RECT  303000.0 655200.0 313200.0 641400.0 ;
      RECT  303000.0 655200.0 313200.0 669000.0 ;
      RECT  303000.0 682800.0 313200.0 669000.0 ;
      RECT  303000.0 682800.0 313200.0 696600.0 ;
      RECT  303000.0 710400.0 313200.0 696600.0 ;
      RECT  303000.0 710400.0 313200.0 724200.0 ;
      RECT  303000.0 738000.0 313200.0 724200.0 ;
      RECT  303000.0 738000.0 313200.0 751800.0 ;
      RECT  303000.0 765600.0 313200.0 751800.0 ;
      RECT  303000.0 765600.0 313200.0 779400.0 ;
      RECT  303000.0 793200.0 313200.0 779400.0 ;
      RECT  303000.0 793200.0 313200.0 807000.0 ;
      RECT  303000.0 820800.0 313200.0 807000.0 ;
      RECT  303000.0 820800.0 313200.0 834600.0 ;
      RECT  303000.0 848400.0 313200.0 834600.0 ;
      RECT  303000.0 848400.0 313200.0 862200.0 ;
      RECT  303000.0 876000.0 313200.0 862200.0 ;
      RECT  303000.0 876000.0 313200.0 889800.0 ;
      RECT  303000.0 903600.0 313200.0 889800.0 ;
      RECT  303000.0 903600.0 313200.0 917400.0 ;
      RECT  303000.0 931200.0 313200.0 917400.0 ;
      RECT  303000.0 931200.0 313200.0 945000.0 ;
      RECT  303000.0 958800.0 313200.0 945000.0 ;
      RECT  303000.0 958800.0 313200.0 972600.0 ;
      RECT  303000.0 986400.0 313200.0 972600.0 ;
      RECT  303000.0 986400.0 313200.0 1000200.0 ;
      RECT  303000.0 1014000.0 313200.0 1000200.0 ;
      RECT  303000.0 1014000.0 313200.0 1027800.0 ;
      RECT  303000.0 1041600.0 313200.0 1027800.0 ;
      RECT  303000.0 1041600.0 313200.0 1055400.0 ;
      RECT  303000.0 1069200.0 313200.0 1055400.0 ;
      RECT  303000.0 1069200.0 313200.0 1083000.0 ;
      RECT  303000.0 1096800.0 313200.0 1083000.0 ;
      RECT  303000.0 1096800.0 313200.0 1110600.0 ;
      RECT  303000.0 1124400.0 313200.0 1110600.0 ;
      RECT  303000.0 1124400.0 313200.0 1138200.0 ;
      RECT  303000.0 1152000.0 313200.0 1138200.0 ;
      RECT  303000.0 1152000.0 313200.0 1165800.0 ;
      RECT  303000.0 1179600.0 313200.0 1165800.0 ;
      RECT  303000.0 1179600.0 313200.0 1193400.0 ;
      RECT  303000.0 1207200.0 313200.0 1193400.0 ;
      RECT  303000.0 1207200.0 313200.0 1221000.0 ;
      RECT  303000.0 1234800.0 313200.0 1221000.0 ;
      RECT  303000.0 1234800.0 313200.0 1248600.0 ;
      RECT  303000.0 1262400.0 313200.0 1248600.0 ;
      RECT  303000.0 1262400.0 313200.0 1276200.0 ;
      RECT  303000.0 1290000.0 313200.0 1276200.0 ;
      RECT  303000.0 1290000.0 313200.0 1303800.0 ;
      RECT  303000.0 1317600.0 313200.0 1303800.0 ;
      RECT  303000.0 1317600.0 313200.0 1331400.0 ;
      RECT  303000.0 1345200.0 313200.0 1331400.0 ;
      RECT  303000.0 1345200.0 313200.0 1359000.0 ;
      RECT  303000.0 1372800.0 313200.0 1359000.0 ;
      RECT  303000.0 1372800.0 313200.0 1386600.0 ;
      RECT  303000.0 1400400.0 313200.0 1386600.0 ;
      RECT  303000.0 1400400.0 313200.0 1414200.0 ;
      RECT  303000.0 1428000.0 313200.0 1414200.0 ;
      RECT  303000.0 1428000.0 313200.0 1441800.0 ;
      RECT  303000.0 1455600.0 313200.0 1441800.0 ;
      RECT  303000.0 1455600.0 313200.0 1469400.0 ;
      RECT  303000.0 1483200.0 313200.0 1469400.0 ;
      RECT  303000.0 1483200.0 313200.0 1497000.0 ;
      RECT  303000.0 1510800.0 313200.0 1497000.0 ;
      RECT  303000.0 1510800.0 313200.0 1524600.0 ;
      RECT  303000.0 1538400.0 313200.0 1524600.0 ;
      RECT  303000.0 1538400.0 313200.0 1552200.0 ;
      RECT  303000.0 1566000.0 313200.0 1552200.0 ;
      RECT  303000.0 1566000.0 313200.0 1579800.0 ;
      RECT  303000.0 1593600.0 313200.0 1579800.0 ;
      RECT  303000.0 1593600.0 313200.0 1607400.0 ;
      RECT  303000.0 1621200.0 313200.0 1607400.0 ;
      RECT  303000.0 1621200.0 313200.0 1635000.0 ;
      RECT  303000.0 1648800.0 313200.0 1635000.0 ;
      RECT  303000.0 1648800.0 313200.0 1662600.0 ;
      RECT  303000.0 1676400.0 313200.0 1662600.0 ;
      RECT  303000.0 1676400.0 313200.0 1690200.0 ;
      RECT  303000.0 1704000.0 313200.0 1690200.0 ;
      RECT  303000.0 1704000.0 313200.0 1717800.0 ;
      RECT  303000.0 1731600.0 313200.0 1717800.0 ;
      RECT  303000.0 1731600.0 313200.0 1745400.0 ;
      RECT  303000.0 1759200.0 313200.0 1745400.0 ;
      RECT  303000.0 1759200.0 313200.0 1773000.0 ;
      RECT  303000.0 1786800.0 313200.0 1773000.0 ;
      RECT  303000.0 1786800.0 313200.0 1800600.0 ;
      RECT  303000.0 1814400.0 313200.0 1800600.0 ;
      RECT  303000.0 1814400.0 313200.0 1828200.0 ;
      RECT  303000.0 1842000.0 313200.0 1828200.0 ;
      RECT  303000.0 1842000.0 313200.0 1855800.0 ;
      RECT  303000.0 1869600.0 313200.0 1855800.0 ;
      RECT  303000.0 1869600.0 313200.0 1883400.0 ;
      RECT  303000.0 1897200.0 313200.0 1883400.0 ;
      RECT  303000.0 1897200.0 313200.0 1911000.0 ;
      RECT  303000.0 1924800.0 313200.0 1911000.0 ;
      RECT  303000.0 1924800.0 313200.0 1938600.0 ;
      RECT  303000.0 1952400.0 313200.0 1938600.0 ;
      RECT  303000.0 1952400.0 313200.0 1966200.0 ;
      RECT  303000.0 1980000.0 313200.0 1966200.0 ;
      RECT  303000.0 1980000.0 313200.0 1993800.0 ;
      RECT  303000.0 2007600.0 313200.0 1993800.0 ;
      RECT  303000.0 2007600.0 313200.0 2021400.0 ;
      RECT  303000.0 2035200.0 313200.0 2021400.0 ;
      RECT  303000.0 2035200.0 313200.0 2049000.0 ;
      RECT  303000.0 2062800.0 313200.0 2049000.0 ;
      RECT  303000.0 2062800.0 313200.0 2076600.0 ;
      RECT  303000.0 2090400.0 313200.0 2076600.0 ;
      RECT  303000.0 2090400.0 313200.0 2104200.0 ;
      RECT  303000.0 2118000.0 313200.0 2104200.0 ;
      RECT  303000.0 2118000.0 313200.0 2131800.0 ;
      RECT  303000.0 2145600.0 313200.0 2131800.0 ;
      RECT  313200.0 379200.0 323400.0 393000.0 ;
      RECT  313200.0 406800.0 323400.0 393000.0 ;
      RECT  313200.0 406800.0 323400.0 420600.0 ;
      RECT  313200.0 434400.0 323400.0 420600.0 ;
      RECT  313200.0 434400.0 323400.0 448200.0 ;
      RECT  313200.0 462000.0 323400.0 448200.0 ;
      RECT  313200.0 462000.0 323400.0 475800.0 ;
      RECT  313200.0 489600.0 323400.0 475800.0 ;
      RECT  313200.0 489600.0 323400.0 503400.0 ;
      RECT  313200.0 517200.0 323400.0 503400.0 ;
      RECT  313200.0 517200.0 323400.0 531000.0 ;
      RECT  313200.0 544800.0 323400.0 531000.0 ;
      RECT  313200.0 544800.0 323400.0 558600.0 ;
      RECT  313200.0 572400.0 323400.0 558600.0 ;
      RECT  313200.0 572400.0 323400.0 586200.0 ;
      RECT  313200.0 600000.0 323400.0 586200.0 ;
      RECT  313200.0 600000.0 323400.0 613800.0 ;
      RECT  313200.0 627600.0 323400.0 613800.0 ;
      RECT  313200.0 627600.0 323400.0 641400.0 ;
      RECT  313200.0 655200.0 323400.0 641400.0 ;
      RECT  313200.0 655200.0 323400.0 669000.0 ;
      RECT  313200.0 682800.0 323400.0 669000.0 ;
      RECT  313200.0 682800.0 323400.0 696600.0 ;
      RECT  313200.0 710400.0 323400.0 696600.0 ;
      RECT  313200.0 710400.0 323400.0 724200.0 ;
      RECT  313200.0 738000.0 323400.0 724200.0 ;
      RECT  313200.0 738000.0 323400.0 751800.0 ;
      RECT  313200.0 765600.0 323400.0 751800.0 ;
      RECT  313200.0 765600.0 323400.0 779400.0 ;
      RECT  313200.0 793200.0 323400.0 779400.0 ;
      RECT  313200.0 793200.0 323400.0 807000.0 ;
      RECT  313200.0 820800.0 323400.0 807000.0 ;
      RECT  313200.0 820800.0 323400.0 834600.0 ;
      RECT  313200.0 848400.0 323400.0 834600.0 ;
      RECT  313200.0 848400.0 323400.0 862200.0 ;
      RECT  313200.0 876000.0 323400.0 862200.0 ;
      RECT  313200.0 876000.0 323400.0 889800.0 ;
      RECT  313200.0 903600.0 323400.0 889800.0 ;
      RECT  313200.0 903600.0 323400.0 917400.0 ;
      RECT  313200.0 931200.0 323400.0 917400.0 ;
      RECT  313200.0 931200.0 323400.0 945000.0 ;
      RECT  313200.0 958800.0 323400.0 945000.0 ;
      RECT  313200.0 958800.0 323400.0 972600.0 ;
      RECT  313200.0 986400.0 323400.0 972600.0 ;
      RECT  313200.0 986400.0 323400.0 1000200.0 ;
      RECT  313200.0 1014000.0 323400.0 1000200.0 ;
      RECT  313200.0 1014000.0 323400.0 1027800.0 ;
      RECT  313200.0 1041600.0 323400.0 1027800.0 ;
      RECT  313200.0 1041600.0 323400.0 1055400.0 ;
      RECT  313200.0 1069200.0 323400.0 1055400.0 ;
      RECT  313200.0 1069200.0 323400.0 1083000.0 ;
      RECT  313200.0 1096800.0 323400.0 1083000.0 ;
      RECT  313200.0 1096800.0 323400.0 1110600.0 ;
      RECT  313200.0 1124400.0 323400.0 1110600.0 ;
      RECT  313200.0 1124400.0 323400.0 1138200.0 ;
      RECT  313200.0 1152000.0 323400.0 1138200.0 ;
      RECT  313200.0 1152000.0 323400.0 1165800.0 ;
      RECT  313200.0 1179600.0 323400.0 1165800.0 ;
      RECT  313200.0 1179600.0 323400.0 1193400.0 ;
      RECT  313200.0 1207200.0 323400.0 1193400.0 ;
      RECT  313200.0 1207200.0 323400.0 1221000.0 ;
      RECT  313200.0 1234800.0 323400.0 1221000.0 ;
      RECT  313200.0 1234800.0 323400.0 1248600.0 ;
      RECT  313200.0 1262400.0 323400.0 1248600.0 ;
      RECT  313200.0 1262400.0 323400.0 1276200.0 ;
      RECT  313200.0 1290000.0 323400.0 1276200.0 ;
      RECT  313200.0 1290000.0 323400.0 1303800.0 ;
      RECT  313200.0 1317600.0 323400.0 1303800.0 ;
      RECT  313200.0 1317600.0 323400.0 1331400.0 ;
      RECT  313200.0 1345200.0 323400.0 1331400.0 ;
      RECT  313200.0 1345200.0 323400.0 1359000.0 ;
      RECT  313200.0 1372800.0 323400.0 1359000.0 ;
      RECT  313200.0 1372800.0 323400.0 1386600.0 ;
      RECT  313200.0 1400400.0 323400.0 1386600.0 ;
      RECT  313200.0 1400400.0 323400.0 1414200.0 ;
      RECT  313200.0 1428000.0 323400.0 1414200.0 ;
      RECT  313200.0 1428000.0 323400.0 1441800.0 ;
      RECT  313200.0 1455600.0 323400.0 1441800.0 ;
      RECT  313200.0 1455600.0 323400.0 1469400.0 ;
      RECT  313200.0 1483200.0 323400.0 1469400.0 ;
      RECT  313200.0 1483200.0 323400.0 1497000.0 ;
      RECT  313200.0 1510800.0 323400.0 1497000.0 ;
      RECT  313200.0 1510800.0 323400.0 1524600.0 ;
      RECT  313200.0 1538400.0 323400.0 1524600.0 ;
      RECT  313200.0 1538400.0 323400.0 1552200.0 ;
      RECT  313200.0 1566000.0 323400.0 1552200.0 ;
      RECT  313200.0 1566000.0 323400.0 1579800.0 ;
      RECT  313200.0 1593600.0 323400.0 1579800.0 ;
      RECT  313200.0 1593600.0 323400.0 1607400.0 ;
      RECT  313200.0 1621200.0 323400.0 1607400.0 ;
      RECT  313200.0 1621200.0 323400.0 1635000.0 ;
      RECT  313200.0 1648800.0 323400.0 1635000.0 ;
      RECT  313200.0 1648800.0 323400.0 1662600.0 ;
      RECT  313200.0 1676400.0 323400.0 1662600.0 ;
      RECT  313200.0 1676400.0 323400.0 1690200.0 ;
      RECT  313200.0 1704000.0 323400.0 1690200.0 ;
      RECT  313200.0 1704000.0 323400.0 1717800.0 ;
      RECT  313200.0 1731600.0 323400.0 1717800.0 ;
      RECT  313200.0 1731600.0 323400.0 1745400.0 ;
      RECT  313200.0 1759200.0 323400.0 1745400.0 ;
      RECT  313200.0 1759200.0 323400.0 1773000.0 ;
      RECT  313200.0 1786800.0 323400.0 1773000.0 ;
      RECT  313200.0 1786800.0 323400.0 1800600.0 ;
      RECT  313200.0 1814400.0 323400.0 1800600.0 ;
      RECT  313200.0 1814400.0 323400.0 1828200.0 ;
      RECT  313200.0 1842000.0 323400.0 1828200.0 ;
      RECT  313200.0 1842000.0 323400.0 1855800.0 ;
      RECT  313200.0 1869600.0 323400.0 1855800.0 ;
      RECT  313200.0 1869600.0 323400.0 1883400.0 ;
      RECT  313200.0 1897200.0 323400.0 1883400.0 ;
      RECT  313200.0 1897200.0 323400.0 1911000.0 ;
      RECT  313200.0 1924800.0 323400.0 1911000.0 ;
      RECT  313200.0 1924800.0 323400.0 1938600.0 ;
      RECT  313200.0 1952400.0 323400.0 1938600.0 ;
      RECT  313200.0 1952400.0 323400.0 1966200.0 ;
      RECT  313200.0 1980000.0 323400.0 1966200.0 ;
      RECT  313200.0 1980000.0 323400.0 1993800.0 ;
      RECT  313200.0 2007600.0 323400.0 1993800.0 ;
      RECT  313200.0 2007600.0 323400.0 2021400.0 ;
      RECT  313200.0 2035200.0 323400.0 2021400.0 ;
      RECT  313200.0 2035200.0 323400.0 2049000.0 ;
      RECT  313200.0 2062800.0 323400.0 2049000.0 ;
      RECT  313200.0 2062800.0 323400.0 2076600.0 ;
      RECT  313200.0 2090400.0 323400.0 2076600.0 ;
      RECT  313200.0 2090400.0 323400.0 2104200.0 ;
      RECT  313200.0 2118000.0 323400.0 2104200.0 ;
      RECT  313200.0 2118000.0 323400.0 2131800.0 ;
      RECT  313200.0 2145600.0 323400.0 2131800.0 ;
      RECT  323400.0 379200.0 333600.0 393000.0 ;
      RECT  323400.0 406800.0 333600.0 393000.0 ;
      RECT  323400.0 406800.0 333600.0 420600.0 ;
      RECT  323400.0 434400.0 333600.0 420600.0 ;
      RECT  323400.0 434400.0 333600.0 448200.0 ;
      RECT  323400.0 462000.0 333600.0 448200.0 ;
      RECT  323400.0 462000.0 333600.0 475800.0 ;
      RECT  323400.0 489600.0 333600.0 475800.0 ;
      RECT  323400.0 489600.0 333600.0 503400.0 ;
      RECT  323400.0 517200.0 333600.0 503400.0 ;
      RECT  323400.0 517200.0 333600.0 531000.0 ;
      RECT  323400.0 544800.0 333600.0 531000.0 ;
      RECT  323400.0 544800.0 333600.0 558600.0 ;
      RECT  323400.0 572400.0 333600.0 558600.0 ;
      RECT  323400.0 572400.0 333600.0 586200.0 ;
      RECT  323400.0 600000.0 333600.0 586200.0 ;
      RECT  323400.0 600000.0 333600.0 613800.0 ;
      RECT  323400.0 627600.0 333600.0 613800.0 ;
      RECT  323400.0 627600.0 333600.0 641400.0 ;
      RECT  323400.0 655200.0 333600.0 641400.0 ;
      RECT  323400.0 655200.0 333600.0 669000.0 ;
      RECT  323400.0 682800.0 333600.0 669000.0 ;
      RECT  323400.0 682800.0 333600.0 696600.0 ;
      RECT  323400.0 710400.0 333600.0 696600.0 ;
      RECT  323400.0 710400.0 333600.0 724200.0 ;
      RECT  323400.0 738000.0 333600.0 724200.0 ;
      RECT  323400.0 738000.0 333600.0 751800.0 ;
      RECT  323400.0 765600.0 333600.0 751800.0 ;
      RECT  323400.0 765600.0 333600.0 779400.0 ;
      RECT  323400.0 793200.0 333600.0 779400.0 ;
      RECT  323400.0 793200.0 333600.0 807000.0 ;
      RECT  323400.0 820800.0 333600.0 807000.0 ;
      RECT  323400.0 820800.0 333600.0 834600.0 ;
      RECT  323400.0 848400.0 333600.0 834600.0 ;
      RECT  323400.0 848400.0 333600.0 862200.0 ;
      RECT  323400.0 876000.0 333600.0 862200.0 ;
      RECT  323400.0 876000.0 333600.0 889800.0 ;
      RECT  323400.0 903600.0 333600.0 889800.0 ;
      RECT  323400.0 903600.0 333600.0 917400.0 ;
      RECT  323400.0 931200.0 333600.0 917400.0 ;
      RECT  323400.0 931200.0 333600.0 945000.0 ;
      RECT  323400.0 958800.0 333600.0 945000.0 ;
      RECT  323400.0 958800.0 333600.0 972600.0 ;
      RECT  323400.0 986400.0 333600.0 972600.0 ;
      RECT  323400.0 986400.0 333600.0 1000200.0 ;
      RECT  323400.0 1014000.0 333600.0 1000200.0 ;
      RECT  323400.0 1014000.0 333600.0 1027800.0 ;
      RECT  323400.0 1041600.0 333600.0 1027800.0 ;
      RECT  323400.0 1041600.0 333600.0 1055400.0 ;
      RECT  323400.0 1069200.0 333600.0 1055400.0 ;
      RECT  323400.0 1069200.0 333600.0 1083000.0 ;
      RECT  323400.0 1096800.0 333600.0 1083000.0 ;
      RECT  323400.0 1096800.0 333600.0 1110600.0 ;
      RECT  323400.0 1124400.0 333600.0 1110600.0 ;
      RECT  323400.0 1124400.0 333600.0 1138200.0 ;
      RECT  323400.0 1152000.0 333600.0 1138200.0 ;
      RECT  323400.0 1152000.0 333600.0 1165800.0 ;
      RECT  323400.0 1179600.0 333600.0 1165800.0 ;
      RECT  323400.0 1179600.0 333600.0 1193400.0 ;
      RECT  323400.0 1207200.0 333600.0 1193400.0 ;
      RECT  323400.0 1207200.0 333600.0 1221000.0 ;
      RECT  323400.0 1234800.0 333600.0 1221000.0 ;
      RECT  323400.0 1234800.0 333600.0 1248600.0 ;
      RECT  323400.0 1262400.0 333600.0 1248600.0 ;
      RECT  323400.0 1262400.0 333600.0 1276200.0 ;
      RECT  323400.0 1290000.0 333600.0 1276200.0 ;
      RECT  323400.0 1290000.0 333600.0 1303800.0 ;
      RECT  323400.0 1317600.0 333600.0 1303800.0 ;
      RECT  323400.0 1317600.0 333600.0 1331400.0 ;
      RECT  323400.0 1345200.0 333600.0 1331400.0 ;
      RECT  323400.0 1345200.0 333600.0 1359000.0 ;
      RECT  323400.0 1372800.0 333600.0 1359000.0 ;
      RECT  323400.0 1372800.0 333600.0 1386600.0 ;
      RECT  323400.0 1400400.0 333600.0 1386600.0 ;
      RECT  323400.0 1400400.0 333600.0 1414200.0 ;
      RECT  323400.0 1428000.0 333600.0 1414200.0 ;
      RECT  323400.0 1428000.0 333600.0 1441800.0 ;
      RECT  323400.0 1455600.0 333600.0 1441800.0 ;
      RECT  323400.0 1455600.0 333600.0 1469400.0 ;
      RECT  323400.0 1483200.0 333600.0 1469400.0 ;
      RECT  323400.0 1483200.0 333600.0 1497000.0 ;
      RECT  323400.0 1510800.0 333600.0 1497000.0 ;
      RECT  323400.0 1510800.0 333600.0 1524600.0 ;
      RECT  323400.0 1538400.0 333600.0 1524600.0 ;
      RECT  323400.0 1538400.0 333600.0 1552200.0 ;
      RECT  323400.0 1566000.0 333600.0 1552200.0 ;
      RECT  323400.0 1566000.0 333600.0 1579800.0 ;
      RECT  323400.0 1593600.0 333600.0 1579800.0 ;
      RECT  323400.0 1593600.0 333600.0 1607400.0 ;
      RECT  323400.0 1621200.0 333600.0 1607400.0 ;
      RECT  323400.0 1621200.0 333600.0 1635000.0 ;
      RECT  323400.0 1648800.0 333600.0 1635000.0 ;
      RECT  323400.0 1648800.0 333600.0 1662600.0 ;
      RECT  323400.0 1676400.0 333600.0 1662600.0 ;
      RECT  323400.0 1676400.0 333600.0 1690200.0 ;
      RECT  323400.0 1704000.0 333600.0 1690200.0 ;
      RECT  323400.0 1704000.0 333600.0 1717800.0 ;
      RECT  323400.0 1731600.0 333600.0 1717800.0 ;
      RECT  323400.0 1731600.0 333600.0 1745400.0 ;
      RECT  323400.0 1759200.0 333600.0 1745400.0 ;
      RECT  323400.0 1759200.0 333600.0 1773000.0 ;
      RECT  323400.0 1786800.0 333600.0 1773000.0 ;
      RECT  323400.0 1786800.0 333600.0 1800600.0 ;
      RECT  323400.0 1814400.0 333600.0 1800600.0 ;
      RECT  323400.0 1814400.0 333600.0 1828200.0 ;
      RECT  323400.0 1842000.0 333600.0 1828200.0 ;
      RECT  323400.0 1842000.0 333600.0 1855800.0 ;
      RECT  323400.0 1869600.0 333600.0 1855800.0 ;
      RECT  323400.0 1869600.0 333600.0 1883400.0 ;
      RECT  323400.0 1897200.0 333600.0 1883400.0 ;
      RECT  323400.0 1897200.0 333600.0 1911000.0 ;
      RECT  323400.0 1924800.0 333600.0 1911000.0 ;
      RECT  323400.0 1924800.0 333600.0 1938600.0 ;
      RECT  323400.0 1952400.0 333600.0 1938600.0 ;
      RECT  323400.0 1952400.0 333600.0 1966200.0 ;
      RECT  323400.0 1980000.0 333600.0 1966200.0 ;
      RECT  323400.0 1980000.0 333600.0 1993800.0 ;
      RECT  323400.0 2007600.0 333600.0 1993800.0 ;
      RECT  323400.0 2007600.0 333600.0 2021400.0 ;
      RECT  323400.0 2035200.0 333600.0 2021400.0 ;
      RECT  323400.0 2035200.0 333600.0 2049000.0 ;
      RECT  323400.0 2062800.0 333600.0 2049000.0 ;
      RECT  323400.0 2062800.0 333600.0 2076600.0 ;
      RECT  323400.0 2090400.0 333600.0 2076600.0 ;
      RECT  323400.0 2090400.0 333600.0 2104200.0 ;
      RECT  323400.0 2118000.0 333600.0 2104200.0 ;
      RECT  323400.0 2118000.0 333600.0 2131800.0 ;
      RECT  323400.0 2145600.0 333600.0 2131800.0 ;
      RECT  333600.0 379200.0 343800.0 393000.0 ;
      RECT  333600.0 406800.0 343800.0 393000.0 ;
      RECT  333600.0 406800.0 343800.0 420600.0 ;
      RECT  333600.0 434400.0 343800.0 420600.0 ;
      RECT  333600.0 434400.0 343800.0 448200.0 ;
      RECT  333600.0 462000.0 343800.0 448200.0 ;
      RECT  333600.0 462000.0 343800.0 475800.0 ;
      RECT  333600.0 489600.0 343800.0 475800.0 ;
      RECT  333600.0 489600.0 343800.0 503400.0 ;
      RECT  333600.0 517200.0 343800.0 503400.0 ;
      RECT  333600.0 517200.0 343800.0 531000.0 ;
      RECT  333600.0 544800.0 343800.0 531000.0 ;
      RECT  333600.0 544800.0 343800.0 558600.0 ;
      RECT  333600.0 572400.0 343800.0 558600.0 ;
      RECT  333600.0 572400.0 343800.0 586200.0 ;
      RECT  333600.0 600000.0 343800.0 586200.0 ;
      RECT  333600.0 600000.0 343800.0 613800.0 ;
      RECT  333600.0 627600.0 343800.0 613800.0 ;
      RECT  333600.0 627600.0 343800.0 641400.0 ;
      RECT  333600.0 655200.0 343800.0 641400.0 ;
      RECT  333600.0 655200.0 343800.0 669000.0 ;
      RECT  333600.0 682800.0 343800.0 669000.0 ;
      RECT  333600.0 682800.0 343800.0 696600.0 ;
      RECT  333600.0 710400.0 343800.0 696600.0 ;
      RECT  333600.0 710400.0 343800.0 724200.0 ;
      RECT  333600.0 738000.0 343800.0 724200.0 ;
      RECT  333600.0 738000.0 343800.0 751800.0 ;
      RECT  333600.0 765600.0 343800.0 751800.0 ;
      RECT  333600.0 765600.0 343800.0 779400.0 ;
      RECT  333600.0 793200.0 343800.0 779400.0 ;
      RECT  333600.0 793200.0 343800.0 807000.0 ;
      RECT  333600.0 820800.0 343800.0 807000.0 ;
      RECT  333600.0 820800.0 343800.0 834600.0 ;
      RECT  333600.0 848400.0 343800.0 834600.0 ;
      RECT  333600.0 848400.0 343800.0 862200.0 ;
      RECT  333600.0 876000.0 343800.0 862200.0 ;
      RECT  333600.0 876000.0 343800.0 889800.0 ;
      RECT  333600.0 903600.0 343800.0 889800.0 ;
      RECT  333600.0 903600.0 343800.0 917400.0 ;
      RECT  333600.0 931200.0 343800.0 917400.0 ;
      RECT  333600.0 931200.0 343800.0 945000.0 ;
      RECT  333600.0 958800.0 343800.0 945000.0 ;
      RECT  333600.0 958800.0 343800.0 972600.0 ;
      RECT  333600.0 986400.0 343800.0 972600.0 ;
      RECT  333600.0 986400.0 343800.0 1000200.0 ;
      RECT  333600.0 1014000.0 343800.0 1000200.0 ;
      RECT  333600.0 1014000.0 343800.0 1027800.0 ;
      RECT  333600.0 1041600.0 343800.0 1027800.0 ;
      RECT  333600.0 1041600.0 343800.0 1055400.0 ;
      RECT  333600.0 1069200.0 343800.0 1055400.0 ;
      RECT  333600.0 1069200.0 343800.0 1083000.0 ;
      RECT  333600.0 1096800.0 343800.0 1083000.0 ;
      RECT  333600.0 1096800.0 343800.0 1110600.0 ;
      RECT  333600.0 1124400.0 343800.0 1110600.0 ;
      RECT  333600.0 1124400.0 343800.0 1138200.0 ;
      RECT  333600.0 1152000.0 343800.0 1138200.0 ;
      RECT  333600.0 1152000.0 343800.0 1165800.0 ;
      RECT  333600.0 1179600.0 343800.0 1165800.0 ;
      RECT  333600.0 1179600.0 343800.0 1193400.0 ;
      RECT  333600.0 1207200.0 343800.0 1193400.0 ;
      RECT  333600.0 1207200.0 343800.0 1221000.0 ;
      RECT  333600.0 1234800.0 343800.0 1221000.0 ;
      RECT  333600.0 1234800.0 343800.0 1248600.0 ;
      RECT  333600.0 1262400.0 343800.0 1248600.0 ;
      RECT  333600.0 1262400.0 343800.0 1276200.0 ;
      RECT  333600.0 1290000.0 343800.0 1276200.0 ;
      RECT  333600.0 1290000.0 343800.0 1303800.0 ;
      RECT  333600.0 1317600.0 343800.0 1303800.0 ;
      RECT  333600.0 1317600.0 343800.0 1331400.0 ;
      RECT  333600.0 1345200.0 343800.0 1331400.0 ;
      RECT  333600.0 1345200.0 343800.0 1359000.0 ;
      RECT  333600.0 1372800.0 343800.0 1359000.0 ;
      RECT  333600.0 1372800.0 343800.0 1386600.0 ;
      RECT  333600.0 1400400.0 343800.0 1386600.0 ;
      RECT  333600.0 1400400.0 343800.0 1414200.0 ;
      RECT  333600.0 1428000.0 343800.0 1414200.0 ;
      RECT  333600.0 1428000.0 343800.0 1441800.0 ;
      RECT  333600.0 1455600.0 343800.0 1441800.0 ;
      RECT  333600.0 1455600.0 343800.0 1469400.0 ;
      RECT  333600.0 1483200.0 343800.0 1469400.0 ;
      RECT  333600.0 1483200.0 343800.0 1497000.0 ;
      RECT  333600.0 1510800.0 343800.0 1497000.0 ;
      RECT  333600.0 1510800.0 343800.0 1524600.0 ;
      RECT  333600.0 1538400.0 343800.0 1524600.0 ;
      RECT  333600.0 1538400.0 343800.0 1552200.0 ;
      RECT  333600.0 1566000.0 343800.0 1552200.0 ;
      RECT  333600.0 1566000.0 343800.0 1579800.0 ;
      RECT  333600.0 1593600.0 343800.0 1579800.0 ;
      RECT  333600.0 1593600.0 343800.0 1607400.0 ;
      RECT  333600.0 1621200.0 343800.0 1607400.0 ;
      RECT  333600.0 1621200.0 343800.0 1635000.0 ;
      RECT  333600.0 1648800.0 343800.0 1635000.0 ;
      RECT  333600.0 1648800.0 343800.0 1662600.0 ;
      RECT  333600.0 1676400.0 343800.0 1662600.0 ;
      RECT  333600.0 1676400.0 343800.0 1690200.0 ;
      RECT  333600.0 1704000.0 343800.0 1690200.0 ;
      RECT  333600.0 1704000.0 343800.0 1717800.0 ;
      RECT  333600.0 1731600.0 343800.0 1717800.0 ;
      RECT  333600.0 1731600.0 343800.0 1745400.0 ;
      RECT  333600.0 1759200.0 343800.0 1745400.0 ;
      RECT  333600.0 1759200.0 343800.0 1773000.0 ;
      RECT  333600.0 1786800.0 343800.0 1773000.0 ;
      RECT  333600.0 1786800.0 343800.0 1800600.0 ;
      RECT  333600.0 1814400.0 343800.0 1800600.0 ;
      RECT  333600.0 1814400.0 343800.0 1828200.0 ;
      RECT  333600.0 1842000.0 343800.0 1828200.0 ;
      RECT  333600.0 1842000.0 343800.0 1855800.0 ;
      RECT  333600.0 1869600.0 343800.0 1855800.0 ;
      RECT  333600.0 1869600.0 343800.0 1883400.0 ;
      RECT  333600.0 1897200.0 343800.0 1883400.0 ;
      RECT  333600.0 1897200.0 343800.0 1911000.0 ;
      RECT  333600.0 1924800.0 343800.0 1911000.0 ;
      RECT  333600.0 1924800.0 343800.0 1938600.0 ;
      RECT  333600.0 1952400.0 343800.0 1938600.0 ;
      RECT  333600.0 1952400.0 343800.0 1966200.0 ;
      RECT  333600.0 1980000.0 343800.0 1966200.0 ;
      RECT  333600.0 1980000.0 343800.0 1993800.0 ;
      RECT  333600.0 2007600.0 343800.0 1993800.0 ;
      RECT  333600.0 2007600.0 343800.0 2021400.0 ;
      RECT  333600.0 2035200.0 343800.0 2021400.0 ;
      RECT  333600.0 2035200.0 343800.0 2049000.0 ;
      RECT  333600.0 2062800.0 343800.0 2049000.0 ;
      RECT  333600.0 2062800.0 343800.0 2076600.0 ;
      RECT  333600.0 2090400.0 343800.0 2076600.0 ;
      RECT  333600.0 2090400.0 343800.0 2104200.0 ;
      RECT  333600.0 2118000.0 343800.0 2104200.0 ;
      RECT  333600.0 2118000.0 343800.0 2131800.0 ;
      RECT  333600.0 2145600.0 343800.0 2131800.0 ;
      RECT  343800.0 379200.0 354000.0 393000.0 ;
      RECT  343800.0 406800.0 354000.0 393000.0 ;
      RECT  343800.0 406800.0 354000.0 420600.0 ;
      RECT  343800.0 434400.0 354000.0 420600.0 ;
      RECT  343800.0 434400.0 354000.0 448200.0 ;
      RECT  343800.0 462000.0 354000.0 448200.0 ;
      RECT  343800.0 462000.0 354000.0 475800.0 ;
      RECT  343800.0 489600.0 354000.0 475800.0 ;
      RECT  343800.0 489600.0 354000.0 503400.0 ;
      RECT  343800.0 517200.0 354000.0 503400.0 ;
      RECT  343800.0 517200.0 354000.0 531000.0 ;
      RECT  343800.0 544800.0 354000.0 531000.0 ;
      RECT  343800.0 544800.0 354000.0 558600.0 ;
      RECT  343800.0 572400.0 354000.0 558600.0 ;
      RECT  343800.0 572400.0 354000.0 586200.0 ;
      RECT  343800.0 600000.0 354000.0 586200.0 ;
      RECT  343800.0 600000.0 354000.0 613800.0 ;
      RECT  343800.0 627600.0 354000.0 613800.0 ;
      RECT  343800.0 627600.0 354000.0 641400.0 ;
      RECT  343800.0 655200.0 354000.0 641400.0 ;
      RECT  343800.0 655200.0 354000.0 669000.0 ;
      RECT  343800.0 682800.0 354000.0 669000.0 ;
      RECT  343800.0 682800.0 354000.0 696600.0 ;
      RECT  343800.0 710400.0 354000.0 696600.0 ;
      RECT  343800.0 710400.0 354000.0 724200.0 ;
      RECT  343800.0 738000.0 354000.0 724200.0 ;
      RECT  343800.0 738000.0 354000.0 751800.0 ;
      RECT  343800.0 765600.0 354000.0 751800.0 ;
      RECT  343800.0 765600.0 354000.0 779400.0 ;
      RECT  343800.0 793200.0 354000.0 779400.0 ;
      RECT  343800.0 793200.0 354000.0 807000.0 ;
      RECT  343800.0 820800.0 354000.0 807000.0 ;
      RECT  343800.0 820800.0 354000.0 834600.0 ;
      RECT  343800.0 848400.0 354000.0 834600.0 ;
      RECT  343800.0 848400.0 354000.0 862200.0 ;
      RECT  343800.0 876000.0 354000.0 862200.0 ;
      RECT  343800.0 876000.0 354000.0 889800.0 ;
      RECT  343800.0 903600.0 354000.0 889800.0 ;
      RECT  343800.0 903600.0 354000.0 917400.0 ;
      RECT  343800.0 931200.0 354000.0 917400.0 ;
      RECT  343800.0 931200.0 354000.0 945000.0 ;
      RECT  343800.0 958800.0 354000.0 945000.0 ;
      RECT  343800.0 958800.0 354000.0 972600.0 ;
      RECT  343800.0 986400.0 354000.0 972600.0 ;
      RECT  343800.0 986400.0 354000.0 1000200.0 ;
      RECT  343800.0 1014000.0 354000.0 1000200.0 ;
      RECT  343800.0 1014000.0 354000.0 1027800.0 ;
      RECT  343800.0 1041600.0 354000.0 1027800.0 ;
      RECT  343800.0 1041600.0 354000.0 1055400.0 ;
      RECT  343800.0 1069200.0 354000.0 1055400.0 ;
      RECT  343800.0 1069200.0 354000.0 1083000.0 ;
      RECT  343800.0 1096800.0 354000.0 1083000.0 ;
      RECT  343800.0 1096800.0 354000.0 1110600.0 ;
      RECT  343800.0 1124400.0 354000.0 1110600.0 ;
      RECT  343800.0 1124400.0 354000.0 1138200.0 ;
      RECT  343800.0 1152000.0 354000.0 1138200.0 ;
      RECT  343800.0 1152000.0 354000.0 1165800.0 ;
      RECT  343800.0 1179600.0 354000.0 1165800.0 ;
      RECT  343800.0 1179600.0 354000.0 1193400.0 ;
      RECT  343800.0 1207200.0 354000.0 1193400.0 ;
      RECT  343800.0 1207200.0 354000.0 1221000.0 ;
      RECT  343800.0 1234800.0 354000.0 1221000.0 ;
      RECT  343800.0 1234800.0 354000.0 1248600.0 ;
      RECT  343800.0 1262400.0 354000.0 1248600.0 ;
      RECT  343800.0 1262400.0 354000.0 1276200.0 ;
      RECT  343800.0 1290000.0 354000.0 1276200.0 ;
      RECT  343800.0 1290000.0 354000.0 1303800.0 ;
      RECT  343800.0 1317600.0 354000.0 1303800.0 ;
      RECT  343800.0 1317600.0 354000.0 1331400.0 ;
      RECT  343800.0 1345200.0 354000.0 1331400.0 ;
      RECT  343800.0 1345200.0 354000.0 1359000.0 ;
      RECT  343800.0 1372800.0 354000.0 1359000.0 ;
      RECT  343800.0 1372800.0 354000.0 1386600.0 ;
      RECT  343800.0 1400400.0 354000.0 1386600.0 ;
      RECT  343800.0 1400400.0 354000.0 1414200.0 ;
      RECT  343800.0 1428000.0 354000.0 1414200.0 ;
      RECT  343800.0 1428000.0 354000.0 1441800.0 ;
      RECT  343800.0 1455600.0 354000.0 1441800.0 ;
      RECT  343800.0 1455600.0 354000.0 1469400.0 ;
      RECT  343800.0 1483200.0 354000.0 1469400.0 ;
      RECT  343800.0 1483200.0 354000.0 1497000.0 ;
      RECT  343800.0 1510800.0 354000.0 1497000.0 ;
      RECT  343800.0 1510800.0 354000.0 1524600.0 ;
      RECT  343800.0 1538400.0 354000.0 1524600.0 ;
      RECT  343800.0 1538400.0 354000.0 1552200.0 ;
      RECT  343800.0 1566000.0 354000.0 1552200.0 ;
      RECT  343800.0 1566000.0 354000.0 1579800.0 ;
      RECT  343800.0 1593600.0 354000.0 1579800.0 ;
      RECT  343800.0 1593600.0 354000.0 1607400.0 ;
      RECT  343800.0 1621200.0 354000.0 1607400.0 ;
      RECT  343800.0 1621200.0 354000.0 1635000.0 ;
      RECT  343800.0 1648800.0 354000.0 1635000.0 ;
      RECT  343800.0 1648800.0 354000.0 1662600.0 ;
      RECT  343800.0 1676400.0 354000.0 1662600.0 ;
      RECT  343800.0 1676400.0 354000.0 1690200.0 ;
      RECT  343800.0 1704000.0 354000.0 1690200.0 ;
      RECT  343800.0 1704000.0 354000.0 1717800.0 ;
      RECT  343800.0 1731600.0 354000.0 1717800.0 ;
      RECT  343800.0 1731600.0 354000.0 1745400.0 ;
      RECT  343800.0 1759200.0 354000.0 1745400.0 ;
      RECT  343800.0 1759200.0 354000.0 1773000.0 ;
      RECT  343800.0 1786800.0 354000.0 1773000.0 ;
      RECT  343800.0 1786800.0 354000.0 1800600.0 ;
      RECT  343800.0 1814400.0 354000.0 1800600.0 ;
      RECT  343800.0 1814400.0 354000.0 1828200.0 ;
      RECT  343800.0 1842000.0 354000.0 1828200.0 ;
      RECT  343800.0 1842000.0 354000.0 1855800.0 ;
      RECT  343800.0 1869600.0 354000.0 1855800.0 ;
      RECT  343800.0 1869600.0 354000.0 1883400.0 ;
      RECT  343800.0 1897200.0 354000.0 1883400.0 ;
      RECT  343800.0 1897200.0 354000.0 1911000.0 ;
      RECT  343800.0 1924800.0 354000.0 1911000.0 ;
      RECT  343800.0 1924800.0 354000.0 1938600.0 ;
      RECT  343800.0 1952400.0 354000.0 1938600.0 ;
      RECT  343800.0 1952400.0 354000.0 1966200.0 ;
      RECT  343800.0 1980000.0 354000.0 1966200.0 ;
      RECT  343800.0 1980000.0 354000.0 1993800.0 ;
      RECT  343800.0 2007600.0 354000.0 1993800.0 ;
      RECT  343800.0 2007600.0 354000.0 2021400.0 ;
      RECT  343800.0 2035200.0 354000.0 2021400.0 ;
      RECT  343800.0 2035200.0 354000.0 2049000.0 ;
      RECT  343800.0 2062800.0 354000.0 2049000.0 ;
      RECT  343800.0 2062800.0 354000.0 2076600.0 ;
      RECT  343800.0 2090400.0 354000.0 2076600.0 ;
      RECT  343800.0 2090400.0 354000.0 2104200.0 ;
      RECT  343800.0 2118000.0 354000.0 2104200.0 ;
      RECT  343800.0 2118000.0 354000.0 2131800.0 ;
      RECT  343800.0 2145600.0 354000.0 2131800.0 ;
      RECT  354000.0 379200.0 364200.0 393000.0 ;
      RECT  354000.0 406800.0 364200.0 393000.0 ;
      RECT  354000.0 406800.0 364200.0 420600.0 ;
      RECT  354000.0 434400.0 364200.0 420600.0 ;
      RECT  354000.0 434400.0 364200.0 448200.0 ;
      RECT  354000.0 462000.0 364200.0 448200.0 ;
      RECT  354000.0 462000.0 364200.0 475800.0 ;
      RECT  354000.0 489600.0 364200.0 475800.0 ;
      RECT  354000.0 489600.0 364200.0 503400.0 ;
      RECT  354000.0 517200.0 364200.0 503400.0 ;
      RECT  354000.0 517200.0 364200.0 531000.0 ;
      RECT  354000.0 544800.0 364200.0 531000.0 ;
      RECT  354000.0 544800.0 364200.0 558600.0 ;
      RECT  354000.0 572400.0 364200.0 558600.0 ;
      RECT  354000.0 572400.0 364200.0 586200.0 ;
      RECT  354000.0 600000.0 364200.0 586200.0 ;
      RECT  354000.0 600000.0 364200.0 613800.0 ;
      RECT  354000.0 627600.0 364200.0 613800.0 ;
      RECT  354000.0 627600.0 364200.0 641400.0 ;
      RECT  354000.0 655200.0 364200.0 641400.0 ;
      RECT  354000.0 655200.0 364200.0 669000.0 ;
      RECT  354000.0 682800.0 364200.0 669000.0 ;
      RECT  354000.0 682800.0 364200.0 696600.0 ;
      RECT  354000.0 710400.0 364200.0 696600.0 ;
      RECT  354000.0 710400.0 364200.0 724200.0 ;
      RECT  354000.0 738000.0 364200.0 724200.0 ;
      RECT  354000.0 738000.0 364200.0 751800.0 ;
      RECT  354000.0 765600.0 364200.0 751800.0 ;
      RECT  354000.0 765600.0 364200.0 779400.0 ;
      RECT  354000.0 793200.0 364200.0 779400.0 ;
      RECT  354000.0 793200.0 364200.0 807000.0 ;
      RECT  354000.0 820800.0 364200.0 807000.0 ;
      RECT  354000.0 820800.0 364200.0 834600.0 ;
      RECT  354000.0 848400.0 364200.0 834600.0 ;
      RECT  354000.0 848400.0 364200.0 862200.0 ;
      RECT  354000.0 876000.0 364200.0 862200.0 ;
      RECT  354000.0 876000.0 364200.0 889800.0 ;
      RECT  354000.0 903600.0 364200.0 889800.0 ;
      RECT  354000.0 903600.0 364200.0 917400.0 ;
      RECT  354000.0 931200.0 364200.0 917400.0 ;
      RECT  354000.0 931200.0 364200.0 945000.0 ;
      RECT  354000.0 958800.0 364200.0 945000.0 ;
      RECT  354000.0 958800.0 364200.0 972600.0 ;
      RECT  354000.0 986400.0 364200.0 972600.0 ;
      RECT  354000.0 986400.0 364200.0 1000200.0 ;
      RECT  354000.0 1014000.0 364200.0 1000200.0 ;
      RECT  354000.0 1014000.0 364200.0 1027800.0 ;
      RECT  354000.0 1041600.0 364200.0 1027800.0 ;
      RECT  354000.0 1041600.0 364200.0 1055400.0 ;
      RECT  354000.0 1069200.0 364200.0 1055400.0 ;
      RECT  354000.0 1069200.0 364200.0 1083000.0 ;
      RECT  354000.0 1096800.0 364200.0 1083000.0 ;
      RECT  354000.0 1096800.0 364200.0 1110600.0 ;
      RECT  354000.0 1124400.0 364200.0 1110600.0 ;
      RECT  354000.0 1124400.0 364200.0 1138200.0 ;
      RECT  354000.0 1152000.0 364200.0 1138200.0 ;
      RECT  354000.0 1152000.0 364200.0 1165800.0 ;
      RECT  354000.0 1179600.0 364200.0 1165800.0 ;
      RECT  354000.0 1179600.0 364200.0 1193400.0 ;
      RECT  354000.0 1207200.0 364200.0 1193400.0 ;
      RECT  354000.0 1207200.0 364200.0 1221000.0 ;
      RECT  354000.0 1234800.0 364200.0 1221000.0 ;
      RECT  354000.0 1234800.0 364200.0 1248600.0 ;
      RECT  354000.0 1262400.0 364200.0 1248600.0 ;
      RECT  354000.0 1262400.0 364200.0 1276200.0 ;
      RECT  354000.0 1290000.0 364200.0 1276200.0 ;
      RECT  354000.0 1290000.0 364200.0 1303800.0 ;
      RECT  354000.0 1317600.0 364200.0 1303800.0 ;
      RECT  354000.0 1317600.0 364200.0 1331400.0 ;
      RECT  354000.0 1345200.0 364200.0 1331400.0 ;
      RECT  354000.0 1345200.0 364200.0 1359000.0 ;
      RECT  354000.0 1372800.0 364200.0 1359000.0 ;
      RECT  354000.0 1372800.0 364200.0 1386600.0 ;
      RECT  354000.0 1400400.0 364200.0 1386600.0 ;
      RECT  354000.0 1400400.0 364200.0 1414200.0 ;
      RECT  354000.0 1428000.0 364200.0 1414200.0 ;
      RECT  354000.0 1428000.0 364200.0 1441800.0 ;
      RECT  354000.0 1455600.0 364200.0 1441800.0 ;
      RECT  354000.0 1455600.0 364200.0 1469400.0 ;
      RECT  354000.0 1483200.0 364200.0 1469400.0 ;
      RECT  354000.0 1483200.0 364200.0 1497000.0 ;
      RECT  354000.0 1510800.0 364200.0 1497000.0 ;
      RECT  354000.0 1510800.0 364200.0 1524600.0 ;
      RECT  354000.0 1538400.0 364200.0 1524600.0 ;
      RECT  354000.0 1538400.0 364200.0 1552200.0 ;
      RECT  354000.0 1566000.0 364200.0 1552200.0 ;
      RECT  354000.0 1566000.0 364200.0 1579800.0 ;
      RECT  354000.0 1593600.0 364200.0 1579800.0 ;
      RECT  354000.0 1593600.0 364200.0 1607400.0 ;
      RECT  354000.0 1621200.0 364200.0 1607400.0 ;
      RECT  354000.0 1621200.0 364200.0 1635000.0 ;
      RECT  354000.0 1648800.0 364200.0 1635000.0 ;
      RECT  354000.0 1648800.0 364200.0 1662600.0 ;
      RECT  354000.0 1676400.0 364200.0 1662600.0 ;
      RECT  354000.0 1676400.0 364200.0 1690200.0 ;
      RECT  354000.0 1704000.0 364200.0 1690200.0 ;
      RECT  354000.0 1704000.0 364200.0 1717800.0 ;
      RECT  354000.0 1731600.0 364200.0 1717800.0 ;
      RECT  354000.0 1731600.0 364200.0 1745400.0 ;
      RECT  354000.0 1759200.0 364200.0 1745400.0 ;
      RECT  354000.0 1759200.0 364200.0 1773000.0 ;
      RECT  354000.0 1786800.0 364200.0 1773000.0 ;
      RECT  354000.0 1786800.0 364200.0 1800600.0 ;
      RECT  354000.0 1814400.0 364200.0 1800600.0 ;
      RECT  354000.0 1814400.0 364200.0 1828200.0 ;
      RECT  354000.0 1842000.0 364200.0 1828200.0 ;
      RECT  354000.0 1842000.0 364200.0 1855800.0 ;
      RECT  354000.0 1869600.0 364200.0 1855800.0 ;
      RECT  354000.0 1869600.0 364200.0 1883400.0 ;
      RECT  354000.0 1897200.0 364200.0 1883400.0 ;
      RECT  354000.0 1897200.0 364200.0 1911000.0 ;
      RECT  354000.0 1924800.0 364200.0 1911000.0 ;
      RECT  354000.0 1924800.0 364200.0 1938600.0 ;
      RECT  354000.0 1952400.0 364200.0 1938600.0 ;
      RECT  354000.0 1952400.0 364200.0 1966200.0 ;
      RECT  354000.0 1980000.0 364200.0 1966200.0 ;
      RECT  354000.0 1980000.0 364200.0 1993800.0 ;
      RECT  354000.0 2007600.0 364200.0 1993800.0 ;
      RECT  354000.0 2007600.0 364200.0 2021400.0 ;
      RECT  354000.0 2035200.0 364200.0 2021400.0 ;
      RECT  354000.0 2035200.0 364200.0 2049000.0 ;
      RECT  354000.0 2062800.0 364200.0 2049000.0 ;
      RECT  354000.0 2062800.0 364200.0 2076600.0 ;
      RECT  354000.0 2090400.0 364200.0 2076600.0 ;
      RECT  354000.0 2090400.0 364200.0 2104200.0 ;
      RECT  354000.0 2118000.0 364200.0 2104200.0 ;
      RECT  354000.0 2118000.0 364200.0 2131800.0 ;
      RECT  354000.0 2145600.0 364200.0 2131800.0 ;
      RECT  364200.0 379200.0 374400.0 393000.0 ;
      RECT  364200.0 406800.0 374400.0 393000.0 ;
      RECT  364200.0 406800.0 374400.0 420600.0 ;
      RECT  364200.0 434400.0 374400.0 420600.0 ;
      RECT  364200.0 434400.0 374400.0 448200.0 ;
      RECT  364200.0 462000.0 374400.0 448200.0 ;
      RECT  364200.0 462000.0 374400.0 475800.0 ;
      RECT  364200.0 489600.0 374400.0 475800.0 ;
      RECT  364200.0 489600.0 374400.0 503400.0 ;
      RECT  364200.0 517200.0 374400.0 503400.0 ;
      RECT  364200.0 517200.0 374400.0 531000.0 ;
      RECT  364200.0 544800.0 374400.0 531000.0 ;
      RECT  364200.0 544800.0 374400.0 558600.0 ;
      RECT  364200.0 572400.0 374400.0 558600.0 ;
      RECT  364200.0 572400.0 374400.0 586200.0 ;
      RECT  364200.0 600000.0 374400.0 586200.0 ;
      RECT  364200.0 600000.0 374400.0 613800.0 ;
      RECT  364200.0 627600.0 374400.0 613800.0 ;
      RECT  364200.0 627600.0 374400.0 641400.0 ;
      RECT  364200.0 655200.0 374400.0 641400.0 ;
      RECT  364200.0 655200.0 374400.0 669000.0 ;
      RECT  364200.0 682800.0 374400.0 669000.0 ;
      RECT  364200.0 682800.0 374400.0 696600.0 ;
      RECT  364200.0 710400.0 374400.0 696600.0 ;
      RECT  364200.0 710400.0 374400.0 724200.0 ;
      RECT  364200.0 738000.0 374400.0 724200.0 ;
      RECT  364200.0 738000.0 374400.0 751800.0 ;
      RECT  364200.0 765600.0 374400.0 751800.0 ;
      RECT  364200.0 765600.0 374400.0 779400.0 ;
      RECT  364200.0 793200.0 374400.0 779400.0 ;
      RECT  364200.0 793200.0 374400.0 807000.0 ;
      RECT  364200.0 820800.0 374400.0 807000.0 ;
      RECT  364200.0 820800.0 374400.0 834600.0 ;
      RECT  364200.0 848400.0 374400.0 834600.0 ;
      RECT  364200.0 848400.0 374400.0 862200.0 ;
      RECT  364200.0 876000.0 374400.0 862200.0 ;
      RECT  364200.0 876000.0 374400.0 889800.0 ;
      RECT  364200.0 903600.0 374400.0 889800.0 ;
      RECT  364200.0 903600.0 374400.0 917400.0 ;
      RECT  364200.0 931200.0 374400.0 917400.0 ;
      RECT  364200.0 931200.0 374400.0 945000.0 ;
      RECT  364200.0 958800.0 374400.0 945000.0 ;
      RECT  364200.0 958800.0 374400.0 972600.0 ;
      RECT  364200.0 986400.0 374400.0 972600.0 ;
      RECT  364200.0 986400.0 374400.0 1000200.0 ;
      RECT  364200.0 1014000.0 374400.0 1000200.0 ;
      RECT  364200.0 1014000.0 374400.0 1027800.0 ;
      RECT  364200.0 1041600.0 374400.0 1027800.0 ;
      RECT  364200.0 1041600.0 374400.0 1055400.0 ;
      RECT  364200.0 1069200.0 374400.0 1055400.0 ;
      RECT  364200.0 1069200.0 374400.0 1083000.0 ;
      RECT  364200.0 1096800.0 374400.0 1083000.0 ;
      RECT  364200.0 1096800.0 374400.0 1110600.0 ;
      RECT  364200.0 1124400.0 374400.0 1110600.0 ;
      RECT  364200.0 1124400.0 374400.0 1138200.0 ;
      RECT  364200.0 1152000.0 374400.0 1138200.0 ;
      RECT  364200.0 1152000.0 374400.0 1165800.0 ;
      RECT  364200.0 1179600.0 374400.0 1165800.0 ;
      RECT  364200.0 1179600.0 374400.0 1193400.0 ;
      RECT  364200.0 1207200.0 374400.0 1193400.0 ;
      RECT  364200.0 1207200.0 374400.0 1221000.0 ;
      RECT  364200.0 1234800.0 374400.0 1221000.0 ;
      RECT  364200.0 1234800.0 374400.0 1248600.0 ;
      RECT  364200.0 1262400.0 374400.0 1248600.0 ;
      RECT  364200.0 1262400.0 374400.0 1276200.0 ;
      RECT  364200.0 1290000.0 374400.0 1276200.0 ;
      RECT  364200.0 1290000.0 374400.0 1303800.0 ;
      RECT  364200.0 1317600.0 374400.0 1303800.0 ;
      RECT  364200.0 1317600.0 374400.0 1331400.0 ;
      RECT  364200.0 1345200.0 374400.0 1331400.0 ;
      RECT  364200.0 1345200.0 374400.0 1359000.0 ;
      RECT  364200.0 1372800.0 374400.0 1359000.0 ;
      RECT  364200.0 1372800.0 374400.0 1386600.0 ;
      RECT  364200.0 1400400.0 374400.0 1386600.0 ;
      RECT  364200.0 1400400.0 374400.0 1414200.0 ;
      RECT  364200.0 1428000.0 374400.0 1414200.0 ;
      RECT  364200.0 1428000.0 374400.0 1441800.0 ;
      RECT  364200.0 1455600.0 374400.0 1441800.0 ;
      RECT  364200.0 1455600.0 374400.0 1469400.0 ;
      RECT  364200.0 1483200.0 374400.0 1469400.0 ;
      RECT  364200.0 1483200.0 374400.0 1497000.0 ;
      RECT  364200.0 1510800.0 374400.0 1497000.0 ;
      RECT  364200.0 1510800.0 374400.0 1524600.0 ;
      RECT  364200.0 1538400.0 374400.0 1524600.0 ;
      RECT  364200.0 1538400.0 374400.0 1552200.0 ;
      RECT  364200.0 1566000.0 374400.0 1552200.0 ;
      RECT  364200.0 1566000.0 374400.0 1579800.0 ;
      RECT  364200.0 1593600.0 374400.0 1579800.0 ;
      RECT  364200.0 1593600.0 374400.0 1607400.0 ;
      RECT  364200.0 1621200.0 374400.0 1607400.0 ;
      RECT  364200.0 1621200.0 374400.0 1635000.0 ;
      RECT  364200.0 1648800.0 374400.0 1635000.0 ;
      RECT  364200.0 1648800.0 374400.0 1662600.0 ;
      RECT  364200.0 1676400.0 374400.0 1662600.0 ;
      RECT  364200.0 1676400.0 374400.0 1690200.0 ;
      RECT  364200.0 1704000.0 374400.0 1690200.0 ;
      RECT  364200.0 1704000.0 374400.0 1717800.0 ;
      RECT  364200.0 1731600.0 374400.0 1717800.0 ;
      RECT  364200.0 1731600.0 374400.0 1745400.0 ;
      RECT  364200.0 1759200.0 374400.0 1745400.0 ;
      RECT  364200.0 1759200.0 374400.0 1773000.0 ;
      RECT  364200.0 1786800.0 374400.0 1773000.0 ;
      RECT  364200.0 1786800.0 374400.0 1800600.0 ;
      RECT  364200.0 1814400.0 374400.0 1800600.0 ;
      RECT  364200.0 1814400.0 374400.0 1828200.0 ;
      RECT  364200.0 1842000.0 374400.0 1828200.0 ;
      RECT  364200.0 1842000.0 374400.0 1855800.0 ;
      RECT  364200.0 1869600.0 374400.0 1855800.0 ;
      RECT  364200.0 1869600.0 374400.0 1883400.0 ;
      RECT  364200.0 1897200.0 374400.0 1883400.0 ;
      RECT  364200.0 1897200.0 374400.0 1911000.0 ;
      RECT  364200.0 1924800.0 374400.0 1911000.0 ;
      RECT  364200.0 1924800.0 374400.0 1938600.0 ;
      RECT  364200.0 1952400.0 374400.0 1938600.0 ;
      RECT  364200.0 1952400.0 374400.0 1966200.0 ;
      RECT  364200.0 1980000.0 374400.0 1966200.0 ;
      RECT  364200.0 1980000.0 374400.0 1993800.0 ;
      RECT  364200.0 2007600.0 374400.0 1993800.0 ;
      RECT  364200.0 2007600.0 374400.0 2021400.0 ;
      RECT  364200.0 2035200.0 374400.0 2021400.0 ;
      RECT  364200.0 2035200.0 374400.0 2049000.0 ;
      RECT  364200.0 2062800.0 374400.0 2049000.0 ;
      RECT  364200.0 2062800.0 374400.0 2076600.0 ;
      RECT  364200.0 2090400.0 374400.0 2076600.0 ;
      RECT  364200.0 2090400.0 374400.0 2104200.0 ;
      RECT  364200.0 2118000.0 374400.0 2104200.0 ;
      RECT  364200.0 2118000.0 374400.0 2131800.0 ;
      RECT  364200.0 2145600.0 374400.0 2131800.0 ;
      RECT  374400.0 379200.0 384600.0 393000.0 ;
      RECT  374400.0 406800.0 384600.0 393000.0 ;
      RECT  374400.0 406800.0 384600.0 420600.0 ;
      RECT  374400.0 434400.0 384600.0 420600.0 ;
      RECT  374400.0 434400.0 384600.0 448200.0 ;
      RECT  374400.0 462000.0 384600.0 448200.0 ;
      RECT  374400.0 462000.0 384600.0 475800.0 ;
      RECT  374400.0 489600.0 384600.0 475800.0 ;
      RECT  374400.0 489600.0 384600.0 503400.0 ;
      RECT  374400.0 517200.0 384600.0 503400.0 ;
      RECT  374400.0 517200.0 384600.0 531000.0 ;
      RECT  374400.0 544800.0 384600.0 531000.0 ;
      RECT  374400.0 544800.0 384600.0 558600.0 ;
      RECT  374400.0 572400.0 384600.0 558600.0 ;
      RECT  374400.0 572400.0 384600.0 586200.0 ;
      RECT  374400.0 600000.0 384600.0 586200.0 ;
      RECT  374400.0 600000.0 384600.0 613800.0 ;
      RECT  374400.0 627600.0 384600.0 613800.0 ;
      RECT  374400.0 627600.0 384600.0 641400.0 ;
      RECT  374400.0 655200.0 384600.0 641400.0 ;
      RECT  374400.0 655200.0 384600.0 669000.0 ;
      RECT  374400.0 682800.0 384600.0 669000.0 ;
      RECT  374400.0 682800.0 384600.0 696600.0 ;
      RECT  374400.0 710400.0 384600.0 696600.0 ;
      RECT  374400.0 710400.0 384600.0 724200.0 ;
      RECT  374400.0 738000.0 384600.0 724200.0 ;
      RECT  374400.0 738000.0 384600.0 751800.0 ;
      RECT  374400.0 765600.0 384600.0 751800.0 ;
      RECT  374400.0 765600.0 384600.0 779400.0 ;
      RECT  374400.0 793200.0 384600.0 779400.0 ;
      RECT  374400.0 793200.0 384600.0 807000.0 ;
      RECT  374400.0 820800.0 384600.0 807000.0 ;
      RECT  374400.0 820800.0 384600.0 834600.0 ;
      RECT  374400.0 848400.0 384600.0 834600.0 ;
      RECT  374400.0 848400.0 384600.0 862200.0 ;
      RECT  374400.0 876000.0 384600.0 862200.0 ;
      RECT  374400.0 876000.0 384600.0 889800.0 ;
      RECT  374400.0 903600.0 384600.0 889800.0 ;
      RECT  374400.0 903600.0 384600.0 917400.0 ;
      RECT  374400.0 931200.0 384600.0 917400.0 ;
      RECT  374400.0 931200.0 384600.0 945000.0 ;
      RECT  374400.0 958800.0 384600.0 945000.0 ;
      RECT  374400.0 958800.0 384600.0 972600.0 ;
      RECT  374400.0 986400.0 384600.0 972600.0 ;
      RECT  374400.0 986400.0 384600.0 1000200.0 ;
      RECT  374400.0 1014000.0 384600.0 1000200.0 ;
      RECT  374400.0 1014000.0 384600.0 1027800.0 ;
      RECT  374400.0 1041600.0 384600.0 1027800.0 ;
      RECT  374400.0 1041600.0 384600.0 1055400.0 ;
      RECT  374400.0 1069200.0 384600.0 1055400.0 ;
      RECT  374400.0 1069200.0 384600.0 1083000.0 ;
      RECT  374400.0 1096800.0 384600.0 1083000.0 ;
      RECT  374400.0 1096800.0 384600.0 1110600.0 ;
      RECT  374400.0 1124400.0 384600.0 1110600.0 ;
      RECT  374400.0 1124400.0 384600.0 1138200.0 ;
      RECT  374400.0 1152000.0 384600.0 1138200.0 ;
      RECT  374400.0 1152000.0 384600.0 1165800.0 ;
      RECT  374400.0 1179600.0 384600.0 1165800.0 ;
      RECT  374400.0 1179600.0 384600.0 1193400.0 ;
      RECT  374400.0 1207200.0 384600.0 1193400.0 ;
      RECT  374400.0 1207200.0 384600.0 1221000.0 ;
      RECT  374400.0 1234800.0 384600.0 1221000.0 ;
      RECT  374400.0 1234800.0 384600.0 1248600.0 ;
      RECT  374400.0 1262400.0 384600.0 1248600.0 ;
      RECT  374400.0 1262400.0 384600.0 1276200.0 ;
      RECT  374400.0 1290000.0 384600.0 1276200.0 ;
      RECT  374400.0 1290000.0 384600.0 1303800.0 ;
      RECT  374400.0 1317600.0 384600.0 1303800.0 ;
      RECT  374400.0 1317600.0 384600.0 1331400.0 ;
      RECT  374400.0 1345200.0 384600.0 1331400.0 ;
      RECT  374400.0 1345200.0 384600.0 1359000.0 ;
      RECT  374400.0 1372800.0 384600.0 1359000.0 ;
      RECT  374400.0 1372800.0 384600.0 1386600.0 ;
      RECT  374400.0 1400400.0 384600.0 1386600.0 ;
      RECT  374400.0 1400400.0 384600.0 1414200.0 ;
      RECT  374400.0 1428000.0 384600.0 1414200.0 ;
      RECT  374400.0 1428000.0 384600.0 1441800.0 ;
      RECT  374400.0 1455600.0 384600.0 1441800.0 ;
      RECT  374400.0 1455600.0 384600.0 1469400.0 ;
      RECT  374400.0 1483200.0 384600.0 1469400.0 ;
      RECT  374400.0 1483200.0 384600.0 1497000.0 ;
      RECT  374400.0 1510800.0 384600.0 1497000.0 ;
      RECT  374400.0 1510800.0 384600.0 1524600.0 ;
      RECT  374400.0 1538400.0 384600.0 1524600.0 ;
      RECT  374400.0 1538400.0 384600.0 1552200.0 ;
      RECT  374400.0 1566000.0 384600.0 1552200.0 ;
      RECT  374400.0 1566000.0 384600.0 1579800.0 ;
      RECT  374400.0 1593600.0 384600.0 1579800.0 ;
      RECT  374400.0 1593600.0 384600.0 1607400.0 ;
      RECT  374400.0 1621200.0 384600.0 1607400.0 ;
      RECT  374400.0 1621200.0 384600.0 1635000.0 ;
      RECT  374400.0 1648800.0 384600.0 1635000.0 ;
      RECT  374400.0 1648800.0 384600.0 1662600.0 ;
      RECT  374400.0 1676400.0 384600.0 1662600.0 ;
      RECT  374400.0 1676400.0 384600.0 1690200.0 ;
      RECT  374400.0 1704000.0 384600.0 1690200.0 ;
      RECT  374400.0 1704000.0 384600.0 1717800.0 ;
      RECT  374400.0 1731600.0 384600.0 1717800.0 ;
      RECT  374400.0 1731600.0 384600.0 1745400.0 ;
      RECT  374400.0 1759200.0 384600.0 1745400.0 ;
      RECT  374400.0 1759200.0 384600.0 1773000.0 ;
      RECT  374400.0 1786800.0 384600.0 1773000.0 ;
      RECT  374400.0 1786800.0 384600.0 1800600.0 ;
      RECT  374400.0 1814400.0 384600.0 1800600.0 ;
      RECT  374400.0 1814400.0 384600.0 1828200.0 ;
      RECT  374400.0 1842000.0 384600.0 1828200.0 ;
      RECT  374400.0 1842000.0 384600.0 1855800.0 ;
      RECT  374400.0 1869600.0 384600.0 1855800.0 ;
      RECT  374400.0 1869600.0 384600.0 1883400.0 ;
      RECT  374400.0 1897200.0 384600.0 1883400.0 ;
      RECT  374400.0 1897200.0 384600.0 1911000.0 ;
      RECT  374400.0 1924800.0 384600.0 1911000.0 ;
      RECT  374400.0 1924800.0 384600.0 1938600.0 ;
      RECT  374400.0 1952400.0 384600.0 1938600.0 ;
      RECT  374400.0 1952400.0 384600.0 1966200.0 ;
      RECT  374400.0 1980000.0 384600.0 1966200.0 ;
      RECT  374400.0 1980000.0 384600.0 1993800.0 ;
      RECT  374400.0 2007600.0 384600.0 1993800.0 ;
      RECT  374400.0 2007600.0 384600.0 2021400.0 ;
      RECT  374400.0 2035200.0 384600.0 2021400.0 ;
      RECT  374400.0 2035200.0 384600.0 2049000.0 ;
      RECT  374400.0 2062800.0 384600.0 2049000.0 ;
      RECT  374400.0 2062800.0 384600.0 2076600.0 ;
      RECT  374400.0 2090400.0 384600.0 2076600.0 ;
      RECT  374400.0 2090400.0 384600.0 2104200.0 ;
      RECT  374400.0 2118000.0 384600.0 2104200.0 ;
      RECT  374400.0 2118000.0 384600.0 2131800.0 ;
      RECT  374400.0 2145600.0 384600.0 2131800.0 ;
      RECT  384600.0 379200.0 394800.0 393000.0 ;
      RECT  384600.0 406800.0 394800.0 393000.0 ;
      RECT  384600.0 406800.0 394800.0 420600.0 ;
      RECT  384600.0 434400.0 394800.0 420600.0 ;
      RECT  384600.0 434400.0 394800.0 448200.0 ;
      RECT  384600.0 462000.0 394800.0 448200.0 ;
      RECT  384600.0 462000.0 394800.0 475800.0 ;
      RECT  384600.0 489600.0 394800.0 475800.0 ;
      RECT  384600.0 489600.0 394800.0 503400.0 ;
      RECT  384600.0 517200.0 394800.0 503400.0 ;
      RECT  384600.0 517200.0 394800.0 531000.0 ;
      RECT  384600.0 544800.0 394800.0 531000.0 ;
      RECT  384600.0 544800.0 394800.0 558600.0 ;
      RECT  384600.0 572400.0 394800.0 558600.0 ;
      RECT  384600.0 572400.0 394800.0 586200.0 ;
      RECT  384600.0 600000.0 394800.0 586200.0 ;
      RECT  384600.0 600000.0 394800.0 613800.0 ;
      RECT  384600.0 627600.0 394800.0 613800.0 ;
      RECT  384600.0 627600.0 394800.0 641400.0 ;
      RECT  384600.0 655200.0 394800.0 641400.0 ;
      RECT  384600.0 655200.0 394800.0 669000.0 ;
      RECT  384600.0 682800.0 394800.0 669000.0 ;
      RECT  384600.0 682800.0 394800.0 696600.0 ;
      RECT  384600.0 710400.0 394800.0 696600.0 ;
      RECT  384600.0 710400.0 394800.0 724200.0 ;
      RECT  384600.0 738000.0 394800.0 724200.0 ;
      RECT  384600.0 738000.0 394800.0 751800.0 ;
      RECT  384600.0 765600.0 394800.0 751800.0 ;
      RECT  384600.0 765600.0 394800.0 779400.0 ;
      RECT  384600.0 793200.0 394800.0 779400.0 ;
      RECT  384600.0 793200.0 394800.0 807000.0 ;
      RECT  384600.0 820800.0 394800.0 807000.0 ;
      RECT  384600.0 820800.0 394800.0 834600.0 ;
      RECT  384600.0 848400.0 394800.0 834600.0 ;
      RECT  384600.0 848400.0 394800.0 862200.0 ;
      RECT  384600.0 876000.0 394800.0 862200.0 ;
      RECT  384600.0 876000.0 394800.0 889800.0 ;
      RECT  384600.0 903600.0 394800.0 889800.0 ;
      RECT  384600.0 903600.0 394800.0 917400.0 ;
      RECT  384600.0 931200.0 394800.0 917400.0 ;
      RECT  384600.0 931200.0 394800.0 945000.0 ;
      RECT  384600.0 958800.0 394800.0 945000.0 ;
      RECT  384600.0 958800.0 394800.0 972600.0 ;
      RECT  384600.0 986400.0 394800.0 972600.0 ;
      RECT  384600.0 986400.0 394800.0 1000200.0 ;
      RECT  384600.0 1014000.0 394800.0 1000200.0 ;
      RECT  384600.0 1014000.0 394800.0 1027800.0 ;
      RECT  384600.0 1041600.0 394800.0 1027800.0 ;
      RECT  384600.0 1041600.0 394800.0 1055400.0 ;
      RECT  384600.0 1069200.0 394800.0 1055400.0 ;
      RECT  384600.0 1069200.0 394800.0 1083000.0 ;
      RECT  384600.0 1096800.0 394800.0 1083000.0 ;
      RECT  384600.0 1096800.0 394800.0 1110600.0 ;
      RECT  384600.0 1124400.0 394800.0 1110600.0 ;
      RECT  384600.0 1124400.0 394800.0 1138200.0 ;
      RECT  384600.0 1152000.0 394800.0 1138200.0 ;
      RECT  384600.0 1152000.0 394800.0 1165800.0 ;
      RECT  384600.0 1179600.0 394800.0 1165800.0 ;
      RECT  384600.0 1179600.0 394800.0 1193400.0 ;
      RECT  384600.0 1207200.0 394800.0 1193400.0 ;
      RECT  384600.0 1207200.0 394800.0 1221000.0 ;
      RECT  384600.0 1234800.0 394800.0 1221000.0 ;
      RECT  384600.0 1234800.0 394800.0 1248600.0 ;
      RECT  384600.0 1262400.0 394800.0 1248600.0 ;
      RECT  384600.0 1262400.0 394800.0 1276200.0 ;
      RECT  384600.0 1290000.0 394800.0 1276200.0 ;
      RECT  384600.0 1290000.0 394800.0 1303800.0 ;
      RECT  384600.0 1317600.0 394800.0 1303800.0 ;
      RECT  384600.0 1317600.0 394800.0 1331400.0 ;
      RECT  384600.0 1345200.0 394800.0 1331400.0 ;
      RECT  384600.0 1345200.0 394800.0 1359000.0 ;
      RECT  384600.0 1372800.0 394800.0 1359000.0 ;
      RECT  384600.0 1372800.0 394800.0 1386600.0 ;
      RECT  384600.0 1400400.0 394800.0 1386600.0 ;
      RECT  384600.0 1400400.0 394800.0 1414200.0 ;
      RECT  384600.0 1428000.0 394800.0 1414200.0 ;
      RECT  384600.0 1428000.0 394800.0 1441800.0 ;
      RECT  384600.0 1455600.0 394800.0 1441800.0 ;
      RECT  384600.0 1455600.0 394800.0 1469400.0 ;
      RECT  384600.0 1483200.0 394800.0 1469400.0 ;
      RECT  384600.0 1483200.0 394800.0 1497000.0 ;
      RECT  384600.0 1510800.0 394800.0 1497000.0 ;
      RECT  384600.0 1510800.0 394800.0 1524600.0 ;
      RECT  384600.0 1538400.0 394800.0 1524600.0 ;
      RECT  384600.0 1538400.0 394800.0 1552200.0 ;
      RECT  384600.0 1566000.0 394800.0 1552200.0 ;
      RECT  384600.0 1566000.0 394800.0 1579800.0 ;
      RECT  384600.0 1593600.0 394800.0 1579800.0 ;
      RECT  384600.0 1593600.0 394800.0 1607400.0 ;
      RECT  384600.0 1621200.0 394800.0 1607400.0 ;
      RECT  384600.0 1621200.0 394800.0 1635000.0 ;
      RECT  384600.0 1648800.0 394800.0 1635000.0 ;
      RECT  384600.0 1648800.0 394800.0 1662600.0 ;
      RECT  384600.0 1676400.0 394800.0 1662600.0 ;
      RECT  384600.0 1676400.0 394800.0 1690200.0 ;
      RECT  384600.0 1704000.0 394800.0 1690200.0 ;
      RECT  384600.0 1704000.0 394800.0 1717800.0 ;
      RECT  384600.0 1731600.0 394800.0 1717800.0 ;
      RECT  384600.0 1731600.0 394800.0 1745400.0 ;
      RECT  384600.0 1759200.0 394800.0 1745400.0 ;
      RECT  384600.0 1759200.0 394800.0 1773000.0 ;
      RECT  384600.0 1786800.0 394800.0 1773000.0 ;
      RECT  384600.0 1786800.0 394800.0 1800600.0 ;
      RECT  384600.0 1814400.0 394800.0 1800600.0 ;
      RECT  384600.0 1814400.0 394800.0 1828200.0 ;
      RECT  384600.0 1842000.0 394800.0 1828200.0 ;
      RECT  384600.0 1842000.0 394800.0 1855800.0 ;
      RECT  384600.0 1869600.0 394800.0 1855800.0 ;
      RECT  384600.0 1869600.0 394800.0 1883400.0 ;
      RECT  384600.0 1897200.0 394800.0 1883400.0 ;
      RECT  384600.0 1897200.0 394800.0 1911000.0 ;
      RECT  384600.0 1924800.0 394800.0 1911000.0 ;
      RECT  384600.0 1924800.0 394800.0 1938600.0 ;
      RECT  384600.0 1952400.0 394800.0 1938600.0 ;
      RECT  384600.0 1952400.0 394800.0 1966200.0 ;
      RECT  384600.0 1980000.0 394800.0 1966200.0 ;
      RECT  384600.0 1980000.0 394800.0 1993800.0 ;
      RECT  384600.0 2007600.0 394800.0 1993800.0 ;
      RECT  384600.0 2007600.0 394800.0 2021400.0 ;
      RECT  384600.0 2035200.0 394800.0 2021400.0 ;
      RECT  384600.0 2035200.0 394800.0 2049000.0 ;
      RECT  384600.0 2062800.0 394800.0 2049000.0 ;
      RECT  384600.0 2062800.0 394800.0 2076600.0 ;
      RECT  384600.0 2090400.0 394800.0 2076600.0 ;
      RECT  384600.0 2090400.0 394800.0 2104200.0 ;
      RECT  384600.0 2118000.0 394800.0 2104200.0 ;
      RECT  384600.0 2118000.0 394800.0 2131800.0 ;
      RECT  384600.0 2145600.0 394800.0 2131800.0 ;
      RECT  394800.0 379200.0 405000.0 393000.0 ;
      RECT  394800.0 406800.0 405000.0 393000.0 ;
      RECT  394800.0 406800.0 405000.0 420600.0 ;
      RECT  394800.0 434400.0 405000.0 420600.0 ;
      RECT  394800.0 434400.0 405000.0 448200.0 ;
      RECT  394800.0 462000.0 405000.0 448200.0 ;
      RECT  394800.0 462000.0 405000.0 475800.0 ;
      RECT  394800.0 489600.0 405000.0 475800.0 ;
      RECT  394800.0 489600.0 405000.0 503400.0 ;
      RECT  394800.0 517200.0 405000.0 503400.0 ;
      RECT  394800.0 517200.0 405000.0 531000.0 ;
      RECT  394800.0 544800.0 405000.0 531000.0 ;
      RECT  394800.0 544800.0 405000.0 558600.0 ;
      RECT  394800.0 572400.0 405000.0 558600.0 ;
      RECT  394800.0 572400.0 405000.0 586200.0 ;
      RECT  394800.0 600000.0 405000.0 586200.0 ;
      RECT  394800.0 600000.0 405000.0 613800.0 ;
      RECT  394800.0 627600.0 405000.0 613800.0 ;
      RECT  394800.0 627600.0 405000.0 641400.0 ;
      RECT  394800.0 655200.0 405000.0 641400.0 ;
      RECT  394800.0 655200.0 405000.0 669000.0 ;
      RECT  394800.0 682800.0 405000.0 669000.0 ;
      RECT  394800.0 682800.0 405000.0 696600.0 ;
      RECT  394800.0 710400.0 405000.0 696600.0 ;
      RECT  394800.0 710400.0 405000.0 724200.0 ;
      RECT  394800.0 738000.0 405000.0 724200.0 ;
      RECT  394800.0 738000.0 405000.0 751800.0 ;
      RECT  394800.0 765600.0 405000.0 751800.0 ;
      RECT  394800.0 765600.0 405000.0 779400.0 ;
      RECT  394800.0 793200.0 405000.0 779400.0 ;
      RECT  394800.0 793200.0 405000.0 807000.0 ;
      RECT  394800.0 820800.0 405000.0 807000.0 ;
      RECT  394800.0 820800.0 405000.0 834600.0 ;
      RECT  394800.0 848400.0 405000.0 834600.0 ;
      RECT  394800.0 848400.0 405000.0 862200.0 ;
      RECT  394800.0 876000.0 405000.0 862200.0 ;
      RECT  394800.0 876000.0 405000.0 889800.0 ;
      RECT  394800.0 903600.0 405000.0 889800.0 ;
      RECT  394800.0 903600.0 405000.0 917400.0 ;
      RECT  394800.0 931200.0 405000.0 917400.0 ;
      RECT  394800.0 931200.0 405000.0 945000.0 ;
      RECT  394800.0 958800.0 405000.0 945000.0 ;
      RECT  394800.0 958800.0 405000.0 972600.0 ;
      RECT  394800.0 986400.0 405000.0 972600.0 ;
      RECT  394800.0 986400.0 405000.0 1000200.0 ;
      RECT  394800.0 1014000.0 405000.0 1000200.0 ;
      RECT  394800.0 1014000.0 405000.0 1027800.0 ;
      RECT  394800.0 1041600.0 405000.0 1027800.0 ;
      RECT  394800.0 1041600.0 405000.0 1055400.0 ;
      RECT  394800.0 1069200.0 405000.0 1055400.0 ;
      RECT  394800.0 1069200.0 405000.0 1083000.0 ;
      RECT  394800.0 1096800.0 405000.0 1083000.0 ;
      RECT  394800.0 1096800.0 405000.0 1110600.0 ;
      RECT  394800.0 1124400.0 405000.0 1110600.0 ;
      RECT  394800.0 1124400.0 405000.0 1138200.0 ;
      RECT  394800.0 1152000.0 405000.0 1138200.0 ;
      RECT  394800.0 1152000.0 405000.0 1165800.0 ;
      RECT  394800.0 1179600.0 405000.0 1165800.0 ;
      RECT  394800.0 1179600.0 405000.0 1193400.0 ;
      RECT  394800.0 1207200.0 405000.0 1193400.0 ;
      RECT  394800.0 1207200.0 405000.0 1221000.0 ;
      RECT  394800.0 1234800.0 405000.0 1221000.0 ;
      RECT  394800.0 1234800.0 405000.0 1248600.0 ;
      RECT  394800.0 1262400.0 405000.0 1248600.0 ;
      RECT  394800.0 1262400.0 405000.0 1276200.0 ;
      RECT  394800.0 1290000.0 405000.0 1276200.0 ;
      RECT  394800.0 1290000.0 405000.0 1303800.0 ;
      RECT  394800.0 1317600.0 405000.0 1303800.0 ;
      RECT  394800.0 1317600.0 405000.0 1331400.0 ;
      RECT  394800.0 1345200.0 405000.0 1331400.0 ;
      RECT  394800.0 1345200.0 405000.0 1359000.0 ;
      RECT  394800.0 1372800.0 405000.0 1359000.0 ;
      RECT  394800.0 1372800.0 405000.0 1386600.0 ;
      RECT  394800.0 1400400.0 405000.0 1386600.0 ;
      RECT  394800.0 1400400.0 405000.0 1414200.0 ;
      RECT  394800.0 1428000.0 405000.0 1414200.0 ;
      RECT  394800.0 1428000.0 405000.0 1441800.0 ;
      RECT  394800.0 1455600.0 405000.0 1441800.0 ;
      RECT  394800.0 1455600.0 405000.0 1469400.0 ;
      RECT  394800.0 1483200.0 405000.0 1469400.0 ;
      RECT  394800.0 1483200.0 405000.0 1497000.0 ;
      RECT  394800.0 1510800.0 405000.0 1497000.0 ;
      RECT  394800.0 1510800.0 405000.0 1524600.0 ;
      RECT  394800.0 1538400.0 405000.0 1524600.0 ;
      RECT  394800.0 1538400.0 405000.0 1552200.0 ;
      RECT  394800.0 1566000.0 405000.0 1552200.0 ;
      RECT  394800.0 1566000.0 405000.0 1579800.0 ;
      RECT  394800.0 1593600.0 405000.0 1579800.0 ;
      RECT  394800.0 1593600.0 405000.0 1607400.0 ;
      RECT  394800.0 1621200.0 405000.0 1607400.0 ;
      RECT  394800.0 1621200.0 405000.0 1635000.0 ;
      RECT  394800.0 1648800.0 405000.0 1635000.0 ;
      RECT  394800.0 1648800.0 405000.0 1662600.0 ;
      RECT  394800.0 1676400.0 405000.0 1662600.0 ;
      RECT  394800.0 1676400.0 405000.0 1690200.0 ;
      RECT  394800.0 1704000.0 405000.0 1690200.0 ;
      RECT  394800.0 1704000.0 405000.0 1717800.0 ;
      RECT  394800.0 1731600.0 405000.0 1717800.0 ;
      RECT  394800.0 1731600.0 405000.0 1745400.0 ;
      RECT  394800.0 1759200.0 405000.0 1745400.0 ;
      RECT  394800.0 1759200.0 405000.0 1773000.0 ;
      RECT  394800.0 1786800.0 405000.0 1773000.0 ;
      RECT  394800.0 1786800.0 405000.0 1800600.0 ;
      RECT  394800.0 1814400.0 405000.0 1800600.0 ;
      RECT  394800.0 1814400.0 405000.0 1828200.0 ;
      RECT  394800.0 1842000.0 405000.0 1828200.0 ;
      RECT  394800.0 1842000.0 405000.0 1855800.0 ;
      RECT  394800.0 1869600.0 405000.0 1855800.0 ;
      RECT  394800.0 1869600.0 405000.0 1883400.0 ;
      RECT  394800.0 1897200.0 405000.0 1883400.0 ;
      RECT  394800.0 1897200.0 405000.0 1911000.0 ;
      RECT  394800.0 1924800.0 405000.0 1911000.0 ;
      RECT  394800.0 1924800.0 405000.0 1938600.0 ;
      RECT  394800.0 1952400.0 405000.0 1938600.0 ;
      RECT  394800.0 1952400.0 405000.0 1966200.0 ;
      RECT  394800.0 1980000.0 405000.0 1966200.0 ;
      RECT  394800.0 1980000.0 405000.0 1993800.0 ;
      RECT  394800.0 2007600.0 405000.0 1993800.0 ;
      RECT  394800.0 2007600.0 405000.0 2021400.0 ;
      RECT  394800.0 2035200.0 405000.0 2021400.0 ;
      RECT  394800.0 2035200.0 405000.0 2049000.0 ;
      RECT  394800.0 2062800.0 405000.0 2049000.0 ;
      RECT  394800.0 2062800.0 405000.0 2076600.0 ;
      RECT  394800.0 2090400.0 405000.0 2076600.0 ;
      RECT  394800.0 2090400.0 405000.0 2104200.0 ;
      RECT  394800.0 2118000.0 405000.0 2104200.0 ;
      RECT  394800.0 2118000.0 405000.0 2131800.0 ;
      RECT  394800.0 2145600.0 405000.0 2131800.0 ;
      RECT  405000.0 379200.0 415200.0 393000.0 ;
      RECT  405000.0 406800.0 415200.0 393000.0 ;
      RECT  405000.0 406800.0 415200.0 420600.0 ;
      RECT  405000.0 434400.0 415200.0 420600.0 ;
      RECT  405000.0 434400.0 415200.0 448200.0 ;
      RECT  405000.0 462000.0 415200.0 448200.0 ;
      RECT  405000.0 462000.0 415200.0 475800.0 ;
      RECT  405000.0 489600.0 415200.0 475800.0 ;
      RECT  405000.0 489600.0 415200.0 503400.0 ;
      RECT  405000.0 517200.0 415200.0 503400.0 ;
      RECT  405000.0 517200.0 415200.0 531000.0 ;
      RECT  405000.0 544800.0 415200.0 531000.0 ;
      RECT  405000.0 544800.0 415200.0 558600.0 ;
      RECT  405000.0 572400.0 415200.0 558600.0 ;
      RECT  405000.0 572400.0 415200.0 586200.0 ;
      RECT  405000.0 600000.0 415200.0 586200.0 ;
      RECT  405000.0 600000.0 415200.0 613800.0 ;
      RECT  405000.0 627600.0 415200.0 613800.0 ;
      RECT  405000.0 627600.0 415200.0 641400.0 ;
      RECT  405000.0 655200.0 415200.0 641400.0 ;
      RECT  405000.0 655200.0 415200.0 669000.0 ;
      RECT  405000.0 682800.0 415200.0 669000.0 ;
      RECT  405000.0 682800.0 415200.0 696600.0 ;
      RECT  405000.0 710400.0 415200.0 696600.0 ;
      RECT  405000.0 710400.0 415200.0 724200.0 ;
      RECT  405000.0 738000.0 415200.0 724200.0 ;
      RECT  405000.0 738000.0 415200.0 751800.0 ;
      RECT  405000.0 765600.0 415200.0 751800.0 ;
      RECT  405000.0 765600.0 415200.0 779400.0 ;
      RECT  405000.0 793200.0 415200.0 779400.0 ;
      RECT  405000.0 793200.0 415200.0 807000.0 ;
      RECT  405000.0 820800.0 415200.0 807000.0 ;
      RECT  405000.0 820800.0 415200.0 834600.0 ;
      RECT  405000.0 848400.0 415200.0 834600.0 ;
      RECT  405000.0 848400.0 415200.0 862200.0 ;
      RECT  405000.0 876000.0 415200.0 862200.0 ;
      RECT  405000.0 876000.0 415200.0 889800.0 ;
      RECT  405000.0 903600.0 415200.0 889800.0 ;
      RECT  405000.0 903600.0 415200.0 917400.0 ;
      RECT  405000.0 931200.0 415200.0 917400.0 ;
      RECT  405000.0 931200.0 415200.0 945000.0 ;
      RECT  405000.0 958800.0 415200.0 945000.0 ;
      RECT  405000.0 958800.0 415200.0 972600.0 ;
      RECT  405000.0 986400.0 415200.0 972600.0 ;
      RECT  405000.0 986400.0 415200.0 1000200.0 ;
      RECT  405000.0 1014000.0 415200.0 1000200.0 ;
      RECT  405000.0 1014000.0 415200.0 1027800.0 ;
      RECT  405000.0 1041600.0 415200.0 1027800.0 ;
      RECT  405000.0 1041600.0 415200.0 1055400.0 ;
      RECT  405000.0 1069200.0 415200.0 1055400.0 ;
      RECT  405000.0 1069200.0 415200.0 1083000.0 ;
      RECT  405000.0 1096800.0 415200.0 1083000.0 ;
      RECT  405000.0 1096800.0 415200.0 1110600.0 ;
      RECT  405000.0 1124400.0 415200.0 1110600.0 ;
      RECT  405000.0 1124400.0 415200.0 1138200.0 ;
      RECT  405000.0 1152000.0 415200.0 1138200.0 ;
      RECT  405000.0 1152000.0 415200.0 1165800.0 ;
      RECT  405000.0 1179600.0 415200.0 1165800.0 ;
      RECT  405000.0 1179600.0 415200.0 1193400.0 ;
      RECT  405000.0 1207200.0 415200.0 1193400.0 ;
      RECT  405000.0 1207200.0 415200.0 1221000.0 ;
      RECT  405000.0 1234800.0 415200.0 1221000.0 ;
      RECT  405000.0 1234800.0 415200.0 1248600.0 ;
      RECT  405000.0 1262400.0 415200.0 1248600.0 ;
      RECT  405000.0 1262400.0 415200.0 1276200.0 ;
      RECT  405000.0 1290000.0 415200.0 1276200.0 ;
      RECT  405000.0 1290000.0 415200.0 1303800.0 ;
      RECT  405000.0 1317600.0 415200.0 1303800.0 ;
      RECT  405000.0 1317600.0 415200.0 1331400.0 ;
      RECT  405000.0 1345200.0 415200.0 1331400.0 ;
      RECT  405000.0 1345200.0 415200.0 1359000.0 ;
      RECT  405000.0 1372800.0 415200.0 1359000.0 ;
      RECT  405000.0 1372800.0 415200.0 1386600.0 ;
      RECT  405000.0 1400400.0 415200.0 1386600.0 ;
      RECT  405000.0 1400400.0 415200.0 1414200.0 ;
      RECT  405000.0 1428000.0 415200.0 1414200.0 ;
      RECT  405000.0 1428000.0 415200.0 1441800.0 ;
      RECT  405000.0 1455600.0 415200.0 1441800.0 ;
      RECT  405000.0 1455600.0 415200.0 1469400.0 ;
      RECT  405000.0 1483200.0 415200.0 1469400.0 ;
      RECT  405000.0 1483200.0 415200.0 1497000.0 ;
      RECT  405000.0 1510800.0 415200.0 1497000.0 ;
      RECT  405000.0 1510800.0 415200.0 1524600.0 ;
      RECT  405000.0 1538400.0 415200.0 1524600.0 ;
      RECT  405000.0 1538400.0 415200.0 1552200.0 ;
      RECT  405000.0 1566000.0 415200.0 1552200.0 ;
      RECT  405000.0 1566000.0 415200.0 1579800.0 ;
      RECT  405000.0 1593600.0 415200.0 1579800.0 ;
      RECT  405000.0 1593600.0 415200.0 1607400.0 ;
      RECT  405000.0 1621200.0 415200.0 1607400.0 ;
      RECT  405000.0 1621200.0 415200.0 1635000.0 ;
      RECT  405000.0 1648800.0 415200.0 1635000.0 ;
      RECT  405000.0 1648800.0 415200.0 1662600.0 ;
      RECT  405000.0 1676400.0 415200.0 1662600.0 ;
      RECT  405000.0 1676400.0 415200.0 1690200.0 ;
      RECT  405000.0 1704000.0 415200.0 1690200.0 ;
      RECT  405000.0 1704000.0 415200.0 1717800.0 ;
      RECT  405000.0 1731600.0 415200.0 1717800.0 ;
      RECT  405000.0 1731600.0 415200.0 1745400.0 ;
      RECT  405000.0 1759200.0 415200.0 1745400.0 ;
      RECT  405000.0 1759200.0 415200.0 1773000.0 ;
      RECT  405000.0 1786800.0 415200.0 1773000.0 ;
      RECT  405000.0 1786800.0 415200.0 1800600.0 ;
      RECT  405000.0 1814400.0 415200.0 1800600.0 ;
      RECT  405000.0 1814400.0 415200.0 1828200.0 ;
      RECT  405000.0 1842000.0 415200.0 1828200.0 ;
      RECT  405000.0 1842000.0 415200.0 1855800.0 ;
      RECT  405000.0 1869600.0 415200.0 1855800.0 ;
      RECT  405000.0 1869600.0 415200.0 1883400.0 ;
      RECT  405000.0 1897200.0 415200.0 1883400.0 ;
      RECT  405000.0 1897200.0 415200.0 1911000.0 ;
      RECT  405000.0 1924800.0 415200.0 1911000.0 ;
      RECT  405000.0 1924800.0 415200.0 1938600.0 ;
      RECT  405000.0 1952400.0 415200.0 1938600.0 ;
      RECT  405000.0 1952400.0 415200.0 1966200.0 ;
      RECT  405000.0 1980000.0 415200.0 1966200.0 ;
      RECT  405000.0 1980000.0 415200.0 1993800.0 ;
      RECT  405000.0 2007600.0 415200.0 1993800.0 ;
      RECT  405000.0 2007600.0 415200.0 2021400.0 ;
      RECT  405000.0 2035200.0 415200.0 2021400.0 ;
      RECT  405000.0 2035200.0 415200.0 2049000.0 ;
      RECT  405000.0 2062800.0 415200.0 2049000.0 ;
      RECT  405000.0 2062800.0 415200.0 2076600.0 ;
      RECT  405000.0 2090400.0 415200.0 2076600.0 ;
      RECT  405000.0 2090400.0 415200.0 2104200.0 ;
      RECT  405000.0 2118000.0 415200.0 2104200.0 ;
      RECT  405000.0 2118000.0 415200.0 2131800.0 ;
      RECT  405000.0 2145600.0 415200.0 2131800.0 ;
      RECT  415200.0 379200.0 425400.0 393000.0 ;
      RECT  415200.0 406800.0 425400.0 393000.0 ;
      RECT  415200.0 406800.0 425400.0 420600.0 ;
      RECT  415200.0 434400.0 425400.0 420600.0 ;
      RECT  415200.0 434400.0 425400.0 448200.0 ;
      RECT  415200.0 462000.0 425400.0 448200.0 ;
      RECT  415200.0 462000.0 425400.0 475800.0 ;
      RECT  415200.0 489600.0 425400.0 475800.0 ;
      RECT  415200.0 489600.0 425400.0 503400.0 ;
      RECT  415200.0 517200.0 425400.0 503400.0 ;
      RECT  415200.0 517200.0 425400.0 531000.0 ;
      RECT  415200.0 544800.0 425400.0 531000.0 ;
      RECT  415200.0 544800.0 425400.0 558600.0 ;
      RECT  415200.0 572400.0 425400.0 558600.0 ;
      RECT  415200.0 572400.0 425400.0 586200.0 ;
      RECT  415200.0 600000.0 425400.0 586200.0 ;
      RECT  415200.0 600000.0 425400.0 613800.0 ;
      RECT  415200.0 627600.0 425400.0 613800.0 ;
      RECT  415200.0 627600.0 425400.0 641400.0 ;
      RECT  415200.0 655200.0 425400.0 641400.0 ;
      RECT  415200.0 655200.0 425400.0 669000.0 ;
      RECT  415200.0 682800.0 425400.0 669000.0 ;
      RECT  415200.0 682800.0 425400.0 696600.0 ;
      RECT  415200.0 710400.0 425400.0 696600.0 ;
      RECT  415200.0 710400.0 425400.0 724200.0 ;
      RECT  415200.0 738000.0 425400.0 724200.0 ;
      RECT  415200.0 738000.0 425400.0 751800.0 ;
      RECT  415200.0 765600.0 425400.0 751800.0 ;
      RECT  415200.0 765600.0 425400.0 779400.0 ;
      RECT  415200.0 793200.0 425400.0 779400.0 ;
      RECT  415200.0 793200.0 425400.0 807000.0 ;
      RECT  415200.0 820800.0 425400.0 807000.0 ;
      RECT  415200.0 820800.0 425400.0 834600.0 ;
      RECT  415200.0 848400.0 425400.0 834600.0 ;
      RECT  415200.0 848400.0 425400.0 862200.0 ;
      RECT  415200.0 876000.0 425400.0 862200.0 ;
      RECT  415200.0 876000.0 425400.0 889800.0 ;
      RECT  415200.0 903600.0 425400.0 889800.0 ;
      RECT  415200.0 903600.0 425400.0 917400.0 ;
      RECT  415200.0 931200.0 425400.0 917400.0 ;
      RECT  415200.0 931200.0 425400.0 945000.0 ;
      RECT  415200.0 958800.0 425400.0 945000.0 ;
      RECT  415200.0 958800.0 425400.0 972600.0 ;
      RECT  415200.0 986400.0 425400.0 972600.0 ;
      RECT  415200.0 986400.0 425400.0 1000200.0 ;
      RECT  415200.0 1014000.0 425400.0 1000200.0 ;
      RECT  415200.0 1014000.0 425400.0 1027800.0 ;
      RECT  415200.0 1041600.0 425400.0 1027800.0 ;
      RECT  415200.0 1041600.0 425400.0 1055400.0 ;
      RECT  415200.0 1069200.0 425400.0 1055400.0 ;
      RECT  415200.0 1069200.0 425400.0 1083000.0 ;
      RECT  415200.0 1096800.0 425400.0 1083000.0 ;
      RECT  415200.0 1096800.0 425400.0 1110600.0 ;
      RECT  415200.0 1124400.0 425400.0 1110600.0 ;
      RECT  415200.0 1124400.0 425400.0 1138200.0 ;
      RECT  415200.0 1152000.0 425400.0 1138200.0 ;
      RECT  415200.0 1152000.0 425400.0 1165800.0 ;
      RECT  415200.0 1179600.0 425400.0 1165800.0 ;
      RECT  415200.0 1179600.0 425400.0 1193400.0 ;
      RECT  415200.0 1207200.0 425400.0 1193400.0 ;
      RECT  415200.0 1207200.0 425400.0 1221000.0 ;
      RECT  415200.0 1234800.0 425400.0 1221000.0 ;
      RECT  415200.0 1234800.0 425400.0 1248600.0 ;
      RECT  415200.0 1262400.0 425400.0 1248600.0 ;
      RECT  415200.0 1262400.0 425400.0 1276200.0 ;
      RECT  415200.0 1290000.0 425400.0 1276200.0 ;
      RECT  415200.0 1290000.0 425400.0 1303800.0 ;
      RECT  415200.0 1317600.0 425400.0 1303800.0 ;
      RECT  415200.0 1317600.0 425400.0 1331400.0 ;
      RECT  415200.0 1345200.0 425400.0 1331400.0 ;
      RECT  415200.0 1345200.0 425400.0 1359000.0 ;
      RECT  415200.0 1372800.0 425400.0 1359000.0 ;
      RECT  415200.0 1372800.0 425400.0 1386600.0 ;
      RECT  415200.0 1400400.0 425400.0 1386600.0 ;
      RECT  415200.0 1400400.0 425400.0 1414200.0 ;
      RECT  415200.0 1428000.0 425400.0 1414200.0 ;
      RECT  415200.0 1428000.0 425400.0 1441800.0 ;
      RECT  415200.0 1455600.0 425400.0 1441800.0 ;
      RECT  415200.0 1455600.0 425400.0 1469400.0 ;
      RECT  415200.0 1483200.0 425400.0 1469400.0 ;
      RECT  415200.0 1483200.0 425400.0 1497000.0 ;
      RECT  415200.0 1510800.0 425400.0 1497000.0 ;
      RECT  415200.0 1510800.0 425400.0 1524600.0 ;
      RECT  415200.0 1538400.0 425400.0 1524600.0 ;
      RECT  415200.0 1538400.0 425400.0 1552200.0 ;
      RECT  415200.0 1566000.0 425400.0 1552200.0 ;
      RECT  415200.0 1566000.0 425400.0 1579800.0 ;
      RECT  415200.0 1593600.0 425400.0 1579800.0 ;
      RECT  415200.0 1593600.0 425400.0 1607400.0 ;
      RECT  415200.0 1621200.0 425400.0 1607400.0 ;
      RECT  415200.0 1621200.0 425400.0 1635000.0 ;
      RECT  415200.0 1648800.0 425400.0 1635000.0 ;
      RECT  415200.0 1648800.0 425400.0 1662600.0 ;
      RECT  415200.0 1676400.0 425400.0 1662600.0 ;
      RECT  415200.0 1676400.0 425400.0 1690200.0 ;
      RECT  415200.0 1704000.0 425400.0 1690200.0 ;
      RECT  415200.0 1704000.0 425400.0 1717800.0 ;
      RECT  415200.0 1731600.0 425400.0 1717800.0 ;
      RECT  415200.0 1731600.0 425400.0 1745400.0 ;
      RECT  415200.0 1759200.0 425400.0 1745400.0 ;
      RECT  415200.0 1759200.0 425400.0 1773000.0 ;
      RECT  415200.0 1786800.0 425400.0 1773000.0 ;
      RECT  415200.0 1786800.0 425400.0 1800600.0 ;
      RECT  415200.0 1814400.0 425400.0 1800600.0 ;
      RECT  415200.0 1814400.0 425400.0 1828200.0 ;
      RECT  415200.0 1842000.0 425400.0 1828200.0 ;
      RECT  415200.0 1842000.0 425400.0 1855800.0 ;
      RECT  415200.0 1869600.0 425400.0 1855800.0 ;
      RECT  415200.0 1869600.0 425400.0 1883400.0 ;
      RECT  415200.0 1897200.0 425400.0 1883400.0 ;
      RECT  415200.0 1897200.0 425400.0 1911000.0 ;
      RECT  415200.0 1924800.0 425400.0 1911000.0 ;
      RECT  415200.0 1924800.0 425400.0 1938600.0 ;
      RECT  415200.0 1952400.0 425400.0 1938600.0 ;
      RECT  415200.0 1952400.0 425400.0 1966200.0 ;
      RECT  415200.0 1980000.0 425400.0 1966200.0 ;
      RECT  415200.0 1980000.0 425400.0 1993800.0 ;
      RECT  415200.0 2007600.0 425400.0 1993800.0 ;
      RECT  415200.0 2007600.0 425400.0 2021400.0 ;
      RECT  415200.0 2035200.0 425400.0 2021400.0 ;
      RECT  415200.0 2035200.0 425400.0 2049000.0 ;
      RECT  415200.0 2062800.0 425400.0 2049000.0 ;
      RECT  415200.0 2062800.0 425400.0 2076600.0 ;
      RECT  415200.0 2090400.0 425400.0 2076600.0 ;
      RECT  415200.0 2090400.0 425400.0 2104200.0 ;
      RECT  415200.0 2118000.0 425400.0 2104200.0 ;
      RECT  415200.0 2118000.0 425400.0 2131800.0 ;
      RECT  415200.0 2145600.0 425400.0 2131800.0 ;
      RECT  425400.0 379200.0 435600.0 393000.0 ;
      RECT  425400.0 406800.0 435600.0 393000.0 ;
      RECT  425400.0 406800.0 435600.0 420600.0 ;
      RECT  425400.0 434400.0 435600.0 420600.0 ;
      RECT  425400.0 434400.0 435600.0 448200.0 ;
      RECT  425400.0 462000.0 435600.0 448200.0 ;
      RECT  425400.0 462000.0 435600.0 475800.0 ;
      RECT  425400.0 489600.0 435600.0 475800.0 ;
      RECT  425400.0 489600.0 435600.0 503400.0 ;
      RECT  425400.0 517200.0 435600.0 503400.0 ;
      RECT  425400.0 517200.0 435600.0 531000.0 ;
      RECT  425400.0 544800.0 435600.0 531000.0 ;
      RECT  425400.0 544800.0 435600.0 558600.0 ;
      RECT  425400.0 572400.0 435600.0 558600.0 ;
      RECT  425400.0 572400.0 435600.0 586200.0 ;
      RECT  425400.0 600000.0 435600.0 586200.0 ;
      RECT  425400.0 600000.0 435600.0 613800.0 ;
      RECT  425400.0 627600.0 435600.0 613800.0 ;
      RECT  425400.0 627600.0 435600.0 641400.0 ;
      RECT  425400.0 655200.0 435600.0 641400.0 ;
      RECT  425400.0 655200.0 435600.0 669000.0 ;
      RECT  425400.0 682800.0 435600.0 669000.0 ;
      RECT  425400.0 682800.0 435600.0 696600.0 ;
      RECT  425400.0 710400.0 435600.0 696600.0 ;
      RECT  425400.0 710400.0 435600.0 724200.0 ;
      RECT  425400.0 738000.0 435600.0 724200.0 ;
      RECT  425400.0 738000.0 435600.0 751800.0 ;
      RECT  425400.0 765600.0 435600.0 751800.0 ;
      RECT  425400.0 765600.0 435600.0 779400.0 ;
      RECT  425400.0 793200.0 435600.0 779400.0 ;
      RECT  425400.0 793200.0 435600.0 807000.0 ;
      RECT  425400.0 820800.0 435600.0 807000.0 ;
      RECT  425400.0 820800.0 435600.0 834600.0 ;
      RECT  425400.0 848400.0 435600.0 834600.0 ;
      RECT  425400.0 848400.0 435600.0 862200.0 ;
      RECT  425400.0 876000.0 435600.0 862200.0 ;
      RECT  425400.0 876000.0 435600.0 889800.0 ;
      RECT  425400.0 903600.0 435600.0 889800.0 ;
      RECT  425400.0 903600.0 435600.0 917400.0 ;
      RECT  425400.0 931200.0 435600.0 917400.0 ;
      RECT  425400.0 931200.0 435600.0 945000.0 ;
      RECT  425400.0 958800.0 435600.0 945000.0 ;
      RECT  425400.0 958800.0 435600.0 972600.0 ;
      RECT  425400.0 986400.0 435600.0 972600.0 ;
      RECT  425400.0 986400.0 435600.0 1000200.0 ;
      RECT  425400.0 1014000.0 435600.0 1000200.0 ;
      RECT  425400.0 1014000.0 435600.0 1027800.0 ;
      RECT  425400.0 1041600.0 435600.0 1027800.0 ;
      RECT  425400.0 1041600.0 435600.0 1055400.0 ;
      RECT  425400.0 1069200.0 435600.0 1055400.0 ;
      RECT  425400.0 1069200.0 435600.0 1083000.0 ;
      RECT  425400.0 1096800.0 435600.0 1083000.0 ;
      RECT  425400.0 1096800.0 435600.0 1110600.0 ;
      RECT  425400.0 1124400.0 435600.0 1110600.0 ;
      RECT  425400.0 1124400.0 435600.0 1138200.0 ;
      RECT  425400.0 1152000.0 435600.0 1138200.0 ;
      RECT  425400.0 1152000.0 435600.0 1165800.0 ;
      RECT  425400.0 1179600.0 435600.0 1165800.0 ;
      RECT  425400.0 1179600.0 435600.0 1193400.0 ;
      RECT  425400.0 1207200.0 435600.0 1193400.0 ;
      RECT  425400.0 1207200.0 435600.0 1221000.0 ;
      RECT  425400.0 1234800.0 435600.0 1221000.0 ;
      RECT  425400.0 1234800.0 435600.0 1248600.0 ;
      RECT  425400.0 1262400.0 435600.0 1248600.0 ;
      RECT  425400.0 1262400.0 435600.0 1276200.0 ;
      RECT  425400.0 1290000.0 435600.0 1276200.0 ;
      RECT  425400.0 1290000.0 435600.0 1303800.0 ;
      RECT  425400.0 1317600.0 435600.0 1303800.0 ;
      RECT  425400.0 1317600.0 435600.0 1331400.0 ;
      RECT  425400.0 1345200.0 435600.0 1331400.0 ;
      RECT  425400.0 1345200.0 435600.0 1359000.0 ;
      RECT  425400.0 1372800.0 435600.0 1359000.0 ;
      RECT  425400.0 1372800.0 435600.0 1386600.0 ;
      RECT  425400.0 1400400.0 435600.0 1386600.0 ;
      RECT  425400.0 1400400.0 435600.0 1414200.0 ;
      RECT  425400.0 1428000.0 435600.0 1414200.0 ;
      RECT  425400.0 1428000.0 435600.0 1441800.0 ;
      RECT  425400.0 1455600.0 435600.0 1441800.0 ;
      RECT  425400.0 1455600.0 435600.0 1469400.0 ;
      RECT  425400.0 1483200.0 435600.0 1469400.0 ;
      RECT  425400.0 1483200.0 435600.0 1497000.0 ;
      RECT  425400.0 1510800.0 435600.0 1497000.0 ;
      RECT  425400.0 1510800.0 435600.0 1524600.0 ;
      RECT  425400.0 1538400.0 435600.0 1524600.0 ;
      RECT  425400.0 1538400.0 435600.0 1552200.0 ;
      RECT  425400.0 1566000.0 435600.0 1552200.0 ;
      RECT  425400.0 1566000.0 435600.0 1579800.0 ;
      RECT  425400.0 1593600.0 435600.0 1579800.0 ;
      RECT  425400.0 1593600.0 435600.0 1607400.0 ;
      RECT  425400.0 1621200.0 435600.0 1607400.0 ;
      RECT  425400.0 1621200.0 435600.0 1635000.0 ;
      RECT  425400.0 1648800.0 435600.0 1635000.0 ;
      RECT  425400.0 1648800.0 435600.0 1662600.0 ;
      RECT  425400.0 1676400.0 435600.0 1662600.0 ;
      RECT  425400.0 1676400.0 435600.0 1690200.0 ;
      RECT  425400.0 1704000.0 435600.0 1690200.0 ;
      RECT  425400.0 1704000.0 435600.0 1717800.0 ;
      RECT  425400.0 1731600.0 435600.0 1717800.0 ;
      RECT  425400.0 1731600.0 435600.0 1745400.0 ;
      RECT  425400.0 1759200.0 435600.0 1745400.0 ;
      RECT  425400.0 1759200.0 435600.0 1773000.0 ;
      RECT  425400.0 1786800.0 435600.0 1773000.0 ;
      RECT  425400.0 1786800.0 435600.0 1800600.0 ;
      RECT  425400.0 1814400.0 435600.0 1800600.0 ;
      RECT  425400.0 1814400.0 435600.0 1828200.0 ;
      RECT  425400.0 1842000.0 435600.0 1828200.0 ;
      RECT  425400.0 1842000.0 435600.0 1855800.0 ;
      RECT  425400.0 1869600.0 435600.0 1855800.0 ;
      RECT  425400.0 1869600.0 435600.0 1883400.0 ;
      RECT  425400.0 1897200.0 435600.0 1883400.0 ;
      RECT  425400.0 1897200.0 435600.0 1911000.0 ;
      RECT  425400.0 1924800.0 435600.0 1911000.0 ;
      RECT  425400.0 1924800.0 435600.0 1938600.0 ;
      RECT  425400.0 1952400.0 435600.0 1938600.0 ;
      RECT  425400.0 1952400.0 435600.0 1966200.0 ;
      RECT  425400.0 1980000.0 435600.0 1966200.0 ;
      RECT  425400.0 1980000.0 435600.0 1993800.0 ;
      RECT  425400.0 2007600.0 435600.0 1993800.0 ;
      RECT  425400.0 2007600.0 435600.0 2021400.0 ;
      RECT  425400.0 2035200.0 435600.0 2021400.0 ;
      RECT  425400.0 2035200.0 435600.0 2049000.0 ;
      RECT  425400.0 2062800.0 435600.0 2049000.0 ;
      RECT  425400.0 2062800.0 435600.0 2076600.0 ;
      RECT  425400.0 2090400.0 435600.0 2076600.0 ;
      RECT  425400.0 2090400.0 435600.0 2104200.0 ;
      RECT  425400.0 2118000.0 435600.0 2104200.0 ;
      RECT  425400.0 2118000.0 435600.0 2131800.0 ;
      RECT  425400.0 2145600.0 435600.0 2131800.0 ;
      RECT  435600.0 379200.0 445800.0 393000.0 ;
      RECT  435600.0 406800.0 445800.0 393000.0 ;
      RECT  435600.0 406800.0 445800.0 420600.0 ;
      RECT  435600.0 434400.0 445800.0 420600.0 ;
      RECT  435600.0 434400.0 445800.0 448200.0 ;
      RECT  435600.0 462000.0 445800.0 448200.0 ;
      RECT  435600.0 462000.0 445800.0 475800.0 ;
      RECT  435600.0 489600.0 445800.0 475800.0 ;
      RECT  435600.0 489600.0 445800.0 503400.0 ;
      RECT  435600.0 517200.0 445800.0 503400.0 ;
      RECT  435600.0 517200.0 445800.0 531000.0 ;
      RECT  435600.0 544800.0 445800.0 531000.0 ;
      RECT  435600.0 544800.0 445800.0 558600.0 ;
      RECT  435600.0 572400.0 445800.0 558600.0 ;
      RECT  435600.0 572400.0 445800.0 586200.0 ;
      RECT  435600.0 600000.0 445800.0 586200.0 ;
      RECT  435600.0 600000.0 445800.0 613800.0 ;
      RECT  435600.0 627600.0 445800.0 613800.0 ;
      RECT  435600.0 627600.0 445800.0 641400.0 ;
      RECT  435600.0 655200.0 445800.0 641400.0 ;
      RECT  435600.0 655200.0 445800.0 669000.0 ;
      RECT  435600.0 682800.0 445800.0 669000.0 ;
      RECT  435600.0 682800.0 445800.0 696600.0 ;
      RECT  435600.0 710400.0 445800.0 696600.0 ;
      RECT  435600.0 710400.0 445800.0 724200.0 ;
      RECT  435600.0 738000.0 445800.0 724200.0 ;
      RECT  435600.0 738000.0 445800.0 751800.0 ;
      RECT  435600.0 765600.0 445800.0 751800.0 ;
      RECT  435600.0 765600.0 445800.0 779400.0 ;
      RECT  435600.0 793200.0 445800.0 779400.0 ;
      RECT  435600.0 793200.0 445800.0 807000.0 ;
      RECT  435600.0 820800.0 445800.0 807000.0 ;
      RECT  435600.0 820800.0 445800.0 834600.0 ;
      RECT  435600.0 848400.0 445800.0 834600.0 ;
      RECT  435600.0 848400.0 445800.0 862200.0 ;
      RECT  435600.0 876000.0 445800.0 862200.0 ;
      RECT  435600.0 876000.0 445800.0 889800.0 ;
      RECT  435600.0 903600.0 445800.0 889800.0 ;
      RECT  435600.0 903600.0 445800.0 917400.0 ;
      RECT  435600.0 931200.0 445800.0 917400.0 ;
      RECT  435600.0 931200.0 445800.0 945000.0 ;
      RECT  435600.0 958800.0 445800.0 945000.0 ;
      RECT  435600.0 958800.0 445800.0 972600.0 ;
      RECT  435600.0 986400.0 445800.0 972600.0 ;
      RECT  435600.0 986400.0 445800.0 1000200.0 ;
      RECT  435600.0 1014000.0 445800.0 1000200.0 ;
      RECT  435600.0 1014000.0 445800.0 1027800.0 ;
      RECT  435600.0 1041600.0 445800.0 1027800.0 ;
      RECT  435600.0 1041600.0 445800.0 1055400.0 ;
      RECT  435600.0 1069200.0 445800.0 1055400.0 ;
      RECT  435600.0 1069200.0 445800.0 1083000.0 ;
      RECT  435600.0 1096800.0 445800.0 1083000.0 ;
      RECT  435600.0 1096800.0 445800.0 1110600.0 ;
      RECT  435600.0 1124400.0 445800.0 1110600.0 ;
      RECT  435600.0 1124400.0 445800.0 1138200.0 ;
      RECT  435600.0 1152000.0 445800.0 1138200.0 ;
      RECT  435600.0 1152000.0 445800.0 1165800.0 ;
      RECT  435600.0 1179600.0 445800.0 1165800.0 ;
      RECT  435600.0 1179600.0 445800.0 1193400.0 ;
      RECT  435600.0 1207200.0 445800.0 1193400.0 ;
      RECT  435600.0 1207200.0 445800.0 1221000.0 ;
      RECT  435600.0 1234800.0 445800.0 1221000.0 ;
      RECT  435600.0 1234800.0 445800.0 1248600.0 ;
      RECT  435600.0 1262400.0 445800.0 1248600.0 ;
      RECT  435600.0 1262400.0 445800.0 1276200.0 ;
      RECT  435600.0 1290000.0 445800.0 1276200.0 ;
      RECT  435600.0 1290000.0 445800.0 1303800.0 ;
      RECT  435600.0 1317600.0 445800.0 1303800.0 ;
      RECT  435600.0 1317600.0 445800.0 1331400.0 ;
      RECT  435600.0 1345200.0 445800.0 1331400.0 ;
      RECT  435600.0 1345200.0 445800.0 1359000.0 ;
      RECT  435600.0 1372800.0 445800.0 1359000.0 ;
      RECT  435600.0 1372800.0 445800.0 1386600.0 ;
      RECT  435600.0 1400400.0 445800.0 1386600.0 ;
      RECT  435600.0 1400400.0 445800.0 1414200.0 ;
      RECT  435600.0 1428000.0 445800.0 1414200.0 ;
      RECT  435600.0 1428000.0 445800.0 1441800.0 ;
      RECT  435600.0 1455600.0 445800.0 1441800.0 ;
      RECT  435600.0 1455600.0 445800.0 1469400.0 ;
      RECT  435600.0 1483200.0 445800.0 1469400.0 ;
      RECT  435600.0 1483200.0 445800.0 1497000.0 ;
      RECT  435600.0 1510800.0 445800.0 1497000.0 ;
      RECT  435600.0 1510800.0 445800.0 1524600.0 ;
      RECT  435600.0 1538400.0 445800.0 1524600.0 ;
      RECT  435600.0 1538400.0 445800.0 1552200.0 ;
      RECT  435600.0 1566000.0 445800.0 1552200.0 ;
      RECT  435600.0 1566000.0 445800.0 1579800.0 ;
      RECT  435600.0 1593600.0 445800.0 1579800.0 ;
      RECT  435600.0 1593600.0 445800.0 1607400.0 ;
      RECT  435600.0 1621200.0 445800.0 1607400.0 ;
      RECT  435600.0 1621200.0 445800.0 1635000.0 ;
      RECT  435600.0 1648800.0 445800.0 1635000.0 ;
      RECT  435600.0 1648800.0 445800.0 1662600.0 ;
      RECT  435600.0 1676400.0 445800.0 1662600.0 ;
      RECT  435600.0 1676400.0 445800.0 1690200.0 ;
      RECT  435600.0 1704000.0 445800.0 1690200.0 ;
      RECT  435600.0 1704000.0 445800.0 1717800.0 ;
      RECT  435600.0 1731600.0 445800.0 1717800.0 ;
      RECT  435600.0 1731600.0 445800.0 1745400.0 ;
      RECT  435600.0 1759200.0 445800.0 1745400.0 ;
      RECT  435600.0 1759200.0 445800.0 1773000.0 ;
      RECT  435600.0 1786800.0 445800.0 1773000.0 ;
      RECT  435600.0 1786800.0 445800.0 1800600.0 ;
      RECT  435600.0 1814400.0 445800.0 1800600.0 ;
      RECT  435600.0 1814400.0 445800.0 1828200.0 ;
      RECT  435600.0 1842000.0 445800.0 1828200.0 ;
      RECT  435600.0 1842000.0 445800.0 1855800.0 ;
      RECT  435600.0 1869600.0 445800.0 1855800.0 ;
      RECT  435600.0 1869600.0 445800.0 1883400.0 ;
      RECT  435600.0 1897200.0 445800.0 1883400.0 ;
      RECT  435600.0 1897200.0 445800.0 1911000.0 ;
      RECT  435600.0 1924800.0 445800.0 1911000.0 ;
      RECT  435600.0 1924800.0 445800.0 1938600.0 ;
      RECT  435600.0 1952400.0 445800.0 1938600.0 ;
      RECT  435600.0 1952400.0 445800.0 1966200.0 ;
      RECT  435600.0 1980000.0 445800.0 1966200.0 ;
      RECT  435600.0 1980000.0 445800.0 1993800.0 ;
      RECT  435600.0 2007600.0 445800.0 1993800.0 ;
      RECT  435600.0 2007600.0 445800.0 2021400.0 ;
      RECT  435600.0 2035200.0 445800.0 2021400.0 ;
      RECT  435600.0 2035200.0 445800.0 2049000.0 ;
      RECT  435600.0 2062800.0 445800.0 2049000.0 ;
      RECT  435600.0 2062800.0 445800.0 2076600.0 ;
      RECT  435600.0 2090400.0 445800.0 2076600.0 ;
      RECT  435600.0 2090400.0 445800.0 2104200.0 ;
      RECT  435600.0 2118000.0 445800.0 2104200.0 ;
      RECT  435600.0 2118000.0 445800.0 2131800.0 ;
      RECT  435600.0 2145600.0 445800.0 2131800.0 ;
      RECT  445800.0 379200.0 456000.0 393000.0 ;
      RECT  445800.0 406800.0 456000.0 393000.0 ;
      RECT  445800.0 406800.0 456000.0 420600.0 ;
      RECT  445800.0 434400.0 456000.0 420600.0 ;
      RECT  445800.0 434400.0 456000.0 448200.0 ;
      RECT  445800.0 462000.0 456000.0 448200.0 ;
      RECT  445800.0 462000.0 456000.0 475800.0 ;
      RECT  445800.0 489600.0 456000.0 475800.0 ;
      RECT  445800.0 489600.0 456000.0 503400.0 ;
      RECT  445800.0 517200.0 456000.0 503400.0 ;
      RECT  445800.0 517200.0 456000.0 531000.0 ;
      RECT  445800.0 544800.0 456000.0 531000.0 ;
      RECT  445800.0 544800.0 456000.0 558600.0 ;
      RECT  445800.0 572400.0 456000.0 558600.0 ;
      RECT  445800.0 572400.0 456000.0 586200.0 ;
      RECT  445800.0 600000.0 456000.0 586200.0 ;
      RECT  445800.0 600000.0 456000.0 613800.0 ;
      RECT  445800.0 627600.0 456000.0 613800.0 ;
      RECT  445800.0 627600.0 456000.0 641400.0 ;
      RECT  445800.0 655200.0 456000.0 641400.0 ;
      RECT  445800.0 655200.0 456000.0 669000.0 ;
      RECT  445800.0 682800.0 456000.0 669000.0 ;
      RECT  445800.0 682800.0 456000.0 696600.0 ;
      RECT  445800.0 710400.0 456000.0 696600.0 ;
      RECT  445800.0 710400.0 456000.0 724200.0 ;
      RECT  445800.0 738000.0 456000.0 724200.0 ;
      RECT  445800.0 738000.0 456000.0 751800.0 ;
      RECT  445800.0 765600.0 456000.0 751800.0 ;
      RECT  445800.0 765600.0 456000.0 779400.0 ;
      RECT  445800.0 793200.0 456000.0 779400.0 ;
      RECT  445800.0 793200.0 456000.0 807000.0 ;
      RECT  445800.0 820800.0 456000.0 807000.0 ;
      RECT  445800.0 820800.0 456000.0 834600.0 ;
      RECT  445800.0 848400.0 456000.0 834600.0 ;
      RECT  445800.0 848400.0 456000.0 862200.0 ;
      RECT  445800.0 876000.0 456000.0 862200.0 ;
      RECT  445800.0 876000.0 456000.0 889800.0 ;
      RECT  445800.0 903600.0 456000.0 889800.0 ;
      RECT  445800.0 903600.0 456000.0 917400.0 ;
      RECT  445800.0 931200.0 456000.0 917400.0 ;
      RECT  445800.0 931200.0 456000.0 945000.0 ;
      RECT  445800.0 958800.0 456000.0 945000.0 ;
      RECT  445800.0 958800.0 456000.0 972600.0 ;
      RECT  445800.0 986400.0 456000.0 972600.0 ;
      RECT  445800.0 986400.0 456000.0 1000200.0 ;
      RECT  445800.0 1014000.0 456000.0 1000200.0 ;
      RECT  445800.0 1014000.0 456000.0 1027800.0 ;
      RECT  445800.0 1041600.0 456000.0 1027800.0 ;
      RECT  445800.0 1041600.0 456000.0 1055400.0 ;
      RECT  445800.0 1069200.0 456000.0 1055400.0 ;
      RECT  445800.0 1069200.0 456000.0 1083000.0 ;
      RECT  445800.0 1096800.0 456000.0 1083000.0 ;
      RECT  445800.0 1096800.0 456000.0 1110600.0 ;
      RECT  445800.0 1124400.0 456000.0 1110600.0 ;
      RECT  445800.0 1124400.0 456000.0 1138200.0 ;
      RECT  445800.0 1152000.0 456000.0 1138200.0 ;
      RECT  445800.0 1152000.0 456000.0 1165800.0 ;
      RECT  445800.0 1179600.0 456000.0 1165800.0 ;
      RECT  445800.0 1179600.0 456000.0 1193400.0 ;
      RECT  445800.0 1207200.0 456000.0 1193400.0 ;
      RECT  445800.0 1207200.0 456000.0 1221000.0 ;
      RECT  445800.0 1234800.0 456000.0 1221000.0 ;
      RECT  445800.0 1234800.0 456000.0 1248600.0 ;
      RECT  445800.0 1262400.0 456000.0 1248600.0 ;
      RECT  445800.0 1262400.0 456000.0 1276200.0 ;
      RECT  445800.0 1290000.0 456000.0 1276200.0 ;
      RECT  445800.0 1290000.0 456000.0 1303800.0 ;
      RECT  445800.0 1317600.0 456000.0 1303800.0 ;
      RECT  445800.0 1317600.0 456000.0 1331400.0 ;
      RECT  445800.0 1345200.0 456000.0 1331400.0 ;
      RECT  445800.0 1345200.0 456000.0 1359000.0 ;
      RECT  445800.0 1372800.0 456000.0 1359000.0 ;
      RECT  445800.0 1372800.0 456000.0 1386600.0 ;
      RECT  445800.0 1400400.0 456000.0 1386600.0 ;
      RECT  445800.0 1400400.0 456000.0 1414200.0 ;
      RECT  445800.0 1428000.0 456000.0 1414200.0 ;
      RECT  445800.0 1428000.0 456000.0 1441800.0 ;
      RECT  445800.0 1455600.0 456000.0 1441800.0 ;
      RECT  445800.0 1455600.0 456000.0 1469400.0 ;
      RECT  445800.0 1483200.0 456000.0 1469400.0 ;
      RECT  445800.0 1483200.0 456000.0 1497000.0 ;
      RECT  445800.0 1510800.0 456000.0 1497000.0 ;
      RECT  445800.0 1510800.0 456000.0 1524600.0 ;
      RECT  445800.0 1538400.0 456000.0 1524600.0 ;
      RECT  445800.0 1538400.0 456000.0 1552200.0 ;
      RECT  445800.0 1566000.0 456000.0 1552200.0 ;
      RECT  445800.0 1566000.0 456000.0 1579800.0 ;
      RECT  445800.0 1593600.0 456000.0 1579800.0 ;
      RECT  445800.0 1593600.0 456000.0 1607400.0 ;
      RECT  445800.0 1621200.0 456000.0 1607400.0 ;
      RECT  445800.0 1621200.0 456000.0 1635000.0 ;
      RECT  445800.0 1648800.0 456000.0 1635000.0 ;
      RECT  445800.0 1648800.0 456000.0 1662600.0 ;
      RECT  445800.0 1676400.0 456000.0 1662600.0 ;
      RECT  445800.0 1676400.0 456000.0 1690200.0 ;
      RECT  445800.0 1704000.0 456000.0 1690200.0 ;
      RECT  445800.0 1704000.0 456000.0 1717800.0 ;
      RECT  445800.0 1731600.0 456000.0 1717800.0 ;
      RECT  445800.0 1731600.0 456000.0 1745400.0 ;
      RECT  445800.0 1759200.0 456000.0 1745400.0 ;
      RECT  445800.0 1759200.0 456000.0 1773000.0 ;
      RECT  445800.0 1786800.0 456000.0 1773000.0 ;
      RECT  445800.0 1786800.0 456000.0 1800600.0 ;
      RECT  445800.0 1814400.0 456000.0 1800600.0 ;
      RECT  445800.0 1814400.0 456000.0 1828200.0 ;
      RECT  445800.0 1842000.0 456000.0 1828200.0 ;
      RECT  445800.0 1842000.0 456000.0 1855800.0 ;
      RECT  445800.0 1869600.0 456000.0 1855800.0 ;
      RECT  445800.0 1869600.0 456000.0 1883400.0 ;
      RECT  445800.0 1897200.0 456000.0 1883400.0 ;
      RECT  445800.0 1897200.0 456000.0 1911000.0 ;
      RECT  445800.0 1924800.0 456000.0 1911000.0 ;
      RECT  445800.0 1924800.0 456000.0 1938600.0 ;
      RECT  445800.0 1952400.0 456000.0 1938600.0 ;
      RECT  445800.0 1952400.0 456000.0 1966200.0 ;
      RECT  445800.0 1980000.0 456000.0 1966200.0 ;
      RECT  445800.0 1980000.0 456000.0 1993800.0 ;
      RECT  445800.0 2007600.0 456000.0 1993800.0 ;
      RECT  445800.0 2007600.0 456000.0 2021400.0 ;
      RECT  445800.0 2035200.0 456000.0 2021400.0 ;
      RECT  445800.0 2035200.0 456000.0 2049000.0 ;
      RECT  445800.0 2062800.0 456000.0 2049000.0 ;
      RECT  445800.0 2062800.0 456000.0 2076600.0 ;
      RECT  445800.0 2090400.0 456000.0 2076600.0 ;
      RECT  445800.0 2090400.0 456000.0 2104200.0 ;
      RECT  445800.0 2118000.0 456000.0 2104200.0 ;
      RECT  445800.0 2118000.0 456000.0 2131800.0 ;
      RECT  445800.0 2145600.0 456000.0 2131800.0 ;
      RECT  456000.0 379200.0 466200.0 393000.0 ;
      RECT  456000.0 406800.0 466200.0 393000.0 ;
      RECT  456000.0 406800.0 466200.0 420600.0 ;
      RECT  456000.0 434400.0 466200.0 420600.0 ;
      RECT  456000.0 434400.0 466200.0 448200.0 ;
      RECT  456000.0 462000.0 466200.0 448200.0 ;
      RECT  456000.0 462000.0 466200.0 475800.0 ;
      RECT  456000.0 489600.0 466200.0 475800.0 ;
      RECT  456000.0 489600.0 466200.0 503400.0 ;
      RECT  456000.0 517200.0 466200.0 503400.0 ;
      RECT  456000.0 517200.0 466200.0 531000.0 ;
      RECT  456000.0 544800.0 466200.0 531000.0 ;
      RECT  456000.0 544800.0 466200.0 558600.0 ;
      RECT  456000.0 572400.0 466200.0 558600.0 ;
      RECT  456000.0 572400.0 466200.0 586200.0 ;
      RECT  456000.0 600000.0 466200.0 586200.0 ;
      RECT  456000.0 600000.0 466200.0 613800.0 ;
      RECT  456000.0 627600.0 466200.0 613800.0 ;
      RECT  456000.0 627600.0 466200.0 641400.0 ;
      RECT  456000.0 655200.0 466200.0 641400.0 ;
      RECT  456000.0 655200.0 466200.0 669000.0 ;
      RECT  456000.0 682800.0 466200.0 669000.0 ;
      RECT  456000.0 682800.0 466200.0 696600.0 ;
      RECT  456000.0 710400.0 466200.0 696600.0 ;
      RECT  456000.0 710400.0 466200.0 724200.0 ;
      RECT  456000.0 738000.0 466200.0 724200.0 ;
      RECT  456000.0 738000.0 466200.0 751800.0 ;
      RECT  456000.0 765600.0 466200.0 751800.0 ;
      RECT  456000.0 765600.0 466200.0 779400.0 ;
      RECT  456000.0 793200.0 466200.0 779400.0 ;
      RECT  456000.0 793200.0 466200.0 807000.0 ;
      RECT  456000.0 820800.0 466200.0 807000.0 ;
      RECT  456000.0 820800.0 466200.0 834600.0 ;
      RECT  456000.0 848400.0 466200.0 834600.0 ;
      RECT  456000.0 848400.0 466200.0 862200.0 ;
      RECT  456000.0 876000.0 466200.0 862200.0 ;
      RECT  456000.0 876000.0 466200.0 889800.0 ;
      RECT  456000.0 903600.0 466200.0 889800.0 ;
      RECT  456000.0 903600.0 466200.0 917400.0 ;
      RECT  456000.0 931200.0 466200.0 917400.0 ;
      RECT  456000.0 931200.0 466200.0 945000.0 ;
      RECT  456000.0 958800.0 466200.0 945000.0 ;
      RECT  456000.0 958800.0 466200.0 972600.0 ;
      RECT  456000.0 986400.0 466200.0 972600.0 ;
      RECT  456000.0 986400.0 466200.0 1000200.0 ;
      RECT  456000.0 1014000.0 466200.0 1000200.0 ;
      RECT  456000.0 1014000.0 466200.0 1027800.0 ;
      RECT  456000.0 1041600.0 466200.0 1027800.0 ;
      RECT  456000.0 1041600.0 466200.0 1055400.0 ;
      RECT  456000.0 1069200.0 466200.0 1055400.0 ;
      RECT  456000.0 1069200.0 466200.0 1083000.0 ;
      RECT  456000.0 1096800.0 466200.0 1083000.0 ;
      RECT  456000.0 1096800.0 466200.0 1110600.0 ;
      RECT  456000.0 1124400.0 466200.0 1110600.0 ;
      RECT  456000.0 1124400.0 466200.0 1138200.0 ;
      RECT  456000.0 1152000.0 466200.0 1138200.0 ;
      RECT  456000.0 1152000.0 466200.0 1165800.0 ;
      RECT  456000.0 1179600.0 466200.0 1165800.0 ;
      RECT  456000.0 1179600.0 466200.0 1193400.0 ;
      RECT  456000.0 1207200.0 466200.0 1193400.0 ;
      RECT  456000.0 1207200.0 466200.0 1221000.0 ;
      RECT  456000.0 1234800.0 466200.0 1221000.0 ;
      RECT  456000.0 1234800.0 466200.0 1248600.0 ;
      RECT  456000.0 1262400.0 466200.0 1248600.0 ;
      RECT  456000.0 1262400.0 466200.0 1276200.0 ;
      RECT  456000.0 1290000.0 466200.0 1276200.0 ;
      RECT  456000.0 1290000.0 466200.0 1303800.0 ;
      RECT  456000.0 1317600.0 466200.0 1303800.0 ;
      RECT  456000.0 1317600.0 466200.0 1331400.0 ;
      RECT  456000.0 1345200.0 466200.0 1331400.0 ;
      RECT  456000.0 1345200.0 466200.0 1359000.0 ;
      RECT  456000.0 1372800.0 466200.0 1359000.0 ;
      RECT  456000.0 1372800.0 466200.0 1386600.0 ;
      RECT  456000.0 1400400.0 466200.0 1386600.0 ;
      RECT  456000.0 1400400.0 466200.0 1414200.0 ;
      RECT  456000.0 1428000.0 466200.0 1414200.0 ;
      RECT  456000.0 1428000.0 466200.0 1441800.0 ;
      RECT  456000.0 1455600.0 466200.0 1441800.0 ;
      RECT  456000.0 1455600.0 466200.0 1469400.0 ;
      RECT  456000.0 1483200.0 466200.0 1469400.0 ;
      RECT  456000.0 1483200.0 466200.0 1497000.0 ;
      RECT  456000.0 1510800.0 466200.0 1497000.0 ;
      RECT  456000.0 1510800.0 466200.0 1524600.0 ;
      RECT  456000.0 1538400.0 466200.0 1524600.0 ;
      RECT  456000.0 1538400.0 466200.0 1552200.0 ;
      RECT  456000.0 1566000.0 466200.0 1552200.0 ;
      RECT  456000.0 1566000.0 466200.0 1579800.0 ;
      RECT  456000.0 1593600.0 466200.0 1579800.0 ;
      RECT  456000.0 1593600.0 466200.0 1607400.0 ;
      RECT  456000.0 1621200.0 466200.0 1607400.0 ;
      RECT  456000.0 1621200.0 466200.0 1635000.0 ;
      RECT  456000.0 1648800.0 466200.0 1635000.0 ;
      RECT  456000.0 1648800.0 466200.0 1662600.0 ;
      RECT  456000.0 1676400.0 466200.0 1662600.0 ;
      RECT  456000.0 1676400.0 466200.0 1690200.0 ;
      RECT  456000.0 1704000.0 466200.0 1690200.0 ;
      RECT  456000.0 1704000.0 466200.0 1717800.0 ;
      RECT  456000.0 1731600.0 466200.0 1717800.0 ;
      RECT  456000.0 1731600.0 466200.0 1745400.0 ;
      RECT  456000.0 1759200.0 466200.0 1745400.0 ;
      RECT  456000.0 1759200.0 466200.0 1773000.0 ;
      RECT  456000.0 1786800.0 466200.0 1773000.0 ;
      RECT  456000.0 1786800.0 466200.0 1800600.0 ;
      RECT  456000.0 1814400.0 466200.0 1800600.0 ;
      RECT  456000.0 1814400.0 466200.0 1828200.0 ;
      RECT  456000.0 1842000.0 466200.0 1828200.0 ;
      RECT  456000.0 1842000.0 466200.0 1855800.0 ;
      RECT  456000.0 1869600.0 466200.0 1855800.0 ;
      RECT  456000.0 1869600.0 466200.0 1883400.0 ;
      RECT  456000.0 1897200.0 466200.0 1883400.0 ;
      RECT  456000.0 1897200.0 466200.0 1911000.0 ;
      RECT  456000.0 1924800.0 466200.0 1911000.0 ;
      RECT  456000.0 1924800.0 466200.0 1938600.0 ;
      RECT  456000.0 1952400.0 466200.0 1938600.0 ;
      RECT  456000.0 1952400.0 466200.0 1966200.0 ;
      RECT  456000.0 1980000.0 466200.0 1966200.0 ;
      RECT  456000.0 1980000.0 466200.0 1993800.0 ;
      RECT  456000.0 2007600.0 466200.0 1993800.0 ;
      RECT  456000.0 2007600.0 466200.0 2021400.0 ;
      RECT  456000.0 2035200.0 466200.0 2021400.0 ;
      RECT  456000.0 2035200.0 466200.0 2049000.0 ;
      RECT  456000.0 2062800.0 466200.0 2049000.0 ;
      RECT  456000.0 2062800.0 466200.0 2076600.0 ;
      RECT  456000.0 2090400.0 466200.0 2076600.0 ;
      RECT  456000.0 2090400.0 466200.0 2104200.0 ;
      RECT  456000.0 2118000.0 466200.0 2104200.0 ;
      RECT  456000.0 2118000.0 466200.0 2131800.0 ;
      RECT  456000.0 2145600.0 466200.0 2131800.0 ;
      RECT  466200.0 379200.0 476400.0 393000.0 ;
      RECT  466200.0 406800.0 476400.0 393000.0 ;
      RECT  466200.0 406800.0 476400.0 420600.0 ;
      RECT  466200.0 434400.0 476400.0 420600.0 ;
      RECT  466200.0 434400.0 476400.0 448200.0 ;
      RECT  466200.0 462000.0 476400.0 448200.0 ;
      RECT  466200.0 462000.0 476400.0 475800.0 ;
      RECT  466200.0 489600.0 476400.0 475800.0 ;
      RECT  466200.0 489600.0 476400.0 503400.0 ;
      RECT  466200.0 517200.0 476400.0 503400.0 ;
      RECT  466200.0 517200.0 476400.0 531000.0 ;
      RECT  466200.0 544800.0 476400.0 531000.0 ;
      RECT  466200.0 544800.0 476400.0 558600.0 ;
      RECT  466200.0 572400.0 476400.0 558600.0 ;
      RECT  466200.0 572400.0 476400.0 586200.0 ;
      RECT  466200.0 600000.0 476400.0 586200.0 ;
      RECT  466200.0 600000.0 476400.0 613800.0 ;
      RECT  466200.0 627600.0 476400.0 613800.0 ;
      RECT  466200.0 627600.0 476400.0 641400.0 ;
      RECT  466200.0 655200.0 476400.0 641400.0 ;
      RECT  466200.0 655200.0 476400.0 669000.0 ;
      RECT  466200.0 682800.0 476400.0 669000.0 ;
      RECT  466200.0 682800.0 476400.0 696600.0 ;
      RECT  466200.0 710400.0 476400.0 696600.0 ;
      RECT  466200.0 710400.0 476400.0 724200.0 ;
      RECT  466200.0 738000.0 476400.0 724200.0 ;
      RECT  466200.0 738000.0 476400.0 751800.0 ;
      RECT  466200.0 765600.0 476400.0 751800.0 ;
      RECT  466200.0 765600.0 476400.0 779400.0 ;
      RECT  466200.0 793200.0 476400.0 779400.0 ;
      RECT  466200.0 793200.0 476400.0 807000.0 ;
      RECT  466200.0 820800.0 476400.0 807000.0 ;
      RECT  466200.0 820800.0 476400.0 834600.0 ;
      RECT  466200.0 848400.0 476400.0 834600.0 ;
      RECT  466200.0 848400.0 476400.0 862200.0 ;
      RECT  466200.0 876000.0 476400.0 862200.0 ;
      RECT  466200.0 876000.0 476400.0 889800.0 ;
      RECT  466200.0 903600.0 476400.0 889800.0 ;
      RECT  466200.0 903600.0 476400.0 917400.0 ;
      RECT  466200.0 931200.0 476400.0 917400.0 ;
      RECT  466200.0 931200.0 476400.0 945000.0 ;
      RECT  466200.0 958800.0 476400.0 945000.0 ;
      RECT  466200.0 958800.0 476400.0 972600.0 ;
      RECT  466200.0 986400.0 476400.0 972600.0 ;
      RECT  466200.0 986400.0 476400.0 1000200.0 ;
      RECT  466200.0 1014000.0 476400.0 1000200.0 ;
      RECT  466200.0 1014000.0 476400.0 1027800.0 ;
      RECT  466200.0 1041600.0 476400.0 1027800.0 ;
      RECT  466200.0 1041600.0 476400.0 1055400.0 ;
      RECT  466200.0 1069200.0 476400.0 1055400.0 ;
      RECT  466200.0 1069200.0 476400.0 1083000.0 ;
      RECT  466200.0 1096800.0 476400.0 1083000.0 ;
      RECT  466200.0 1096800.0 476400.0 1110600.0 ;
      RECT  466200.0 1124400.0 476400.0 1110600.0 ;
      RECT  466200.0 1124400.0 476400.0 1138200.0 ;
      RECT  466200.0 1152000.0 476400.0 1138200.0 ;
      RECT  466200.0 1152000.0 476400.0 1165800.0 ;
      RECT  466200.0 1179600.0 476400.0 1165800.0 ;
      RECT  466200.0 1179600.0 476400.0 1193400.0 ;
      RECT  466200.0 1207200.0 476400.0 1193400.0 ;
      RECT  466200.0 1207200.0 476400.0 1221000.0 ;
      RECT  466200.0 1234800.0 476400.0 1221000.0 ;
      RECT  466200.0 1234800.0 476400.0 1248600.0 ;
      RECT  466200.0 1262400.0 476400.0 1248600.0 ;
      RECT  466200.0 1262400.0 476400.0 1276200.0 ;
      RECT  466200.0 1290000.0 476400.0 1276200.0 ;
      RECT  466200.0 1290000.0 476400.0 1303800.0 ;
      RECT  466200.0 1317600.0 476400.0 1303800.0 ;
      RECT  466200.0 1317600.0 476400.0 1331400.0 ;
      RECT  466200.0 1345200.0 476400.0 1331400.0 ;
      RECT  466200.0 1345200.0 476400.0 1359000.0 ;
      RECT  466200.0 1372800.0 476400.0 1359000.0 ;
      RECT  466200.0 1372800.0 476400.0 1386600.0 ;
      RECT  466200.0 1400400.0 476400.0 1386600.0 ;
      RECT  466200.0 1400400.0 476400.0 1414200.0 ;
      RECT  466200.0 1428000.0 476400.0 1414200.0 ;
      RECT  466200.0 1428000.0 476400.0 1441800.0 ;
      RECT  466200.0 1455600.0 476400.0 1441800.0 ;
      RECT  466200.0 1455600.0 476400.0 1469400.0 ;
      RECT  466200.0 1483200.0 476400.0 1469400.0 ;
      RECT  466200.0 1483200.0 476400.0 1497000.0 ;
      RECT  466200.0 1510800.0 476400.0 1497000.0 ;
      RECT  466200.0 1510800.0 476400.0 1524600.0 ;
      RECT  466200.0 1538400.0 476400.0 1524600.0 ;
      RECT  466200.0 1538400.0 476400.0 1552200.0 ;
      RECT  466200.0 1566000.0 476400.0 1552200.0 ;
      RECT  466200.0 1566000.0 476400.0 1579800.0 ;
      RECT  466200.0 1593600.0 476400.0 1579800.0 ;
      RECT  466200.0 1593600.0 476400.0 1607400.0 ;
      RECT  466200.0 1621200.0 476400.0 1607400.0 ;
      RECT  466200.0 1621200.0 476400.0 1635000.0 ;
      RECT  466200.0 1648800.0 476400.0 1635000.0 ;
      RECT  466200.0 1648800.0 476400.0 1662600.0 ;
      RECT  466200.0 1676400.0 476400.0 1662600.0 ;
      RECT  466200.0 1676400.0 476400.0 1690200.0 ;
      RECT  466200.0 1704000.0 476400.0 1690200.0 ;
      RECT  466200.0 1704000.0 476400.0 1717800.0 ;
      RECT  466200.0 1731600.0 476400.0 1717800.0 ;
      RECT  466200.0 1731600.0 476400.0 1745400.0 ;
      RECT  466200.0 1759200.0 476400.0 1745400.0 ;
      RECT  466200.0 1759200.0 476400.0 1773000.0 ;
      RECT  466200.0 1786800.0 476400.0 1773000.0 ;
      RECT  466200.0 1786800.0 476400.0 1800600.0 ;
      RECT  466200.0 1814400.0 476400.0 1800600.0 ;
      RECT  466200.0 1814400.0 476400.0 1828200.0 ;
      RECT  466200.0 1842000.0 476400.0 1828200.0 ;
      RECT  466200.0 1842000.0 476400.0 1855800.0 ;
      RECT  466200.0 1869600.0 476400.0 1855800.0 ;
      RECT  466200.0 1869600.0 476400.0 1883400.0 ;
      RECT  466200.0 1897200.0 476400.0 1883400.0 ;
      RECT  466200.0 1897200.0 476400.0 1911000.0 ;
      RECT  466200.0 1924800.0 476400.0 1911000.0 ;
      RECT  466200.0 1924800.0 476400.0 1938600.0 ;
      RECT  466200.0 1952400.0 476400.0 1938600.0 ;
      RECT  466200.0 1952400.0 476400.0 1966200.0 ;
      RECT  466200.0 1980000.0 476400.0 1966200.0 ;
      RECT  466200.0 1980000.0 476400.0 1993800.0 ;
      RECT  466200.0 2007600.0 476400.0 1993800.0 ;
      RECT  466200.0 2007600.0 476400.0 2021400.0 ;
      RECT  466200.0 2035200.0 476400.0 2021400.0 ;
      RECT  466200.0 2035200.0 476400.0 2049000.0 ;
      RECT  466200.0 2062800.0 476400.0 2049000.0 ;
      RECT  466200.0 2062800.0 476400.0 2076600.0 ;
      RECT  466200.0 2090400.0 476400.0 2076600.0 ;
      RECT  466200.0 2090400.0 476400.0 2104200.0 ;
      RECT  466200.0 2118000.0 476400.0 2104200.0 ;
      RECT  466200.0 2118000.0 476400.0 2131800.0 ;
      RECT  466200.0 2145600.0 476400.0 2131800.0 ;
      RECT  476400.0 379200.0 486600.0 393000.0 ;
      RECT  476400.0 406800.0 486600.0 393000.0 ;
      RECT  476400.0 406800.0 486600.0 420600.0 ;
      RECT  476400.0 434400.0 486600.0 420600.0 ;
      RECT  476400.0 434400.0 486600.0 448200.0 ;
      RECT  476400.0 462000.0 486600.0 448200.0 ;
      RECT  476400.0 462000.0 486600.0 475800.0 ;
      RECT  476400.0 489600.0 486600.0 475800.0 ;
      RECT  476400.0 489600.0 486600.0 503400.0 ;
      RECT  476400.0 517200.0 486600.0 503400.0 ;
      RECT  476400.0 517200.0 486600.0 531000.0 ;
      RECT  476400.0 544800.0 486600.0 531000.0 ;
      RECT  476400.0 544800.0 486600.0 558600.0 ;
      RECT  476400.0 572400.0 486600.0 558600.0 ;
      RECT  476400.0 572400.0 486600.0 586200.0 ;
      RECT  476400.0 600000.0 486600.0 586200.0 ;
      RECT  476400.0 600000.0 486600.0 613800.0 ;
      RECT  476400.0 627600.0 486600.0 613800.0 ;
      RECT  476400.0 627600.0 486600.0 641400.0 ;
      RECT  476400.0 655200.0 486600.0 641400.0 ;
      RECT  476400.0 655200.0 486600.0 669000.0 ;
      RECT  476400.0 682800.0 486600.0 669000.0 ;
      RECT  476400.0 682800.0 486600.0 696600.0 ;
      RECT  476400.0 710400.0 486600.0 696600.0 ;
      RECT  476400.0 710400.0 486600.0 724200.0 ;
      RECT  476400.0 738000.0 486600.0 724200.0 ;
      RECT  476400.0 738000.0 486600.0 751800.0 ;
      RECT  476400.0 765600.0 486600.0 751800.0 ;
      RECT  476400.0 765600.0 486600.0 779400.0 ;
      RECT  476400.0 793200.0 486600.0 779400.0 ;
      RECT  476400.0 793200.0 486600.0 807000.0 ;
      RECT  476400.0 820800.0 486600.0 807000.0 ;
      RECT  476400.0 820800.0 486600.0 834600.0 ;
      RECT  476400.0 848400.0 486600.0 834600.0 ;
      RECT  476400.0 848400.0 486600.0 862200.0 ;
      RECT  476400.0 876000.0 486600.0 862200.0 ;
      RECT  476400.0 876000.0 486600.0 889800.0 ;
      RECT  476400.0 903600.0 486600.0 889800.0 ;
      RECT  476400.0 903600.0 486600.0 917400.0 ;
      RECT  476400.0 931200.0 486600.0 917400.0 ;
      RECT  476400.0 931200.0 486600.0 945000.0 ;
      RECT  476400.0 958800.0 486600.0 945000.0 ;
      RECT  476400.0 958800.0 486600.0 972600.0 ;
      RECT  476400.0 986400.0 486600.0 972600.0 ;
      RECT  476400.0 986400.0 486600.0 1000200.0 ;
      RECT  476400.0 1014000.0 486600.0 1000200.0 ;
      RECT  476400.0 1014000.0 486600.0 1027800.0 ;
      RECT  476400.0 1041600.0 486600.0 1027800.0 ;
      RECT  476400.0 1041600.0 486600.0 1055400.0 ;
      RECT  476400.0 1069200.0 486600.0 1055400.0 ;
      RECT  476400.0 1069200.0 486600.0 1083000.0 ;
      RECT  476400.0 1096800.0 486600.0 1083000.0 ;
      RECT  476400.0 1096800.0 486600.0 1110600.0 ;
      RECT  476400.0 1124400.0 486600.0 1110600.0 ;
      RECT  476400.0 1124400.0 486600.0 1138200.0 ;
      RECT  476400.0 1152000.0 486600.0 1138200.0 ;
      RECT  476400.0 1152000.0 486600.0 1165800.0 ;
      RECT  476400.0 1179600.0 486600.0 1165800.0 ;
      RECT  476400.0 1179600.0 486600.0 1193400.0 ;
      RECT  476400.0 1207200.0 486600.0 1193400.0 ;
      RECT  476400.0 1207200.0 486600.0 1221000.0 ;
      RECT  476400.0 1234800.0 486600.0 1221000.0 ;
      RECT  476400.0 1234800.0 486600.0 1248600.0 ;
      RECT  476400.0 1262400.0 486600.0 1248600.0 ;
      RECT  476400.0 1262400.0 486600.0 1276200.0 ;
      RECT  476400.0 1290000.0 486600.0 1276200.0 ;
      RECT  476400.0 1290000.0 486600.0 1303800.0 ;
      RECT  476400.0 1317600.0 486600.0 1303800.0 ;
      RECT  476400.0 1317600.0 486600.0 1331400.0 ;
      RECT  476400.0 1345200.0 486600.0 1331400.0 ;
      RECT  476400.0 1345200.0 486600.0 1359000.0 ;
      RECT  476400.0 1372800.0 486600.0 1359000.0 ;
      RECT  476400.0 1372800.0 486600.0 1386600.0 ;
      RECT  476400.0 1400400.0 486600.0 1386600.0 ;
      RECT  476400.0 1400400.0 486600.0 1414200.0 ;
      RECT  476400.0 1428000.0 486600.0 1414200.0 ;
      RECT  476400.0 1428000.0 486600.0 1441800.0 ;
      RECT  476400.0 1455600.0 486600.0 1441800.0 ;
      RECT  476400.0 1455600.0 486600.0 1469400.0 ;
      RECT  476400.0 1483200.0 486600.0 1469400.0 ;
      RECT  476400.0 1483200.0 486600.0 1497000.0 ;
      RECT  476400.0 1510800.0 486600.0 1497000.0 ;
      RECT  476400.0 1510800.0 486600.0 1524600.0 ;
      RECT  476400.0 1538400.0 486600.0 1524600.0 ;
      RECT  476400.0 1538400.0 486600.0 1552200.0 ;
      RECT  476400.0 1566000.0 486600.0 1552200.0 ;
      RECT  476400.0 1566000.0 486600.0 1579800.0 ;
      RECT  476400.0 1593600.0 486600.0 1579800.0 ;
      RECT  476400.0 1593600.0 486600.0 1607400.0 ;
      RECT  476400.0 1621200.0 486600.0 1607400.0 ;
      RECT  476400.0 1621200.0 486600.0 1635000.0 ;
      RECT  476400.0 1648800.0 486600.0 1635000.0 ;
      RECT  476400.0 1648800.0 486600.0 1662600.0 ;
      RECT  476400.0 1676400.0 486600.0 1662600.0 ;
      RECT  476400.0 1676400.0 486600.0 1690200.0 ;
      RECT  476400.0 1704000.0 486600.0 1690200.0 ;
      RECT  476400.0 1704000.0 486600.0 1717800.0 ;
      RECT  476400.0 1731600.0 486600.0 1717800.0 ;
      RECT  476400.0 1731600.0 486600.0 1745400.0 ;
      RECT  476400.0 1759200.0 486600.0 1745400.0 ;
      RECT  476400.0 1759200.0 486600.0 1773000.0 ;
      RECT  476400.0 1786800.0 486600.0 1773000.0 ;
      RECT  476400.0 1786800.0 486600.0 1800600.0 ;
      RECT  476400.0 1814400.0 486600.0 1800600.0 ;
      RECT  476400.0 1814400.0 486600.0 1828200.0 ;
      RECT  476400.0 1842000.0 486600.0 1828200.0 ;
      RECT  476400.0 1842000.0 486600.0 1855800.0 ;
      RECT  476400.0 1869600.0 486600.0 1855800.0 ;
      RECT  476400.0 1869600.0 486600.0 1883400.0 ;
      RECT  476400.0 1897200.0 486600.0 1883400.0 ;
      RECT  476400.0 1897200.0 486600.0 1911000.0 ;
      RECT  476400.0 1924800.0 486600.0 1911000.0 ;
      RECT  476400.0 1924800.0 486600.0 1938600.0 ;
      RECT  476400.0 1952400.0 486600.0 1938600.0 ;
      RECT  476400.0 1952400.0 486600.0 1966200.0 ;
      RECT  476400.0 1980000.0 486600.0 1966200.0 ;
      RECT  476400.0 1980000.0 486600.0 1993800.0 ;
      RECT  476400.0 2007600.0 486600.0 1993800.0 ;
      RECT  476400.0 2007600.0 486600.0 2021400.0 ;
      RECT  476400.0 2035200.0 486600.0 2021400.0 ;
      RECT  476400.0 2035200.0 486600.0 2049000.0 ;
      RECT  476400.0 2062800.0 486600.0 2049000.0 ;
      RECT  476400.0 2062800.0 486600.0 2076600.0 ;
      RECT  476400.0 2090400.0 486600.0 2076600.0 ;
      RECT  476400.0 2090400.0 486600.0 2104200.0 ;
      RECT  476400.0 2118000.0 486600.0 2104200.0 ;
      RECT  476400.0 2118000.0 486600.0 2131800.0 ;
      RECT  476400.0 2145600.0 486600.0 2131800.0 ;
      RECT  486600.0 379200.0 496800.0 393000.0 ;
      RECT  486600.0 406800.0 496800.0 393000.0 ;
      RECT  486600.0 406800.0 496800.0 420600.0 ;
      RECT  486600.0 434400.0 496800.0 420600.0 ;
      RECT  486600.0 434400.0 496800.0 448200.0 ;
      RECT  486600.0 462000.0 496800.0 448200.0 ;
      RECT  486600.0 462000.0 496800.0 475800.0 ;
      RECT  486600.0 489600.0 496800.0 475800.0 ;
      RECT  486600.0 489600.0 496800.0 503400.0 ;
      RECT  486600.0 517200.0 496800.0 503400.0 ;
      RECT  486600.0 517200.0 496800.0 531000.0 ;
      RECT  486600.0 544800.0 496800.0 531000.0 ;
      RECT  486600.0 544800.0 496800.0 558600.0 ;
      RECT  486600.0 572400.0 496800.0 558600.0 ;
      RECT  486600.0 572400.0 496800.0 586200.0 ;
      RECT  486600.0 600000.0 496800.0 586200.0 ;
      RECT  486600.0 600000.0 496800.0 613800.0 ;
      RECT  486600.0 627600.0 496800.0 613800.0 ;
      RECT  486600.0 627600.0 496800.0 641400.0 ;
      RECT  486600.0 655200.0 496800.0 641400.0 ;
      RECT  486600.0 655200.0 496800.0 669000.0 ;
      RECT  486600.0 682800.0 496800.0 669000.0 ;
      RECT  486600.0 682800.0 496800.0 696600.0 ;
      RECT  486600.0 710400.0 496800.0 696600.0 ;
      RECT  486600.0 710400.0 496800.0 724200.0 ;
      RECT  486600.0 738000.0 496800.0 724200.0 ;
      RECT  486600.0 738000.0 496800.0 751800.0 ;
      RECT  486600.0 765600.0 496800.0 751800.0 ;
      RECT  486600.0 765600.0 496800.0 779400.0 ;
      RECT  486600.0 793200.0 496800.0 779400.0 ;
      RECT  486600.0 793200.0 496800.0 807000.0 ;
      RECT  486600.0 820800.0 496800.0 807000.0 ;
      RECT  486600.0 820800.0 496800.0 834600.0 ;
      RECT  486600.0 848400.0 496800.0 834600.0 ;
      RECT  486600.0 848400.0 496800.0 862200.0 ;
      RECT  486600.0 876000.0 496800.0 862200.0 ;
      RECT  486600.0 876000.0 496800.0 889800.0 ;
      RECT  486600.0 903600.0 496800.0 889800.0 ;
      RECT  486600.0 903600.0 496800.0 917400.0 ;
      RECT  486600.0 931200.0 496800.0 917400.0 ;
      RECT  486600.0 931200.0 496800.0 945000.0 ;
      RECT  486600.0 958800.0 496800.0 945000.0 ;
      RECT  486600.0 958800.0 496800.0 972600.0 ;
      RECT  486600.0 986400.0 496800.0 972600.0 ;
      RECT  486600.0 986400.0 496800.0 1000200.0 ;
      RECT  486600.0 1014000.0 496800.0 1000200.0 ;
      RECT  486600.0 1014000.0 496800.0 1027800.0 ;
      RECT  486600.0 1041600.0 496800.0 1027800.0 ;
      RECT  486600.0 1041600.0 496800.0 1055400.0 ;
      RECT  486600.0 1069200.0 496800.0 1055400.0 ;
      RECT  486600.0 1069200.0 496800.0 1083000.0 ;
      RECT  486600.0 1096800.0 496800.0 1083000.0 ;
      RECT  486600.0 1096800.0 496800.0 1110600.0 ;
      RECT  486600.0 1124400.0 496800.0 1110600.0 ;
      RECT  486600.0 1124400.0 496800.0 1138200.0 ;
      RECT  486600.0 1152000.0 496800.0 1138200.0 ;
      RECT  486600.0 1152000.0 496800.0 1165800.0 ;
      RECT  486600.0 1179600.0 496800.0 1165800.0 ;
      RECT  486600.0 1179600.0 496800.0 1193400.0 ;
      RECT  486600.0 1207200.0 496800.0 1193400.0 ;
      RECT  486600.0 1207200.0 496800.0 1221000.0 ;
      RECT  486600.0 1234800.0 496800.0 1221000.0 ;
      RECT  486600.0 1234800.0 496800.0 1248600.0 ;
      RECT  486600.0 1262400.0 496800.0 1248600.0 ;
      RECT  486600.0 1262400.0 496800.0 1276200.0 ;
      RECT  486600.0 1290000.0 496800.0 1276200.0 ;
      RECT  486600.0 1290000.0 496800.0 1303800.0 ;
      RECT  486600.0 1317600.0 496800.0 1303800.0 ;
      RECT  486600.0 1317600.0 496800.0 1331400.0 ;
      RECT  486600.0 1345200.0 496800.0 1331400.0 ;
      RECT  486600.0 1345200.0 496800.0 1359000.0 ;
      RECT  486600.0 1372800.0 496800.0 1359000.0 ;
      RECT  486600.0 1372800.0 496800.0 1386600.0 ;
      RECT  486600.0 1400400.0 496800.0 1386600.0 ;
      RECT  486600.0 1400400.0 496800.0 1414200.0 ;
      RECT  486600.0 1428000.0 496800.0 1414200.0 ;
      RECT  486600.0 1428000.0 496800.0 1441800.0 ;
      RECT  486600.0 1455600.0 496800.0 1441800.0 ;
      RECT  486600.0 1455600.0 496800.0 1469400.0 ;
      RECT  486600.0 1483200.0 496800.0 1469400.0 ;
      RECT  486600.0 1483200.0 496800.0 1497000.0 ;
      RECT  486600.0 1510800.0 496800.0 1497000.0 ;
      RECT  486600.0 1510800.0 496800.0 1524600.0 ;
      RECT  486600.0 1538400.0 496800.0 1524600.0 ;
      RECT  486600.0 1538400.0 496800.0 1552200.0 ;
      RECT  486600.0 1566000.0 496800.0 1552200.0 ;
      RECT  486600.0 1566000.0 496800.0 1579800.0 ;
      RECT  486600.0 1593600.0 496800.0 1579800.0 ;
      RECT  486600.0 1593600.0 496800.0 1607400.0 ;
      RECT  486600.0 1621200.0 496800.0 1607400.0 ;
      RECT  486600.0 1621200.0 496800.0 1635000.0 ;
      RECT  486600.0 1648800.0 496800.0 1635000.0 ;
      RECT  486600.0 1648800.0 496800.0 1662600.0 ;
      RECT  486600.0 1676400.0 496800.0 1662600.0 ;
      RECT  486600.0 1676400.0 496800.0 1690200.0 ;
      RECT  486600.0 1704000.0 496800.0 1690200.0 ;
      RECT  486600.0 1704000.0 496800.0 1717800.0 ;
      RECT  486600.0 1731600.0 496800.0 1717800.0 ;
      RECT  486600.0 1731600.0 496800.0 1745400.0 ;
      RECT  486600.0 1759200.0 496800.0 1745400.0 ;
      RECT  486600.0 1759200.0 496800.0 1773000.0 ;
      RECT  486600.0 1786800.0 496800.0 1773000.0 ;
      RECT  486600.0 1786800.0 496800.0 1800600.0 ;
      RECT  486600.0 1814400.0 496800.0 1800600.0 ;
      RECT  486600.0 1814400.0 496800.0 1828200.0 ;
      RECT  486600.0 1842000.0 496800.0 1828200.0 ;
      RECT  486600.0 1842000.0 496800.0 1855800.0 ;
      RECT  486600.0 1869600.0 496800.0 1855800.0 ;
      RECT  486600.0 1869600.0 496800.0 1883400.0 ;
      RECT  486600.0 1897200.0 496800.0 1883400.0 ;
      RECT  486600.0 1897200.0 496800.0 1911000.0 ;
      RECT  486600.0 1924800.0 496800.0 1911000.0 ;
      RECT  486600.0 1924800.0 496800.0 1938600.0 ;
      RECT  486600.0 1952400.0 496800.0 1938600.0 ;
      RECT  486600.0 1952400.0 496800.0 1966200.0 ;
      RECT  486600.0 1980000.0 496800.0 1966200.0 ;
      RECT  486600.0 1980000.0 496800.0 1993800.0 ;
      RECT  486600.0 2007600.0 496800.0 1993800.0 ;
      RECT  486600.0 2007600.0 496800.0 2021400.0 ;
      RECT  486600.0 2035200.0 496800.0 2021400.0 ;
      RECT  486600.0 2035200.0 496800.0 2049000.0 ;
      RECT  486600.0 2062800.0 496800.0 2049000.0 ;
      RECT  486600.0 2062800.0 496800.0 2076600.0 ;
      RECT  486600.0 2090400.0 496800.0 2076600.0 ;
      RECT  486600.0 2090400.0 496800.0 2104200.0 ;
      RECT  486600.0 2118000.0 496800.0 2104200.0 ;
      RECT  486600.0 2118000.0 496800.0 2131800.0 ;
      RECT  486600.0 2145600.0 496800.0 2131800.0 ;
      RECT  496800.0 379200.0 507000.0 393000.0 ;
      RECT  496800.0 406800.0 507000.0 393000.0 ;
      RECT  496800.0 406800.0 507000.0 420600.0 ;
      RECT  496800.0 434400.0 507000.0 420600.0 ;
      RECT  496800.0 434400.0 507000.0 448200.0 ;
      RECT  496800.0 462000.0 507000.0 448200.0 ;
      RECT  496800.0 462000.0 507000.0 475800.0 ;
      RECT  496800.0 489600.0 507000.0 475800.0 ;
      RECT  496800.0 489600.0 507000.0 503400.0 ;
      RECT  496800.0 517200.0 507000.0 503400.0 ;
      RECT  496800.0 517200.0 507000.0 531000.0 ;
      RECT  496800.0 544800.0 507000.0 531000.0 ;
      RECT  496800.0 544800.0 507000.0 558600.0 ;
      RECT  496800.0 572400.0 507000.0 558600.0 ;
      RECT  496800.0 572400.0 507000.0 586200.0 ;
      RECT  496800.0 600000.0 507000.0 586200.0 ;
      RECT  496800.0 600000.0 507000.0 613800.0 ;
      RECT  496800.0 627600.0 507000.0 613800.0 ;
      RECT  496800.0 627600.0 507000.0 641400.0 ;
      RECT  496800.0 655200.0 507000.0 641400.0 ;
      RECT  496800.0 655200.0 507000.0 669000.0 ;
      RECT  496800.0 682800.0 507000.0 669000.0 ;
      RECT  496800.0 682800.0 507000.0 696600.0 ;
      RECT  496800.0 710400.0 507000.0 696600.0 ;
      RECT  496800.0 710400.0 507000.0 724200.0 ;
      RECT  496800.0 738000.0 507000.0 724200.0 ;
      RECT  496800.0 738000.0 507000.0 751800.0 ;
      RECT  496800.0 765600.0 507000.0 751800.0 ;
      RECT  496800.0 765600.0 507000.0 779400.0 ;
      RECT  496800.0 793200.0 507000.0 779400.0 ;
      RECT  496800.0 793200.0 507000.0 807000.0 ;
      RECT  496800.0 820800.0 507000.0 807000.0 ;
      RECT  496800.0 820800.0 507000.0 834600.0 ;
      RECT  496800.0 848400.0 507000.0 834600.0 ;
      RECT  496800.0 848400.0 507000.0 862200.0 ;
      RECT  496800.0 876000.0 507000.0 862200.0 ;
      RECT  496800.0 876000.0 507000.0 889800.0 ;
      RECT  496800.0 903600.0 507000.0 889800.0 ;
      RECT  496800.0 903600.0 507000.0 917400.0 ;
      RECT  496800.0 931200.0 507000.0 917400.0 ;
      RECT  496800.0 931200.0 507000.0 945000.0 ;
      RECT  496800.0 958800.0 507000.0 945000.0 ;
      RECT  496800.0 958800.0 507000.0 972600.0 ;
      RECT  496800.0 986400.0 507000.0 972600.0 ;
      RECT  496800.0 986400.0 507000.0 1000200.0 ;
      RECT  496800.0 1014000.0 507000.0 1000200.0 ;
      RECT  496800.0 1014000.0 507000.0 1027800.0 ;
      RECT  496800.0 1041600.0 507000.0 1027800.0 ;
      RECT  496800.0 1041600.0 507000.0 1055400.0 ;
      RECT  496800.0 1069200.0 507000.0 1055400.0 ;
      RECT  496800.0 1069200.0 507000.0 1083000.0 ;
      RECT  496800.0 1096800.0 507000.0 1083000.0 ;
      RECT  496800.0 1096800.0 507000.0 1110600.0 ;
      RECT  496800.0 1124400.0 507000.0 1110600.0 ;
      RECT  496800.0 1124400.0 507000.0 1138200.0 ;
      RECT  496800.0 1152000.0 507000.0 1138200.0 ;
      RECT  496800.0 1152000.0 507000.0 1165800.0 ;
      RECT  496800.0 1179600.0 507000.0 1165800.0 ;
      RECT  496800.0 1179600.0 507000.0 1193400.0 ;
      RECT  496800.0 1207200.0 507000.0 1193400.0 ;
      RECT  496800.0 1207200.0 507000.0 1221000.0 ;
      RECT  496800.0 1234800.0 507000.0 1221000.0 ;
      RECT  496800.0 1234800.0 507000.0 1248600.0 ;
      RECT  496800.0 1262400.0 507000.0 1248600.0 ;
      RECT  496800.0 1262400.0 507000.0 1276200.0 ;
      RECT  496800.0 1290000.0 507000.0 1276200.0 ;
      RECT  496800.0 1290000.0 507000.0 1303800.0 ;
      RECT  496800.0 1317600.0 507000.0 1303800.0 ;
      RECT  496800.0 1317600.0 507000.0 1331400.0 ;
      RECT  496800.0 1345200.0 507000.0 1331400.0 ;
      RECT  496800.0 1345200.0 507000.0 1359000.0 ;
      RECT  496800.0 1372800.0 507000.0 1359000.0 ;
      RECT  496800.0 1372800.0 507000.0 1386600.0 ;
      RECT  496800.0 1400400.0 507000.0 1386600.0 ;
      RECT  496800.0 1400400.0 507000.0 1414200.0 ;
      RECT  496800.0 1428000.0 507000.0 1414200.0 ;
      RECT  496800.0 1428000.0 507000.0 1441800.0 ;
      RECT  496800.0 1455600.0 507000.0 1441800.0 ;
      RECT  496800.0 1455600.0 507000.0 1469400.0 ;
      RECT  496800.0 1483200.0 507000.0 1469400.0 ;
      RECT  496800.0 1483200.0 507000.0 1497000.0 ;
      RECT  496800.0 1510800.0 507000.0 1497000.0 ;
      RECT  496800.0 1510800.0 507000.0 1524600.0 ;
      RECT  496800.0 1538400.0 507000.0 1524600.0 ;
      RECT  496800.0 1538400.0 507000.0 1552200.0 ;
      RECT  496800.0 1566000.0 507000.0 1552200.0 ;
      RECT  496800.0 1566000.0 507000.0 1579800.0 ;
      RECT  496800.0 1593600.0 507000.0 1579800.0 ;
      RECT  496800.0 1593600.0 507000.0 1607400.0 ;
      RECT  496800.0 1621200.0 507000.0 1607400.0 ;
      RECT  496800.0 1621200.0 507000.0 1635000.0 ;
      RECT  496800.0 1648800.0 507000.0 1635000.0 ;
      RECT  496800.0 1648800.0 507000.0 1662600.0 ;
      RECT  496800.0 1676400.0 507000.0 1662600.0 ;
      RECT  496800.0 1676400.0 507000.0 1690200.0 ;
      RECT  496800.0 1704000.0 507000.0 1690200.0 ;
      RECT  496800.0 1704000.0 507000.0 1717800.0 ;
      RECT  496800.0 1731600.0 507000.0 1717800.0 ;
      RECT  496800.0 1731600.0 507000.0 1745400.0 ;
      RECT  496800.0 1759200.0 507000.0 1745400.0 ;
      RECT  496800.0 1759200.0 507000.0 1773000.0 ;
      RECT  496800.0 1786800.0 507000.0 1773000.0 ;
      RECT  496800.0 1786800.0 507000.0 1800600.0 ;
      RECT  496800.0 1814400.0 507000.0 1800600.0 ;
      RECT  496800.0 1814400.0 507000.0 1828200.0 ;
      RECT  496800.0 1842000.0 507000.0 1828200.0 ;
      RECT  496800.0 1842000.0 507000.0 1855800.0 ;
      RECT  496800.0 1869600.0 507000.0 1855800.0 ;
      RECT  496800.0 1869600.0 507000.0 1883400.0 ;
      RECT  496800.0 1897200.0 507000.0 1883400.0 ;
      RECT  496800.0 1897200.0 507000.0 1911000.0 ;
      RECT  496800.0 1924800.0 507000.0 1911000.0 ;
      RECT  496800.0 1924800.0 507000.0 1938600.0 ;
      RECT  496800.0 1952400.0 507000.0 1938600.0 ;
      RECT  496800.0 1952400.0 507000.0 1966200.0 ;
      RECT  496800.0 1980000.0 507000.0 1966200.0 ;
      RECT  496800.0 1980000.0 507000.0 1993800.0 ;
      RECT  496800.0 2007600.0 507000.0 1993800.0 ;
      RECT  496800.0 2007600.0 507000.0 2021400.0 ;
      RECT  496800.0 2035200.0 507000.0 2021400.0 ;
      RECT  496800.0 2035200.0 507000.0 2049000.0 ;
      RECT  496800.0 2062800.0 507000.0 2049000.0 ;
      RECT  496800.0 2062800.0 507000.0 2076600.0 ;
      RECT  496800.0 2090400.0 507000.0 2076600.0 ;
      RECT  496800.0 2090400.0 507000.0 2104200.0 ;
      RECT  496800.0 2118000.0 507000.0 2104200.0 ;
      RECT  496800.0 2118000.0 507000.0 2131800.0 ;
      RECT  496800.0 2145600.0 507000.0 2131800.0 ;
      RECT  507000.0 379200.0 517200.0 393000.0 ;
      RECT  507000.0 406800.0 517200.0 393000.0 ;
      RECT  507000.0 406800.0 517200.0 420600.0 ;
      RECT  507000.0 434400.0 517200.0 420600.0 ;
      RECT  507000.0 434400.0 517200.0 448200.0 ;
      RECT  507000.0 462000.0 517200.0 448200.0 ;
      RECT  507000.0 462000.0 517200.0 475800.0 ;
      RECT  507000.0 489600.0 517200.0 475800.0 ;
      RECT  507000.0 489600.0 517200.0 503400.0 ;
      RECT  507000.0 517200.0 517200.0 503400.0 ;
      RECT  507000.0 517200.0 517200.0 531000.0 ;
      RECT  507000.0 544800.0 517200.0 531000.0 ;
      RECT  507000.0 544800.0 517200.0 558600.0 ;
      RECT  507000.0 572400.0 517200.0 558600.0 ;
      RECT  507000.0 572400.0 517200.0 586200.0 ;
      RECT  507000.0 600000.0 517200.0 586200.0 ;
      RECT  507000.0 600000.0 517200.0 613800.0 ;
      RECT  507000.0 627600.0 517200.0 613800.0 ;
      RECT  507000.0 627600.0 517200.0 641400.0 ;
      RECT  507000.0 655200.0 517200.0 641400.0 ;
      RECT  507000.0 655200.0 517200.0 669000.0 ;
      RECT  507000.0 682800.0 517200.0 669000.0 ;
      RECT  507000.0 682800.0 517200.0 696600.0 ;
      RECT  507000.0 710400.0 517200.0 696600.0 ;
      RECT  507000.0 710400.0 517200.0 724200.0 ;
      RECT  507000.0 738000.0 517200.0 724200.0 ;
      RECT  507000.0 738000.0 517200.0 751800.0 ;
      RECT  507000.0 765600.0 517200.0 751800.0 ;
      RECT  507000.0 765600.0 517200.0 779400.0 ;
      RECT  507000.0 793200.0 517200.0 779400.0 ;
      RECT  507000.0 793200.0 517200.0 807000.0 ;
      RECT  507000.0 820800.0 517200.0 807000.0 ;
      RECT  507000.0 820800.0 517200.0 834600.0 ;
      RECT  507000.0 848400.0 517200.0 834600.0 ;
      RECT  507000.0 848400.0 517200.0 862200.0 ;
      RECT  507000.0 876000.0 517200.0 862200.0 ;
      RECT  507000.0 876000.0 517200.0 889800.0 ;
      RECT  507000.0 903600.0 517200.0 889800.0 ;
      RECT  507000.0 903600.0 517200.0 917400.0 ;
      RECT  507000.0 931200.0 517200.0 917400.0 ;
      RECT  507000.0 931200.0 517200.0 945000.0 ;
      RECT  507000.0 958800.0 517200.0 945000.0 ;
      RECT  507000.0 958800.0 517200.0 972600.0 ;
      RECT  507000.0 986400.0 517200.0 972600.0 ;
      RECT  507000.0 986400.0 517200.0 1000200.0 ;
      RECT  507000.0 1014000.0 517200.0 1000200.0 ;
      RECT  507000.0 1014000.0 517200.0 1027800.0 ;
      RECT  507000.0 1041600.0 517200.0 1027800.0 ;
      RECT  507000.0 1041600.0 517200.0 1055400.0 ;
      RECT  507000.0 1069200.0 517200.0 1055400.0 ;
      RECT  507000.0 1069200.0 517200.0 1083000.0 ;
      RECT  507000.0 1096800.0 517200.0 1083000.0 ;
      RECT  507000.0 1096800.0 517200.0 1110600.0 ;
      RECT  507000.0 1124400.0 517200.0 1110600.0 ;
      RECT  507000.0 1124400.0 517200.0 1138200.0 ;
      RECT  507000.0 1152000.0 517200.0 1138200.0 ;
      RECT  507000.0 1152000.0 517200.0 1165800.0 ;
      RECT  507000.0 1179600.0 517200.0 1165800.0 ;
      RECT  507000.0 1179600.0 517200.0 1193400.0 ;
      RECT  507000.0 1207200.0 517200.0 1193400.0 ;
      RECT  507000.0 1207200.0 517200.0 1221000.0 ;
      RECT  507000.0 1234800.0 517200.0 1221000.0 ;
      RECT  507000.0 1234800.0 517200.0 1248600.0 ;
      RECT  507000.0 1262400.0 517200.0 1248600.0 ;
      RECT  507000.0 1262400.0 517200.0 1276200.0 ;
      RECT  507000.0 1290000.0 517200.0 1276200.0 ;
      RECT  507000.0 1290000.0 517200.0 1303800.0 ;
      RECT  507000.0 1317600.0 517200.0 1303800.0 ;
      RECT  507000.0 1317600.0 517200.0 1331400.0 ;
      RECT  507000.0 1345200.0 517200.0 1331400.0 ;
      RECT  507000.0 1345200.0 517200.0 1359000.0 ;
      RECT  507000.0 1372800.0 517200.0 1359000.0 ;
      RECT  507000.0 1372800.0 517200.0 1386600.0 ;
      RECT  507000.0 1400400.0 517200.0 1386600.0 ;
      RECT  507000.0 1400400.0 517200.0 1414200.0 ;
      RECT  507000.0 1428000.0 517200.0 1414200.0 ;
      RECT  507000.0 1428000.0 517200.0 1441800.0 ;
      RECT  507000.0 1455600.0 517200.0 1441800.0 ;
      RECT  507000.0 1455600.0 517200.0 1469400.0 ;
      RECT  507000.0 1483200.0 517200.0 1469400.0 ;
      RECT  507000.0 1483200.0 517200.0 1497000.0 ;
      RECT  507000.0 1510800.0 517200.0 1497000.0 ;
      RECT  507000.0 1510800.0 517200.0 1524600.0 ;
      RECT  507000.0 1538400.0 517200.0 1524600.0 ;
      RECT  507000.0 1538400.0 517200.0 1552200.0 ;
      RECT  507000.0 1566000.0 517200.0 1552200.0 ;
      RECT  507000.0 1566000.0 517200.0 1579800.0 ;
      RECT  507000.0 1593600.0 517200.0 1579800.0 ;
      RECT  507000.0 1593600.0 517200.0 1607400.0 ;
      RECT  507000.0 1621200.0 517200.0 1607400.0 ;
      RECT  507000.0 1621200.0 517200.0 1635000.0 ;
      RECT  507000.0 1648800.0 517200.0 1635000.0 ;
      RECT  507000.0 1648800.0 517200.0 1662600.0 ;
      RECT  507000.0 1676400.0 517200.0 1662600.0 ;
      RECT  507000.0 1676400.0 517200.0 1690200.0 ;
      RECT  507000.0 1704000.0 517200.0 1690200.0 ;
      RECT  507000.0 1704000.0 517200.0 1717800.0 ;
      RECT  507000.0 1731600.0 517200.0 1717800.0 ;
      RECT  507000.0 1731600.0 517200.0 1745400.0 ;
      RECT  507000.0 1759200.0 517200.0 1745400.0 ;
      RECT  507000.0 1759200.0 517200.0 1773000.0 ;
      RECT  507000.0 1786800.0 517200.0 1773000.0 ;
      RECT  507000.0 1786800.0 517200.0 1800600.0 ;
      RECT  507000.0 1814400.0 517200.0 1800600.0 ;
      RECT  507000.0 1814400.0 517200.0 1828200.0 ;
      RECT  507000.0 1842000.0 517200.0 1828200.0 ;
      RECT  507000.0 1842000.0 517200.0 1855800.0 ;
      RECT  507000.0 1869600.0 517200.0 1855800.0 ;
      RECT  507000.0 1869600.0 517200.0 1883400.0 ;
      RECT  507000.0 1897200.0 517200.0 1883400.0 ;
      RECT  507000.0 1897200.0 517200.0 1911000.0 ;
      RECT  507000.0 1924800.0 517200.0 1911000.0 ;
      RECT  507000.0 1924800.0 517200.0 1938600.0 ;
      RECT  507000.0 1952400.0 517200.0 1938600.0 ;
      RECT  507000.0 1952400.0 517200.0 1966200.0 ;
      RECT  507000.0 1980000.0 517200.0 1966200.0 ;
      RECT  507000.0 1980000.0 517200.0 1993800.0 ;
      RECT  507000.0 2007600.0 517200.0 1993800.0 ;
      RECT  507000.0 2007600.0 517200.0 2021400.0 ;
      RECT  507000.0 2035200.0 517200.0 2021400.0 ;
      RECT  507000.0 2035200.0 517200.0 2049000.0 ;
      RECT  507000.0 2062800.0 517200.0 2049000.0 ;
      RECT  507000.0 2062800.0 517200.0 2076600.0 ;
      RECT  507000.0 2090400.0 517200.0 2076600.0 ;
      RECT  507000.0 2090400.0 517200.0 2104200.0 ;
      RECT  507000.0 2118000.0 517200.0 2104200.0 ;
      RECT  507000.0 2118000.0 517200.0 2131800.0 ;
      RECT  507000.0 2145600.0 517200.0 2131800.0 ;
      RECT  517200.0 379200.0 527400.0 393000.0 ;
      RECT  517200.0 406800.0 527400.0 393000.0 ;
      RECT  517200.0 406800.0 527400.0 420600.0 ;
      RECT  517200.0 434400.0 527400.0 420600.0 ;
      RECT  517200.0 434400.0 527400.0 448200.0 ;
      RECT  517200.0 462000.0 527400.0 448200.0 ;
      RECT  517200.0 462000.0 527400.0 475800.0 ;
      RECT  517200.0 489600.0 527400.0 475800.0 ;
      RECT  517200.0 489600.0 527400.0 503400.0 ;
      RECT  517200.0 517200.0 527400.0 503400.0 ;
      RECT  517200.0 517200.0 527400.0 531000.0 ;
      RECT  517200.0 544800.0 527400.0 531000.0 ;
      RECT  517200.0 544800.0 527400.0 558600.0 ;
      RECT  517200.0 572400.0 527400.0 558600.0 ;
      RECT  517200.0 572400.0 527400.0 586200.0 ;
      RECT  517200.0 600000.0 527400.0 586200.0 ;
      RECT  517200.0 600000.0 527400.0 613800.0 ;
      RECT  517200.0 627600.0 527400.0 613800.0 ;
      RECT  517200.0 627600.0 527400.0 641400.0 ;
      RECT  517200.0 655200.0 527400.0 641400.0 ;
      RECT  517200.0 655200.0 527400.0 669000.0 ;
      RECT  517200.0 682800.0 527400.0 669000.0 ;
      RECT  517200.0 682800.0 527400.0 696600.0 ;
      RECT  517200.0 710400.0 527400.0 696600.0 ;
      RECT  517200.0 710400.0 527400.0 724200.0 ;
      RECT  517200.0 738000.0 527400.0 724200.0 ;
      RECT  517200.0 738000.0 527400.0 751800.0 ;
      RECT  517200.0 765600.0 527400.0 751800.0 ;
      RECT  517200.0 765600.0 527400.0 779400.0 ;
      RECT  517200.0 793200.0 527400.0 779400.0 ;
      RECT  517200.0 793200.0 527400.0 807000.0 ;
      RECT  517200.0 820800.0 527400.0 807000.0 ;
      RECT  517200.0 820800.0 527400.0 834600.0 ;
      RECT  517200.0 848400.0 527400.0 834600.0 ;
      RECT  517200.0 848400.0 527400.0 862200.0 ;
      RECT  517200.0 876000.0 527400.0 862200.0 ;
      RECT  517200.0 876000.0 527400.0 889800.0 ;
      RECT  517200.0 903600.0 527400.0 889800.0 ;
      RECT  517200.0 903600.0 527400.0 917400.0 ;
      RECT  517200.0 931200.0 527400.0 917400.0 ;
      RECT  517200.0 931200.0 527400.0 945000.0 ;
      RECT  517200.0 958800.0 527400.0 945000.0 ;
      RECT  517200.0 958800.0 527400.0 972600.0 ;
      RECT  517200.0 986400.0 527400.0 972600.0 ;
      RECT  517200.0 986400.0 527400.0 1000200.0 ;
      RECT  517200.0 1014000.0 527400.0 1000200.0 ;
      RECT  517200.0 1014000.0 527400.0 1027800.0 ;
      RECT  517200.0 1041600.0 527400.0 1027800.0 ;
      RECT  517200.0 1041600.0 527400.0 1055400.0 ;
      RECT  517200.0 1069200.0 527400.0 1055400.0 ;
      RECT  517200.0 1069200.0 527400.0 1083000.0 ;
      RECT  517200.0 1096800.0 527400.0 1083000.0 ;
      RECT  517200.0 1096800.0 527400.0 1110600.0 ;
      RECT  517200.0 1124400.0 527400.0 1110600.0 ;
      RECT  517200.0 1124400.0 527400.0 1138200.0 ;
      RECT  517200.0 1152000.0 527400.0 1138200.0 ;
      RECT  517200.0 1152000.0 527400.0 1165800.0 ;
      RECT  517200.0 1179600.0 527400.0 1165800.0 ;
      RECT  517200.0 1179600.0 527400.0 1193400.0 ;
      RECT  517200.0 1207200.0 527400.0 1193400.0 ;
      RECT  517200.0 1207200.0 527400.0 1221000.0 ;
      RECT  517200.0 1234800.0 527400.0 1221000.0 ;
      RECT  517200.0 1234800.0 527400.0 1248600.0 ;
      RECT  517200.0 1262400.0 527400.0 1248600.0 ;
      RECT  517200.0 1262400.0 527400.0 1276200.0 ;
      RECT  517200.0 1290000.0 527400.0 1276200.0 ;
      RECT  517200.0 1290000.0 527400.0 1303800.0 ;
      RECT  517200.0 1317600.0 527400.0 1303800.0 ;
      RECT  517200.0 1317600.0 527400.0 1331400.0 ;
      RECT  517200.0 1345200.0 527400.0 1331400.0 ;
      RECT  517200.0 1345200.0 527400.0 1359000.0 ;
      RECT  517200.0 1372800.0 527400.0 1359000.0 ;
      RECT  517200.0 1372800.0 527400.0 1386600.0 ;
      RECT  517200.0 1400400.0 527400.0 1386600.0 ;
      RECT  517200.0 1400400.0 527400.0 1414200.0 ;
      RECT  517200.0 1428000.0 527400.0 1414200.0 ;
      RECT  517200.0 1428000.0 527400.0 1441800.0 ;
      RECT  517200.0 1455600.0 527400.0 1441800.0 ;
      RECT  517200.0 1455600.0 527400.0 1469400.0 ;
      RECT  517200.0 1483200.0 527400.0 1469400.0 ;
      RECT  517200.0 1483200.0 527400.0 1497000.0 ;
      RECT  517200.0 1510800.0 527400.0 1497000.0 ;
      RECT  517200.0 1510800.0 527400.0 1524600.0 ;
      RECT  517200.0 1538400.0 527400.0 1524600.0 ;
      RECT  517200.0 1538400.0 527400.0 1552200.0 ;
      RECT  517200.0 1566000.0 527400.0 1552200.0 ;
      RECT  517200.0 1566000.0 527400.0 1579800.0 ;
      RECT  517200.0 1593600.0 527400.0 1579800.0 ;
      RECT  517200.0 1593600.0 527400.0 1607400.0 ;
      RECT  517200.0 1621200.0 527400.0 1607400.0 ;
      RECT  517200.0 1621200.0 527400.0 1635000.0 ;
      RECT  517200.0 1648800.0 527400.0 1635000.0 ;
      RECT  517200.0 1648800.0 527400.0 1662600.0 ;
      RECT  517200.0 1676400.0 527400.0 1662600.0 ;
      RECT  517200.0 1676400.0 527400.0 1690200.0 ;
      RECT  517200.0 1704000.0 527400.0 1690200.0 ;
      RECT  517200.0 1704000.0 527400.0 1717800.0 ;
      RECT  517200.0 1731600.0 527400.0 1717800.0 ;
      RECT  517200.0 1731600.0 527400.0 1745400.0 ;
      RECT  517200.0 1759200.0 527400.0 1745400.0 ;
      RECT  517200.0 1759200.0 527400.0 1773000.0 ;
      RECT  517200.0 1786800.0 527400.0 1773000.0 ;
      RECT  517200.0 1786800.0 527400.0 1800600.0 ;
      RECT  517200.0 1814400.0 527400.0 1800600.0 ;
      RECT  517200.0 1814400.0 527400.0 1828200.0 ;
      RECT  517200.0 1842000.0 527400.0 1828200.0 ;
      RECT  517200.0 1842000.0 527400.0 1855800.0 ;
      RECT  517200.0 1869600.0 527400.0 1855800.0 ;
      RECT  517200.0 1869600.0 527400.0 1883400.0 ;
      RECT  517200.0 1897200.0 527400.0 1883400.0 ;
      RECT  517200.0 1897200.0 527400.0 1911000.0 ;
      RECT  517200.0 1924800.0 527400.0 1911000.0 ;
      RECT  517200.0 1924800.0 527400.0 1938600.0 ;
      RECT  517200.0 1952400.0 527400.0 1938600.0 ;
      RECT  517200.0 1952400.0 527400.0 1966200.0 ;
      RECT  517200.0 1980000.0 527400.0 1966200.0 ;
      RECT  517200.0 1980000.0 527400.0 1993800.0 ;
      RECT  517200.0 2007600.0 527400.0 1993800.0 ;
      RECT  517200.0 2007600.0 527400.0 2021400.0 ;
      RECT  517200.0 2035200.0 527400.0 2021400.0 ;
      RECT  517200.0 2035200.0 527400.0 2049000.0 ;
      RECT  517200.0 2062800.0 527400.0 2049000.0 ;
      RECT  517200.0 2062800.0 527400.0 2076600.0 ;
      RECT  517200.0 2090400.0 527400.0 2076600.0 ;
      RECT  517200.0 2090400.0 527400.0 2104200.0 ;
      RECT  517200.0 2118000.0 527400.0 2104200.0 ;
      RECT  517200.0 2118000.0 527400.0 2131800.0 ;
      RECT  517200.0 2145600.0 527400.0 2131800.0 ;
      RECT  527400.0 379200.0 537600.0 393000.0 ;
      RECT  527400.0 406800.0 537600.0 393000.0 ;
      RECT  527400.0 406800.0 537600.0 420600.0 ;
      RECT  527400.0 434400.0 537600.0 420600.0 ;
      RECT  527400.0 434400.0 537600.0 448200.0 ;
      RECT  527400.0 462000.0 537600.0 448200.0 ;
      RECT  527400.0 462000.0 537600.0 475800.0 ;
      RECT  527400.0 489600.0 537600.0 475800.0 ;
      RECT  527400.0 489600.0 537600.0 503400.0 ;
      RECT  527400.0 517200.0 537600.0 503400.0 ;
      RECT  527400.0 517200.0 537600.0 531000.0 ;
      RECT  527400.0 544800.0 537600.0 531000.0 ;
      RECT  527400.0 544800.0 537600.0 558600.0 ;
      RECT  527400.0 572400.0 537600.0 558600.0 ;
      RECT  527400.0 572400.0 537600.0 586200.0 ;
      RECT  527400.0 600000.0 537600.0 586200.0 ;
      RECT  527400.0 600000.0 537600.0 613800.0 ;
      RECT  527400.0 627600.0 537600.0 613800.0 ;
      RECT  527400.0 627600.0 537600.0 641400.0 ;
      RECT  527400.0 655200.0 537600.0 641400.0 ;
      RECT  527400.0 655200.0 537600.0 669000.0 ;
      RECT  527400.0 682800.0 537600.0 669000.0 ;
      RECT  527400.0 682800.0 537600.0 696600.0 ;
      RECT  527400.0 710400.0 537600.0 696600.0 ;
      RECT  527400.0 710400.0 537600.0 724200.0 ;
      RECT  527400.0 738000.0 537600.0 724200.0 ;
      RECT  527400.0 738000.0 537600.0 751800.0 ;
      RECT  527400.0 765600.0 537600.0 751800.0 ;
      RECT  527400.0 765600.0 537600.0 779400.0 ;
      RECT  527400.0 793200.0 537600.0 779400.0 ;
      RECT  527400.0 793200.0 537600.0 807000.0 ;
      RECT  527400.0 820800.0 537600.0 807000.0 ;
      RECT  527400.0 820800.0 537600.0 834600.0 ;
      RECT  527400.0 848400.0 537600.0 834600.0 ;
      RECT  527400.0 848400.0 537600.0 862200.0 ;
      RECT  527400.0 876000.0 537600.0 862200.0 ;
      RECT  527400.0 876000.0 537600.0 889800.0 ;
      RECT  527400.0 903600.0 537600.0 889800.0 ;
      RECT  527400.0 903600.0 537600.0 917400.0 ;
      RECT  527400.0 931200.0 537600.0 917400.0 ;
      RECT  527400.0 931200.0 537600.0 945000.0 ;
      RECT  527400.0 958800.0 537600.0 945000.0 ;
      RECT  527400.0 958800.0 537600.0 972600.0 ;
      RECT  527400.0 986400.0 537600.0 972600.0 ;
      RECT  527400.0 986400.0 537600.0 1000200.0 ;
      RECT  527400.0 1014000.0 537600.0 1000200.0 ;
      RECT  527400.0 1014000.0 537600.0 1027800.0 ;
      RECT  527400.0 1041600.0 537600.0 1027800.0 ;
      RECT  527400.0 1041600.0 537600.0 1055400.0 ;
      RECT  527400.0 1069200.0 537600.0 1055400.0 ;
      RECT  527400.0 1069200.0 537600.0 1083000.0 ;
      RECT  527400.0 1096800.0 537600.0 1083000.0 ;
      RECT  527400.0 1096800.0 537600.0 1110600.0 ;
      RECT  527400.0 1124400.0 537600.0 1110600.0 ;
      RECT  527400.0 1124400.0 537600.0 1138200.0 ;
      RECT  527400.0 1152000.0 537600.0 1138200.0 ;
      RECT  527400.0 1152000.0 537600.0 1165800.0 ;
      RECT  527400.0 1179600.0 537600.0 1165800.0 ;
      RECT  527400.0 1179600.0 537600.0 1193400.0 ;
      RECT  527400.0 1207200.0 537600.0 1193400.0 ;
      RECT  527400.0 1207200.0 537600.0 1221000.0 ;
      RECT  527400.0 1234800.0 537600.0 1221000.0 ;
      RECT  527400.0 1234800.0 537600.0 1248600.0 ;
      RECT  527400.0 1262400.0 537600.0 1248600.0 ;
      RECT  527400.0 1262400.0 537600.0 1276200.0 ;
      RECT  527400.0 1290000.0 537600.0 1276200.0 ;
      RECT  527400.0 1290000.0 537600.0 1303800.0 ;
      RECT  527400.0 1317600.0 537600.0 1303800.0 ;
      RECT  527400.0 1317600.0 537600.0 1331400.0 ;
      RECT  527400.0 1345200.0 537600.0 1331400.0 ;
      RECT  527400.0 1345200.0 537600.0 1359000.0 ;
      RECT  527400.0 1372800.0 537600.0 1359000.0 ;
      RECT  527400.0 1372800.0 537600.0 1386600.0 ;
      RECT  527400.0 1400400.0 537600.0 1386600.0 ;
      RECT  527400.0 1400400.0 537600.0 1414200.0 ;
      RECT  527400.0 1428000.0 537600.0 1414200.0 ;
      RECT  527400.0 1428000.0 537600.0 1441800.0 ;
      RECT  527400.0 1455600.0 537600.0 1441800.0 ;
      RECT  527400.0 1455600.0 537600.0 1469400.0 ;
      RECT  527400.0 1483200.0 537600.0 1469400.0 ;
      RECT  527400.0 1483200.0 537600.0 1497000.0 ;
      RECT  527400.0 1510800.0 537600.0 1497000.0 ;
      RECT  527400.0 1510800.0 537600.0 1524600.0 ;
      RECT  527400.0 1538400.0 537600.0 1524600.0 ;
      RECT  527400.0 1538400.0 537600.0 1552200.0 ;
      RECT  527400.0 1566000.0 537600.0 1552200.0 ;
      RECT  527400.0 1566000.0 537600.0 1579800.0 ;
      RECT  527400.0 1593600.0 537600.0 1579800.0 ;
      RECT  527400.0 1593600.0 537600.0 1607400.0 ;
      RECT  527400.0 1621200.0 537600.0 1607400.0 ;
      RECT  527400.0 1621200.0 537600.0 1635000.0 ;
      RECT  527400.0 1648800.0 537600.0 1635000.0 ;
      RECT  527400.0 1648800.0 537600.0 1662600.0 ;
      RECT  527400.0 1676400.0 537600.0 1662600.0 ;
      RECT  527400.0 1676400.0 537600.0 1690200.0 ;
      RECT  527400.0 1704000.0 537600.0 1690200.0 ;
      RECT  527400.0 1704000.0 537600.0 1717800.0 ;
      RECT  527400.0 1731600.0 537600.0 1717800.0 ;
      RECT  527400.0 1731600.0 537600.0 1745400.0 ;
      RECT  527400.0 1759200.0 537600.0 1745400.0 ;
      RECT  527400.0 1759200.0 537600.0 1773000.0 ;
      RECT  527400.0 1786800.0 537600.0 1773000.0 ;
      RECT  527400.0 1786800.0 537600.0 1800600.0 ;
      RECT  527400.0 1814400.0 537600.0 1800600.0 ;
      RECT  527400.0 1814400.0 537600.0 1828200.0 ;
      RECT  527400.0 1842000.0 537600.0 1828200.0 ;
      RECT  527400.0 1842000.0 537600.0 1855800.0 ;
      RECT  527400.0 1869600.0 537600.0 1855800.0 ;
      RECT  527400.0 1869600.0 537600.0 1883400.0 ;
      RECT  527400.0 1897200.0 537600.0 1883400.0 ;
      RECT  527400.0 1897200.0 537600.0 1911000.0 ;
      RECT  527400.0 1924800.0 537600.0 1911000.0 ;
      RECT  527400.0 1924800.0 537600.0 1938600.0 ;
      RECT  527400.0 1952400.0 537600.0 1938600.0 ;
      RECT  527400.0 1952400.0 537600.0 1966200.0 ;
      RECT  527400.0 1980000.0 537600.0 1966200.0 ;
      RECT  527400.0 1980000.0 537600.0 1993800.0 ;
      RECT  527400.0 2007600.0 537600.0 1993800.0 ;
      RECT  527400.0 2007600.0 537600.0 2021400.0 ;
      RECT  527400.0 2035200.0 537600.0 2021400.0 ;
      RECT  527400.0 2035200.0 537600.0 2049000.0 ;
      RECT  527400.0 2062800.0 537600.0 2049000.0 ;
      RECT  527400.0 2062800.0 537600.0 2076600.0 ;
      RECT  527400.0 2090400.0 537600.0 2076600.0 ;
      RECT  527400.0 2090400.0 537600.0 2104200.0 ;
      RECT  527400.0 2118000.0 537600.0 2104200.0 ;
      RECT  527400.0 2118000.0 537600.0 2131800.0 ;
      RECT  527400.0 2145600.0 537600.0 2131800.0 ;
      RECT  537600.0 379200.0 547800.0 393000.0 ;
      RECT  537600.0 406800.0 547800.0 393000.0 ;
      RECT  537600.0 406800.0 547800.0 420600.0 ;
      RECT  537600.0 434400.0 547800.0 420600.0 ;
      RECT  537600.0 434400.0 547800.0 448200.0 ;
      RECT  537600.0 462000.0 547800.0 448200.0 ;
      RECT  537600.0 462000.0 547800.0 475800.0 ;
      RECT  537600.0 489600.0 547800.0 475800.0 ;
      RECT  537600.0 489600.0 547800.0 503400.0 ;
      RECT  537600.0 517200.0 547800.0 503400.0 ;
      RECT  537600.0 517200.0 547800.0 531000.0 ;
      RECT  537600.0 544800.0 547800.0 531000.0 ;
      RECT  537600.0 544800.0 547800.0 558600.0 ;
      RECT  537600.0 572400.0 547800.0 558600.0 ;
      RECT  537600.0 572400.0 547800.0 586200.0 ;
      RECT  537600.0 600000.0 547800.0 586200.0 ;
      RECT  537600.0 600000.0 547800.0 613800.0 ;
      RECT  537600.0 627600.0 547800.0 613800.0 ;
      RECT  537600.0 627600.0 547800.0 641400.0 ;
      RECT  537600.0 655200.0 547800.0 641400.0 ;
      RECT  537600.0 655200.0 547800.0 669000.0 ;
      RECT  537600.0 682800.0 547800.0 669000.0 ;
      RECT  537600.0 682800.0 547800.0 696600.0 ;
      RECT  537600.0 710400.0 547800.0 696600.0 ;
      RECT  537600.0 710400.0 547800.0 724200.0 ;
      RECT  537600.0 738000.0 547800.0 724200.0 ;
      RECT  537600.0 738000.0 547800.0 751800.0 ;
      RECT  537600.0 765600.0 547800.0 751800.0 ;
      RECT  537600.0 765600.0 547800.0 779400.0 ;
      RECT  537600.0 793200.0 547800.0 779400.0 ;
      RECT  537600.0 793200.0 547800.0 807000.0 ;
      RECT  537600.0 820800.0 547800.0 807000.0 ;
      RECT  537600.0 820800.0 547800.0 834600.0 ;
      RECT  537600.0 848400.0 547800.0 834600.0 ;
      RECT  537600.0 848400.0 547800.0 862200.0 ;
      RECT  537600.0 876000.0 547800.0 862200.0 ;
      RECT  537600.0 876000.0 547800.0 889800.0 ;
      RECT  537600.0 903600.0 547800.0 889800.0 ;
      RECT  537600.0 903600.0 547800.0 917400.0 ;
      RECT  537600.0 931200.0 547800.0 917400.0 ;
      RECT  537600.0 931200.0 547800.0 945000.0 ;
      RECT  537600.0 958800.0 547800.0 945000.0 ;
      RECT  537600.0 958800.0 547800.0 972600.0 ;
      RECT  537600.0 986400.0 547800.0 972600.0 ;
      RECT  537600.0 986400.0 547800.0 1000200.0 ;
      RECT  537600.0 1014000.0 547800.0 1000200.0 ;
      RECT  537600.0 1014000.0 547800.0 1027800.0 ;
      RECT  537600.0 1041600.0 547800.0 1027800.0 ;
      RECT  537600.0 1041600.0 547800.0 1055400.0 ;
      RECT  537600.0 1069200.0 547800.0 1055400.0 ;
      RECT  537600.0 1069200.0 547800.0 1083000.0 ;
      RECT  537600.0 1096800.0 547800.0 1083000.0 ;
      RECT  537600.0 1096800.0 547800.0 1110600.0 ;
      RECT  537600.0 1124400.0 547800.0 1110600.0 ;
      RECT  537600.0 1124400.0 547800.0 1138200.0 ;
      RECT  537600.0 1152000.0 547800.0 1138200.0 ;
      RECT  537600.0 1152000.0 547800.0 1165800.0 ;
      RECT  537600.0 1179600.0 547800.0 1165800.0 ;
      RECT  537600.0 1179600.0 547800.0 1193400.0 ;
      RECT  537600.0 1207200.0 547800.0 1193400.0 ;
      RECT  537600.0 1207200.0 547800.0 1221000.0 ;
      RECT  537600.0 1234800.0 547800.0 1221000.0 ;
      RECT  537600.0 1234800.0 547800.0 1248600.0 ;
      RECT  537600.0 1262400.0 547800.0 1248600.0 ;
      RECT  537600.0 1262400.0 547800.0 1276200.0 ;
      RECT  537600.0 1290000.0 547800.0 1276200.0 ;
      RECT  537600.0 1290000.0 547800.0 1303800.0 ;
      RECT  537600.0 1317600.0 547800.0 1303800.0 ;
      RECT  537600.0 1317600.0 547800.0 1331400.0 ;
      RECT  537600.0 1345200.0 547800.0 1331400.0 ;
      RECT  537600.0 1345200.0 547800.0 1359000.0 ;
      RECT  537600.0 1372800.0 547800.0 1359000.0 ;
      RECT  537600.0 1372800.0 547800.0 1386600.0 ;
      RECT  537600.0 1400400.0 547800.0 1386600.0 ;
      RECT  537600.0 1400400.0 547800.0 1414200.0 ;
      RECT  537600.0 1428000.0 547800.0 1414200.0 ;
      RECT  537600.0 1428000.0 547800.0 1441800.0 ;
      RECT  537600.0 1455600.0 547800.0 1441800.0 ;
      RECT  537600.0 1455600.0 547800.0 1469400.0 ;
      RECT  537600.0 1483200.0 547800.0 1469400.0 ;
      RECT  537600.0 1483200.0 547800.0 1497000.0 ;
      RECT  537600.0 1510800.0 547800.0 1497000.0 ;
      RECT  537600.0 1510800.0 547800.0 1524600.0 ;
      RECT  537600.0 1538400.0 547800.0 1524600.0 ;
      RECT  537600.0 1538400.0 547800.0 1552200.0 ;
      RECT  537600.0 1566000.0 547800.0 1552200.0 ;
      RECT  537600.0 1566000.0 547800.0 1579800.0 ;
      RECT  537600.0 1593600.0 547800.0 1579800.0 ;
      RECT  537600.0 1593600.0 547800.0 1607400.0 ;
      RECT  537600.0 1621200.0 547800.0 1607400.0 ;
      RECT  537600.0 1621200.0 547800.0 1635000.0 ;
      RECT  537600.0 1648800.0 547800.0 1635000.0 ;
      RECT  537600.0 1648800.0 547800.0 1662600.0 ;
      RECT  537600.0 1676400.0 547800.0 1662600.0 ;
      RECT  537600.0 1676400.0 547800.0 1690200.0 ;
      RECT  537600.0 1704000.0 547800.0 1690200.0 ;
      RECT  537600.0 1704000.0 547800.0 1717800.0 ;
      RECT  537600.0 1731600.0 547800.0 1717800.0 ;
      RECT  537600.0 1731600.0 547800.0 1745400.0 ;
      RECT  537600.0 1759200.0 547800.0 1745400.0 ;
      RECT  537600.0 1759200.0 547800.0 1773000.0 ;
      RECT  537600.0 1786800.0 547800.0 1773000.0 ;
      RECT  537600.0 1786800.0 547800.0 1800600.0 ;
      RECT  537600.0 1814400.0 547800.0 1800600.0 ;
      RECT  537600.0 1814400.0 547800.0 1828200.0 ;
      RECT  537600.0 1842000.0 547800.0 1828200.0 ;
      RECT  537600.0 1842000.0 547800.0 1855800.0 ;
      RECT  537600.0 1869600.0 547800.0 1855800.0 ;
      RECT  537600.0 1869600.0 547800.0 1883400.0 ;
      RECT  537600.0 1897200.0 547800.0 1883400.0 ;
      RECT  537600.0 1897200.0 547800.0 1911000.0 ;
      RECT  537600.0 1924800.0 547800.0 1911000.0 ;
      RECT  537600.0 1924800.0 547800.0 1938600.0 ;
      RECT  537600.0 1952400.0 547800.0 1938600.0 ;
      RECT  537600.0 1952400.0 547800.0 1966200.0 ;
      RECT  537600.0 1980000.0 547800.0 1966200.0 ;
      RECT  537600.0 1980000.0 547800.0 1993800.0 ;
      RECT  537600.0 2007600.0 547800.0 1993800.0 ;
      RECT  537600.0 2007600.0 547800.0 2021400.0 ;
      RECT  537600.0 2035200.0 547800.0 2021400.0 ;
      RECT  537600.0 2035200.0 547800.0 2049000.0 ;
      RECT  537600.0 2062800.0 547800.0 2049000.0 ;
      RECT  537600.0 2062800.0 547800.0 2076600.0 ;
      RECT  537600.0 2090400.0 547800.0 2076600.0 ;
      RECT  537600.0 2090400.0 547800.0 2104200.0 ;
      RECT  537600.0 2118000.0 547800.0 2104200.0 ;
      RECT  537600.0 2118000.0 547800.0 2131800.0 ;
      RECT  537600.0 2145600.0 547800.0 2131800.0 ;
      RECT  547800.0 379200.0 558000.0 393000.0 ;
      RECT  547800.0 406800.0 558000.0 393000.0 ;
      RECT  547800.0 406800.0 558000.0 420600.0 ;
      RECT  547800.0 434400.0 558000.0 420600.0 ;
      RECT  547800.0 434400.0 558000.0 448200.0 ;
      RECT  547800.0 462000.0 558000.0 448200.0 ;
      RECT  547800.0 462000.0 558000.0 475800.0 ;
      RECT  547800.0 489600.0 558000.0 475800.0 ;
      RECT  547800.0 489600.0 558000.0 503400.0 ;
      RECT  547800.0 517200.0 558000.0 503400.0 ;
      RECT  547800.0 517200.0 558000.0 531000.0 ;
      RECT  547800.0 544800.0 558000.0 531000.0 ;
      RECT  547800.0 544800.0 558000.0 558600.0 ;
      RECT  547800.0 572400.0 558000.0 558600.0 ;
      RECT  547800.0 572400.0 558000.0 586200.0 ;
      RECT  547800.0 600000.0 558000.0 586200.0 ;
      RECT  547800.0 600000.0 558000.0 613800.0 ;
      RECT  547800.0 627600.0 558000.0 613800.0 ;
      RECT  547800.0 627600.0 558000.0 641400.0 ;
      RECT  547800.0 655200.0 558000.0 641400.0 ;
      RECT  547800.0 655200.0 558000.0 669000.0 ;
      RECT  547800.0 682800.0 558000.0 669000.0 ;
      RECT  547800.0 682800.0 558000.0 696600.0 ;
      RECT  547800.0 710400.0 558000.0 696600.0 ;
      RECT  547800.0 710400.0 558000.0 724200.0 ;
      RECT  547800.0 738000.0 558000.0 724200.0 ;
      RECT  547800.0 738000.0 558000.0 751800.0 ;
      RECT  547800.0 765600.0 558000.0 751800.0 ;
      RECT  547800.0 765600.0 558000.0 779400.0 ;
      RECT  547800.0 793200.0 558000.0 779400.0 ;
      RECT  547800.0 793200.0 558000.0 807000.0 ;
      RECT  547800.0 820800.0 558000.0 807000.0 ;
      RECT  547800.0 820800.0 558000.0 834600.0 ;
      RECT  547800.0 848400.0 558000.0 834600.0 ;
      RECT  547800.0 848400.0 558000.0 862200.0 ;
      RECT  547800.0 876000.0 558000.0 862200.0 ;
      RECT  547800.0 876000.0 558000.0 889800.0 ;
      RECT  547800.0 903600.0 558000.0 889800.0 ;
      RECT  547800.0 903600.0 558000.0 917400.0 ;
      RECT  547800.0 931200.0 558000.0 917400.0 ;
      RECT  547800.0 931200.0 558000.0 945000.0 ;
      RECT  547800.0 958800.0 558000.0 945000.0 ;
      RECT  547800.0 958800.0 558000.0 972600.0 ;
      RECT  547800.0 986400.0 558000.0 972600.0 ;
      RECT  547800.0 986400.0 558000.0 1000200.0 ;
      RECT  547800.0 1014000.0 558000.0 1000200.0 ;
      RECT  547800.0 1014000.0 558000.0 1027800.0 ;
      RECT  547800.0 1041600.0 558000.0 1027800.0 ;
      RECT  547800.0 1041600.0 558000.0 1055400.0 ;
      RECT  547800.0 1069200.0 558000.0 1055400.0 ;
      RECT  547800.0 1069200.0 558000.0 1083000.0 ;
      RECT  547800.0 1096800.0 558000.0 1083000.0 ;
      RECT  547800.0 1096800.0 558000.0 1110600.0 ;
      RECT  547800.0 1124400.0 558000.0 1110600.0 ;
      RECT  547800.0 1124400.0 558000.0 1138200.0 ;
      RECT  547800.0 1152000.0 558000.0 1138200.0 ;
      RECT  547800.0 1152000.0 558000.0 1165800.0 ;
      RECT  547800.0 1179600.0 558000.0 1165800.0 ;
      RECT  547800.0 1179600.0 558000.0 1193400.0 ;
      RECT  547800.0 1207200.0 558000.0 1193400.0 ;
      RECT  547800.0 1207200.0 558000.0 1221000.0 ;
      RECT  547800.0 1234800.0 558000.0 1221000.0 ;
      RECT  547800.0 1234800.0 558000.0 1248600.0 ;
      RECT  547800.0 1262400.0 558000.0 1248600.0 ;
      RECT  547800.0 1262400.0 558000.0 1276200.0 ;
      RECT  547800.0 1290000.0 558000.0 1276200.0 ;
      RECT  547800.0 1290000.0 558000.0 1303800.0 ;
      RECT  547800.0 1317600.0 558000.0 1303800.0 ;
      RECT  547800.0 1317600.0 558000.0 1331400.0 ;
      RECT  547800.0 1345200.0 558000.0 1331400.0 ;
      RECT  547800.0 1345200.0 558000.0 1359000.0 ;
      RECT  547800.0 1372800.0 558000.0 1359000.0 ;
      RECT  547800.0 1372800.0 558000.0 1386600.0 ;
      RECT  547800.0 1400400.0 558000.0 1386600.0 ;
      RECT  547800.0 1400400.0 558000.0 1414200.0 ;
      RECT  547800.0 1428000.0 558000.0 1414200.0 ;
      RECT  547800.0 1428000.0 558000.0 1441800.0 ;
      RECT  547800.0 1455600.0 558000.0 1441800.0 ;
      RECT  547800.0 1455600.0 558000.0 1469400.0 ;
      RECT  547800.0 1483200.0 558000.0 1469400.0 ;
      RECT  547800.0 1483200.0 558000.0 1497000.0 ;
      RECT  547800.0 1510800.0 558000.0 1497000.0 ;
      RECT  547800.0 1510800.0 558000.0 1524600.0 ;
      RECT  547800.0 1538400.0 558000.0 1524600.0 ;
      RECT  547800.0 1538400.0 558000.0 1552200.0 ;
      RECT  547800.0 1566000.0 558000.0 1552200.0 ;
      RECT  547800.0 1566000.0 558000.0 1579800.0 ;
      RECT  547800.0 1593600.0 558000.0 1579800.0 ;
      RECT  547800.0 1593600.0 558000.0 1607400.0 ;
      RECT  547800.0 1621200.0 558000.0 1607400.0 ;
      RECT  547800.0 1621200.0 558000.0 1635000.0 ;
      RECT  547800.0 1648800.0 558000.0 1635000.0 ;
      RECT  547800.0 1648800.0 558000.0 1662600.0 ;
      RECT  547800.0 1676400.0 558000.0 1662600.0 ;
      RECT  547800.0 1676400.0 558000.0 1690200.0 ;
      RECT  547800.0 1704000.0 558000.0 1690200.0 ;
      RECT  547800.0 1704000.0 558000.0 1717800.0 ;
      RECT  547800.0 1731600.0 558000.0 1717800.0 ;
      RECT  547800.0 1731600.0 558000.0 1745400.0 ;
      RECT  547800.0 1759200.0 558000.0 1745400.0 ;
      RECT  547800.0 1759200.0 558000.0 1773000.0 ;
      RECT  547800.0 1786800.0 558000.0 1773000.0 ;
      RECT  547800.0 1786800.0 558000.0 1800600.0 ;
      RECT  547800.0 1814400.0 558000.0 1800600.0 ;
      RECT  547800.0 1814400.0 558000.0 1828200.0 ;
      RECT  547800.0 1842000.0 558000.0 1828200.0 ;
      RECT  547800.0 1842000.0 558000.0 1855800.0 ;
      RECT  547800.0 1869600.0 558000.0 1855800.0 ;
      RECT  547800.0 1869600.0 558000.0 1883400.0 ;
      RECT  547800.0 1897200.0 558000.0 1883400.0 ;
      RECT  547800.0 1897200.0 558000.0 1911000.0 ;
      RECT  547800.0 1924800.0 558000.0 1911000.0 ;
      RECT  547800.0 1924800.0 558000.0 1938600.0 ;
      RECT  547800.0 1952400.0 558000.0 1938600.0 ;
      RECT  547800.0 1952400.0 558000.0 1966200.0 ;
      RECT  547800.0 1980000.0 558000.0 1966200.0 ;
      RECT  547800.0 1980000.0 558000.0 1993800.0 ;
      RECT  547800.0 2007600.0 558000.0 1993800.0 ;
      RECT  547800.0 2007600.0 558000.0 2021400.0 ;
      RECT  547800.0 2035200.0 558000.0 2021400.0 ;
      RECT  547800.0 2035200.0 558000.0 2049000.0 ;
      RECT  547800.0 2062800.0 558000.0 2049000.0 ;
      RECT  547800.0 2062800.0 558000.0 2076600.0 ;
      RECT  547800.0 2090400.0 558000.0 2076600.0 ;
      RECT  547800.0 2090400.0 558000.0 2104200.0 ;
      RECT  547800.0 2118000.0 558000.0 2104200.0 ;
      RECT  547800.0 2118000.0 558000.0 2131800.0 ;
      RECT  547800.0 2145600.0 558000.0 2131800.0 ;
      RECT  558000.0 379200.0 568200.0 393000.0 ;
      RECT  558000.0 406800.0 568200.0 393000.0 ;
      RECT  558000.0 406800.0 568200.0 420600.0 ;
      RECT  558000.0 434400.0 568200.0 420600.0 ;
      RECT  558000.0 434400.0 568200.0 448200.0 ;
      RECT  558000.0 462000.0 568200.0 448200.0 ;
      RECT  558000.0 462000.0 568200.0 475800.0 ;
      RECT  558000.0 489600.0 568200.0 475800.0 ;
      RECT  558000.0 489600.0 568200.0 503400.0 ;
      RECT  558000.0 517200.0 568200.0 503400.0 ;
      RECT  558000.0 517200.0 568200.0 531000.0 ;
      RECT  558000.0 544800.0 568200.0 531000.0 ;
      RECT  558000.0 544800.0 568200.0 558600.0 ;
      RECT  558000.0 572400.0 568200.0 558600.0 ;
      RECT  558000.0 572400.0 568200.0 586200.0 ;
      RECT  558000.0 600000.0 568200.0 586200.0 ;
      RECT  558000.0 600000.0 568200.0 613800.0 ;
      RECT  558000.0 627600.0 568200.0 613800.0 ;
      RECT  558000.0 627600.0 568200.0 641400.0 ;
      RECT  558000.0 655200.0 568200.0 641400.0 ;
      RECT  558000.0 655200.0 568200.0 669000.0 ;
      RECT  558000.0 682800.0 568200.0 669000.0 ;
      RECT  558000.0 682800.0 568200.0 696600.0 ;
      RECT  558000.0 710400.0 568200.0 696600.0 ;
      RECT  558000.0 710400.0 568200.0 724200.0 ;
      RECT  558000.0 738000.0 568200.0 724200.0 ;
      RECT  558000.0 738000.0 568200.0 751800.0 ;
      RECT  558000.0 765600.0 568200.0 751800.0 ;
      RECT  558000.0 765600.0 568200.0 779400.0 ;
      RECT  558000.0 793200.0 568200.0 779400.0 ;
      RECT  558000.0 793200.0 568200.0 807000.0 ;
      RECT  558000.0 820800.0 568200.0 807000.0 ;
      RECT  558000.0 820800.0 568200.0 834600.0 ;
      RECT  558000.0 848400.0 568200.0 834600.0 ;
      RECT  558000.0 848400.0 568200.0 862200.0 ;
      RECT  558000.0 876000.0 568200.0 862200.0 ;
      RECT  558000.0 876000.0 568200.0 889800.0 ;
      RECT  558000.0 903600.0 568200.0 889800.0 ;
      RECT  558000.0 903600.0 568200.0 917400.0 ;
      RECT  558000.0 931200.0 568200.0 917400.0 ;
      RECT  558000.0 931200.0 568200.0 945000.0 ;
      RECT  558000.0 958800.0 568200.0 945000.0 ;
      RECT  558000.0 958800.0 568200.0 972600.0 ;
      RECT  558000.0 986400.0 568200.0 972600.0 ;
      RECT  558000.0 986400.0 568200.0 1000200.0 ;
      RECT  558000.0 1014000.0 568200.0 1000200.0 ;
      RECT  558000.0 1014000.0 568200.0 1027800.0 ;
      RECT  558000.0 1041600.0 568200.0 1027800.0 ;
      RECT  558000.0 1041600.0 568200.0 1055400.0 ;
      RECT  558000.0 1069200.0 568200.0 1055400.0 ;
      RECT  558000.0 1069200.0 568200.0 1083000.0 ;
      RECT  558000.0 1096800.0 568200.0 1083000.0 ;
      RECT  558000.0 1096800.0 568200.0 1110600.0 ;
      RECT  558000.0 1124400.0 568200.0 1110600.0 ;
      RECT  558000.0 1124400.0 568200.0 1138200.0 ;
      RECT  558000.0 1152000.0 568200.0 1138200.0 ;
      RECT  558000.0 1152000.0 568200.0 1165800.0 ;
      RECT  558000.0 1179600.0 568200.0 1165800.0 ;
      RECT  558000.0 1179600.0 568200.0 1193400.0 ;
      RECT  558000.0 1207200.0 568200.0 1193400.0 ;
      RECT  558000.0 1207200.0 568200.0 1221000.0 ;
      RECT  558000.0 1234800.0 568200.0 1221000.0 ;
      RECT  558000.0 1234800.0 568200.0 1248600.0 ;
      RECT  558000.0 1262400.0 568200.0 1248600.0 ;
      RECT  558000.0 1262400.0 568200.0 1276200.0 ;
      RECT  558000.0 1290000.0 568200.0 1276200.0 ;
      RECT  558000.0 1290000.0 568200.0 1303800.0 ;
      RECT  558000.0 1317600.0 568200.0 1303800.0 ;
      RECT  558000.0 1317600.0 568200.0 1331400.0 ;
      RECT  558000.0 1345200.0 568200.0 1331400.0 ;
      RECT  558000.0 1345200.0 568200.0 1359000.0 ;
      RECT  558000.0 1372800.0 568200.0 1359000.0 ;
      RECT  558000.0 1372800.0 568200.0 1386600.0 ;
      RECT  558000.0 1400400.0 568200.0 1386600.0 ;
      RECT  558000.0 1400400.0 568200.0 1414200.0 ;
      RECT  558000.0 1428000.0 568200.0 1414200.0 ;
      RECT  558000.0 1428000.0 568200.0 1441800.0 ;
      RECT  558000.0 1455600.0 568200.0 1441800.0 ;
      RECT  558000.0 1455600.0 568200.0 1469400.0 ;
      RECT  558000.0 1483200.0 568200.0 1469400.0 ;
      RECT  558000.0 1483200.0 568200.0 1497000.0 ;
      RECT  558000.0 1510800.0 568200.0 1497000.0 ;
      RECT  558000.0 1510800.0 568200.0 1524600.0 ;
      RECT  558000.0 1538400.0 568200.0 1524600.0 ;
      RECT  558000.0 1538400.0 568200.0 1552200.0 ;
      RECT  558000.0 1566000.0 568200.0 1552200.0 ;
      RECT  558000.0 1566000.0 568200.0 1579800.0 ;
      RECT  558000.0 1593600.0 568200.0 1579800.0 ;
      RECT  558000.0 1593600.0 568200.0 1607400.0 ;
      RECT  558000.0 1621200.0 568200.0 1607400.0 ;
      RECT  558000.0 1621200.0 568200.0 1635000.0 ;
      RECT  558000.0 1648800.0 568200.0 1635000.0 ;
      RECT  558000.0 1648800.0 568200.0 1662600.0 ;
      RECT  558000.0 1676400.0 568200.0 1662600.0 ;
      RECT  558000.0 1676400.0 568200.0 1690200.0 ;
      RECT  558000.0 1704000.0 568200.0 1690200.0 ;
      RECT  558000.0 1704000.0 568200.0 1717800.0 ;
      RECT  558000.0 1731600.0 568200.0 1717800.0 ;
      RECT  558000.0 1731600.0 568200.0 1745400.0 ;
      RECT  558000.0 1759200.0 568200.0 1745400.0 ;
      RECT  558000.0 1759200.0 568200.0 1773000.0 ;
      RECT  558000.0 1786800.0 568200.0 1773000.0 ;
      RECT  558000.0 1786800.0 568200.0 1800600.0 ;
      RECT  558000.0 1814400.0 568200.0 1800600.0 ;
      RECT  558000.0 1814400.0 568200.0 1828200.0 ;
      RECT  558000.0 1842000.0 568200.0 1828200.0 ;
      RECT  558000.0 1842000.0 568200.0 1855800.0 ;
      RECT  558000.0 1869600.0 568200.0 1855800.0 ;
      RECT  558000.0 1869600.0 568200.0 1883400.0 ;
      RECT  558000.0 1897200.0 568200.0 1883400.0 ;
      RECT  558000.0 1897200.0 568200.0 1911000.0 ;
      RECT  558000.0 1924800.0 568200.0 1911000.0 ;
      RECT  558000.0 1924800.0 568200.0 1938600.0 ;
      RECT  558000.0 1952400.0 568200.0 1938600.0 ;
      RECT  558000.0 1952400.0 568200.0 1966200.0 ;
      RECT  558000.0 1980000.0 568200.0 1966200.0 ;
      RECT  558000.0 1980000.0 568200.0 1993800.0 ;
      RECT  558000.0 2007600.0 568200.0 1993800.0 ;
      RECT  558000.0 2007600.0 568200.0 2021400.0 ;
      RECT  558000.0 2035200.0 568200.0 2021400.0 ;
      RECT  558000.0 2035200.0 568200.0 2049000.0 ;
      RECT  558000.0 2062800.0 568200.0 2049000.0 ;
      RECT  558000.0 2062800.0 568200.0 2076600.0 ;
      RECT  558000.0 2090400.0 568200.0 2076600.0 ;
      RECT  558000.0 2090400.0 568200.0 2104200.0 ;
      RECT  558000.0 2118000.0 568200.0 2104200.0 ;
      RECT  558000.0 2118000.0 568200.0 2131800.0 ;
      RECT  558000.0 2145600.0 568200.0 2131800.0 ;
      RECT  568200.0 379200.0 578400.0 393000.0 ;
      RECT  568200.0 406800.0 578400.0 393000.0 ;
      RECT  568200.0 406800.0 578400.0 420600.0 ;
      RECT  568200.0 434400.0 578400.0 420600.0 ;
      RECT  568200.0 434400.0 578400.0 448200.0 ;
      RECT  568200.0 462000.0 578400.0 448200.0 ;
      RECT  568200.0 462000.0 578400.0 475800.0 ;
      RECT  568200.0 489600.0 578400.0 475800.0 ;
      RECT  568200.0 489600.0 578400.0 503400.0 ;
      RECT  568200.0 517200.0 578400.0 503400.0 ;
      RECT  568200.0 517200.0 578400.0 531000.0 ;
      RECT  568200.0 544800.0 578400.0 531000.0 ;
      RECT  568200.0 544800.0 578400.0 558600.0 ;
      RECT  568200.0 572400.0 578400.0 558600.0 ;
      RECT  568200.0 572400.0 578400.0 586200.0 ;
      RECT  568200.0 600000.0 578400.0 586200.0 ;
      RECT  568200.0 600000.0 578400.0 613800.0 ;
      RECT  568200.0 627600.0 578400.0 613800.0 ;
      RECT  568200.0 627600.0 578400.0 641400.0 ;
      RECT  568200.0 655200.0 578400.0 641400.0 ;
      RECT  568200.0 655200.0 578400.0 669000.0 ;
      RECT  568200.0 682800.0 578400.0 669000.0 ;
      RECT  568200.0 682800.0 578400.0 696600.0 ;
      RECT  568200.0 710400.0 578400.0 696600.0 ;
      RECT  568200.0 710400.0 578400.0 724200.0 ;
      RECT  568200.0 738000.0 578400.0 724200.0 ;
      RECT  568200.0 738000.0 578400.0 751800.0 ;
      RECT  568200.0 765600.0 578400.0 751800.0 ;
      RECT  568200.0 765600.0 578400.0 779400.0 ;
      RECT  568200.0 793200.0 578400.0 779400.0 ;
      RECT  568200.0 793200.0 578400.0 807000.0 ;
      RECT  568200.0 820800.0 578400.0 807000.0 ;
      RECT  568200.0 820800.0 578400.0 834600.0 ;
      RECT  568200.0 848400.0 578400.0 834600.0 ;
      RECT  568200.0 848400.0 578400.0 862200.0 ;
      RECT  568200.0 876000.0 578400.0 862200.0 ;
      RECT  568200.0 876000.0 578400.0 889800.0 ;
      RECT  568200.0 903600.0 578400.0 889800.0 ;
      RECT  568200.0 903600.0 578400.0 917400.0 ;
      RECT  568200.0 931200.0 578400.0 917400.0 ;
      RECT  568200.0 931200.0 578400.0 945000.0 ;
      RECT  568200.0 958800.0 578400.0 945000.0 ;
      RECT  568200.0 958800.0 578400.0 972600.0 ;
      RECT  568200.0 986400.0 578400.0 972600.0 ;
      RECT  568200.0 986400.0 578400.0 1000200.0 ;
      RECT  568200.0 1014000.0 578400.0 1000200.0 ;
      RECT  568200.0 1014000.0 578400.0 1027800.0 ;
      RECT  568200.0 1041600.0 578400.0 1027800.0 ;
      RECT  568200.0 1041600.0 578400.0 1055400.0 ;
      RECT  568200.0 1069200.0 578400.0 1055400.0 ;
      RECT  568200.0 1069200.0 578400.0 1083000.0 ;
      RECT  568200.0 1096800.0 578400.0 1083000.0 ;
      RECT  568200.0 1096800.0 578400.0 1110600.0 ;
      RECT  568200.0 1124400.0 578400.0 1110600.0 ;
      RECT  568200.0 1124400.0 578400.0 1138200.0 ;
      RECT  568200.0 1152000.0 578400.0 1138200.0 ;
      RECT  568200.0 1152000.0 578400.0 1165800.0 ;
      RECT  568200.0 1179600.0 578400.0 1165800.0 ;
      RECT  568200.0 1179600.0 578400.0 1193400.0 ;
      RECT  568200.0 1207200.0 578400.0 1193400.0 ;
      RECT  568200.0 1207200.0 578400.0 1221000.0 ;
      RECT  568200.0 1234800.0 578400.0 1221000.0 ;
      RECT  568200.0 1234800.0 578400.0 1248600.0 ;
      RECT  568200.0 1262400.0 578400.0 1248600.0 ;
      RECT  568200.0 1262400.0 578400.0 1276200.0 ;
      RECT  568200.0 1290000.0 578400.0 1276200.0 ;
      RECT  568200.0 1290000.0 578400.0 1303800.0 ;
      RECT  568200.0 1317600.0 578400.0 1303800.0 ;
      RECT  568200.0 1317600.0 578400.0 1331400.0 ;
      RECT  568200.0 1345200.0 578400.0 1331400.0 ;
      RECT  568200.0 1345200.0 578400.0 1359000.0 ;
      RECT  568200.0 1372800.0 578400.0 1359000.0 ;
      RECT  568200.0 1372800.0 578400.0 1386600.0 ;
      RECT  568200.0 1400400.0 578400.0 1386600.0 ;
      RECT  568200.0 1400400.0 578400.0 1414200.0 ;
      RECT  568200.0 1428000.0 578400.0 1414200.0 ;
      RECT  568200.0 1428000.0 578400.0 1441800.0 ;
      RECT  568200.0 1455600.0 578400.0 1441800.0 ;
      RECT  568200.0 1455600.0 578400.0 1469400.0 ;
      RECT  568200.0 1483200.0 578400.0 1469400.0 ;
      RECT  568200.0 1483200.0 578400.0 1497000.0 ;
      RECT  568200.0 1510800.0 578400.0 1497000.0 ;
      RECT  568200.0 1510800.0 578400.0 1524600.0 ;
      RECT  568200.0 1538400.0 578400.0 1524600.0 ;
      RECT  568200.0 1538400.0 578400.0 1552200.0 ;
      RECT  568200.0 1566000.0 578400.0 1552200.0 ;
      RECT  568200.0 1566000.0 578400.0 1579800.0 ;
      RECT  568200.0 1593600.0 578400.0 1579800.0 ;
      RECT  568200.0 1593600.0 578400.0 1607400.0 ;
      RECT  568200.0 1621200.0 578400.0 1607400.0 ;
      RECT  568200.0 1621200.0 578400.0 1635000.0 ;
      RECT  568200.0 1648800.0 578400.0 1635000.0 ;
      RECT  568200.0 1648800.0 578400.0 1662600.0 ;
      RECT  568200.0 1676400.0 578400.0 1662600.0 ;
      RECT  568200.0 1676400.0 578400.0 1690200.0 ;
      RECT  568200.0 1704000.0 578400.0 1690200.0 ;
      RECT  568200.0 1704000.0 578400.0 1717800.0 ;
      RECT  568200.0 1731600.0 578400.0 1717800.0 ;
      RECT  568200.0 1731600.0 578400.0 1745400.0 ;
      RECT  568200.0 1759200.0 578400.0 1745400.0 ;
      RECT  568200.0 1759200.0 578400.0 1773000.0 ;
      RECT  568200.0 1786800.0 578400.0 1773000.0 ;
      RECT  568200.0 1786800.0 578400.0 1800600.0 ;
      RECT  568200.0 1814400.0 578400.0 1800600.0 ;
      RECT  568200.0 1814400.0 578400.0 1828200.0 ;
      RECT  568200.0 1842000.0 578400.0 1828200.0 ;
      RECT  568200.0 1842000.0 578400.0 1855800.0 ;
      RECT  568200.0 1869600.0 578400.0 1855800.0 ;
      RECT  568200.0 1869600.0 578400.0 1883400.0 ;
      RECT  568200.0 1897200.0 578400.0 1883400.0 ;
      RECT  568200.0 1897200.0 578400.0 1911000.0 ;
      RECT  568200.0 1924800.0 578400.0 1911000.0 ;
      RECT  568200.0 1924800.0 578400.0 1938600.0 ;
      RECT  568200.0 1952400.0 578400.0 1938600.0 ;
      RECT  568200.0 1952400.0 578400.0 1966200.0 ;
      RECT  568200.0 1980000.0 578400.0 1966200.0 ;
      RECT  568200.0 1980000.0 578400.0 1993800.0 ;
      RECT  568200.0 2007600.0 578400.0 1993800.0 ;
      RECT  568200.0 2007600.0 578400.0 2021400.0 ;
      RECT  568200.0 2035200.0 578400.0 2021400.0 ;
      RECT  568200.0 2035200.0 578400.0 2049000.0 ;
      RECT  568200.0 2062800.0 578400.0 2049000.0 ;
      RECT  568200.0 2062800.0 578400.0 2076600.0 ;
      RECT  568200.0 2090400.0 578400.0 2076600.0 ;
      RECT  568200.0 2090400.0 578400.0 2104200.0 ;
      RECT  568200.0 2118000.0 578400.0 2104200.0 ;
      RECT  568200.0 2118000.0 578400.0 2131800.0 ;
      RECT  568200.0 2145600.0 578400.0 2131800.0 ;
      RECT  578400.0 379200.0 588600.0 393000.0 ;
      RECT  578400.0 406800.0 588600.0 393000.0 ;
      RECT  578400.0 406800.0 588600.0 420600.0 ;
      RECT  578400.0 434400.0 588600.0 420600.0 ;
      RECT  578400.0 434400.0 588600.0 448200.0 ;
      RECT  578400.0 462000.0 588600.0 448200.0 ;
      RECT  578400.0 462000.0 588600.0 475800.0 ;
      RECT  578400.0 489600.0 588600.0 475800.0 ;
      RECT  578400.0 489600.0 588600.0 503400.0 ;
      RECT  578400.0 517200.0 588600.0 503400.0 ;
      RECT  578400.0 517200.0 588600.0 531000.0 ;
      RECT  578400.0 544800.0 588600.0 531000.0 ;
      RECT  578400.0 544800.0 588600.0 558600.0 ;
      RECT  578400.0 572400.0 588600.0 558600.0 ;
      RECT  578400.0 572400.0 588600.0 586200.0 ;
      RECT  578400.0 600000.0 588600.0 586200.0 ;
      RECT  578400.0 600000.0 588600.0 613800.0 ;
      RECT  578400.0 627600.0 588600.0 613800.0 ;
      RECT  578400.0 627600.0 588600.0 641400.0 ;
      RECT  578400.0 655200.0 588600.0 641400.0 ;
      RECT  578400.0 655200.0 588600.0 669000.0 ;
      RECT  578400.0 682800.0 588600.0 669000.0 ;
      RECT  578400.0 682800.0 588600.0 696600.0 ;
      RECT  578400.0 710400.0 588600.0 696600.0 ;
      RECT  578400.0 710400.0 588600.0 724200.0 ;
      RECT  578400.0 738000.0 588600.0 724200.0 ;
      RECT  578400.0 738000.0 588600.0 751800.0 ;
      RECT  578400.0 765600.0 588600.0 751800.0 ;
      RECT  578400.0 765600.0 588600.0 779400.0 ;
      RECT  578400.0 793200.0 588600.0 779400.0 ;
      RECT  578400.0 793200.0 588600.0 807000.0 ;
      RECT  578400.0 820800.0 588600.0 807000.0 ;
      RECT  578400.0 820800.0 588600.0 834600.0 ;
      RECT  578400.0 848400.0 588600.0 834600.0 ;
      RECT  578400.0 848400.0 588600.0 862200.0 ;
      RECT  578400.0 876000.0 588600.0 862200.0 ;
      RECT  578400.0 876000.0 588600.0 889800.0 ;
      RECT  578400.0 903600.0 588600.0 889800.0 ;
      RECT  578400.0 903600.0 588600.0 917400.0 ;
      RECT  578400.0 931200.0 588600.0 917400.0 ;
      RECT  578400.0 931200.0 588600.0 945000.0 ;
      RECT  578400.0 958800.0 588600.0 945000.0 ;
      RECT  578400.0 958800.0 588600.0 972600.0 ;
      RECT  578400.0 986400.0 588600.0 972600.0 ;
      RECT  578400.0 986400.0 588600.0 1000200.0 ;
      RECT  578400.0 1014000.0 588600.0 1000200.0 ;
      RECT  578400.0 1014000.0 588600.0 1027800.0 ;
      RECT  578400.0 1041600.0 588600.0 1027800.0 ;
      RECT  578400.0 1041600.0 588600.0 1055400.0 ;
      RECT  578400.0 1069200.0 588600.0 1055400.0 ;
      RECT  578400.0 1069200.0 588600.0 1083000.0 ;
      RECT  578400.0 1096800.0 588600.0 1083000.0 ;
      RECT  578400.0 1096800.0 588600.0 1110600.0 ;
      RECT  578400.0 1124400.0 588600.0 1110600.0 ;
      RECT  578400.0 1124400.0 588600.0 1138200.0 ;
      RECT  578400.0 1152000.0 588600.0 1138200.0 ;
      RECT  578400.0 1152000.0 588600.0 1165800.0 ;
      RECT  578400.0 1179600.0 588600.0 1165800.0 ;
      RECT  578400.0 1179600.0 588600.0 1193400.0 ;
      RECT  578400.0 1207200.0 588600.0 1193400.0 ;
      RECT  578400.0 1207200.0 588600.0 1221000.0 ;
      RECT  578400.0 1234800.0 588600.0 1221000.0 ;
      RECT  578400.0 1234800.0 588600.0 1248600.0 ;
      RECT  578400.0 1262400.0 588600.0 1248600.0 ;
      RECT  578400.0 1262400.0 588600.0 1276200.0 ;
      RECT  578400.0 1290000.0 588600.0 1276200.0 ;
      RECT  578400.0 1290000.0 588600.0 1303800.0 ;
      RECT  578400.0 1317600.0 588600.0 1303800.0 ;
      RECT  578400.0 1317600.0 588600.0 1331400.0 ;
      RECT  578400.0 1345200.0 588600.0 1331400.0 ;
      RECT  578400.0 1345200.0 588600.0 1359000.0 ;
      RECT  578400.0 1372800.0 588600.0 1359000.0 ;
      RECT  578400.0 1372800.0 588600.0 1386600.0 ;
      RECT  578400.0 1400400.0 588600.0 1386600.0 ;
      RECT  578400.0 1400400.0 588600.0 1414200.0 ;
      RECT  578400.0 1428000.0 588600.0 1414200.0 ;
      RECT  578400.0 1428000.0 588600.0 1441800.0 ;
      RECT  578400.0 1455600.0 588600.0 1441800.0 ;
      RECT  578400.0 1455600.0 588600.0 1469400.0 ;
      RECT  578400.0 1483200.0 588600.0 1469400.0 ;
      RECT  578400.0 1483200.0 588600.0 1497000.0 ;
      RECT  578400.0 1510800.0 588600.0 1497000.0 ;
      RECT  578400.0 1510800.0 588600.0 1524600.0 ;
      RECT  578400.0 1538400.0 588600.0 1524600.0 ;
      RECT  578400.0 1538400.0 588600.0 1552200.0 ;
      RECT  578400.0 1566000.0 588600.0 1552200.0 ;
      RECT  578400.0 1566000.0 588600.0 1579800.0 ;
      RECT  578400.0 1593600.0 588600.0 1579800.0 ;
      RECT  578400.0 1593600.0 588600.0 1607400.0 ;
      RECT  578400.0 1621200.0 588600.0 1607400.0 ;
      RECT  578400.0 1621200.0 588600.0 1635000.0 ;
      RECT  578400.0 1648800.0 588600.0 1635000.0 ;
      RECT  578400.0 1648800.0 588600.0 1662600.0 ;
      RECT  578400.0 1676400.0 588600.0 1662600.0 ;
      RECT  578400.0 1676400.0 588600.0 1690200.0 ;
      RECT  578400.0 1704000.0 588600.0 1690200.0 ;
      RECT  578400.0 1704000.0 588600.0 1717800.0 ;
      RECT  578400.0 1731600.0 588600.0 1717800.0 ;
      RECT  578400.0 1731600.0 588600.0 1745400.0 ;
      RECT  578400.0 1759200.0 588600.0 1745400.0 ;
      RECT  578400.0 1759200.0 588600.0 1773000.0 ;
      RECT  578400.0 1786800.0 588600.0 1773000.0 ;
      RECT  578400.0 1786800.0 588600.0 1800600.0 ;
      RECT  578400.0 1814400.0 588600.0 1800600.0 ;
      RECT  578400.0 1814400.0 588600.0 1828200.0 ;
      RECT  578400.0 1842000.0 588600.0 1828200.0 ;
      RECT  578400.0 1842000.0 588600.0 1855800.0 ;
      RECT  578400.0 1869600.0 588600.0 1855800.0 ;
      RECT  578400.0 1869600.0 588600.0 1883400.0 ;
      RECT  578400.0 1897200.0 588600.0 1883400.0 ;
      RECT  578400.0 1897200.0 588600.0 1911000.0 ;
      RECT  578400.0 1924800.0 588600.0 1911000.0 ;
      RECT  578400.0 1924800.0 588600.0 1938600.0 ;
      RECT  578400.0 1952400.0 588600.0 1938600.0 ;
      RECT  578400.0 1952400.0 588600.0 1966200.0 ;
      RECT  578400.0 1980000.0 588600.0 1966200.0 ;
      RECT  578400.0 1980000.0 588600.0 1993800.0 ;
      RECT  578400.0 2007600.0 588600.0 1993800.0 ;
      RECT  578400.0 2007600.0 588600.0 2021400.0 ;
      RECT  578400.0 2035200.0 588600.0 2021400.0 ;
      RECT  578400.0 2035200.0 588600.0 2049000.0 ;
      RECT  578400.0 2062800.0 588600.0 2049000.0 ;
      RECT  578400.0 2062800.0 588600.0 2076600.0 ;
      RECT  578400.0 2090400.0 588600.0 2076600.0 ;
      RECT  578400.0 2090400.0 588600.0 2104200.0 ;
      RECT  578400.0 2118000.0 588600.0 2104200.0 ;
      RECT  578400.0 2118000.0 588600.0 2131800.0 ;
      RECT  578400.0 2145600.0 588600.0 2131800.0 ;
      RECT  588600.0 379200.0 598800.0 393000.0 ;
      RECT  588600.0 406800.0 598800.0 393000.0 ;
      RECT  588600.0 406800.0 598800.0 420600.0 ;
      RECT  588600.0 434400.0 598800.0 420600.0 ;
      RECT  588600.0 434400.0 598800.0 448200.0 ;
      RECT  588600.0 462000.0 598800.0 448200.0 ;
      RECT  588600.0 462000.0 598800.0 475800.0 ;
      RECT  588600.0 489600.0 598800.0 475800.0 ;
      RECT  588600.0 489600.0 598800.0 503400.0 ;
      RECT  588600.0 517200.0 598800.0 503400.0 ;
      RECT  588600.0 517200.0 598800.0 531000.0 ;
      RECT  588600.0 544800.0 598800.0 531000.0 ;
      RECT  588600.0 544800.0 598800.0 558600.0 ;
      RECT  588600.0 572400.0 598800.0 558600.0 ;
      RECT  588600.0 572400.0 598800.0 586200.0 ;
      RECT  588600.0 600000.0 598800.0 586200.0 ;
      RECT  588600.0 600000.0 598800.0 613800.0 ;
      RECT  588600.0 627600.0 598800.0 613800.0 ;
      RECT  588600.0 627600.0 598800.0 641400.0 ;
      RECT  588600.0 655200.0 598800.0 641400.0 ;
      RECT  588600.0 655200.0 598800.0 669000.0 ;
      RECT  588600.0 682800.0 598800.0 669000.0 ;
      RECT  588600.0 682800.0 598800.0 696600.0 ;
      RECT  588600.0 710400.0 598800.0 696600.0 ;
      RECT  588600.0 710400.0 598800.0 724200.0 ;
      RECT  588600.0 738000.0 598800.0 724200.0 ;
      RECT  588600.0 738000.0 598800.0 751800.0 ;
      RECT  588600.0 765600.0 598800.0 751800.0 ;
      RECT  588600.0 765600.0 598800.0 779400.0 ;
      RECT  588600.0 793200.0 598800.0 779400.0 ;
      RECT  588600.0 793200.0 598800.0 807000.0 ;
      RECT  588600.0 820800.0 598800.0 807000.0 ;
      RECT  588600.0 820800.0 598800.0 834600.0 ;
      RECT  588600.0 848400.0 598800.0 834600.0 ;
      RECT  588600.0 848400.0 598800.0 862200.0 ;
      RECT  588600.0 876000.0 598800.0 862200.0 ;
      RECT  588600.0 876000.0 598800.0 889800.0 ;
      RECT  588600.0 903600.0 598800.0 889800.0 ;
      RECT  588600.0 903600.0 598800.0 917400.0 ;
      RECT  588600.0 931200.0 598800.0 917400.0 ;
      RECT  588600.0 931200.0 598800.0 945000.0 ;
      RECT  588600.0 958800.0 598800.0 945000.0 ;
      RECT  588600.0 958800.0 598800.0 972600.0 ;
      RECT  588600.0 986400.0 598800.0 972600.0 ;
      RECT  588600.0 986400.0 598800.0 1000200.0 ;
      RECT  588600.0 1014000.0 598800.0 1000200.0 ;
      RECT  588600.0 1014000.0 598800.0 1027800.0 ;
      RECT  588600.0 1041600.0 598800.0 1027800.0 ;
      RECT  588600.0 1041600.0 598800.0 1055400.0 ;
      RECT  588600.0 1069200.0 598800.0 1055400.0 ;
      RECT  588600.0 1069200.0 598800.0 1083000.0 ;
      RECT  588600.0 1096800.0 598800.0 1083000.0 ;
      RECT  588600.0 1096800.0 598800.0 1110600.0 ;
      RECT  588600.0 1124400.0 598800.0 1110600.0 ;
      RECT  588600.0 1124400.0 598800.0 1138200.0 ;
      RECT  588600.0 1152000.0 598800.0 1138200.0 ;
      RECT  588600.0 1152000.0 598800.0 1165800.0 ;
      RECT  588600.0 1179600.0 598800.0 1165800.0 ;
      RECT  588600.0 1179600.0 598800.0 1193400.0 ;
      RECT  588600.0 1207200.0 598800.0 1193400.0 ;
      RECT  588600.0 1207200.0 598800.0 1221000.0 ;
      RECT  588600.0 1234800.0 598800.0 1221000.0 ;
      RECT  588600.0 1234800.0 598800.0 1248600.0 ;
      RECT  588600.0 1262400.0 598800.0 1248600.0 ;
      RECT  588600.0 1262400.0 598800.0 1276200.0 ;
      RECT  588600.0 1290000.0 598800.0 1276200.0 ;
      RECT  588600.0 1290000.0 598800.0 1303800.0 ;
      RECT  588600.0 1317600.0 598800.0 1303800.0 ;
      RECT  588600.0 1317600.0 598800.0 1331400.0 ;
      RECT  588600.0 1345200.0 598800.0 1331400.0 ;
      RECT  588600.0 1345200.0 598800.0 1359000.0 ;
      RECT  588600.0 1372800.0 598800.0 1359000.0 ;
      RECT  588600.0 1372800.0 598800.0 1386600.0 ;
      RECT  588600.0 1400400.0 598800.0 1386600.0 ;
      RECT  588600.0 1400400.0 598800.0 1414200.0 ;
      RECT  588600.0 1428000.0 598800.0 1414200.0 ;
      RECT  588600.0 1428000.0 598800.0 1441800.0 ;
      RECT  588600.0 1455600.0 598800.0 1441800.0 ;
      RECT  588600.0 1455600.0 598800.0 1469400.0 ;
      RECT  588600.0 1483200.0 598800.0 1469400.0 ;
      RECT  588600.0 1483200.0 598800.0 1497000.0 ;
      RECT  588600.0 1510800.0 598800.0 1497000.0 ;
      RECT  588600.0 1510800.0 598800.0 1524600.0 ;
      RECT  588600.0 1538400.0 598800.0 1524600.0 ;
      RECT  588600.0 1538400.0 598800.0 1552200.0 ;
      RECT  588600.0 1566000.0 598800.0 1552200.0 ;
      RECT  588600.0 1566000.0 598800.0 1579800.0 ;
      RECT  588600.0 1593600.0 598800.0 1579800.0 ;
      RECT  588600.0 1593600.0 598800.0 1607400.0 ;
      RECT  588600.0 1621200.0 598800.0 1607400.0 ;
      RECT  588600.0 1621200.0 598800.0 1635000.0 ;
      RECT  588600.0 1648800.0 598800.0 1635000.0 ;
      RECT  588600.0 1648800.0 598800.0 1662600.0 ;
      RECT  588600.0 1676400.0 598800.0 1662600.0 ;
      RECT  588600.0 1676400.0 598800.0 1690200.0 ;
      RECT  588600.0 1704000.0 598800.0 1690200.0 ;
      RECT  588600.0 1704000.0 598800.0 1717800.0 ;
      RECT  588600.0 1731600.0 598800.0 1717800.0 ;
      RECT  588600.0 1731600.0 598800.0 1745400.0 ;
      RECT  588600.0 1759200.0 598800.0 1745400.0 ;
      RECT  588600.0 1759200.0 598800.0 1773000.0 ;
      RECT  588600.0 1786800.0 598800.0 1773000.0 ;
      RECT  588600.0 1786800.0 598800.0 1800600.0 ;
      RECT  588600.0 1814400.0 598800.0 1800600.0 ;
      RECT  588600.0 1814400.0 598800.0 1828200.0 ;
      RECT  588600.0 1842000.0 598800.0 1828200.0 ;
      RECT  588600.0 1842000.0 598800.0 1855800.0 ;
      RECT  588600.0 1869600.0 598800.0 1855800.0 ;
      RECT  588600.0 1869600.0 598800.0 1883400.0 ;
      RECT  588600.0 1897200.0 598800.0 1883400.0 ;
      RECT  588600.0 1897200.0 598800.0 1911000.0 ;
      RECT  588600.0 1924800.0 598800.0 1911000.0 ;
      RECT  588600.0 1924800.0 598800.0 1938600.0 ;
      RECT  588600.0 1952400.0 598800.0 1938600.0 ;
      RECT  588600.0 1952400.0 598800.0 1966200.0 ;
      RECT  588600.0 1980000.0 598800.0 1966200.0 ;
      RECT  588600.0 1980000.0 598800.0 1993800.0 ;
      RECT  588600.0 2007600.0 598800.0 1993800.0 ;
      RECT  588600.0 2007600.0 598800.0 2021400.0 ;
      RECT  588600.0 2035200.0 598800.0 2021400.0 ;
      RECT  588600.0 2035200.0 598800.0 2049000.0 ;
      RECT  588600.0 2062800.0 598800.0 2049000.0 ;
      RECT  588600.0 2062800.0 598800.0 2076600.0 ;
      RECT  588600.0 2090400.0 598800.0 2076600.0 ;
      RECT  588600.0 2090400.0 598800.0 2104200.0 ;
      RECT  588600.0 2118000.0 598800.0 2104200.0 ;
      RECT  588600.0 2118000.0 598800.0 2131800.0 ;
      RECT  588600.0 2145600.0 598800.0 2131800.0 ;
      RECT  598800.0 379200.0 609000.0 393000.0 ;
      RECT  598800.0 406800.0 609000.0 393000.0 ;
      RECT  598800.0 406800.0 609000.0 420600.0 ;
      RECT  598800.0 434400.0 609000.0 420600.0 ;
      RECT  598800.0 434400.0 609000.0 448200.0 ;
      RECT  598800.0 462000.0 609000.0 448200.0 ;
      RECT  598800.0 462000.0 609000.0 475800.0 ;
      RECT  598800.0 489600.0 609000.0 475800.0 ;
      RECT  598800.0 489600.0 609000.0 503400.0 ;
      RECT  598800.0 517200.0 609000.0 503400.0 ;
      RECT  598800.0 517200.0 609000.0 531000.0 ;
      RECT  598800.0 544800.0 609000.0 531000.0 ;
      RECT  598800.0 544800.0 609000.0 558600.0 ;
      RECT  598800.0 572400.0 609000.0 558600.0 ;
      RECT  598800.0 572400.0 609000.0 586200.0 ;
      RECT  598800.0 600000.0 609000.0 586200.0 ;
      RECT  598800.0 600000.0 609000.0 613800.0 ;
      RECT  598800.0 627600.0 609000.0 613800.0 ;
      RECT  598800.0 627600.0 609000.0 641400.0 ;
      RECT  598800.0 655200.0 609000.0 641400.0 ;
      RECT  598800.0 655200.0 609000.0 669000.0 ;
      RECT  598800.0 682800.0 609000.0 669000.0 ;
      RECT  598800.0 682800.0 609000.0 696600.0 ;
      RECT  598800.0 710400.0 609000.0 696600.0 ;
      RECT  598800.0 710400.0 609000.0 724200.0 ;
      RECT  598800.0 738000.0 609000.0 724200.0 ;
      RECT  598800.0 738000.0 609000.0 751800.0 ;
      RECT  598800.0 765600.0 609000.0 751800.0 ;
      RECT  598800.0 765600.0 609000.0 779400.0 ;
      RECT  598800.0 793200.0 609000.0 779400.0 ;
      RECT  598800.0 793200.0 609000.0 807000.0 ;
      RECT  598800.0 820800.0 609000.0 807000.0 ;
      RECT  598800.0 820800.0 609000.0 834600.0 ;
      RECT  598800.0 848400.0 609000.0 834600.0 ;
      RECT  598800.0 848400.0 609000.0 862200.0 ;
      RECT  598800.0 876000.0 609000.0 862200.0 ;
      RECT  598800.0 876000.0 609000.0 889800.0 ;
      RECT  598800.0 903600.0 609000.0 889800.0 ;
      RECT  598800.0 903600.0 609000.0 917400.0 ;
      RECT  598800.0 931200.0 609000.0 917400.0 ;
      RECT  598800.0 931200.0 609000.0 945000.0 ;
      RECT  598800.0 958800.0 609000.0 945000.0 ;
      RECT  598800.0 958800.0 609000.0 972600.0 ;
      RECT  598800.0 986400.0 609000.0 972600.0 ;
      RECT  598800.0 986400.0 609000.0 1000200.0 ;
      RECT  598800.0 1014000.0 609000.0 1000200.0 ;
      RECT  598800.0 1014000.0 609000.0 1027800.0 ;
      RECT  598800.0 1041600.0 609000.0 1027800.0 ;
      RECT  598800.0 1041600.0 609000.0 1055400.0 ;
      RECT  598800.0 1069200.0 609000.0 1055400.0 ;
      RECT  598800.0 1069200.0 609000.0 1083000.0 ;
      RECT  598800.0 1096800.0 609000.0 1083000.0 ;
      RECT  598800.0 1096800.0 609000.0 1110600.0 ;
      RECT  598800.0 1124400.0 609000.0 1110600.0 ;
      RECT  598800.0 1124400.0 609000.0 1138200.0 ;
      RECT  598800.0 1152000.0 609000.0 1138200.0 ;
      RECT  598800.0 1152000.0 609000.0 1165800.0 ;
      RECT  598800.0 1179600.0 609000.0 1165800.0 ;
      RECT  598800.0 1179600.0 609000.0 1193400.0 ;
      RECT  598800.0 1207200.0 609000.0 1193400.0 ;
      RECT  598800.0 1207200.0 609000.0 1221000.0 ;
      RECT  598800.0 1234800.0 609000.0 1221000.0 ;
      RECT  598800.0 1234800.0 609000.0 1248600.0 ;
      RECT  598800.0 1262400.0 609000.0 1248600.0 ;
      RECT  598800.0 1262400.0 609000.0 1276200.0 ;
      RECT  598800.0 1290000.0 609000.0 1276200.0 ;
      RECT  598800.0 1290000.0 609000.0 1303800.0 ;
      RECT  598800.0 1317600.0 609000.0 1303800.0 ;
      RECT  598800.0 1317600.0 609000.0 1331400.0 ;
      RECT  598800.0 1345200.0 609000.0 1331400.0 ;
      RECT  598800.0 1345200.0 609000.0 1359000.0 ;
      RECT  598800.0 1372800.0 609000.0 1359000.0 ;
      RECT  598800.0 1372800.0 609000.0 1386600.0 ;
      RECT  598800.0 1400400.0 609000.0 1386600.0 ;
      RECT  598800.0 1400400.0 609000.0 1414200.0 ;
      RECT  598800.0 1428000.0 609000.0 1414200.0 ;
      RECT  598800.0 1428000.0 609000.0 1441800.0 ;
      RECT  598800.0 1455600.0 609000.0 1441800.0 ;
      RECT  598800.0 1455600.0 609000.0 1469400.0 ;
      RECT  598800.0 1483200.0 609000.0 1469400.0 ;
      RECT  598800.0 1483200.0 609000.0 1497000.0 ;
      RECT  598800.0 1510800.0 609000.0 1497000.0 ;
      RECT  598800.0 1510800.0 609000.0 1524600.0 ;
      RECT  598800.0 1538400.0 609000.0 1524600.0 ;
      RECT  598800.0 1538400.0 609000.0 1552200.0 ;
      RECT  598800.0 1566000.0 609000.0 1552200.0 ;
      RECT  598800.0 1566000.0 609000.0 1579800.0 ;
      RECT  598800.0 1593600.0 609000.0 1579800.0 ;
      RECT  598800.0 1593600.0 609000.0 1607400.0 ;
      RECT  598800.0 1621200.0 609000.0 1607400.0 ;
      RECT  598800.0 1621200.0 609000.0 1635000.0 ;
      RECT  598800.0 1648800.0 609000.0 1635000.0 ;
      RECT  598800.0 1648800.0 609000.0 1662600.0 ;
      RECT  598800.0 1676400.0 609000.0 1662600.0 ;
      RECT  598800.0 1676400.0 609000.0 1690200.0 ;
      RECT  598800.0 1704000.0 609000.0 1690200.0 ;
      RECT  598800.0 1704000.0 609000.0 1717800.0 ;
      RECT  598800.0 1731600.0 609000.0 1717800.0 ;
      RECT  598800.0 1731600.0 609000.0 1745400.0 ;
      RECT  598800.0 1759200.0 609000.0 1745400.0 ;
      RECT  598800.0 1759200.0 609000.0 1773000.0 ;
      RECT  598800.0 1786800.0 609000.0 1773000.0 ;
      RECT  598800.0 1786800.0 609000.0 1800600.0 ;
      RECT  598800.0 1814400.0 609000.0 1800600.0 ;
      RECT  598800.0 1814400.0 609000.0 1828200.0 ;
      RECT  598800.0 1842000.0 609000.0 1828200.0 ;
      RECT  598800.0 1842000.0 609000.0 1855800.0 ;
      RECT  598800.0 1869600.0 609000.0 1855800.0 ;
      RECT  598800.0 1869600.0 609000.0 1883400.0 ;
      RECT  598800.0 1897200.0 609000.0 1883400.0 ;
      RECT  598800.0 1897200.0 609000.0 1911000.0 ;
      RECT  598800.0 1924800.0 609000.0 1911000.0 ;
      RECT  598800.0 1924800.0 609000.0 1938600.0 ;
      RECT  598800.0 1952400.0 609000.0 1938600.0 ;
      RECT  598800.0 1952400.0 609000.0 1966200.0 ;
      RECT  598800.0 1980000.0 609000.0 1966200.0 ;
      RECT  598800.0 1980000.0 609000.0 1993800.0 ;
      RECT  598800.0 2007600.0 609000.0 1993800.0 ;
      RECT  598800.0 2007600.0 609000.0 2021400.0 ;
      RECT  598800.0 2035200.0 609000.0 2021400.0 ;
      RECT  598800.0 2035200.0 609000.0 2049000.0 ;
      RECT  598800.0 2062800.0 609000.0 2049000.0 ;
      RECT  598800.0 2062800.0 609000.0 2076600.0 ;
      RECT  598800.0 2090400.0 609000.0 2076600.0 ;
      RECT  598800.0 2090400.0 609000.0 2104200.0 ;
      RECT  598800.0 2118000.0 609000.0 2104200.0 ;
      RECT  598800.0 2118000.0 609000.0 2131800.0 ;
      RECT  598800.0 2145600.0 609000.0 2131800.0 ;
      RECT  609000.0 379200.0 619200.0 393000.0 ;
      RECT  609000.0 406800.0 619200.0 393000.0 ;
      RECT  609000.0 406800.0 619200.0 420600.0 ;
      RECT  609000.0 434400.0 619200.0 420600.0 ;
      RECT  609000.0 434400.0 619200.0 448200.0 ;
      RECT  609000.0 462000.0 619200.0 448200.0 ;
      RECT  609000.0 462000.0 619200.0 475800.0 ;
      RECT  609000.0 489600.0 619200.0 475800.0 ;
      RECT  609000.0 489600.0 619200.0 503400.0 ;
      RECT  609000.0 517200.0 619200.0 503400.0 ;
      RECT  609000.0 517200.0 619200.0 531000.0 ;
      RECT  609000.0 544800.0 619200.0 531000.0 ;
      RECT  609000.0 544800.0 619200.0 558600.0 ;
      RECT  609000.0 572400.0 619200.0 558600.0 ;
      RECT  609000.0 572400.0 619200.0 586200.0 ;
      RECT  609000.0 600000.0 619200.0 586200.0 ;
      RECT  609000.0 600000.0 619200.0 613800.0 ;
      RECT  609000.0 627600.0 619200.0 613800.0 ;
      RECT  609000.0 627600.0 619200.0 641400.0 ;
      RECT  609000.0 655200.0 619200.0 641400.0 ;
      RECT  609000.0 655200.0 619200.0 669000.0 ;
      RECT  609000.0 682800.0 619200.0 669000.0 ;
      RECT  609000.0 682800.0 619200.0 696600.0 ;
      RECT  609000.0 710400.0 619200.0 696600.0 ;
      RECT  609000.0 710400.0 619200.0 724200.0 ;
      RECT  609000.0 738000.0 619200.0 724200.0 ;
      RECT  609000.0 738000.0 619200.0 751800.0 ;
      RECT  609000.0 765600.0 619200.0 751800.0 ;
      RECT  609000.0 765600.0 619200.0 779400.0 ;
      RECT  609000.0 793200.0 619200.0 779400.0 ;
      RECT  609000.0 793200.0 619200.0 807000.0 ;
      RECT  609000.0 820800.0 619200.0 807000.0 ;
      RECT  609000.0 820800.0 619200.0 834600.0 ;
      RECT  609000.0 848400.0 619200.0 834600.0 ;
      RECT  609000.0 848400.0 619200.0 862200.0 ;
      RECT  609000.0 876000.0 619200.0 862200.0 ;
      RECT  609000.0 876000.0 619200.0 889800.0 ;
      RECT  609000.0 903600.0 619200.0 889800.0 ;
      RECT  609000.0 903600.0 619200.0 917400.0 ;
      RECT  609000.0 931200.0 619200.0 917400.0 ;
      RECT  609000.0 931200.0 619200.0 945000.0 ;
      RECT  609000.0 958800.0 619200.0 945000.0 ;
      RECT  609000.0 958800.0 619200.0 972600.0 ;
      RECT  609000.0 986400.0 619200.0 972600.0 ;
      RECT  609000.0 986400.0 619200.0 1000200.0 ;
      RECT  609000.0 1014000.0 619200.0 1000200.0 ;
      RECT  609000.0 1014000.0 619200.0 1027800.0 ;
      RECT  609000.0 1041600.0 619200.0 1027800.0 ;
      RECT  609000.0 1041600.0 619200.0 1055400.0 ;
      RECT  609000.0 1069200.0 619200.0 1055400.0 ;
      RECT  609000.0 1069200.0 619200.0 1083000.0 ;
      RECT  609000.0 1096800.0 619200.0 1083000.0 ;
      RECT  609000.0 1096800.0 619200.0 1110600.0 ;
      RECT  609000.0 1124400.0 619200.0 1110600.0 ;
      RECT  609000.0 1124400.0 619200.0 1138200.0 ;
      RECT  609000.0 1152000.0 619200.0 1138200.0 ;
      RECT  609000.0 1152000.0 619200.0 1165800.0 ;
      RECT  609000.0 1179600.0 619200.0 1165800.0 ;
      RECT  609000.0 1179600.0 619200.0 1193400.0 ;
      RECT  609000.0 1207200.0 619200.0 1193400.0 ;
      RECT  609000.0 1207200.0 619200.0 1221000.0 ;
      RECT  609000.0 1234800.0 619200.0 1221000.0 ;
      RECT  609000.0 1234800.0 619200.0 1248600.0 ;
      RECT  609000.0 1262400.0 619200.0 1248600.0 ;
      RECT  609000.0 1262400.0 619200.0 1276200.0 ;
      RECT  609000.0 1290000.0 619200.0 1276200.0 ;
      RECT  609000.0 1290000.0 619200.0 1303800.0 ;
      RECT  609000.0 1317600.0 619200.0 1303800.0 ;
      RECT  609000.0 1317600.0 619200.0 1331400.0 ;
      RECT  609000.0 1345200.0 619200.0 1331400.0 ;
      RECT  609000.0 1345200.0 619200.0 1359000.0 ;
      RECT  609000.0 1372800.0 619200.0 1359000.0 ;
      RECT  609000.0 1372800.0 619200.0 1386600.0 ;
      RECT  609000.0 1400400.0 619200.0 1386600.0 ;
      RECT  609000.0 1400400.0 619200.0 1414200.0 ;
      RECT  609000.0 1428000.0 619200.0 1414200.0 ;
      RECT  609000.0 1428000.0 619200.0 1441800.0 ;
      RECT  609000.0 1455600.0 619200.0 1441800.0 ;
      RECT  609000.0 1455600.0 619200.0 1469400.0 ;
      RECT  609000.0 1483200.0 619200.0 1469400.0 ;
      RECT  609000.0 1483200.0 619200.0 1497000.0 ;
      RECT  609000.0 1510800.0 619200.0 1497000.0 ;
      RECT  609000.0 1510800.0 619200.0 1524600.0 ;
      RECT  609000.0 1538400.0 619200.0 1524600.0 ;
      RECT  609000.0 1538400.0 619200.0 1552200.0 ;
      RECT  609000.0 1566000.0 619200.0 1552200.0 ;
      RECT  609000.0 1566000.0 619200.0 1579800.0 ;
      RECT  609000.0 1593600.0 619200.0 1579800.0 ;
      RECT  609000.0 1593600.0 619200.0 1607400.0 ;
      RECT  609000.0 1621200.0 619200.0 1607400.0 ;
      RECT  609000.0 1621200.0 619200.0 1635000.0 ;
      RECT  609000.0 1648800.0 619200.0 1635000.0 ;
      RECT  609000.0 1648800.0 619200.0 1662600.0 ;
      RECT  609000.0 1676400.0 619200.0 1662600.0 ;
      RECT  609000.0 1676400.0 619200.0 1690200.0 ;
      RECT  609000.0 1704000.0 619200.0 1690200.0 ;
      RECT  609000.0 1704000.0 619200.0 1717800.0 ;
      RECT  609000.0 1731600.0 619200.0 1717800.0 ;
      RECT  609000.0 1731600.0 619200.0 1745400.0 ;
      RECT  609000.0 1759200.0 619200.0 1745400.0 ;
      RECT  609000.0 1759200.0 619200.0 1773000.0 ;
      RECT  609000.0 1786800.0 619200.0 1773000.0 ;
      RECT  609000.0 1786800.0 619200.0 1800600.0 ;
      RECT  609000.0 1814400.0 619200.0 1800600.0 ;
      RECT  609000.0 1814400.0 619200.0 1828200.0 ;
      RECT  609000.0 1842000.0 619200.0 1828200.0 ;
      RECT  609000.0 1842000.0 619200.0 1855800.0 ;
      RECT  609000.0 1869600.0 619200.0 1855800.0 ;
      RECT  609000.0 1869600.0 619200.0 1883400.0 ;
      RECT  609000.0 1897200.0 619200.0 1883400.0 ;
      RECT  609000.0 1897200.0 619200.0 1911000.0 ;
      RECT  609000.0 1924800.0 619200.0 1911000.0 ;
      RECT  609000.0 1924800.0 619200.0 1938600.0 ;
      RECT  609000.0 1952400.0 619200.0 1938600.0 ;
      RECT  609000.0 1952400.0 619200.0 1966200.0 ;
      RECT  609000.0 1980000.0 619200.0 1966200.0 ;
      RECT  609000.0 1980000.0 619200.0 1993800.0 ;
      RECT  609000.0 2007600.0 619200.0 1993800.0 ;
      RECT  609000.0 2007600.0 619200.0 2021400.0 ;
      RECT  609000.0 2035200.0 619200.0 2021400.0 ;
      RECT  609000.0 2035200.0 619200.0 2049000.0 ;
      RECT  609000.0 2062800.0 619200.0 2049000.0 ;
      RECT  609000.0 2062800.0 619200.0 2076600.0 ;
      RECT  609000.0 2090400.0 619200.0 2076600.0 ;
      RECT  609000.0 2090400.0 619200.0 2104200.0 ;
      RECT  609000.0 2118000.0 619200.0 2104200.0 ;
      RECT  609000.0 2118000.0 619200.0 2131800.0 ;
      RECT  609000.0 2145600.0 619200.0 2131800.0 ;
      RECT  619200.0 379200.0 629400.0 393000.0 ;
      RECT  619200.0 406800.0 629400.0 393000.0 ;
      RECT  619200.0 406800.0 629400.0 420600.0 ;
      RECT  619200.0 434400.0 629400.0 420600.0 ;
      RECT  619200.0 434400.0 629400.0 448200.0 ;
      RECT  619200.0 462000.0 629400.0 448200.0 ;
      RECT  619200.0 462000.0 629400.0 475800.0 ;
      RECT  619200.0 489600.0 629400.0 475800.0 ;
      RECT  619200.0 489600.0 629400.0 503400.0 ;
      RECT  619200.0 517200.0 629400.0 503400.0 ;
      RECT  619200.0 517200.0 629400.0 531000.0 ;
      RECT  619200.0 544800.0 629400.0 531000.0 ;
      RECT  619200.0 544800.0 629400.0 558600.0 ;
      RECT  619200.0 572400.0 629400.0 558600.0 ;
      RECT  619200.0 572400.0 629400.0 586200.0 ;
      RECT  619200.0 600000.0 629400.0 586200.0 ;
      RECT  619200.0 600000.0 629400.0 613800.0 ;
      RECT  619200.0 627600.0 629400.0 613800.0 ;
      RECT  619200.0 627600.0 629400.0 641400.0 ;
      RECT  619200.0 655200.0 629400.0 641400.0 ;
      RECT  619200.0 655200.0 629400.0 669000.0 ;
      RECT  619200.0 682800.0 629400.0 669000.0 ;
      RECT  619200.0 682800.0 629400.0 696600.0 ;
      RECT  619200.0 710400.0 629400.0 696600.0 ;
      RECT  619200.0 710400.0 629400.0 724200.0 ;
      RECT  619200.0 738000.0 629400.0 724200.0 ;
      RECT  619200.0 738000.0 629400.0 751800.0 ;
      RECT  619200.0 765600.0 629400.0 751800.0 ;
      RECT  619200.0 765600.0 629400.0 779400.0 ;
      RECT  619200.0 793200.0 629400.0 779400.0 ;
      RECT  619200.0 793200.0 629400.0 807000.0 ;
      RECT  619200.0 820800.0 629400.0 807000.0 ;
      RECT  619200.0 820800.0 629400.0 834600.0 ;
      RECT  619200.0 848400.0 629400.0 834600.0 ;
      RECT  619200.0 848400.0 629400.0 862200.0 ;
      RECT  619200.0 876000.0 629400.0 862200.0 ;
      RECT  619200.0 876000.0 629400.0 889800.0 ;
      RECT  619200.0 903600.0 629400.0 889800.0 ;
      RECT  619200.0 903600.0 629400.0 917400.0 ;
      RECT  619200.0 931200.0 629400.0 917400.0 ;
      RECT  619200.0 931200.0 629400.0 945000.0 ;
      RECT  619200.0 958800.0 629400.0 945000.0 ;
      RECT  619200.0 958800.0 629400.0 972600.0 ;
      RECT  619200.0 986400.0 629400.0 972600.0 ;
      RECT  619200.0 986400.0 629400.0 1000200.0 ;
      RECT  619200.0 1014000.0 629400.0 1000200.0 ;
      RECT  619200.0 1014000.0 629400.0 1027800.0 ;
      RECT  619200.0 1041600.0 629400.0 1027800.0 ;
      RECT  619200.0 1041600.0 629400.0 1055400.0 ;
      RECT  619200.0 1069200.0 629400.0 1055400.0 ;
      RECT  619200.0 1069200.0 629400.0 1083000.0 ;
      RECT  619200.0 1096800.0 629400.0 1083000.0 ;
      RECT  619200.0 1096800.0 629400.0 1110600.0 ;
      RECT  619200.0 1124400.0 629400.0 1110600.0 ;
      RECT  619200.0 1124400.0 629400.0 1138200.0 ;
      RECT  619200.0 1152000.0 629400.0 1138200.0 ;
      RECT  619200.0 1152000.0 629400.0 1165800.0 ;
      RECT  619200.0 1179600.0 629400.0 1165800.0 ;
      RECT  619200.0 1179600.0 629400.0 1193400.0 ;
      RECT  619200.0 1207200.0 629400.0 1193400.0 ;
      RECT  619200.0 1207200.0 629400.0 1221000.0 ;
      RECT  619200.0 1234800.0 629400.0 1221000.0 ;
      RECT  619200.0 1234800.0 629400.0 1248600.0 ;
      RECT  619200.0 1262400.0 629400.0 1248600.0 ;
      RECT  619200.0 1262400.0 629400.0 1276200.0 ;
      RECT  619200.0 1290000.0 629400.0 1276200.0 ;
      RECT  619200.0 1290000.0 629400.0 1303800.0 ;
      RECT  619200.0 1317600.0 629400.0 1303800.0 ;
      RECT  619200.0 1317600.0 629400.0 1331400.0 ;
      RECT  619200.0 1345200.0 629400.0 1331400.0 ;
      RECT  619200.0 1345200.0 629400.0 1359000.0 ;
      RECT  619200.0 1372800.0 629400.0 1359000.0 ;
      RECT  619200.0 1372800.0 629400.0 1386600.0 ;
      RECT  619200.0 1400400.0 629400.0 1386600.0 ;
      RECT  619200.0 1400400.0 629400.0 1414200.0 ;
      RECT  619200.0 1428000.0 629400.0 1414200.0 ;
      RECT  619200.0 1428000.0 629400.0 1441800.0 ;
      RECT  619200.0 1455600.0 629400.0 1441800.0 ;
      RECT  619200.0 1455600.0 629400.0 1469400.0 ;
      RECT  619200.0 1483200.0 629400.0 1469400.0 ;
      RECT  619200.0 1483200.0 629400.0 1497000.0 ;
      RECT  619200.0 1510800.0 629400.0 1497000.0 ;
      RECT  619200.0 1510800.0 629400.0 1524600.0 ;
      RECT  619200.0 1538400.0 629400.0 1524600.0 ;
      RECT  619200.0 1538400.0 629400.0 1552200.0 ;
      RECT  619200.0 1566000.0 629400.0 1552200.0 ;
      RECT  619200.0 1566000.0 629400.0 1579800.0 ;
      RECT  619200.0 1593600.0 629400.0 1579800.0 ;
      RECT  619200.0 1593600.0 629400.0 1607400.0 ;
      RECT  619200.0 1621200.0 629400.0 1607400.0 ;
      RECT  619200.0 1621200.0 629400.0 1635000.0 ;
      RECT  619200.0 1648800.0 629400.0 1635000.0 ;
      RECT  619200.0 1648800.0 629400.0 1662600.0 ;
      RECT  619200.0 1676400.0 629400.0 1662600.0 ;
      RECT  619200.0 1676400.0 629400.0 1690200.0 ;
      RECT  619200.0 1704000.0 629400.0 1690200.0 ;
      RECT  619200.0 1704000.0 629400.0 1717800.0 ;
      RECT  619200.0 1731600.0 629400.0 1717800.0 ;
      RECT  619200.0 1731600.0 629400.0 1745400.0 ;
      RECT  619200.0 1759200.0 629400.0 1745400.0 ;
      RECT  619200.0 1759200.0 629400.0 1773000.0 ;
      RECT  619200.0 1786800.0 629400.0 1773000.0 ;
      RECT  619200.0 1786800.0 629400.0 1800600.0 ;
      RECT  619200.0 1814400.0 629400.0 1800600.0 ;
      RECT  619200.0 1814400.0 629400.0 1828200.0 ;
      RECT  619200.0 1842000.0 629400.0 1828200.0 ;
      RECT  619200.0 1842000.0 629400.0 1855800.0 ;
      RECT  619200.0 1869600.0 629400.0 1855800.0 ;
      RECT  619200.0 1869600.0 629400.0 1883400.0 ;
      RECT  619200.0 1897200.0 629400.0 1883400.0 ;
      RECT  619200.0 1897200.0 629400.0 1911000.0 ;
      RECT  619200.0 1924800.0 629400.0 1911000.0 ;
      RECT  619200.0 1924800.0 629400.0 1938600.0 ;
      RECT  619200.0 1952400.0 629400.0 1938600.0 ;
      RECT  619200.0 1952400.0 629400.0 1966200.0 ;
      RECT  619200.0 1980000.0 629400.0 1966200.0 ;
      RECT  619200.0 1980000.0 629400.0 1993800.0 ;
      RECT  619200.0 2007600.0 629400.0 1993800.0 ;
      RECT  619200.0 2007600.0 629400.0 2021400.0 ;
      RECT  619200.0 2035200.0 629400.0 2021400.0 ;
      RECT  619200.0 2035200.0 629400.0 2049000.0 ;
      RECT  619200.0 2062800.0 629400.0 2049000.0 ;
      RECT  619200.0 2062800.0 629400.0 2076600.0 ;
      RECT  619200.0 2090400.0 629400.0 2076600.0 ;
      RECT  619200.0 2090400.0 629400.0 2104200.0 ;
      RECT  619200.0 2118000.0 629400.0 2104200.0 ;
      RECT  619200.0 2118000.0 629400.0 2131800.0 ;
      RECT  619200.0 2145600.0 629400.0 2131800.0 ;
      RECT  629400.0 379200.0 639600.0 393000.0 ;
      RECT  629400.0 406800.0 639600.0 393000.0 ;
      RECT  629400.0 406800.0 639600.0 420600.0 ;
      RECT  629400.0 434400.0 639600.0 420600.0 ;
      RECT  629400.0 434400.0 639600.0 448200.0 ;
      RECT  629400.0 462000.0 639600.0 448200.0 ;
      RECT  629400.0 462000.0 639600.0 475800.0 ;
      RECT  629400.0 489600.0 639600.0 475800.0 ;
      RECT  629400.0 489600.0 639600.0 503400.0 ;
      RECT  629400.0 517200.0 639600.0 503400.0 ;
      RECT  629400.0 517200.0 639600.0 531000.0 ;
      RECT  629400.0 544800.0 639600.0 531000.0 ;
      RECT  629400.0 544800.0 639600.0 558600.0 ;
      RECT  629400.0 572400.0 639600.0 558600.0 ;
      RECT  629400.0 572400.0 639600.0 586200.0 ;
      RECT  629400.0 600000.0 639600.0 586200.0 ;
      RECT  629400.0 600000.0 639600.0 613800.0 ;
      RECT  629400.0 627600.0 639600.0 613800.0 ;
      RECT  629400.0 627600.0 639600.0 641400.0 ;
      RECT  629400.0 655200.0 639600.0 641400.0 ;
      RECT  629400.0 655200.0 639600.0 669000.0 ;
      RECT  629400.0 682800.0 639600.0 669000.0 ;
      RECT  629400.0 682800.0 639600.0 696600.0 ;
      RECT  629400.0 710400.0 639600.0 696600.0 ;
      RECT  629400.0 710400.0 639600.0 724200.0 ;
      RECT  629400.0 738000.0 639600.0 724200.0 ;
      RECT  629400.0 738000.0 639600.0 751800.0 ;
      RECT  629400.0 765600.0 639600.0 751800.0 ;
      RECT  629400.0 765600.0 639600.0 779400.0 ;
      RECT  629400.0 793200.0 639600.0 779400.0 ;
      RECT  629400.0 793200.0 639600.0 807000.0 ;
      RECT  629400.0 820800.0 639600.0 807000.0 ;
      RECT  629400.0 820800.0 639600.0 834600.0 ;
      RECT  629400.0 848400.0 639600.0 834600.0 ;
      RECT  629400.0 848400.0 639600.0 862200.0 ;
      RECT  629400.0 876000.0 639600.0 862200.0 ;
      RECT  629400.0 876000.0 639600.0 889800.0 ;
      RECT  629400.0 903600.0 639600.0 889800.0 ;
      RECT  629400.0 903600.0 639600.0 917400.0 ;
      RECT  629400.0 931200.0 639600.0 917400.0 ;
      RECT  629400.0 931200.0 639600.0 945000.0 ;
      RECT  629400.0 958800.0 639600.0 945000.0 ;
      RECT  629400.0 958800.0 639600.0 972600.0 ;
      RECT  629400.0 986400.0 639600.0 972600.0 ;
      RECT  629400.0 986400.0 639600.0 1000200.0 ;
      RECT  629400.0 1014000.0 639600.0 1000200.0 ;
      RECT  629400.0 1014000.0 639600.0 1027800.0 ;
      RECT  629400.0 1041600.0 639600.0 1027800.0 ;
      RECT  629400.0 1041600.0 639600.0 1055400.0 ;
      RECT  629400.0 1069200.0 639600.0 1055400.0 ;
      RECT  629400.0 1069200.0 639600.0 1083000.0 ;
      RECT  629400.0 1096800.0 639600.0 1083000.0 ;
      RECT  629400.0 1096800.0 639600.0 1110600.0 ;
      RECT  629400.0 1124400.0 639600.0 1110600.0 ;
      RECT  629400.0 1124400.0 639600.0 1138200.0 ;
      RECT  629400.0 1152000.0 639600.0 1138200.0 ;
      RECT  629400.0 1152000.0 639600.0 1165800.0 ;
      RECT  629400.0 1179600.0 639600.0 1165800.0 ;
      RECT  629400.0 1179600.0 639600.0 1193400.0 ;
      RECT  629400.0 1207200.0 639600.0 1193400.0 ;
      RECT  629400.0 1207200.0 639600.0 1221000.0 ;
      RECT  629400.0 1234800.0 639600.0 1221000.0 ;
      RECT  629400.0 1234800.0 639600.0 1248600.0 ;
      RECT  629400.0 1262400.0 639600.0 1248600.0 ;
      RECT  629400.0 1262400.0 639600.0 1276200.0 ;
      RECT  629400.0 1290000.0 639600.0 1276200.0 ;
      RECT  629400.0 1290000.0 639600.0 1303800.0 ;
      RECT  629400.0 1317600.0 639600.0 1303800.0 ;
      RECT  629400.0 1317600.0 639600.0 1331400.0 ;
      RECT  629400.0 1345200.0 639600.0 1331400.0 ;
      RECT  629400.0 1345200.0 639600.0 1359000.0 ;
      RECT  629400.0 1372800.0 639600.0 1359000.0 ;
      RECT  629400.0 1372800.0 639600.0 1386600.0 ;
      RECT  629400.0 1400400.0 639600.0 1386600.0 ;
      RECT  629400.0 1400400.0 639600.0 1414200.0 ;
      RECT  629400.0 1428000.0 639600.0 1414200.0 ;
      RECT  629400.0 1428000.0 639600.0 1441800.0 ;
      RECT  629400.0 1455600.0 639600.0 1441800.0 ;
      RECT  629400.0 1455600.0 639600.0 1469400.0 ;
      RECT  629400.0 1483200.0 639600.0 1469400.0 ;
      RECT  629400.0 1483200.0 639600.0 1497000.0 ;
      RECT  629400.0 1510800.0 639600.0 1497000.0 ;
      RECT  629400.0 1510800.0 639600.0 1524600.0 ;
      RECT  629400.0 1538400.0 639600.0 1524600.0 ;
      RECT  629400.0 1538400.0 639600.0 1552200.0 ;
      RECT  629400.0 1566000.0 639600.0 1552200.0 ;
      RECT  629400.0 1566000.0 639600.0 1579800.0 ;
      RECT  629400.0 1593600.0 639600.0 1579800.0 ;
      RECT  629400.0 1593600.0 639600.0 1607400.0 ;
      RECT  629400.0 1621200.0 639600.0 1607400.0 ;
      RECT  629400.0 1621200.0 639600.0 1635000.0 ;
      RECT  629400.0 1648800.0 639600.0 1635000.0 ;
      RECT  629400.0 1648800.0 639600.0 1662600.0 ;
      RECT  629400.0 1676400.0 639600.0 1662600.0 ;
      RECT  629400.0 1676400.0 639600.0 1690200.0 ;
      RECT  629400.0 1704000.0 639600.0 1690200.0 ;
      RECT  629400.0 1704000.0 639600.0 1717800.0 ;
      RECT  629400.0 1731600.0 639600.0 1717800.0 ;
      RECT  629400.0 1731600.0 639600.0 1745400.0 ;
      RECT  629400.0 1759200.0 639600.0 1745400.0 ;
      RECT  629400.0 1759200.0 639600.0 1773000.0 ;
      RECT  629400.0 1786800.0 639600.0 1773000.0 ;
      RECT  629400.0 1786800.0 639600.0 1800600.0 ;
      RECT  629400.0 1814400.0 639600.0 1800600.0 ;
      RECT  629400.0 1814400.0 639600.0 1828200.0 ;
      RECT  629400.0 1842000.0 639600.0 1828200.0 ;
      RECT  629400.0 1842000.0 639600.0 1855800.0 ;
      RECT  629400.0 1869600.0 639600.0 1855800.0 ;
      RECT  629400.0 1869600.0 639600.0 1883400.0 ;
      RECT  629400.0 1897200.0 639600.0 1883400.0 ;
      RECT  629400.0 1897200.0 639600.0 1911000.0 ;
      RECT  629400.0 1924800.0 639600.0 1911000.0 ;
      RECT  629400.0 1924800.0 639600.0 1938600.0 ;
      RECT  629400.0 1952400.0 639600.0 1938600.0 ;
      RECT  629400.0 1952400.0 639600.0 1966200.0 ;
      RECT  629400.0 1980000.0 639600.0 1966200.0 ;
      RECT  629400.0 1980000.0 639600.0 1993800.0 ;
      RECT  629400.0 2007600.0 639600.0 1993800.0 ;
      RECT  629400.0 2007600.0 639600.0 2021400.0 ;
      RECT  629400.0 2035200.0 639600.0 2021400.0 ;
      RECT  629400.0 2035200.0 639600.0 2049000.0 ;
      RECT  629400.0 2062800.0 639600.0 2049000.0 ;
      RECT  629400.0 2062800.0 639600.0 2076600.0 ;
      RECT  629400.0 2090400.0 639600.0 2076600.0 ;
      RECT  629400.0 2090400.0 639600.0 2104200.0 ;
      RECT  629400.0 2118000.0 639600.0 2104200.0 ;
      RECT  629400.0 2118000.0 639600.0 2131800.0 ;
      RECT  629400.0 2145600.0 639600.0 2131800.0 ;
      RECT  639600.0 379200.0 649800.0 393000.0 ;
      RECT  639600.0 406800.0 649800.0 393000.0 ;
      RECT  639600.0 406800.0 649800.0 420600.0 ;
      RECT  639600.0 434400.0 649800.0 420600.0 ;
      RECT  639600.0 434400.0 649800.0 448200.0 ;
      RECT  639600.0 462000.0 649800.0 448200.0 ;
      RECT  639600.0 462000.0 649800.0 475800.0 ;
      RECT  639600.0 489600.0 649800.0 475800.0 ;
      RECT  639600.0 489600.0 649800.0 503400.0 ;
      RECT  639600.0 517200.0 649800.0 503400.0 ;
      RECT  639600.0 517200.0 649800.0 531000.0 ;
      RECT  639600.0 544800.0 649800.0 531000.0 ;
      RECT  639600.0 544800.0 649800.0 558600.0 ;
      RECT  639600.0 572400.0 649800.0 558600.0 ;
      RECT  639600.0 572400.0 649800.0 586200.0 ;
      RECT  639600.0 600000.0 649800.0 586200.0 ;
      RECT  639600.0 600000.0 649800.0 613800.0 ;
      RECT  639600.0 627600.0 649800.0 613800.0 ;
      RECT  639600.0 627600.0 649800.0 641400.0 ;
      RECT  639600.0 655200.0 649800.0 641400.0 ;
      RECT  639600.0 655200.0 649800.0 669000.0 ;
      RECT  639600.0 682800.0 649800.0 669000.0 ;
      RECT  639600.0 682800.0 649800.0 696600.0 ;
      RECT  639600.0 710400.0 649800.0 696600.0 ;
      RECT  639600.0 710400.0 649800.0 724200.0 ;
      RECT  639600.0 738000.0 649800.0 724200.0 ;
      RECT  639600.0 738000.0 649800.0 751800.0 ;
      RECT  639600.0 765600.0 649800.0 751800.0 ;
      RECT  639600.0 765600.0 649800.0 779400.0 ;
      RECT  639600.0 793200.0 649800.0 779400.0 ;
      RECT  639600.0 793200.0 649800.0 807000.0 ;
      RECT  639600.0 820800.0 649800.0 807000.0 ;
      RECT  639600.0 820800.0 649800.0 834600.0 ;
      RECT  639600.0 848400.0 649800.0 834600.0 ;
      RECT  639600.0 848400.0 649800.0 862200.0 ;
      RECT  639600.0 876000.0 649800.0 862200.0 ;
      RECT  639600.0 876000.0 649800.0 889800.0 ;
      RECT  639600.0 903600.0 649800.0 889800.0 ;
      RECT  639600.0 903600.0 649800.0 917400.0 ;
      RECT  639600.0 931200.0 649800.0 917400.0 ;
      RECT  639600.0 931200.0 649800.0 945000.0 ;
      RECT  639600.0 958800.0 649800.0 945000.0 ;
      RECT  639600.0 958800.0 649800.0 972600.0 ;
      RECT  639600.0 986400.0 649800.0 972600.0 ;
      RECT  639600.0 986400.0 649800.0 1000200.0 ;
      RECT  639600.0 1014000.0 649800.0 1000200.0 ;
      RECT  639600.0 1014000.0 649800.0 1027800.0 ;
      RECT  639600.0 1041600.0 649800.0 1027800.0 ;
      RECT  639600.0 1041600.0 649800.0 1055400.0 ;
      RECT  639600.0 1069200.0 649800.0 1055400.0 ;
      RECT  639600.0 1069200.0 649800.0 1083000.0 ;
      RECT  639600.0 1096800.0 649800.0 1083000.0 ;
      RECT  639600.0 1096800.0 649800.0 1110600.0 ;
      RECT  639600.0 1124400.0 649800.0 1110600.0 ;
      RECT  639600.0 1124400.0 649800.0 1138200.0 ;
      RECT  639600.0 1152000.0 649800.0 1138200.0 ;
      RECT  639600.0 1152000.0 649800.0 1165800.0 ;
      RECT  639600.0 1179600.0 649800.0 1165800.0 ;
      RECT  639600.0 1179600.0 649800.0 1193400.0 ;
      RECT  639600.0 1207200.0 649800.0 1193400.0 ;
      RECT  639600.0 1207200.0 649800.0 1221000.0 ;
      RECT  639600.0 1234800.0 649800.0 1221000.0 ;
      RECT  639600.0 1234800.0 649800.0 1248600.0 ;
      RECT  639600.0 1262400.0 649800.0 1248600.0 ;
      RECT  639600.0 1262400.0 649800.0 1276200.0 ;
      RECT  639600.0 1290000.0 649800.0 1276200.0 ;
      RECT  639600.0 1290000.0 649800.0 1303800.0 ;
      RECT  639600.0 1317600.0 649800.0 1303800.0 ;
      RECT  639600.0 1317600.0 649800.0 1331400.0 ;
      RECT  639600.0 1345200.0 649800.0 1331400.0 ;
      RECT  639600.0 1345200.0 649800.0 1359000.0 ;
      RECT  639600.0 1372800.0 649800.0 1359000.0 ;
      RECT  639600.0 1372800.0 649800.0 1386600.0 ;
      RECT  639600.0 1400400.0 649800.0 1386600.0 ;
      RECT  639600.0 1400400.0 649800.0 1414200.0 ;
      RECT  639600.0 1428000.0 649800.0 1414200.0 ;
      RECT  639600.0 1428000.0 649800.0 1441800.0 ;
      RECT  639600.0 1455600.0 649800.0 1441800.0 ;
      RECT  639600.0 1455600.0 649800.0 1469400.0 ;
      RECT  639600.0 1483200.0 649800.0 1469400.0 ;
      RECT  639600.0 1483200.0 649800.0 1497000.0 ;
      RECT  639600.0 1510800.0 649800.0 1497000.0 ;
      RECT  639600.0 1510800.0 649800.0 1524600.0 ;
      RECT  639600.0 1538400.0 649800.0 1524600.0 ;
      RECT  639600.0 1538400.0 649800.0 1552200.0 ;
      RECT  639600.0 1566000.0 649800.0 1552200.0 ;
      RECT  639600.0 1566000.0 649800.0 1579800.0 ;
      RECT  639600.0 1593600.0 649800.0 1579800.0 ;
      RECT  639600.0 1593600.0 649800.0 1607400.0 ;
      RECT  639600.0 1621200.0 649800.0 1607400.0 ;
      RECT  639600.0 1621200.0 649800.0 1635000.0 ;
      RECT  639600.0 1648800.0 649800.0 1635000.0 ;
      RECT  639600.0 1648800.0 649800.0 1662600.0 ;
      RECT  639600.0 1676400.0 649800.0 1662600.0 ;
      RECT  639600.0 1676400.0 649800.0 1690200.0 ;
      RECT  639600.0 1704000.0 649800.0 1690200.0 ;
      RECT  639600.0 1704000.0 649800.0 1717800.0 ;
      RECT  639600.0 1731600.0 649800.0 1717800.0 ;
      RECT  639600.0 1731600.0 649800.0 1745400.0 ;
      RECT  639600.0 1759200.0 649800.0 1745400.0 ;
      RECT  639600.0 1759200.0 649800.0 1773000.0 ;
      RECT  639600.0 1786800.0 649800.0 1773000.0 ;
      RECT  639600.0 1786800.0 649800.0 1800600.0 ;
      RECT  639600.0 1814400.0 649800.0 1800600.0 ;
      RECT  639600.0 1814400.0 649800.0 1828200.0 ;
      RECT  639600.0 1842000.0 649800.0 1828200.0 ;
      RECT  639600.0 1842000.0 649800.0 1855800.0 ;
      RECT  639600.0 1869600.0 649800.0 1855800.0 ;
      RECT  639600.0 1869600.0 649800.0 1883400.0 ;
      RECT  639600.0 1897200.0 649800.0 1883400.0 ;
      RECT  639600.0 1897200.0 649800.0 1911000.0 ;
      RECT  639600.0 1924800.0 649800.0 1911000.0 ;
      RECT  639600.0 1924800.0 649800.0 1938600.0 ;
      RECT  639600.0 1952400.0 649800.0 1938600.0 ;
      RECT  639600.0 1952400.0 649800.0 1966200.0 ;
      RECT  639600.0 1980000.0 649800.0 1966200.0 ;
      RECT  639600.0 1980000.0 649800.0 1993800.0 ;
      RECT  639600.0 2007600.0 649800.0 1993800.0 ;
      RECT  639600.0 2007600.0 649800.0 2021400.0 ;
      RECT  639600.0 2035200.0 649800.0 2021400.0 ;
      RECT  639600.0 2035200.0 649800.0 2049000.0 ;
      RECT  639600.0 2062800.0 649800.0 2049000.0 ;
      RECT  639600.0 2062800.0 649800.0 2076600.0 ;
      RECT  639600.0 2090400.0 649800.0 2076600.0 ;
      RECT  639600.0 2090400.0 649800.0 2104200.0 ;
      RECT  639600.0 2118000.0 649800.0 2104200.0 ;
      RECT  639600.0 2118000.0 649800.0 2131800.0 ;
      RECT  639600.0 2145600.0 649800.0 2131800.0 ;
      RECT  649800.0 379200.0 660000.0 393000.0 ;
      RECT  649800.0 406800.0 660000.0 393000.0 ;
      RECT  649800.0 406800.0 660000.0 420600.0 ;
      RECT  649800.0 434400.0 660000.0 420600.0 ;
      RECT  649800.0 434400.0 660000.0 448200.0 ;
      RECT  649800.0 462000.0 660000.0 448200.0 ;
      RECT  649800.0 462000.0 660000.0 475800.0 ;
      RECT  649800.0 489600.0 660000.0 475800.0 ;
      RECT  649800.0 489600.0 660000.0 503400.0 ;
      RECT  649800.0 517200.0 660000.0 503400.0 ;
      RECT  649800.0 517200.0 660000.0 531000.0 ;
      RECT  649800.0 544800.0 660000.0 531000.0 ;
      RECT  649800.0 544800.0 660000.0 558600.0 ;
      RECT  649800.0 572400.0 660000.0 558600.0 ;
      RECT  649800.0 572400.0 660000.0 586200.0 ;
      RECT  649800.0 600000.0 660000.0 586200.0 ;
      RECT  649800.0 600000.0 660000.0 613800.0 ;
      RECT  649800.0 627600.0 660000.0 613800.0 ;
      RECT  649800.0 627600.0 660000.0 641400.0 ;
      RECT  649800.0 655200.0 660000.0 641400.0 ;
      RECT  649800.0 655200.0 660000.0 669000.0 ;
      RECT  649800.0 682800.0 660000.0 669000.0 ;
      RECT  649800.0 682800.0 660000.0 696600.0 ;
      RECT  649800.0 710400.0 660000.0 696600.0 ;
      RECT  649800.0 710400.0 660000.0 724200.0 ;
      RECT  649800.0 738000.0 660000.0 724200.0 ;
      RECT  649800.0 738000.0 660000.0 751800.0 ;
      RECT  649800.0 765600.0 660000.0 751800.0 ;
      RECT  649800.0 765600.0 660000.0 779400.0 ;
      RECT  649800.0 793200.0 660000.0 779400.0 ;
      RECT  649800.0 793200.0 660000.0 807000.0 ;
      RECT  649800.0 820800.0 660000.0 807000.0 ;
      RECT  649800.0 820800.0 660000.0 834600.0 ;
      RECT  649800.0 848400.0 660000.0 834600.0 ;
      RECT  649800.0 848400.0 660000.0 862200.0 ;
      RECT  649800.0 876000.0 660000.0 862200.0 ;
      RECT  649800.0 876000.0 660000.0 889800.0 ;
      RECT  649800.0 903600.0 660000.0 889800.0 ;
      RECT  649800.0 903600.0 660000.0 917400.0 ;
      RECT  649800.0 931200.0 660000.0 917400.0 ;
      RECT  649800.0 931200.0 660000.0 945000.0 ;
      RECT  649800.0 958800.0 660000.0 945000.0 ;
      RECT  649800.0 958800.0 660000.0 972600.0 ;
      RECT  649800.0 986400.0 660000.0 972600.0 ;
      RECT  649800.0 986400.0 660000.0 1000200.0 ;
      RECT  649800.0 1014000.0 660000.0 1000200.0 ;
      RECT  649800.0 1014000.0 660000.0 1027800.0 ;
      RECT  649800.0 1041600.0 660000.0 1027800.0 ;
      RECT  649800.0 1041600.0 660000.0 1055400.0 ;
      RECT  649800.0 1069200.0 660000.0 1055400.0 ;
      RECT  649800.0 1069200.0 660000.0 1083000.0 ;
      RECT  649800.0 1096800.0 660000.0 1083000.0 ;
      RECT  649800.0 1096800.0 660000.0 1110600.0 ;
      RECT  649800.0 1124400.0 660000.0 1110600.0 ;
      RECT  649800.0 1124400.0 660000.0 1138200.0 ;
      RECT  649800.0 1152000.0 660000.0 1138200.0 ;
      RECT  649800.0 1152000.0 660000.0 1165800.0 ;
      RECT  649800.0 1179600.0 660000.0 1165800.0 ;
      RECT  649800.0 1179600.0 660000.0 1193400.0 ;
      RECT  649800.0 1207200.0 660000.0 1193400.0 ;
      RECT  649800.0 1207200.0 660000.0 1221000.0 ;
      RECT  649800.0 1234800.0 660000.0 1221000.0 ;
      RECT  649800.0 1234800.0 660000.0 1248600.0 ;
      RECT  649800.0 1262400.0 660000.0 1248600.0 ;
      RECT  649800.0 1262400.0 660000.0 1276200.0 ;
      RECT  649800.0 1290000.0 660000.0 1276200.0 ;
      RECT  649800.0 1290000.0 660000.0 1303800.0 ;
      RECT  649800.0 1317600.0 660000.0 1303800.0 ;
      RECT  649800.0 1317600.0 660000.0 1331400.0 ;
      RECT  649800.0 1345200.0 660000.0 1331400.0 ;
      RECT  649800.0 1345200.0 660000.0 1359000.0 ;
      RECT  649800.0 1372800.0 660000.0 1359000.0 ;
      RECT  649800.0 1372800.0 660000.0 1386600.0 ;
      RECT  649800.0 1400400.0 660000.0 1386600.0 ;
      RECT  649800.0 1400400.0 660000.0 1414200.0 ;
      RECT  649800.0 1428000.0 660000.0 1414200.0 ;
      RECT  649800.0 1428000.0 660000.0 1441800.0 ;
      RECT  649800.0 1455600.0 660000.0 1441800.0 ;
      RECT  649800.0 1455600.0 660000.0 1469400.0 ;
      RECT  649800.0 1483200.0 660000.0 1469400.0 ;
      RECT  649800.0 1483200.0 660000.0 1497000.0 ;
      RECT  649800.0 1510800.0 660000.0 1497000.0 ;
      RECT  649800.0 1510800.0 660000.0 1524600.0 ;
      RECT  649800.0 1538400.0 660000.0 1524600.0 ;
      RECT  649800.0 1538400.0 660000.0 1552200.0 ;
      RECT  649800.0 1566000.0 660000.0 1552200.0 ;
      RECT  649800.0 1566000.0 660000.0 1579800.0 ;
      RECT  649800.0 1593600.0 660000.0 1579800.0 ;
      RECT  649800.0 1593600.0 660000.0 1607400.0 ;
      RECT  649800.0 1621200.0 660000.0 1607400.0 ;
      RECT  649800.0 1621200.0 660000.0 1635000.0 ;
      RECT  649800.0 1648800.0 660000.0 1635000.0 ;
      RECT  649800.0 1648800.0 660000.0 1662600.0 ;
      RECT  649800.0 1676400.0 660000.0 1662600.0 ;
      RECT  649800.0 1676400.0 660000.0 1690200.0 ;
      RECT  649800.0 1704000.0 660000.0 1690200.0 ;
      RECT  649800.0 1704000.0 660000.0 1717800.0 ;
      RECT  649800.0 1731600.0 660000.0 1717800.0 ;
      RECT  649800.0 1731600.0 660000.0 1745400.0 ;
      RECT  649800.0 1759200.0 660000.0 1745400.0 ;
      RECT  649800.0 1759200.0 660000.0 1773000.0 ;
      RECT  649800.0 1786800.0 660000.0 1773000.0 ;
      RECT  649800.0 1786800.0 660000.0 1800600.0 ;
      RECT  649800.0 1814400.0 660000.0 1800600.0 ;
      RECT  649800.0 1814400.0 660000.0 1828200.0 ;
      RECT  649800.0 1842000.0 660000.0 1828200.0 ;
      RECT  649800.0 1842000.0 660000.0 1855800.0 ;
      RECT  649800.0 1869600.0 660000.0 1855800.0 ;
      RECT  649800.0 1869600.0 660000.0 1883400.0 ;
      RECT  649800.0 1897200.0 660000.0 1883400.0 ;
      RECT  649800.0 1897200.0 660000.0 1911000.0 ;
      RECT  649800.0 1924800.0 660000.0 1911000.0 ;
      RECT  649800.0 1924800.0 660000.0 1938600.0 ;
      RECT  649800.0 1952400.0 660000.0 1938600.0 ;
      RECT  649800.0 1952400.0 660000.0 1966200.0 ;
      RECT  649800.0 1980000.0 660000.0 1966200.0 ;
      RECT  649800.0 1980000.0 660000.0 1993800.0 ;
      RECT  649800.0 2007600.0 660000.0 1993800.0 ;
      RECT  649800.0 2007600.0 660000.0 2021400.0 ;
      RECT  649800.0 2035200.0 660000.0 2021400.0 ;
      RECT  649800.0 2035200.0 660000.0 2049000.0 ;
      RECT  649800.0 2062800.0 660000.0 2049000.0 ;
      RECT  649800.0 2062800.0 660000.0 2076600.0 ;
      RECT  649800.0 2090400.0 660000.0 2076600.0 ;
      RECT  649800.0 2090400.0 660000.0 2104200.0 ;
      RECT  649800.0 2118000.0 660000.0 2104200.0 ;
      RECT  649800.0 2118000.0 660000.0 2131800.0 ;
      RECT  649800.0 2145600.0 660000.0 2131800.0 ;
      RECT  660000.0 379200.0 670200.0 393000.0 ;
      RECT  660000.0 406800.0 670200.0 393000.0 ;
      RECT  660000.0 406800.0 670200.0 420600.0 ;
      RECT  660000.0 434400.0 670200.0 420600.0 ;
      RECT  660000.0 434400.0 670200.0 448200.0 ;
      RECT  660000.0 462000.0 670200.0 448200.0 ;
      RECT  660000.0 462000.0 670200.0 475800.0 ;
      RECT  660000.0 489600.0 670200.0 475800.0 ;
      RECT  660000.0 489600.0 670200.0 503400.0 ;
      RECT  660000.0 517200.0 670200.0 503400.0 ;
      RECT  660000.0 517200.0 670200.0 531000.0 ;
      RECT  660000.0 544800.0 670200.0 531000.0 ;
      RECT  660000.0 544800.0 670200.0 558600.0 ;
      RECT  660000.0 572400.0 670200.0 558600.0 ;
      RECT  660000.0 572400.0 670200.0 586200.0 ;
      RECT  660000.0 600000.0 670200.0 586200.0 ;
      RECT  660000.0 600000.0 670200.0 613800.0 ;
      RECT  660000.0 627600.0 670200.0 613800.0 ;
      RECT  660000.0 627600.0 670200.0 641400.0 ;
      RECT  660000.0 655200.0 670200.0 641400.0 ;
      RECT  660000.0 655200.0 670200.0 669000.0 ;
      RECT  660000.0 682800.0 670200.0 669000.0 ;
      RECT  660000.0 682800.0 670200.0 696600.0 ;
      RECT  660000.0 710400.0 670200.0 696600.0 ;
      RECT  660000.0 710400.0 670200.0 724200.0 ;
      RECT  660000.0 738000.0 670200.0 724200.0 ;
      RECT  660000.0 738000.0 670200.0 751800.0 ;
      RECT  660000.0 765600.0 670200.0 751800.0 ;
      RECT  660000.0 765600.0 670200.0 779400.0 ;
      RECT  660000.0 793200.0 670200.0 779400.0 ;
      RECT  660000.0 793200.0 670200.0 807000.0 ;
      RECT  660000.0 820800.0 670200.0 807000.0 ;
      RECT  660000.0 820800.0 670200.0 834600.0 ;
      RECT  660000.0 848400.0 670200.0 834600.0 ;
      RECT  660000.0 848400.0 670200.0 862200.0 ;
      RECT  660000.0 876000.0 670200.0 862200.0 ;
      RECT  660000.0 876000.0 670200.0 889800.0 ;
      RECT  660000.0 903600.0 670200.0 889800.0 ;
      RECT  660000.0 903600.0 670200.0 917400.0 ;
      RECT  660000.0 931200.0 670200.0 917400.0 ;
      RECT  660000.0 931200.0 670200.0 945000.0 ;
      RECT  660000.0 958800.0 670200.0 945000.0 ;
      RECT  660000.0 958800.0 670200.0 972600.0 ;
      RECT  660000.0 986400.0 670200.0 972600.0 ;
      RECT  660000.0 986400.0 670200.0 1000200.0 ;
      RECT  660000.0 1014000.0 670200.0 1000200.0 ;
      RECT  660000.0 1014000.0 670200.0 1027800.0 ;
      RECT  660000.0 1041600.0 670200.0 1027800.0 ;
      RECT  660000.0 1041600.0 670200.0 1055400.0 ;
      RECT  660000.0 1069200.0 670200.0 1055400.0 ;
      RECT  660000.0 1069200.0 670200.0 1083000.0 ;
      RECT  660000.0 1096800.0 670200.0 1083000.0 ;
      RECT  660000.0 1096800.0 670200.0 1110600.0 ;
      RECT  660000.0 1124400.0 670200.0 1110600.0 ;
      RECT  660000.0 1124400.0 670200.0 1138200.0 ;
      RECT  660000.0 1152000.0 670200.0 1138200.0 ;
      RECT  660000.0 1152000.0 670200.0 1165800.0 ;
      RECT  660000.0 1179600.0 670200.0 1165800.0 ;
      RECT  660000.0 1179600.0 670200.0 1193400.0 ;
      RECT  660000.0 1207200.0 670200.0 1193400.0 ;
      RECT  660000.0 1207200.0 670200.0 1221000.0 ;
      RECT  660000.0 1234800.0 670200.0 1221000.0 ;
      RECT  660000.0 1234800.0 670200.0 1248600.0 ;
      RECT  660000.0 1262400.0 670200.0 1248600.0 ;
      RECT  660000.0 1262400.0 670200.0 1276200.0 ;
      RECT  660000.0 1290000.0 670200.0 1276200.0 ;
      RECT  660000.0 1290000.0 670200.0 1303800.0 ;
      RECT  660000.0 1317600.0 670200.0 1303800.0 ;
      RECT  660000.0 1317600.0 670200.0 1331400.0 ;
      RECT  660000.0 1345200.0 670200.0 1331400.0 ;
      RECT  660000.0 1345200.0 670200.0 1359000.0 ;
      RECT  660000.0 1372800.0 670200.0 1359000.0 ;
      RECT  660000.0 1372800.0 670200.0 1386600.0 ;
      RECT  660000.0 1400400.0 670200.0 1386600.0 ;
      RECT  660000.0 1400400.0 670200.0 1414200.0 ;
      RECT  660000.0 1428000.0 670200.0 1414200.0 ;
      RECT  660000.0 1428000.0 670200.0 1441800.0 ;
      RECT  660000.0 1455600.0 670200.0 1441800.0 ;
      RECT  660000.0 1455600.0 670200.0 1469400.0 ;
      RECT  660000.0 1483200.0 670200.0 1469400.0 ;
      RECT  660000.0 1483200.0 670200.0 1497000.0 ;
      RECT  660000.0 1510800.0 670200.0 1497000.0 ;
      RECT  660000.0 1510800.0 670200.0 1524600.0 ;
      RECT  660000.0 1538400.0 670200.0 1524600.0 ;
      RECT  660000.0 1538400.0 670200.0 1552200.0 ;
      RECT  660000.0 1566000.0 670200.0 1552200.0 ;
      RECT  660000.0 1566000.0 670200.0 1579800.0 ;
      RECT  660000.0 1593600.0 670200.0 1579800.0 ;
      RECT  660000.0 1593600.0 670200.0 1607400.0 ;
      RECT  660000.0 1621200.0 670200.0 1607400.0 ;
      RECT  660000.0 1621200.0 670200.0 1635000.0 ;
      RECT  660000.0 1648800.0 670200.0 1635000.0 ;
      RECT  660000.0 1648800.0 670200.0 1662600.0 ;
      RECT  660000.0 1676400.0 670200.0 1662600.0 ;
      RECT  660000.0 1676400.0 670200.0 1690200.0 ;
      RECT  660000.0 1704000.0 670200.0 1690200.0 ;
      RECT  660000.0 1704000.0 670200.0 1717800.0 ;
      RECT  660000.0 1731600.0 670200.0 1717800.0 ;
      RECT  660000.0 1731600.0 670200.0 1745400.0 ;
      RECT  660000.0 1759200.0 670200.0 1745400.0 ;
      RECT  660000.0 1759200.0 670200.0 1773000.0 ;
      RECT  660000.0 1786800.0 670200.0 1773000.0 ;
      RECT  660000.0 1786800.0 670200.0 1800600.0 ;
      RECT  660000.0 1814400.0 670200.0 1800600.0 ;
      RECT  660000.0 1814400.0 670200.0 1828200.0 ;
      RECT  660000.0 1842000.0 670200.0 1828200.0 ;
      RECT  660000.0 1842000.0 670200.0 1855800.0 ;
      RECT  660000.0 1869600.0 670200.0 1855800.0 ;
      RECT  660000.0 1869600.0 670200.0 1883400.0 ;
      RECT  660000.0 1897200.0 670200.0 1883400.0 ;
      RECT  660000.0 1897200.0 670200.0 1911000.0 ;
      RECT  660000.0 1924800.0 670200.0 1911000.0 ;
      RECT  660000.0 1924800.0 670200.0 1938600.0 ;
      RECT  660000.0 1952400.0 670200.0 1938600.0 ;
      RECT  660000.0 1952400.0 670200.0 1966200.0 ;
      RECT  660000.0 1980000.0 670200.0 1966200.0 ;
      RECT  660000.0 1980000.0 670200.0 1993800.0 ;
      RECT  660000.0 2007600.0 670200.0 1993800.0 ;
      RECT  660000.0 2007600.0 670200.0 2021400.0 ;
      RECT  660000.0 2035200.0 670200.0 2021400.0 ;
      RECT  660000.0 2035200.0 670200.0 2049000.0 ;
      RECT  660000.0 2062800.0 670200.0 2049000.0 ;
      RECT  660000.0 2062800.0 670200.0 2076600.0 ;
      RECT  660000.0 2090400.0 670200.0 2076600.0 ;
      RECT  660000.0 2090400.0 670200.0 2104200.0 ;
      RECT  660000.0 2118000.0 670200.0 2104200.0 ;
      RECT  660000.0 2118000.0 670200.0 2131800.0 ;
      RECT  660000.0 2145600.0 670200.0 2131800.0 ;
      RECT  670200.0 379200.0 680400.0 393000.0 ;
      RECT  670200.0 406800.0 680400.0 393000.0 ;
      RECT  670200.0 406800.0 680400.0 420600.0 ;
      RECT  670200.0 434400.0 680400.0 420600.0 ;
      RECT  670200.0 434400.0 680400.0 448200.0 ;
      RECT  670200.0 462000.0 680400.0 448200.0 ;
      RECT  670200.0 462000.0 680400.0 475800.0 ;
      RECT  670200.0 489600.0 680400.0 475800.0 ;
      RECT  670200.0 489600.0 680400.0 503400.0 ;
      RECT  670200.0 517200.0 680400.0 503400.0 ;
      RECT  670200.0 517200.0 680400.0 531000.0 ;
      RECT  670200.0 544800.0 680400.0 531000.0 ;
      RECT  670200.0 544800.0 680400.0 558600.0 ;
      RECT  670200.0 572400.0 680400.0 558600.0 ;
      RECT  670200.0 572400.0 680400.0 586200.0 ;
      RECT  670200.0 600000.0 680400.0 586200.0 ;
      RECT  670200.0 600000.0 680400.0 613800.0 ;
      RECT  670200.0 627600.0 680400.0 613800.0 ;
      RECT  670200.0 627600.0 680400.0 641400.0 ;
      RECT  670200.0 655200.0 680400.0 641400.0 ;
      RECT  670200.0 655200.0 680400.0 669000.0 ;
      RECT  670200.0 682800.0 680400.0 669000.0 ;
      RECT  670200.0 682800.0 680400.0 696600.0 ;
      RECT  670200.0 710400.0 680400.0 696600.0 ;
      RECT  670200.0 710400.0 680400.0 724200.0 ;
      RECT  670200.0 738000.0 680400.0 724200.0 ;
      RECT  670200.0 738000.0 680400.0 751800.0 ;
      RECT  670200.0 765600.0 680400.0 751800.0 ;
      RECT  670200.0 765600.0 680400.0 779400.0 ;
      RECT  670200.0 793200.0 680400.0 779400.0 ;
      RECT  670200.0 793200.0 680400.0 807000.0 ;
      RECT  670200.0 820800.0 680400.0 807000.0 ;
      RECT  670200.0 820800.0 680400.0 834600.0 ;
      RECT  670200.0 848400.0 680400.0 834600.0 ;
      RECT  670200.0 848400.0 680400.0 862200.0 ;
      RECT  670200.0 876000.0 680400.0 862200.0 ;
      RECT  670200.0 876000.0 680400.0 889800.0 ;
      RECT  670200.0 903600.0 680400.0 889800.0 ;
      RECT  670200.0 903600.0 680400.0 917400.0 ;
      RECT  670200.0 931200.0 680400.0 917400.0 ;
      RECT  670200.0 931200.0 680400.0 945000.0 ;
      RECT  670200.0 958800.0 680400.0 945000.0 ;
      RECT  670200.0 958800.0 680400.0 972600.0 ;
      RECT  670200.0 986400.0 680400.0 972600.0 ;
      RECT  670200.0 986400.0 680400.0 1000200.0 ;
      RECT  670200.0 1014000.0 680400.0 1000200.0 ;
      RECT  670200.0 1014000.0 680400.0 1027800.0 ;
      RECT  670200.0 1041600.0 680400.0 1027800.0 ;
      RECT  670200.0 1041600.0 680400.0 1055400.0 ;
      RECT  670200.0 1069200.0 680400.0 1055400.0 ;
      RECT  670200.0 1069200.0 680400.0 1083000.0 ;
      RECT  670200.0 1096800.0 680400.0 1083000.0 ;
      RECT  670200.0 1096800.0 680400.0 1110600.0 ;
      RECT  670200.0 1124400.0 680400.0 1110600.0 ;
      RECT  670200.0 1124400.0 680400.0 1138200.0 ;
      RECT  670200.0 1152000.0 680400.0 1138200.0 ;
      RECT  670200.0 1152000.0 680400.0 1165800.0 ;
      RECT  670200.0 1179600.0 680400.0 1165800.0 ;
      RECT  670200.0 1179600.0 680400.0 1193400.0 ;
      RECT  670200.0 1207200.0 680400.0 1193400.0 ;
      RECT  670200.0 1207200.0 680400.0 1221000.0 ;
      RECT  670200.0 1234800.0 680400.0 1221000.0 ;
      RECT  670200.0 1234800.0 680400.0 1248600.0 ;
      RECT  670200.0 1262400.0 680400.0 1248600.0 ;
      RECT  670200.0 1262400.0 680400.0 1276200.0 ;
      RECT  670200.0 1290000.0 680400.0 1276200.0 ;
      RECT  670200.0 1290000.0 680400.0 1303800.0 ;
      RECT  670200.0 1317600.0 680400.0 1303800.0 ;
      RECT  670200.0 1317600.0 680400.0 1331400.0 ;
      RECT  670200.0 1345200.0 680400.0 1331400.0 ;
      RECT  670200.0 1345200.0 680400.0 1359000.0 ;
      RECT  670200.0 1372800.0 680400.0 1359000.0 ;
      RECT  670200.0 1372800.0 680400.0 1386600.0 ;
      RECT  670200.0 1400400.0 680400.0 1386600.0 ;
      RECT  670200.0 1400400.0 680400.0 1414200.0 ;
      RECT  670200.0 1428000.0 680400.0 1414200.0 ;
      RECT  670200.0 1428000.0 680400.0 1441800.0 ;
      RECT  670200.0 1455600.0 680400.0 1441800.0 ;
      RECT  670200.0 1455600.0 680400.0 1469400.0 ;
      RECT  670200.0 1483200.0 680400.0 1469400.0 ;
      RECT  670200.0 1483200.0 680400.0 1497000.0 ;
      RECT  670200.0 1510800.0 680400.0 1497000.0 ;
      RECT  670200.0 1510800.0 680400.0 1524600.0 ;
      RECT  670200.0 1538400.0 680400.0 1524600.0 ;
      RECT  670200.0 1538400.0 680400.0 1552200.0 ;
      RECT  670200.0 1566000.0 680400.0 1552200.0 ;
      RECT  670200.0 1566000.0 680400.0 1579800.0 ;
      RECT  670200.0 1593600.0 680400.0 1579800.0 ;
      RECT  670200.0 1593600.0 680400.0 1607400.0 ;
      RECT  670200.0 1621200.0 680400.0 1607400.0 ;
      RECT  670200.0 1621200.0 680400.0 1635000.0 ;
      RECT  670200.0 1648800.0 680400.0 1635000.0 ;
      RECT  670200.0 1648800.0 680400.0 1662600.0 ;
      RECT  670200.0 1676400.0 680400.0 1662600.0 ;
      RECT  670200.0 1676400.0 680400.0 1690200.0 ;
      RECT  670200.0 1704000.0 680400.0 1690200.0 ;
      RECT  670200.0 1704000.0 680400.0 1717800.0 ;
      RECT  670200.0 1731600.0 680400.0 1717800.0 ;
      RECT  670200.0 1731600.0 680400.0 1745400.0 ;
      RECT  670200.0 1759200.0 680400.0 1745400.0 ;
      RECT  670200.0 1759200.0 680400.0 1773000.0 ;
      RECT  670200.0 1786800.0 680400.0 1773000.0 ;
      RECT  670200.0 1786800.0 680400.0 1800600.0 ;
      RECT  670200.0 1814400.0 680400.0 1800600.0 ;
      RECT  670200.0 1814400.0 680400.0 1828200.0 ;
      RECT  670200.0 1842000.0 680400.0 1828200.0 ;
      RECT  670200.0 1842000.0 680400.0 1855800.0 ;
      RECT  670200.0 1869600.0 680400.0 1855800.0 ;
      RECT  670200.0 1869600.0 680400.0 1883400.0 ;
      RECT  670200.0 1897200.0 680400.0 1883400.0 ;
      RECT  670200.0 1897200.0 680400.0 1911000.0 ;
      RECT  670200.0 1924800.0 680400.0 1911000.0 ;
      RECT  670200.0 1924800.0 680400.0 1938600.0 ;
      RECT  670200.0 1952400.0 680400.0 1938600.0 ;
      RECT  670200.0 1952400.0 680400.0 1966200.0 ;
      RECT  670200.0 1980000.0 680400.0 1966200.0 ;
      RECT  670200.0 1980000.0 680400.0 1993800.0 ;
      RECT  670200.0 2007600.0 680400.0 1993800.0 ;
      RECT  670200.0 2007600.0 680400.0 2021400.0 ;
      RECT  670200.0 2035200.0 680400.0 2021400.0 ;
      RECT  670200.0 2035200.0 680400.0 2049000.0 ;
      RECT  670200.0 2062800.0 680400.0 2049000.0 ;
      RECT  670200.0 2062800.0 680400.0 2076600.0 ;
      RECT  670200.0 2090400.0 680400.0 2076600.0 ;
      RECT  670200.0 2090400.0 680400.0 2104200.0 ;
      RECT  670200.0 2118000.0 680400.0 2104200.0 ;
      RECT  670200.0 2118000.0 680400.0 2131800.0 ;
      RECT  670200.0 2145600.0 680400.0 2131800.0 ;
      RECT  680400.0 379200.0 690600.0 393000.0 ;
      RECT  680400.0 406800.0 690600.0 393000.0 ;
      RECT  680400.0 406800.0 690600.0 420600.0 ;
      RECT  680400.0 434400.0 690600.0 420600.0 ;
      RECT  680400.0 434400.0 690600.0 448200.0 ;
      RECT  680400.0 462000.0 690600.0 448200.0 ;
      RECT  680400.0 462000.0 690600.0 475800.0 ;
      RECT  680400.0 489600.0 690600.0 475800.0 ;
      RECT  680400.0 489600.0 690600.0 503400.0 ;
      RECT  680400.0 517200.0 690600.0 503400.0 ;
      RECT  680400.0 517200.0 690600.0 531000.0 ;
      RECT  680400.0 544800.0 690600.0 531000.0 ;
      RECT  680400.0 544800.0 690600.0 558600.0 ;
      RECT  680400.0 572400.0 690600.0 558600.0 ;
      RECT  680400.0 572400.0 690600.0 586200.0 ;
      RECT  680400.0 600000.0 690600.0 586200.0 ;
      RECT  680400.0 600000.0 690600.0 613800.0 ;
      RECT  680400.0 627600.0 690600.0 613800.0 ;
      RECT  680400.0 627600.0 690600.0 641400.0 ;
      RECT  680400.0 655200.0 690600.0 641400.0 ;
      RECT  680400.0 655200.0 690600.0 669000.0 ;
      RECT  680400.0 682800.0 690600.0 669000.0 ;
      RECT  680400.0 682800.0 690600.0 696600.0 ;
      RECT  680400.0 710400.0 690600.0 696600.0 ;
      RECT  680400.0 710400.0 690600.0 724200.0 ;
      RECT  680400.0 738000.0 690600.0 724200.0 ;
      RECT  680400.0 738000.0 690600.0 751800.0 ;
      RECT  680400.0 765600.0 690600.0 751800.0 ;
      RECT  680400.0 765600.0 690600.0 779400.0 ;
      RECT  680400.0 793200.0 690600.0 779400.0 ;
      RECT  680400.0 793200.0 690600.0 807000.0 ;
      RECT  680400.0 820800.0 690600.0 807000.0 ;
      RECT  680400.0 820800.0 690600.0 834600.0 ;
      RECT  680400.0 848400.0 690600.0 834600.0 ;
      RECT  680400.0 848400.0 690600.0 862200.0 ;
      RECT  680400.0 876000.0 690600.0 862200.0 ;
      RECT  680400.0 876000.0 690600.0 889800.0 ;
      RECT  680400.0 903600.0 690600.0 889800.0 ;
      RECT  680400.0 903600.0 690600.0 917400.0 ;
      RECT  680400.0 931200.0 690600.0 917400.0 ;
      RECT  680400.0 931200.0 690600.0 945000.0 ;
      RECT  680400.0 958800.0 690600.0 945000.0 ;
      RECT  680400.0 958800.0 690600.0 972600.0 ;
      RECT  680400.0 986400.0 690600.0 972600.0 ;
      RECT  680400.0 986400.0 690600.0 1000200.0 ;
      RECT  680400.0 1014000.0 690600.0 1000200.0 ;
      RECT  680400.0 1014000.0 690600.0 1027800.0 ;
      RECT  680400.0 1041600.0 690600.0 1027800.0 ;
      RECT  680400.0 1041600.0 690600.0 1055400.0 ;
      RECT  680400.0 1069200.0 690600.0 1055400.0 ;
      RECT  680400.0 1069200.0 690600.0 1083000.0 ;
      RECT  680400.0 1096800.0 690600.0 1083000.0 ;
      RECT  680400.0 1096800.0 690600.0 1110600.0 ;
      RECT  680400.0 1124400.0 690600.0 1110600.0 ;
      RECT  680400.0 1124400.0 690600.0 1138200.0 ;
      RECT  680400.0 1152000.0 690600.0 1138200.0 ;
      RECT  680400.0 1152000.0 690600.0 1165800.0 ;
      RECT  680400.0 1179600.0 690600.0 1165800.0 ;
      RECT  680400.0 1179600.0 690600.0 1193400.0 ;
      RECT  680400.0 1207200.0 690600.0 1193400.0 ;
      RECT  680400.0 1207200.0 690600.0 1221000.0 ;
      RECT  680400.0 1234800.0 690600.0 1221000.0 ;
      RECT  680400.0 1234800.0 690600.0 1248600.0 ;
      RECT  680400.0 1262400.0 690600.0 1248600.0 ;
      RECT  680400.0 1262400.0 690600.0 1276200.0 ;
      RECT  680400.0 1290000.0 690600.0 1276200.0 ;
      RECT  680400.0 1290000.0 690600.0 1303800.0 ;
      RECT  680400.0 1317600.0 690600.0 1303800.0 ;
      RECT  680400.0 1317600.0 690600.0 1331400.0 ;
      RECT  680400.0 1345200.0 690600.0 1331400.0 ;
      RECT  680400.0 1345200.0 690600.0 1359000.0 ;
      RECT  680400.0 1372800.0 690600.0 1359000.0 ;
      RECT  680400.0 1372800.0 690600.0 1386600.0 ;
      RECT  680400.0 1400400.0 690600.0 1386600.0 ;
      RECT  680400.0 1400400.0 690600.0 1414200.0 ;
      RECT  680400.0 1428000.0 690600.0 1414200.0 ;
      RECT  680400.0 1428000.0 690600.0 1441800.0 ;
      RECT  680400.0 1455600.0 690600.0 1441800.0 ;
      RECT  680400.0 1455600.0 690600.0 1469400.0 ;
      RECT  680400.0 1483200.0 690600.0 1469400.0 ;
      RECT  680400.0 1483200.0 690600.0 1497000.0 ;
      RECT  680400.0 1510800.0 690600.0 1497000.0 ;
      RECT  680400.0 1510800.0 690600.0 1524600.0 ;
      RECT  680400.0 1538400.0 690600.0 1524600.0 ;
      RECT  680400.0 1538400.0 690600.0 1552200.0 ;
      RECT  680400.0 1566000.0 690600.0 1552200.0 ;
      RECT  680400.0 1566000.0 690600.0 1579800.0 ;
      RECT  680400.0 1593600.0 690600.0 1579800.0 ;
      RECT  680400.0 1593600.0 690600.0 1607400.0 ;
      RECT  680400.0 1621200.0 690600.0 1607400.0 ;
      RECT  680400.0 1621200.0 690600.0 1635000.0 ;
      RECT  680400.0 1648800.0 690600.0 1635000.0 ;
      RECT  680400.0 1648800.0 690600.0 1662600.0 ;
      RECT  680400.0 1676400.0 690600.0 1662600.0 ;
      RECT  680400.0 1676400.0 690600.0 1690200.0 ;
      RECT  680400.0 1704000.0 690600.0 1690200.0 ;
      RECT  680400.0 1704000.0 690600.0 1717800.0 ;
      RECT  680400.0 1731600.0 690600.0 1717800.0 ;
      RECT  680400.0 1731600.0 690600.0 1745400.0 ;
      RECT  680400.0 1759200.0 690600.0 1745400.0 ;
      RECT  680400.0 1759200.0 690600.0 1773000.0 ;
      RECT  680400.0 1786800.0 690600.0 1773000.0 ;
      RECT  680400.0 1786800.0 690600.0 1800600.0 ;
      RECT  680400.0 1814400.0 690600.0 1800600.0 ;
      RECT  680400.0 1814400.0 690600.0 1828200.0 ;
      RECT  680400.0 1842000.0 690600.0 1828200.0 ;
      RECT  680400.0 1842000.0 690600.0 1855800.0 ;
      RECT  680400.0 1869600.0 690600.0 1855800.0 ;
      RECT  680400.0 1869600.0 690600.0 1883400.0 ;
      RECT  680400.0 1897200.0 690600.0 1883400.0 ;
      RECT  680400.0 1897200.0 690600.0 1911000.0 ;
      RECT  680400.0 1924800.0 690600.0 1911000.0 ;
      RECT  680400.0 1924800.0 690600.0 1938600.0 ;
      RECT  680400.0 1952400.0 690600.0 1938600.0 ;
      RECT  680400.0 1952400.0 690600.0 1966200.0 ;
      RECT  680400.0 1980000.0 690600.0 1966200.0 ;
      RECT  680400.0 1980000.0 690600.0 1993800.0 ;
      RECT  680400.0 2007600.0 690600.0 1993800.0 ;
      RECT  680400.0 2007600.0 690600.0 2021400.0 ;
      RECT  680400.0 2035200.0 690600.0 2021400.0 ;
      RECT  680400.0 2035200.0 690600.0 2049000.0 ;
      RECT  680400.0 2062800.0 690600.0 2049000.0 ;
      RECT  680400.0 2062800.0 690600.0 2076600.0 ;
      RECT  680400.0 2090400.0 690600.0 2076600.0 ;
      RECT  680400.0 2090400.0 690600.0 2104200.0 ;
      RECT  680400.0 2118000.0 690600.0 2104200.0 ;
      RECT  680400.0 2118000.0 690600.0 2131800.0 ;
      RECT  680400.0 2145600.0 690600.0 2131800.0 ;
      RECT  690600.0 379200.0 700800.0 393000.0 ;
      RECT  690600.0 406800.0 700800.0 393000.0 ;
      RECT  690600.0 406800.0 700800.0 420600.0 ;
      RECT  690600.0 434400.0 700800.0 420600.0 ;
      RECT  690600.0 434400.0 700800.0 448200.0 ;
      RECT  690600.0 462000.0 700800.0 448200.0 ;
      RECT  690600.0 462000.0 700800.0 475800.0 ;
      RECT  690600.0 489600.0 700800.0 475800.0 ;
      RECT  690600.0 489600.0 700800.0 503400.0 ;
      RECT  690600.0 517200.0 700800.0 503400.0 ;
      RECT  690600.0 517200.0 700800.0 531000.0 ;
      RECT  690600.0 544800.0 700800.0 531000.0 ;
      RECT  690600.0 544800.0 700800.0 558600.0 ;
      RECT  690600.0 572400.0 700800.0 558600.0 ;
      RECT  690600.0 572400.0 700800.0 586200.0 ;
      RECT  690600.0 600000.0 700800.0 586200.0 ;
      RECT  690600.0 600000.0 700800.0 613800.0 ;
      RECT  690600.0 627600.0 700800.0 613800.0 ;
      RECT  690600.0 627600.0 700800.0 641400.0 ;
      RECT  690600.0 655200.0 700800.0 641400.0 ;
      RECT  690600.0 655200.0 700800.0 669000.0 ;
      RECT  690600.0 682800.0 700800.0 669000.0 ;
      RECT  690600.0 682800.0 700800.0 696600.0 ;
      RECT  690600.0 710400.0 700800.0 696600.0 ;
      RECT  690600.0 710400.0 700800.0 724200.0 ;
      RECT  690600.0 738000.0 700800.0 724200.0 ;
      RECT  690600.0 738000.0 700800.0 751800.0 ;
      RECT  690600.0 765600.0 700800.0 751800.0 ;
      RECT  690600.0 765600.0 700800.0 779400.0 ;
      RECT  690600.0 793200.0 700800.0 779400.0 ;
      RECT  690600.0 793200.0 700800.0 807000.0 ;
      RECT  690600.0 820800.0 700800.0 807000.0 ;
      RECT  690600.0 820800.0 700800.0 834600.0 ;
      RECT  690600.0 848400.0 700800.0 834600.0 ;
      RECT  690600.0 848400.0 700800.0 862200.0 ;
      RECT  690600.0 876000.0 700800.0 862200.0 ;
      RECT  690600.0 876000.0 700800.0 889800.0 ;
      RECT  690600.0 903600.0 700800.0 889800.0 ;
      RECT  690600.0 903600.0 700800.0 917400.0 ;
      RECT  690600.0 931200.0 700800.0 917400.0 ;
      RECT  690600.0 931200.0 700800.0 945000.0 ;
      RECT  690600.0 958800.0 700800.0 945000.0 ;
      RECT  690600.0 958800.0 700800.0 972600.0 ;
      RECT  690600.0 986400.0 700800.0 972600.0 ;
      RECT  690600.0 986400.0 700800.0 1000200.0 ;
      RECT  690600.0 1014000.0 700800.0 1000200.0 ;
      RECT  690600.0 1014000.0 700800.0 1027800.0 ;
      RECT  690600.0 1041600.0 700800.0 1027800.0 ;
      RECT  690600.0 1041600.0 700800.0 1055400.0 ;
      RECT  690600.0 1069200.0 700800.0 1055400.0 ;
      RECT  690600.0 1069200.0 700800.0 1083000.0 ;
      RECT  690600.0 1096800.0 700800.0 1083000.0 ;
      RECT  690600.0 1096800.0 700800.0 1110600.0 ;
      RECT  690600.0 1124400.0 700800.0 1110600.0 ;
      RECT  690600.0 1124400.0 700800.0 1138200.0 ;
      RECT  690600.0 1152000.0 700800.0 1138200.0 ;
      RECT  690600.0 1152000.0 700800.0 1165800.0 ;
      RECT  690600.0 1179600.0 700800.0 1165800.0 ;
      RECT  690600.0 1179600.0 700800.0 1193400.0 ;
      RECT  690600.0 1207200.0 700800.0 1193400.0 ;
      RECT  690600.0 1207200.0 700800.0 1221000.0 ;
      RECT  690600.0 1234800.0 700800.0 1221000.0 ;
      RECT  690600.0 1234800.0 700800.0 1248600.0 ;
      RECT  690600.0 1262400.0 700800.0 1248600.0 ;
      RECT  690600.0 1262400.0 700800.0 1276200.0 ;
      RECT  690600.0 1290000.0 700800.0 1276200.0 ;
      RECT  690600.0 1290000.0 700800.0 1303800.0 ;
      RECT  690600.0 1317600.0 700800.0 1303800.0 ;
      RECT  690600.0 1317600.0 700800.0 1331400.0 ;
      RECT  690600.0 1345200.0 700800.0 1331400.0 ;
      RECT  690600.0 1345200.0 700800.0 1359000.0 ;
      RECT  690600.0 1372800.0 700800.0 1359000.0 ;
      RECT  690600.0 1372800.0 700800.0 1386600.0 ;
      RECT  690600.0 1400400.0 700800.0 1386600.0 ;
      RECT  690600.0 1400400.0 700800.0 1414200.0 ;
      RECT  690600.0 1428000.0 700800.0 1414200.0 ;
      RECT  690600.0 1428000.0 700800.0 1441800.0 ;
      RECT  690600.0 1455600.0 700800.0 1441800.0 ;
      RECT  690600.0 1455600.0 700800.0 1469400.0 ;
      RECT  690600.0 1483200.0 700800.0 1469400.0 ;
      RECT  690600.0 1483200.0 700800.0 1497000.0 ;
      RECT  690600.0 1510800.0 700800.0 1497000.0 ;
      RECT  690600.0 1510800.0 700800.0 1524600.0 ;
      RECT  690600.0 1538400.0 700800.0 1524600.0 ;
      RECT  690600.0 1538400.0 700800.0 1552200.0 ;
      RECT  690600.0 1566000.0 700800.0 1552200.0 ;
      RECT  690600.0 1566000.0 700800.0 1579800.0 ;
      RECT  690600.0 1593600.0 700800.0 1579800.0 ;
      RECT  690600.0 1593600.0 700800.0 1607400.0 ;
      RECT  690600.0 1621200.0 700800.0 1607400.0 ;
      RECT  690600.0 1621200.0 700800.0 1635000.0 ;
      RECT  690600.0 1648800.0 700800.0 1635000.0 ;
      RECT  690600.0 1648800.0 700800.0 1662600.0 ;
      RECT  690600.0 1676400.0 700800.0 1662600.0 ;
      RECT  690600.0 1676400.0 700800.0 1690200.0 ;
      RECT  690600.0 1704000.0 700800.0 1690200.0 ;
      RECT  690600.0 1704000.0 700800.0 1717800.0 ;
      RECT  690600.0 1731600.0 700800.0 1717800.0 ;
      RECT  690600.0 1731600.0 700800.0 1745400.0 ;
      RECT  690600.0 1759200.0 700800.0 1745400.0 ;
      RECT  690600.0 1759200.0 700800.0 1773000.0 ;
      RECT  690600.0 1786800.0 700800.0 1773000.0 ;
      RECT  690600.0 1786800.0 700800.0 1800600.0 ;
      RECT  690600.0 1814400.0 700800.0 1800600.0 ;
      RECT  690600.0 1814400.0 700800.0 1828200.0 ;
      RECT  690600.0 1842000.0 700800.0 1828200.0 ;
      RECT  690600.0 1842000.0 700800.0 1855800.0 ;
      RECT  690600.0 1869600.0 700800.0 1855800.0 ;
      RECT  690600.0 1869600.0 700800.0 1883400.0 ;
      RECT  690600.0 1897200.0 700800.0 1883400.0 ;
      RECT  690600.0 1897200.0 700800.0 1911000.0 ;
      RECT  690600.0 1924800.0 700800.0 1911000.0 ;
      RECT  690600.0 1924800.0 700800.0 1938600.0 ;
      RECT  690600.0 1952400.0 700800.0 1938600.0 ;
      RECT  690600.0 1952400.0 700800.0 1966200.0 ;
      RECT  690600.0 1980000.0 700800.0 1966200.0 ;
      RECT  690600.0 1980000.0 700800.0 1993800.0 ;
      RECT  690600.0 2007600.0 700800.0 1993800.0 ;
      RECT  690600.0 2007600.0 700800.0 2021400.0 ;
      RECT  690600.0 2035200.0 700800.0 2021400.0 ;
      RECT  690600.0 2035200.0 700800.0 2049000.0 ;
      RECT  690600.0 2062800.0 700800.0 2049000.0 ;
      RECT  690600.0 2062800.0 700800.0 2076600.0 ;
      RECT  690600.0 2090400.0 700800.0 2076600.0 ;
      RECT  690600.0 2090400.0 700800.0 2104200.0 ;
      RECT  690600.0 2118000.0 700800.0 2104200.0 ;
      RECT  690600.0 2118000.0 700800.0 2131800.0 ;
      RECT  690600.0 2145600.0 700800.0 2131800.0 ;
      RECT  700800.0 379200.0 711000.0 393000.0 ;
      RECT  700800.0 406800.0 711000.0 393000.0 ;
      RECT  700800.0 406800.0 711000.0 420600.0 ;
      RECT  700800.0 434400.0 711000.0 420600.0 ;
      RECT  700800.0 434400.0 711000.0 448200.0 ;
      RECT  700800.0 462000.0 711000.0 448200.0 ;
      RECT  700800.0 462000.0 711000.0 475800.0 ;
      RECT  700800.0 489600.0 711000.0 475800.0 ;
      RECT  700800.0 489600.0 711000.0 503400.0 ;
      RECT  700800.0 517200.0 711000.0 503400.0 ;
      RECT  700800.0 517200.0 711000.0 531000.0 ;
      RECT  700800.0 544800.0 711000.0 531000.0 ;
      RECT  700800.0 544800.0 711000.0 558600.0 ;
      RECT  700800.0 572400.0 711000.0 558600.0 ;
      RECT  700800.0 572400.0 711000.0 586200.0 ;
      RECT  700800.0 600000.0 711000.0 586200.0 ;
      RECT  700800.0 600000.0 711000.0 613800.0 ;
      RECT  700800.0 627600.0 711000.0 613800.0 ;
      RECT  700800.0 627600.0 711000.0 641400.0 ;
      RECT  700800.0 655200.0 711000.0 641400.0 ;
      RECT  700800.0 655200.0 711000.0 669000.0 ;
      RECT  700800.0 682800.0 711000.0 669000.0 ;
      RECT  700800.0 682800.0 711000.0 696600.0 ;
      RECT  700800.0 710400.0 711000.0 696600.0 ;
      RECT  700800.0 710400.0 711000.0 724200.0 ;
      RECT  700800.0 738000.0 711000.0 724200.0 ;
      RECT  700800.0 738000.0 711000.0 751800.0 ;
      RECT  700800.0 765600.0 711000.0 751800.0 ;
      RECT  700800.0 765600.0 711000.0 779400.0 ;
      RECT  700800.0 793200.0 711000.0 779400.0 ;
      RECT  700800.0 793200.0 711000.0 807000.0 ;
      RECT  700800.0 820800.0 711000.0 807000.0 ;
      RECT  700800.0 820800.0 711000.0 834600.0 ;
      RECT  700800.0 848400.0 711000.0 834600.0 ;
      RECT  700800.0 848400.0 711000.0 862200.0 ;
      RECT  700800.0 876000.0 711000.0 862200.0 ;
      RECT  700800.0 876000.0 711000.0 889800.0 ;
      RECT  700800.0 903600.0 711000.0 889800.0 ;
      RECT  700800.0 903600.0 711000.0 917400.0 ;
      RECT  700800.0 931200.0 711000.0 917400.0 ;
      RECT  700800.0 931200.0 711000.0 945000.0 ;
      RECT  700800.0 958800.0 711000.0 945000.0 ;
      RECT  700800.0 958800.0 711000.0 972600.0 ;
      RECT  700800.0 986400.0 711000.0 972600.0 ;
      RECT  700800.0 986400.0 711000.0 1000200.0 ;
      RECT  700800.0 1014000.0 711000.0 1000200.0 ;
      RECT  700800.0 1014000.0 711000.0 1027800.0 ;
      RECT  700800.0 1041600.0 711000.0 1027800.0 ;
      RECT  700800.0 1041600.0 711000.0 1055400.0 ;
      RECT  700800.0 1069200.0 711000.0 1055400.0 ;
      RECT  700800.0 1069200.0 711000.0 1083000.0 ;
      RECT  700800.0 1096800.0 711000.0 1083000.0 ;
      RECT  700800.0 1096800.0 711000.0 1110600.0 ;
      RECT  700800.0 1124400.0 711000.0 1110600.0 ;
      RECT  700800.0 1124400.0 711000.0 1138200.0 ;
      RECT  700800.0 1152000.0 711000.0 1138200.0 ;
      RECT  700800.0 1152000.0 711000.0 1165800.0 ;
      RECT  700800.0 1179600.0 711000.0 1165800.0 ;
      RECT  700800.0 1179600.0 711000.0 1193400.0 ;
      RECT  700800.0 1207200.0 711000.0 1193400.0 ;
      RECT  700800.0 1207200.0 711000.0 1221000.0 ;
      RECT  700800.0 1234800.0 711000.0 1221000.0 ;
      RECT  700800.0 1234800.0 711000.0 1248600.0 ;
      RECT  700800.0 1262400.0 711000.0 1248600.0 ;
      RECT  700800.0 1262400.0 711000.0 1276200.0 ;
      RECT  700800.0 1290000.0 711000.0 1276200.0 ;
      RECT  700800.0 1290000.0 711000.0 1303800.0 ;
      RECT  700800.0 1317600.0 711000.0 1303800.0 ;
      RECT  700800.0 1317600.0 711000.0 1331400.0 ;
      RECT  700800.0 1345200.0 711000.0 1331400.0 ;
      RECT  700800.0 1345200.0 711000.0 1359000.0 ;
      RECT  700800.0 1372800.0 711000.0 1359000.0 ;
      RECT  700800.0 1372800.0 711000.0 1386600.0 ;
      RECT  700800.0 1400400.0 711000.0 1386600.0 ;
      RECT  700800.0 1400400.0 711000.0 1414200.0 ;
      RECT  700800.0 1428000.0 711000.0 1414200.0 ;
      RECT  700800.0 1428000.0 711000.0 1441800.0 ;
      RECT  700800.0 1455600.0 711000.0 1441800.0 ;
      RECT  700800.0 1455600.0 711000.0 1469400.0 ;
      RECT  700800.0 1483200.0 711000.0 1469400.0 ;
      RECT  700800.0 1483200.0 711000.0 1497000.0 ;
      RECT  700800.0 1510800.0 711000.0 1497000.0 ;
      RECT  700800.0 1510800.0 711000.0 1524600.0 ;
      RECT  700800.0 1538400.0 711000.0 1524600.0 ;
      RECT  700800.0 1538400.0 711000.0 1552200.0 ;
      RECT  700800.0 1566000.0 711000.0 1552200.0 ;
      RECT  700800.0 1566000.0 711000.0 1579800.0 ;
      RECT  700800.0 1593600.0 711000.0 1579800.0 ;
      RECT  700800.0 1593600.0 711000.0 1607400.0 ;
      RECT  700800.0 1621200.0 711000.0 1607400.0 ;
      RECT  700800.0 1621200.0 711000.0 1635000.0 ;
      RECT  700800.0 1648800.0 711000.0 1635000.0 ;
      RECT  700800.0 1648800.0 711000.0 1662600.0 ;
      RECT  700800.0 1676400.0 711000.0 1662600.0 ;
      RECT  700800.0 1676400.0 711000.0 1690200.0 ;
      RECT  700800.0 1704000.0 711000.0 1690200.0 ;
      RECT  700800.0 1704000.0 711000.0 1717800.0 ;
      RECT  700800.0 1731600.0 711000.0 1717800.0 ;
      RECT  700800.0 1731600.0 711000.0 1745400.0 ;
      RECT  700800.0 1759200.0 711000.0 1745400.0 ;
      RECT  700800.0 1759200.0 711000.0 1773000.0 ;
      RECT  700800.0 1786800.0 711000.0 1773000.0 ;
      RECT  700800.0 1786800.0 711000.0 1800600.0 ;
      RECT  700800.0 1814400.0 711000.0 1800600.0 ;
      RECT  700800.0 1814400.0 711000.0 1828200.0 ;
      RECT  700800.0 1842000.0 711000.0 1828200.0 ;
      RECT  700800.0 1842000.0 711000.0 1855800.0 ;
      RECT  700800.0 1869600.0 711000.0 1855800.0 ;
      RECT  700800.0 1869600.0 711000.0 1883400.0 ;
      RECT  700800.0 1897200.0 711000.0 1883400.0 ;
      RECT  700800.0 1897200.0 711000.0 1911000.0 ;
      RECT  700800.0 1924800.0 711000.0 1911000.0 ;
      RECT  700800.0 1924800.0 711000.0 1938600.0 ;
      RECT  700800.0 1952400.0 711000.0 1938600.0 ;
      RECT  700800.0 1952400.0 711000.0 1966200.0 ;
      RECT  700800.0 1980000.0 711000.0 1966200.0 ;
      RECT  700800.0 1980000.0 711000.0 1993800.0 ;
      RECT  700800.0 2007600.0 711000.0 1993800.0 ;
      RECT  700800.0 2007600.0 711000.0 2021400.0 ;
      RECT  700800.0 2035200.0 711000.0 2021400.0 ;
      RECT  700800.0 2035200.0 711000.0 2049000.0 ;
      RECT  700800.0 2062800.0 711000.0 2049000.0 ;
      RECT  700800.0 2062800.0 711000.0 2076600.0 ;
      RECT  700800.0 2090400.0 711000.0 2076600.0 ;
      RECT  700800.0 2090400.0 711000.0 2104200.0 ;
      RECT  700800.0 2118000.0 711000.0 2104200.0 ;
      RECT  700800.0 2118000.0 711000.0 2131800.0 ;
      RECT  700800.0 2145600.0 711000.0 2131800.0 ;
      RECT  711000.0 379200.0 721200.0 393000.0 ;
      RECT  711000.0 406800.0 721200.0 393000.0 ;
      RECT  711000.0 406800.0 721200.0 420600.0 ;
      RECT  711000.0 434400.0 721200.0 420600.0 ;
      RECT  711000.0 434400.0 721200.0 448200.0 ;
      RECT  711000.0 462000.0 721200.0 448200.0 ;
      RECT  711000.0 462000.0 721200.0 475800.0 ;
      RECT  711000.0 489600.0 721200.0 475800.0 ;
      RECT  711000.0 489600.0 721200.0 503400.0 ;
      RECT  711000.0 517200.0 721200.0 503400.0 ;
      RECT  711000.0 517200.0 721200.0 531000.0 ;
      RECT  711000.0 544800.0 721200.0 531000.0 ;
      RECT  711000.0 544800.0 721200.0 558600.0 ;
      RECT  711000.0 572400.0 721200.0 558600.0 ;
      RECT  711000.0 572400.0 721200.0 586200.0 ;
      RECT  711000.0 600000.0 721200.0 586200.0 ;
      RECT  711000.0 600000.0 721200.0 613800.0 ;
      RECT  711000.0 627600.0 721200.0 613800.0 ;
      RECT  711000.0 627600.0 721200.0 641400.0 ;
      RECT  711000.0 655200.0 721200.0 641400.0 ;
      RECT  711000.0 655200.0 721200.0 669000.0 ;
      RECT  711000.0 682800.0 721200.0 669000.0 ;
      RECT  711000.0 682800.0 721200.0 696600.0 ;
      RECT  711000.0 710400.0 721200.0 696600.0 ;
      RECT  711000.0 710400.0 721200.0 724200.0 ;
      RECT  711000.0 738000.0 721200.0 724200.0 ;
      RECT  711000.0 738000.0 721200.0 751800.0 ;
      RECT  711000.0 765600.0 721200.0 751800.0 ;
      RECT  711000.0 765600.0 721200.0 779400.0 ;
      RECT  711000.0 793200.0 721200.0 779400.0 ;
      RECT  711000.0 793200.0 721200.0 807000.0 ;
      RECT  711000.0 820800.0 721200.0 807000.0 ;
      RECT  711000.0 820800.0 721200.0 834600.0 ;
      RECT  711000.0 848400.0 721200.0 834600.0 ;
      RECT  711000.0 848400.0 721200.0 862200.0 ;
      RECT  711000.0 876000.0 721200.0 862200.0 ;
      RECT  711000.0 876000.0 721200.0 889800.0 ;
      RECT  711000.0 903600.0 721200.0 889800.0 ;
      RECT  711000.0 903600.0 721200.0 917400.0 ;
      RECT  711000.0 931200.0 721200.0 917400.0 ;
      RECT  711000.0 931200.0 721200.0 945000.0 ;
      RECT  711000.0 958800.0 721200.0 945000.0 ;
      RECT  711000.0 958800.0 721200.0 972600.0 ;
      RECT  711000.0 986400.0 721200.0 972600.0 ;
      RECT  711000.0 986400.0 721200.0 1000200.0 ;
      RECT  711000.0 1014000.0 721200.0 1000200.0 ;
      RECT  711000.0 1014000.0 721200.0 1027800.0 ;
      RECT  711000.0 1041600.0 721200.0 1027800.0 ;
      RECT  711000.0 1041600.0 721200.0 1055400.0 ;
      RECT  711000.0 1069200.0 721200.0 1055400.0 ;
      RECT  711000.0 1069200.0 721200.0 1083000.0 ;
      RECT  711000.0 1096800.0 721200.0 1083000.0 ;
      RECT  711000.0 1096800.0 721200.0 1110600.0 ;
      RECT  711000.0 1124400.0 721200.0 1110600.0 ;
      RECT  711000.0 1124400.0 721200.0 1138200.0 ;
      RECT  711000.0 1152000.0 721200.0 1138200.0 ;
      RECT  711000.0 1152000.0 721200.0 1165800.0 ;
      RECT  711000.0 1179600.0 721200.0 1165800.0 ;
      RECT  711000.0 1179600.0 721200.0 1193400.0 ;
      RECT  711000.0 1207200.0 721200.0 1193400.0 ;
      RECT  711000.0 1207200.0 721200.0 1221000.0 ;
      RECT  711000.0 1234800.0 721200.0 1221000.0 ;
      RECT  711000.0 1234800.0 721200.0 1248600.0 ;
      RECT  711000.0 1262400.0 721200.0 1248600.0 ;
      RECT  711000.0 1262400.0 721200.0 1276200.0 ;
      RECT  711000.0 1290000.0 721200.0 1276200.0 ;
      RECT  711000.0 1290000.0 721200.0 1303800.0 ;
      RECT  711000.0 1317600.0 721200.0 1303800.0 ;
      RECT  711000.0 1317600.0 721200.0 1331400.0 ;
      RECT  711000.0 1345200.0 721200.0 1331400.0 ;
      RECT  711000.0 1345200.0 721200.0 1359000.0 ;
      RECT  711000.0 1372800.0 721200.0 1359000.0 ;
      RECT  711000.0 1372800.0 721200.0 1386600.0 ;
      RECT  711000.0 1400400.0 721200.0 1386600.0 ;
      RECT  711000.0 1400400.0 721200.0 1414200.0 ;
      RECT  711000.0 1428000.0 721200.0 1414200.0 ;
      RECT  711000.0 1428000.0 721200.0 1441800.0 ;
      RECT  711000.0 1455600.0 721200.0 1441800.0 ;
      RECT  711000.0 1455600.0 721200.0 1469400.0 ;
      RECT  711000.0 1483200.0 721200.0 1469400.0 ;
      RECT  711000.0 1483200.0 721200.0 1497000.0 ;
      RECT  711000.0 1510800.0 721200.0 1497000.0 ;
      RECT  711000.0 1510800.0 721200.0 1524600.0 ;
      RECT  711000.0 1538400.0 721200.0 1524600.0 ;
      RECT  711000.0 1538400.0 721200.0 1552200.0 ;
      RECT  711000.0 1566000.0 721200.0 1552200.0 ;
      RECT  711000.0 1566000.0 721200.0 1579800.0 ;
      RECT  711000.0 1593600.0 721200.0 1579800.0 ;
      RECT  711000.0 1593600.0 721200.0 1607400.0 ;
      RECT  711000.0 1621200.0 721200.0 1607400.0 ;
      RECT  711000.0 1621200.0 721200.0 1635000.0 ;
      RECT  711000.0 1648800.0 721200.0 1635000.0 ;
      RECT  711000.0 1648800.0 721200.0 1662600.0 ;
      RECT  711000.0 1676400.0 721200.0 1662600.0 ;
      RECT  711000.0 1676400.0 721200.0 1690200.0 ;
      RECT  711000.0 1704000.0 721200.0 1690200.0 ;
      RECT  711000.0 1704000.0 721200.0 1717800.0 ;
      RECT  711000.0 1731600.0 721200.0 1717800.0 ;
      RECT  711000.0 1731600.0 721200.0 1745400.0 ;
      RECT  711000.0 1759200.0 721200.0 1745400.0 ;
      RECT  711000.0 1759200.0 721200.0 1773000.0 ;
      RECT  711000.0 1786800.0 721200.0 1773000.0 ;
      RECT  711000.0 1786800.0 721200.0 1800600.0 ;
      RECT  711000.0 1814400.0 721200.0 1800600.0 ;
      RECT  711000.0 1814400.0 721200.0 1828200.0 ;
      RECT  711000.0 1842000.0 721200.0 1828200.0 ;
      RECT  711000.0 1842000.0 721200.0 1855800.0 ;
      RECT  711000.0 1869600.0 721200.0 1855800.0 ;
      RECT  711000.0 1869600.0 721200.0 1883400.0 ;
      RECT  711000.0 1897200.0 721200.0 1883400.0 ;
      RECT  711000.0 1897200.0 721200.0 1911000.0 ;
      RECT  711000.0 1924800.0 721200.0 1911000.0 ;
      RECT  711000.0 1924800.0 721200.0 1938600.0 ;
      RECT  711000.0 1952400.0 721200.0 1938600.0 ;
      RECT  711000.0 1952400.0 721200.0 1966200.0 ;
      RECT  711000.0 1980000.0 721200.0 1966200.0 ;
      RECT  711000.0 1980000.0 721200.0 1993800.0 ;
      RECT  711000.0 2007600.0 721200.0 1993800.0 ;
      RECT  711000.0 2007600.0 721200.0 2021400.0 ;
      RECT  711000.0 2035200.0 721200.0 2021400.0 ;
      RECT  711000.0 2035200.0 721200.0 2049000.0 ;
      RECT  711000.0 2062800.0 721200.0 2049000.0 ;
      RECT  711000.0 2062800.0 721200.0 2076600.0 ;
      RECT  711000.0 2090400.0 721200.0 2076600.0 ;
      RECT  711000.0 2090400.0 721200.0 2104200.0 ;
      RECT  711000.0 2118000.0 721200.0 2104200.0 ;
      RECT  711000.0 2118000.0 721200.0 2131800.0 ;
      RECT  711000.0 2145600.0 721200.0 2131800.0 ;
      RECT  721200.0 379200.0 731400.0 393000.0 ;
      RECT  721200.0 406800.0 731400.0 393000.0 ;
      RECT  721200.0 406800.0 731400.0 420600.0 ;
      RECT  721200.0 434400.0 731400.0 420600.0 ;
      RECT  721200.0 434400.0 731400.0 448200.0 ;
      RECT  721200.0 462000.0 731400.0 448200.0 ;
      RECT  721200.0 462000.0 731400.0 475800.0 ;
      RECT  721200.0 489600.0 731400.0 475800.0 ;
      RECT  721200.0 489600.0 731400.0 503400.0 ;
      RECT  721200.0 517200.0 731400.0 503400.0 ;
      RECT  721200.0 517200.0 731400.0 531000.0 ;
      RECT  721200.0 544800.0 731400.0 531000.0 ;
      RECT  721200.0 544800.0 731400.0 558600.0 ;
      RECT  721200.0 572400.0 731400.0 558600.0 ;
      RECT  721200.0 572400.0 731400.0 586200.0 ;
      RECT  721200.0 600000.0 731400.0 586200.0 ;
      RECT  721200.0 600000.0 731400.0 613800.0 ;
      RECT  721200.0 627600.0 731400.0 613800.0 ;
      RECT  721200.0 627600.0 731400.0 641400.0 ;
      RECT  721200.0 655200.0 731400.0 641400.0 ;
      RECT  721200.0 655200.0 731400.0 669000.0 ;
      RECT  721200.0 682800.0 731400.0 669000.0 ;
      RECT  721200.0 682800.0 731400.0 696600.0 ;
      RECT  721200.0 710400.0 731400.0 696600.0 ;
      RECT  721200.0 710400.0 731400.0 724200.0 ;
      RECT  721200.0 738000.0 731400.0 724200.0 ;
      RECT  721200.0 738000.0 731400.0 751800.0 ;
      RECT  721200.0 765600.0 731400.0 751800.0 ;
      RECT  721200.0 765600.0 731400.0 779400.0 ;
      RECT  721200.0 793200.0 731400.0 779400.0 ;
      RECT  721200.0 793200.0 731400.0 807000.0 ;
      RECT  721200.0 820800.0 731400.0 807000.0 ;
      RECT  721200.0 820800.0 731400.0 834600.0 ;
      RECT  721200.0 848400.0 731400.0 834600.0 ;
      RECT  721200.0 848400.0 731400.0 862200.0 ;
      RECT  721200.0 876000.0 731400.0 862200.0 ;
      RECT  721200.0 876000.0 731400.0 889800.0 ;
      RECT  721200.0 903600.0 731400.0 889800.0 ;
      RECT  721200.0 903600.0 731400.0 917400.0 ;
      RECT  721200.0 931200.0 731400.0 917400.0 ;
      RECT  721200.0 931200.0 731400.0 945000.0 ;
      RECT  721200.0 958800.0 731400.0 945000.0 ;
      RECT  721200.0 958800.0 731400.0 972600.0 ;
      RECT  721200.0 986400.0 731400.0 972600.0 ;
      RECT  721200.0 986400.0 731400.0 1000200.0 ;
      RECT  721200.0 1014000.0 731400.0 1000200.0 ;
      RECT  721200.0 1014000.0 731400.0 1027800.0 ;
      RECT  721200.0 1041600.0 731400.0 1027800.0 ;
      RECT  721200.0 1041600.0 731400.0 1055400.0 ;
      RECT  721200.0 1069200.0 731400.0 1055400.0 ;
      RECT  721200.0 1069200.0 731400.0 1083000.0 ;
      RECT  721200.0 1096800.0 731400.0 1083000.0 ;
      RECT  721200.0 1096800.0 731400.0 1110600.0 ;
      RECT  721200.0 1124400.0 731400.0 1110600.0 ;
      RECT  721200.0 1124400.0 731400.0 1138200.0 ;
      RECT  721200.0 1152000.0 731400.0 1138200.0 ;
      RECT  721200.0 1152000.0 731400.0 1165800.0 ;
      RECT  721200.0 1179600.0 731400.0 1165800.0 ;
      RECT  721200.0 1179600.0 731400.0 1193400.0 ;
      RECT  721200.0 1207200.0 731400.0 1193400.0 ;
      RECT  721200.0 1207200.0 731400.0 1221000.0 ;
      RECT  721200.0 1234800.0 731400.0 1221000.0 ;
      RECT  721200.0 1234800.0 731400.0 1248600.0 ;
      RECT  721200.0 1262400.0 731400.0 1248600.0 ;
      RECT  721200.0 1262400.0 731400.0 1276200.0 ;
      RECT  721200.0 1290000.0 731400.0 1276200.0 ;
      RECT  721200.0 1290000.0 731400.0 1303800.0 ;
      RECT  721200.0 1317600.0 731400.0 1303800.0 ;
      RECT  721200.0 1317600.0 731400.0 1331400.0 ;
      RECT  721200.0 1345200.0 731400.0 1331400.0 ;
      RECT  721200.0 1345200.0 731400.0 1359000.0 ;
      RECT  721200.0 1372800.0 731400.0 1359000.0 ;
      RECT  721200.0 1372800.0 731400.0 1386600.0 ;
      RECT  721200.0 1400400.0 731400.0 1386600.0 ;
      RECT  721200.0 1400400.0 731400.0 1414200.0 ;
      RECT  721200.0 1428000.0 731400.0 1414200.0 ;
      RECT  721200.0 1428000.0 731400.0 1441800.0 ;
      RECT  721200.0 1455600.0 731400.0 1441800.0 ;
      RECT  721200.0 1455600.0 731400.0 1469400.0 ;
      RECT  721200.0 1483200.0 731400.0 1469400.0 ;
      RECT  721200.0 1483200.0 731400.0 1497000.0 ;
      RECT  721200.0 1510800.0 731400.0 1497000.0 ;
      RECT  721200.0 1510800.0 731400.0 1524600.0 ;
      RECT  721200.0 1538400.0 731400.0 1524600.0 ;
      RECT  721200.0 1538400.0 731400.0 1552200.0 ;
      RECT  721200.0 1566000.0 731400.0 1552200.0 ;
      RECT  721200.0 1566000.0 731400.0 1579800.0 ;
      RECT  721200.0 1593600.0 731400.0 1579800.0 ;
      RECT  721200.0 1593600.0 731400.0 1607400.0 ;
      RECT  721200.0 1621200.0 731400.0 1607400.0 ;
      RECT  721200.0 1621200.0 731400.0 1635000.0 ;
      RECT  721200.0 1648800.0 731400.0 1635000.0 ;
      RECT  721200.0 1648800.0 731400.0 1662600.0 ;
      RECT  721200.0 1676400.0 731400.0 1662600.0 ;
      RECT  721200.0 1676400.0 731400.0 1690200.0 ;
      RECT  721200.0 1704000.0 731400.0 1690200.0 ;
      RECT  721200.0 1704000.0 731400.0 1717800.0 ;
      RECT  721200.0 1731600.0 731400.0 1717800.0 ;
      RECT  721200.0 1731600.0 731400.0 1745400.0 ;
      RECT  721200.0 1759200.0 731400.0 1745400.0 ;
      RECT  721200.0 1759200.0 731400.0 1773000.0 ;
      RECT  721200.0 1786800.0 731400.0 1773000.0 ;
      RECT  721200.0 1786800.0 731400.0 1800600.0 ;
      RECT  721200.0 1814400.0 731400.0 1800600.0 ;
      RECT  721200.0 1814400.0 731400.0 1828200.0 ;
      RECT  721200.0 1842000.0 731400.0 1828200.0 ;
      RECT  721200.0 1842000.0 731400.0 1855800.0 ;
      RECT  721200.0 1869600.0 731400.0 1855800.0 ;
      RECT  721200.0 1869600.0 731400.0 1883400.0 ;
      RECT  721200.0 1897200.0 731400.0 1883400.0 ;
      RECT  721200.0 1897200.0 731400.0 1911000.0 ;
      RECT  721200.0 1924800.0 731400.0 1911000.0 ;
      RECT  721200.0 1924800.0 731400.0 1938600.0 ;
      RECT  721200.0 1952400.0 731400.0 1938600.0 ;
      RECT  721200.0 1952400.0 731400.0 1966200.0 ;
      RECT  721200.0 1980000.0 731400.0 1966200.0 ;
      RECT  721200.0 1980000.0 731400.0 1993800.0 ;
      RECT  721200.0 2007600.0 731400.0 1993800.0 ;
      RECT  721200.0 2007600.0 731400.0 2021400.0 ;
      RECT  721200.0 2035200.0 731400.0 2021400.0 ;
      RECT  721200.0 2035200.0 731400.0 2049000.0 ;
      RECT  721200.0 2062800.0 731400.0 2049000.0 ;
      RECT  721200.0 2062800.0 731400.0 2076600.0 ;
      RECT  721200.0 2090400.0 731400.0 2076600.0 ;
      RECT  721200.0 2090400.0 731400.0 2104200.0 ;
      RECT  721200.0 2118000.0 731400.0 2104200.0 ;
      RECT  721200.0 2118000.0 731400.0 2131800.0 ;
      RECT  721200.0 2145600.0 731400.0 2131800.0 ;
      RECT  731400.0 379200.0 741600.0 393000.0 ;
      RECT  731400.0 406800.0 741600.0 393000.0 ;
      RECT  731400.0 406800.0 741600.0 420600.0 ;
      RECT  731400.0 434400.0 741600.0 420600.0 ;
      RECT  731400.0 434400.0 741600.0 448200.0 ;
      RECT  731400.0 462000.0 741600.0 448200.0 ;
      RECT  731400.0 462000.0 741600.0 475800.0 ;
      RECT  731400.0 489600.0 741600.0 475800.0 ;
      RECT  731400.0 489600.0 741600.0 503400.0 ;
      RECT  731400.0 517200.0 741600.0 503400.0 ;
      RECT  731400.0 517200.0 741600.0 531000.0 ;
      RECT  731400.0 544800.0 741600.0 531000.0 ;
      RECT  731400.0 544800.0 741600.0 558600.0 ;
      RECT  731400.0 572400.0 741600.0 558600.0 ;
      RECT  731400.0 572400.0 741600.0 586200.0 ;
      RECT  731400.0 600000.0 741600.0 586200.0 ;
      RECT  731400.0 600000.0 741600.0 613800.0 ;
      RECT  731400.0 627600.0 741600.0 613800.0 ;
      RECT  731400.0 627600.0 741600.0 641400.0 ;
      RECT  731400.0 655200.0 741600.0 641400.0 ;
      RECT  731400.0 655200.0 741600.0 669000.0 ;
      RECT  731400.0 682800.0 741600.0 669000.0 ;
      RECT  731400.0 682800.0 741600.0 696600.0 ;
      RECT  731400.0 710400.0 741600.0 696600.0 ;
      RECT  731400.0 710400.0 741600.0 724200.0 ;
      RECT  731400.0 738000.0 741600.0 724200.0 ;
      RECT  731400.0 738000.0 741600.0 751800.0 ;
      RECT  731400.0 765600.0 741600.0 751800.0 ;
      RECT  731400.0 765600.0 741600.0 779400.0 ;
      RECT  731400.0 793200.0 741600.0 779400.0 ;
      RECT  731400.0 793200.0 741600.0 807000.0 ;
      RECT  731400.0 820800.0 741600.0 807000.0 ;
      RECT  731400.0 820800.0 741600.0 834600.0 ;
      RECT  731400.0 848400.0 741600.0 834600.0 ;
      RECT  731400.0 848400.0 741600.0 862200.0 ;
      RECT  731400.0 876000.0 741600.0 862200.0 ;
      RECT  731400.0 876000.0 741600.0 889800.0 ;
      RECT  731400.0 903600.0 741600.0 889800.0 ;
      RECT  731400.0 903600.0 741600.0 917400.0 ;
      RECT  731400.0 931200.0 741600.0 917400.0 ;
      RECT  731400.0 931200.0 741600.0 945000.0 ;
      RECT  731400.0 958800.0 741600.0 945000.0 ;
      RECT  731400.0 958800.0 741600.0 972600.0 ;
      RECT  731400.0 986400.0 741600.0 972600.0 ;
      RECT  731400.0 986400.0 741600.0 1000200.0 ;
      RECT  731400.0 1014000.0 741600.0 1000200.0 ;
      RECT  731400.0 1014000.0 741600.0 1027800.0 ;
      RECT  731400.0 1041600.0 741600.0 1027800.0 ;
      RECT  731400.0 1041600.0 741600.0 1055400.0 ;
      RECT  731400.0 1069200.0 741600.0 1055400.0 ;
      RECT  731400.0 1069200.0 741600.0 1083000.0 ;
      RECT  731400.0 1096800.0 741600.0 1083000.0 ;
      RECT  731400.0 1096800.0 741600.0 1110600.0 ;
      RECT  731400.0 1124400.0 741600.0 1110600.0 ;
      RECT  731400.0 1124400.0 741600.0 1138200.0 ;
      RECT  731400.0 1152000.0 741600.0 1138200.0 ;
      RECT  731400.0 1152000.0 741600.0 1165800.0 ;
      RECT  731400.0 1179600.0 741600.0 1165800.0 ;
      RECT  731400.0 1179600.0 741600.0 1193400.0 ;
      RECT  731400.0 1207200.0 741600.0 1193400.0 ;
      RECT  731400.0 1207200.0 741600.0 1221000.0 ;
      RECT  731400.0 1234800.0 741600.0 1221000.0 ;
      RECT  731400.0 1234800.0 741600.0 1248600.0 ;
      RECT  731400.0 1262400.0 741600.0 1248600.0 ;
      RECT  731400.0 1262400.0 741600.0 1276200.0 ;
      RECT  731400.0 1290000.0 741600.0 1276200.0 ;
      RECT  731400.0 1290000.0 741600.0 1303800.0 ;
      RECT  731400.0 1317600.0 741600.0 1303800.0 ;
      RECT  731400.0 1317600.0 741600.0 1331400.0 ;
      RECT  731400.0 1345200.0 741600.0 1331400.0 ;
      RECT  731400.0 1345200.0 741600.0 1359000.0 ;
      RECT  731400.0 1372800.0 741600.0 1359000.0 ;
      RECT  731400.0 1372800.0 741600.0 1386600.0 ;
      RECT  731400.0 1400400.0 741600.0 1386600.0 ;
      RECT  731400.0 1400400.0 741600.0 1414200.0 ;
      RECT  731400.0 1428000.0 741600.0 1414200.0 ;
      RECT  731400.0 1428000.0 741600.0 1441800.0 ;
      RECT  731400.0 1455600.0 741600.0 1441800.0 ;
      RECT  731400.0 1455600.0 741600.0 1469400.0 ;
      RECT  731400.0 1483200.0 741600.0 1469400.0 ;
      RECT  731400.0 1483200.0 741600.0 1497000.0 ;
      RECT  731400.0 1510800.0 741600.0 1497000.0 ;
      RECT  731400.0 1510800.0 741600.0 1524600.0 ;
      RECT  731400.0 1538400.0 741600.0 1524600.0 ;
      RECT  731400.0 1538400.0 741600.0 1552200.0 ;
      RECT  731400.0 1566000.0 741600.0 1552200.0 ;
      RECT  731400.0 1566000.0 741600.0 1579800.0 ;
      RECT  731400.0 1593600.0 741600.0 1579800.0 ;
      RECT  731400.0 1593600.0 741600.0 1607400.0 ;
      RECT  731400.0 1621200.0 741600.0 1607400.0 ;
      RECT  731400.0 1621200.0 741600.0 1635000.0 ;
      RECT  731400.0 1648800.0 741600.0 1635000.0 ;
      RECT  731400.0 1648800.0 741600.0 1662600.0 ;
      RECT  731400.0 1676400.0 741600.0 1662600.0 ;
      RECT  731400.0 1676400.0 741600.0 1690200.0 ;
      RECT  731400.0 1704000.0 741600.0 1690200.0 ;
      RECT  731400.0 1704000.0 741600.0 1717800.0 ;
      RECT  731400.0 1731600.0 741600.0 1717800.0 ;
      RECT  731400.0 1731600.0 741600.0 1745400.0 ;
      RECT  731400.0 1759200.0 741600.0 1745400.0 ;
      RECT  731400.0 1759200.0 741600.0 1773000.0 ;
      RECT  731400.0 1786800.0 741600.0 1773000.0 ;
      RECT  731400.0 1786800.0 741600.0 1800600.0 ;
      RECT  731400.0 1814400.0 741600.0 1800600.0 ;
      RECT  731400.0 1814400.0 741600.0 1828200.0 ;
      RECT  731400.0 1842000.0 741600.0 1828200.0 ;
      RECT  731400.0 1842000.0 741600.0 1855800.0 ;
      RECT  731400.0 1869600.0 741600.0 1855800.0 ;
      RECT  731400.0 1869600.0 741600.0 1883400.0 ;
      RECT  731400.0 1897200.0 741600.0 1883400.0 ;
      RECT  731400.0 1897200.0 741600.0 1911000.0 ;
      RECT  731400.0 1924800.0 741600.0 1911000.0 ;
      RECT  731400.0 1924800.0 741600.0 1938600.0 ;
      RECT  731400.0 1952400.0 741600.0 1938600.0 ;
      RECT  731400.0 1952400.0 741600.0 1966200.0 ;
      RECT  731400.0 1980000.0 741600.0 1966200.0 ;
      RECT  731400.0 1980000.0 741600.0 1993800.0 ;
      RECT  731400.0 2007600.0 741600.0 1993800.0 ;
      RECT  731400.0 2007600.0 741600.0 2021400.0 ;
      RECT  731400.0 2035200.0 741600.0 2021400.0 ;
      RECT  731400.0 2035200.0 741600.0 2049000.0 ;
      RECT  731400.0 2062800.0 741600.0 2049000.0 ;
      RECT  731400.0 2062800.0 741600.0 2076600.0 ;
      RECT  731400.0 2090400.0 741600.0 2076600.0 ;
      RECT  731400.0 2090400.0 741600.0 2104200.0 ;
      RECT  731400.0 2118000.0 741600.0 2104200.0 ;
      RECT  731400.0 2118000.0 741600.0 2131800.0 ;
      RECT  731400.0 2145600.0 741600.0 2131800.0 ;
      RECT  741600.0 379200.0 751800.0 393000.0 ;
      RECT  741600.0 406800.0 751800.0 393000.0 ;
      RECT  741600.0 406800.0 751800.0 420600.0 ;
      RECT  741600.0 434400.0 751800.0 420600.0 ;
      RECT  741600.0 434400.0 751800.0 448200.0 ;
      RECT  741600.0 462000.0 751800.0 448200.0 ;
      RECT  741600.0 462000.0 751800.0 475800.0 ;
      RECT  741600.0 489600.0 751800.0 475800.0 ;
      RECT  741600.0 489600.0 751800.0 503400.0 ;
      RECT  741600.0 517200.0 751800.0 503400.0 ;
      RECT  741600.0 517200.0 751800.0 531000.0 ;
      RECT  741600.0 544800.0 751800.0 531000.0 ;
      RECT  741600.0 544800.0 751800.0 558600.0 ;
      RECT  741600.0 572400.0 751800.0 558600.0 ;
      RECT  741600.0 572400.0 751800.0 586200.0 ;
      RECT  741600.0 600000.0 751800.0 586200.0 ;
      RECT  741600.0 600000.0 751800.0 613800.0 ;
      RECT  741600.0 627600.0 751800.0 613800.0 ;
      RECT  741600.0 627600.0 751800.0 641400.0 ;
      RECT  741600.0 655200.0 751800.0 641400.0 ;
      RECT  741600.0 655200.0 751800.0 669000.0 ;
      RECT  741600.0 682800.0 751800.0 669000.0 ;
      RECT  741600.0 682800.0 751800.0 696600.0 ;
      RECT  741600.0 710400.0 751800.0 696600.0 ;
      RECT  741600.0 710400.0 751800.0 724200.0 ;
      RECT  741600.0 738000.0 751800.0 724200.0 ;
      RECT  741600.0 738000.0 751800.0 751800.0 ;
      RECT  741600.0 765600.0 751800.0 751800.0 ;
      RECT  741600.0 765600.0 751800.0 779400.0 ;
      RECT  741600.0 793200.0 751800.0 779400.0 ;
      RECT  741600.0 793200.0 751800.0 807000.0 ;
      RECT  741600.0 820800.0 751800.0 807000.0 ;
      RECT  741600.0 820800.0 751800.0 834600.0 ;
      RECT  741600.0 848400.0 751800.0 834600.0 ;
      RECT  741600.0 848400.0 751800.0 862200.0 ;
      RECT  741600.0 876000.0 751800.0 862200.0 ;
      RECT  741600.0 876000.0 751800.0 889800.0 ;
      RECT  741600.0 903600.0 751800.0 889800.0 ;
      RECT  741600.0 903600.0 751800.0 917400.0 ;
      RECT  741600.0 931200.0 751800.0 917400.0 ;
      RECT  741600.0 931200.0 751800.0 945000.0 ;
      RECT  741600.0 958800.0 751800.0 945000.0 ;
      RECT  741600.0 958800.0 751800.0 972600.0 ;
      RECT  741600.0 986400.0 751800.0 972600.0 ;
      RECT  741600.0 986400.0 751800.0 1000200.0 ;
      RECT  741600.0 1014000.0 751800.0 1000200.0 ;
      RECT  741600.0 1014000.0 751800.0 1027800.0 ;
      RECT  741600.0 1041600.0 751800.0 1027800.0 ;
      RECT  741600.0 1041600.0 751800.0 1055400.0 ;
      RECT  741600.0 1069200.0 751800.0 1055400.0 ;
      RECT  741600.0 1069200.0 751800.0 1083000.0 ;
      RECT  741600.0 1096800.0 751800.0 1083000.0 ;
      RECT  741600.0 1096800.0 751800.0 1110600.0 ;
      RECT  741600.0 1124400.0 751800.0 1110600.0 ;
      RECT  741600.0 1124400.0 751800.0 1138200.0 ;
      RECT  741600.0 1152000.0 751800.0 1138200.0 ;
      RECT  741600.0 1152000.0 751800.0 1165800.0 ;
      RECT  741600.0 1179600.0 751800.0 1165800.0 ;
      RECT  741600.0 1179600.0 751800.0 1193400.0 ;
      RECT  741600.0 1207200.0 751800.0 1193400.0 ;
      RECT  741600.0 1207200.0 751800.0 1221000.0 ;
      RECT  741600.0 1234800.0 751800.0 1221000.0 ;
      RECT  741600.0 1234800.0 751800.0 1248600.0 ;
      RECT  741600.0 1262400.0 751800.0 1248600.0 ;
      RECT  741600.0 1262400.0 751800.0 1276200.0 ;
      RECT  741600.0 1290000.0 751800.0 1276200.0 ;
      RECT  741600.0 1290000.0 751800.0 1303800.0 ;
      RECT  741600.0 1317600.0 751800.0 1303800.0 ;
      RECT  741600.0 1317600.0 751800.0 1331400.0 ;
      RECT  741600.0 1345200.0 751800.0 1331400.0 ;
      RECT  741600.0 1345200.0 751800.0 1359000.0 ;
      RECT  741600.0 1372800.0 751800.0 1359000.0 ;
      RECT  741600.0 1372800.0 751800.0 1386600.0 ;
      RECT  741600.0 1400400.0 751800.0 1386600.0 ;
      RECT  741600.0 1400400.0 751800.0 1414200.0 ;
      RECT  741600.0 1428000.0 751800.0 1414200.0 ;
      RECT  741600.0 1428000.0 751800.0 1441800.0 ;
      RECT  741600.0 1455600.0 751800.0 1441800.0 ;
      RECT  741600.0 1455600.0 751800.0 1469400.0 ;
      RECT  741600.0 1483200.0 751800.0 1469400.0 ;
      RECT  741600.0 1483200.0 751800.0 1497000.0 ;
      RECT  741600.0 1510800.0 751800.0 1497000.0 ;
      RECT  741600.0 1510800.0 751800.0 1524600.0 ;
      RECT  741600.0 1538400.0 751800.0 1524600.0 ;
      RECT  741600.0 1538400.0 751800.0 1552200.0 ;
      RECT  741600.0 1566000.0 751800.0 1552200.0 ;
      RECT  741600.0 1566000.0 751800.0 1579800.0 ;
      RECT  741600.0 1593600.0 751800.0 1579800.0 ;
      RECT  741600.0 1593600.0 751800.0 1607400.0 ;
      RECT  741600.0 1621200.0 751800.0 1607400.0 ;
      RECT  741600.0 1621200.0 751800.0 1635000.0 ;
      RECT  741600.0 1648800.0 751800.0 1635000.0 ;
      RECT  741600.0 1648800.0 751800.0 1662600.0 ;
      RECT  741600.0 1676400.0 751800.0 1662600.0 ;
      RECT  741600.0 1676400.0 751800.0 1690200.0 ;
      RECT  741600.0 1704000.0 751800.0 1690200.0 ;
      RECT  741600.0 1704000.0 751800.0 1717800.0 ;
      RECT  741600.0 1731600.0 751800.0 1717800.0 ;
      RECT  741600.0 1731600.0 751800.0 1745400.0 ;
      RECT  741600.0 1759200.0 751800.0 1745400.0 ;
      RECT  741600.0 1759200.0 751800.0 1773000.0 ;
      RECT  741600.0 1786800.0 751800.0 1773000.0 ;
      RECT  741600.0 1786800.0 751800.0 1800600.0 ;
      RECT  741600.0 1814400.0 751800.0 1800600.0 ;
      RECT  741600.0 1814400.0 751800.0 1828200.0 ;
      RECT  741600.0 1842000.0 751800.0 1828200.0 ;
      RECT  741600.0 1842000.0 751800.0 1855800.0 ;
      RECT  741600.0 1869600.0 751800.0 1855800.0 ;
      RECT  741600.0 1869600.0 751800.0 1883400.0 ;
      RECT  741600.0 1897200.0 751800.0 1883400.0 ;
      RECT  741600.0 1897200.0 751800.0 1911000.0 ;
      RECT  741600.0 1924800.0 751800.0 1911000.0 ;
      RECT  741600.0 1924800.0 751800.0 1938600.0 ;
      RECT  741600.0 1952400.0 751800.0 1938600.0 ;
      RECT  741600.0 1952400.0 751800.0 1966200.0 ;
      RECT  741600.0 1980000.0 751800.0 1966200.0 ;
      RECT  741600.0 1980000.0 751800.0 1993800.0 ;
      RECT  741600.0 2007600.0 751800.0 1993800.0 ;
      RECT  741600.0 2007600.0 751800.0 2021400.0 ;
      RECT  741600.0 2035200.0 751800.0 2021400.0 ;
      RECT  741600.0 2035200.0 751800.0 2049000.0 ;
      RECT  741600.0 2062800.0 751800.0 2049000.0 ;
      RECT  741600.0 2062800.0 751800.0 2076600.0 ;
      RECT  741600.0 2090400.0 751800.0 2076600.0 ;
      RECT  741600.0 2090400.0 751800.0 2104200.0 ;
      RECT  741600.0 2118000.0 751800.0 2104200.0 ;
      RECT  741600.0 2118000.0 751800.0 2131800.0 ;
      RECT  741600.0 2145600.0 751800.0 2131800.0 ;
      RECT  751800.0 379200.0 762000.0 393000.0 ;
      RECT  751800.0 406800.0 762000.0 393000.0 ;
      RECT  751800.0 406800.0 762000.0 420600.0 ;
      RECT  751800.0 434400.0 762000.0 420600.0 ;
      RECT  751800.0 434400.0 762000.0 448200.0 ;
      RECT  751800.0 462000.0 762000.0 448200.0 ;
      RECT  751800.0 462000.0 762000.0 475800.0 ;
      RECT  751800.0 489600.0 762000.0 475800.0 ;
      RECT  751800.0 489600.0 762000.0 503400.0 ;
      RECT  751800.0 517200.0 762000.0 503400.0 ;
      RECT  751800.0 517200.0 762000.0 531000.0 ;
      RECT  751800.0 544800.0 762000.0 531000.0 ;
      RECT  751800.0 544800.0 762000.0 558600.0 ;
      RECT  751800.0 572400.0 762000.0 558600.0 ;
      RECT  751800.0 572400.0 762000.0 586200.0 ;
      RECT  751800.0 600000.0 762000.0 586200.0 ;
      RECT  751800.0 600000.0 762000.0 613800.0 ;
      RECT  751800.0 627600.0 762000.0 613800.0 ;
      RECT  751800.0 627600.0 762000.0 641400.0 ;
      RECT  751800.0 655200.0 762000.0 641400.0 ;
      RECT  751800.0 655200.0 762000.0 669000.0 ;
      RECT  751800.0 682800.0 762000.0 669000.0 ;
      RECT  751800.0 682800.0 762000.0 696600.0 ;
      RECT  751800.0 710400.0 762000.0 696600.0 ;
      RECT  751800.0 710400.0 762000.0 724200.0 ;
      RECT  751800.0 738000.0 762000.0 724200.0 ;
      RECT  751800.0 738000.0 762000.0 751800.0 ;
      RECT  751800.0 765600.0 762000.0 751800.0 ;
      RECT  751800.0 765600.0 762000.0 779400.0 ;
      RECT  751800.0 793200.0 762000.0 779400.0 ;
      RECT  751800.0 793200.0 762000.0 807000.0 ;
      RECT  751800.0 820800.0 762000.0 807000.0 ;
      RECT  751800.0 820800.0 762000.0 834600.0 ;
      RECT  751800.0 848400.0 762000.0 834600.0 ;
      RECT  751800.0 848400.0 762000.0 862200.0 ;
      RECT  751800.0 876000.0 762000.0 862200.0 ;
      RECT  751800.0 876000.0 762000.0 889800.0 ;
      RECT  751800.0 903600.0 762000.0 889800.0 ;
      RECT  751800.0 903600.0 762000.0 917400.0 ;
      RECT  751800.0 931200.0 762000.0 917400.0 ;
      RECT  751800.0 931200.0 762000.0 945000.0 ;
      RECT  751800.0 958800.0 762000.0 945000.0 ;
      RECT  751800.0 958800.0 762000.0 972600.0 ;
      RECT  751800.0 986400.0 762000.0 972600.0 ;
      RECT  751800.0 986400.0 762000.0 1000200.0 ;
      RECT  751800.0 1014000.0 762000.0 1000200.0 ;
      RECT  751800.0 1014000.0 762000.0 1027800.0 ;
      RECT  751800.0 1041600.0 762000.0 1027800.0 ;
      RECT  751800.0 1041600.0 762000.0 1055400.0 ;
      RECT  751800.0 1069200.0 762000.0 1055400.0 ;
      RECT  751800.0 1069200.0 762000.0 1083000.0 ;
      RECT  751800.0 1096800.0 762000.0 1083000.0 ;
      RECT  751800.0 1096800.0 762000.0 1110600.0 ;
      RECT  751800.0 1124400.0 762000.0 1110600.0 ;
      RECT  751800.0 1124400.0 762000.0 1138200.0 ;
      RECT  751800.0 1152000.0 762000.0 1138200.0 ;
      RECT  751800.0 1152000.0 762000.0 1165800.0 ;
      RECT  751800.0 1179600.0 762000.0 1165800.0 ;
      RECT  751800.0 1179600.0 762000.0 1193400.0 ;
      RECT  751800.0 1207200.0 762000.0 1193400.0 ;
      RECT  751800.0 1207200.0 762000.0 1221000.0 ;
      RECT  751800.0 1234800.0 762000.0 1221000.0 ;
      RECT  751800.0 1234800.0 762000.0 1248600.0 ;
      RECT  751800.0 1262400.0 762000.0 1248600.0 ;
      RECT  751800.0 1262400.0 762000.0 1276200.0 ;
      RECT  751800.0 1290000.0 762000.0 1276200.0 ;
      RECT  751800.0 1290000.0 762000.0 1303800.0 ;
      RECT  751800.0 1317600.0 762000.0 1303800.0 ;
      RECT  751800.0 1317600.0 762000.0 1331400.0 ;
      RECT  751800.0 1345200.0 762000.0 1331400.0 ;
      RECT  751800.0 1345200.0 762000.0 1359000.0 ;
      RECT  751800.0 1372800.0 762000.0 1359000.0 ;
      RECT  751800.0 1372800.0 762000.0 1386600.0 ;
      RECT  751800.0 1400400.0 762000.0 1386600.0 ;
      RECT  751800.0 1400400.0 762000.0 1414200.0 ;
      RECT  751800.0 1428000.0 762000.0 1414200.0 ;
      RECT  751800.0 1428000.0 762000.0 1441800.0 ;
      RECT  751800.0 1455600.0 762000.0 1441800.0 ;
      RECT  751800.0 1455600.0 762000.0 1469400.0 ;
      RECT  751800.0 1483200.0 762000.0 1469400.0 ;
      RECT  751800.0 1483200.0 762000.0 1497000.0 ;
      RECT  751800.0 1510800.0 762000.0 1497000.0 ;
      RECT  751800.0 1510800.0 762000.0 1524600.0 ;
      RECT  751800.0 1538400.0 762000.0 1524600.0 ;
      RECT  751800.0 1538400.0 762000.0 1552200.0 ;
      RECT  751800.0 1566000.0 762000.0 1552200.0 ;
      RECT  751800.0 1566000.0 762000.0 1579800.0 ;
      RECT  751800.0 1593600.0 762000.0 1579800.0 ;
      RECT  751800.0 1593600.0 762000.0 1607400.0 ;
      RECT  751800.0 1621200.0 762000.0 1607400.0 ;
      RECT  751800.0 1621200.0 762000.0 1635000.0 ;
      RECT  751800.0 1648800.0 762000.0 1635000.0 ;
      RECT  751800.0 1648800.0 762000.0 1662600.0 ;
      RECT  751800.0 1676400.0 762000.0 1662600.0 ;
      RECT  751800.0 1676400.0 762000.0 1690200.0 ;
      RECT  751800.0 1704000.0 762000.0 1690200.0 ;
      RECT  751800.0 1704000.0 762000.0 1717800.0 ;
      RECT  751800.0 1731600.0 762000.0 1717800.0 ;
      RECT  751800.0 1731600.0 762000.0 1745400.0 ;
      RECT  751800.0 1759200.0 762000.0 1745400.0 ;
      RECT  751800.0 1759200.0 762000.0 1773000.0 ;
      RECT  751800.0 1786800.0 762000.0 1773000.0 ;
      RECT  751800.0 1786800.0 762000.0 1800600.0 ;
      RECT  751800.0 1814400.0 762000.0 1800600.0 ;
      RECT  751800.0 1814400.0 762000.0 1828200.0 ;
      RECT  751800.0 1842000.0 762000.0 1828200.0 ;
      RECT  751800.0 1842000.0 762000.0 1855800.0 ;
      RECT  751800.0 1869600.0 762000.0 1855800.0 ;
      RECT  751800.0 1869600.0 762000.0 1883400.0 ;
      RECT  751800.0 1897200.0 762000.0 1883400.0 ;
      RECT  751800.0 1897200.0 762000.0 1911000.0 ;
      RECT  751800.0 1924800.0 762000.0 1911000.0 ;
      RECT  751800.0 1924800.0 762000.0 1938600.0 ;
      RECT  751800.0 1952400.0 762000.0 1938600.0 ;
      RECT  751800.0 1952400.0 762000.0 1966200.0 ;
      RECT  751800.0 1980000.0 762000.0 1966200.0 ;
      RECT  751800.0 1980000.0 762000.0 1993800.0 ;
      RECT  751800.0 2007600.0 762000.0 1993800.0 ;
      RECT  751800.0 2007600.0 762000.0 2021400.0 ;
      RECT  751800.0 2035200.0 762000.0 2021400.0 ;
      RECT  751800.0 2035200.0 762000.0 2049000.0 ;
      RECT  751800.0 2062800.0 762000.0 2049000.0 ;
      RECT  751800.0 2062800.0 762000.0 2076600.0 ;
      RECT  751800.0 2090400.0 762000.0 2076600.0 ;
      RECT  751800.0 2090400.0 762000.0 2104200.0 ;
      RECT  751800.0 2118000.0 762000.0 2104200.0 ;
      RECT  751800.0 2118000.0 762000.0 2131800.0 ;
      RECT  751800.0 2145600.0 762000.0 2131800.0 ;
      RECT  762000.0 379200.0 772200.0 393000.0 ;
      RECT  762000.0 406800.0 772200.0 393000.0 ;
      RECT  762000.0 406800.0 772200.0 420600.0 ;
      RECT  762000.0 434400.0 772200.0 420600.0 ;
      RECT  762000.0 434400.0 772200.0 448200.0 ;
      RECT  762000.0 462000.0 772200.0 448200.0 ;
      RECT  762000.0 462000.0 772200.0 475800.0 ;
      RECT  762000.0 489600.0 772200.0 475800.0 ;
      RECT  762000.0 489600.0 772200.0 503400.0 ;
      RECT  762000.0 517200.0 772200.0 503400.0 ;
      RECT  762000.0 517200.0 772200.0 531000.0 ;
      RECT  762000.0 544800.0 772200.0 531000.0 ;
      RECT  762000.0 544800.0 772200.0 558600.0 ;
      RECT  762000.0 572400.0 772200.0 558600.0 ;
      RECT  762000.0 572400.0 772200.0 586200.0 ;
      RECT  762000.0 600000.0 772200.0 586200.0 ;
      RECT  762000.0 600000.0 772200.0 613800.0 ;
      RECT  762000.0 627600.0 772200.0 613800.0 ;
      RECT  762000.0 627600.0 772200.0 641400.0 ;
      RECT  762000.0 655200.0 772200.0 641400.0 ;
      RECT  762000.0 655200.0 772200.0 669000.0 ;
      RECT  762000.0 682800.0 772200.0 669000.0 ;
      RECT  762000.0 682800.0 772200.0 696600.0 ;
      RECT  762000.0 710400.0 772200.0 696600.0 ;
      RECT  762000.0 710400.0 772200.0 724200.0 ;
      RECT  762000.0 738000.0 772200.0 724200.0 ;
      RECT  762000.0 738000.0 772200.0 751800.0 ;
      RECT  762000.0 765600.0 772200.0 751800.0 ;
      RECT  762000.0 765600.0 772200.0 779400.0 ;
      RECT  762000.0 793200.0 772200.0 779400.0 ;
      RECT  762000.0 793200.0 772200.0 807000.0 ;
      RECT  762000.0 820800.0 772200.0 807000.0 ;
      RECT  762000.0 820800.0 772200.0 834600.0 ;
      RECT  762000.0 848400.0 772200.0 834600.0 ;
      RECT  762000.0 848400.0 772200.0 862200.0 ;
      RECT  762000.0 876000.0 772200.0 862200.0 ;
      RECT  762000.0 876000.0 772200.0 889800.0 ;
      RECT  762000.0 903600.0 772200.0 889800.0 ;
      RECT  762000.0 903600.0 772200.0 917400.0 ;
      RECT  762000.0 931200.0 772200.0 917400.0 ;
      RECT  762000.0 931200.0 772200.0 945000.0 ;
      RECT  762000.0 958800.0 772200.0 945000.0 ;
      RECT  762000.0 958800.0 772200.0 972600.0 ;
      RECT  762000.0 986400.0 772200.0 972600.0 ;
      RECT  762000.0 986400.0 772200.0 1000200.0 ;
      RECT  762000.0 1014000.0 772200.0 1000200.0 ;
      RECT  762000.0 1014000.0 772200.0 1027800.0 ;
      RECT  762000.0 1041600.0 772200.0 1027800.0 ;
      RECT  762000.0 1041600.0 772200.0 1055400.0 ;
      RECT  762000.0 1069200.0 772200.0 1055400.0 ;
      RECT  762000.0 1069200.0 772200.0 1083000.0 ;
      RECT  762000.0 1096800.0 772200.0 1083000.0 ;
      RECT  762000.0 1096800.0 772200.0 1110600.0 ;
      RECT  762000.0 1124400.0 772200.0 1110600.0 ;
      RECT  762000.0 1124400.0 772200.0 1138200.0 ;
      RECT  762000.0 1152000.0 772200.0 1138200.0 ;
      RECT  762000.0 1152000.0 772200.0 1165800.0 ;
      RECT  762000.0 1179600.0 772200.0 1165800.0 ;
      RECT  762000.0 1179600.0 772200.0 1193400.0 ;
      RECT  762000.0 1207200.0 772200.0 1193400.0 ;
      RECT  762000.0 1207200.0 772200.0 1221000.0 ;
      RECT  762000.0 1234800.0 772200.0 1221000.0 ;
      RECT  762000.0 1234800.0 772200.0 1248600.0 ;
      RECT  762000.0 1262400.0 772200.0 1248600.0 ;
      RECT  762000.0 1262400.0 772200.0 1276200.0 ;
      RECT  762000.0 1290000.0 772200.0 1276200.0 ;
      RECT  762000.0 1290000.0 772200.0 1303800.0 ;
      RECT  762000.0 1317600.0 772200.0 1303800.0 ;
      RECT  762000.0 1317600.0 772200.0 1331400.0 ;
      RECT  762000.0 1345200.0 772200.0 1331400.0 ;
      RECT  762000.0 1345200.0 772200.0 1359000.0 ;
      RECT  762000.0 1372800.0 772200.0 1359000.0 ;
      RECT  762000.0 1372800.0 772200.0 1386600.0 ;
      RECT  762000.0 1400400.0 772200.0 1386600.0 ;
      RECT  762000.0 1400400.0 772200.0 1414200.0 ;
      RECT  762000.0 1428000.0 772200.0 1414200.0 ;
      RECT  762000.0 1428000.0 772200.0 1441800.0 ;
      RECT  762000.0 1455600.0 772200.0 1441800.0 ;
      RECT  762000.0 1455600.0 772200.0 1469400.0 ;
      RECT  762000.0 1483200.0 772200.0 1469400.0 ;
      RECT  762000.0 1483200.0 772200.0 1497000.0 ;
      RECT  762000.0 1510800.0 772200.0 1497000.0 ;
      RECT  762000.0 1510800.0 772200.0 1524600.0 ;
      RECT  762000.0 1538400.0 772200.0 1524600.0 ;
      RECT  762000.0 1538400.0 772200.0 1552200.0 ;
      RECT  762000.0 1566000.0 772200.0 1552200.0 ;
      RECT  762000.0 1566000.0 772200.0 1579800.0 ;
      RECT  762000.0 1593600.0 772200.0 1579800.0 ;
      RECT  762000.0 1593600.0 772200.0 1607400.0 ;
      RECT  762000.0 1621200.0 772200.0 1607400.0 ;
      RECT  762000.0 1621200.0 772200.0 1635000.0 ;
      RECT  762000.0 1648800.0 772200.0 1635000.0 ;
      RECT  762000.0 1648800.0 772200.0 1662600.0 ;
      RECT  762000.0 1676400.0 772200.0 1662600.0 ;
      RECT  762000.0 1676400.0 772200.0 1690200.0 ;
      RECT  762000.0 1704000.0 772200.0 1690200.0 ;
      RECT  762000.0 1704000.0 772200.0 1717800.0 ;
      RECT  762000.0 1731600.0 772200.0 1717800.0 ;
      RECT  762000.0 1731600.0 772200.0 1745400.0 ;
      RECT  762000.0 1759200.0 772200.0 1745400.0 ;
      RECT  762000.0 1759200.0 772200.0 1773000.0 ;
      RECT  762000.0 1786800.0 772200.0 1773000.0 ;
      RECT  762000.0 1786800.0 772200.0 1800600.0 ;
      RECT  762000.0 1814400.0 772200.0 1800600.0 ;
      RECT  762000.0 1814400.0 772200.0 1828200.0 ;
      RECT  762000.0 1842000.0 772200.0 1828200.0 ;
      RECT  762000.0 1842000.0 772200.0 1855800.0 ;
      RECT  762000.0 1869600.0 772200.0 1855800.0 ;
      RECT  762000.0 1869600.0 772200.0 1883400.0 ;
      RECT  762000.0 1897200.0 772200.0 1883400.0 ;
      RECT  762000.0 1897200.0 772200.0 1911000.0 ;
      RECT  762000.0 1924800.0 772200.0 1911000.0 ;
      RECT  762000.0 1924800.0 772200.0 1938600.0 ;
      RECT  762000.0 1952400.0 772200.0 1938600.0 ;
      RECT  762000.0 1952400.0 772200.0 1966200.0 ;
      RECT  762000.0 1980000.0 772200.0 1966200.0 ;
      RECT  762000.0 1980000.0 772200.0 1993800.0 ;
      RECT  762000.0 2007600.0 772200.0 1993800.0 ;
      RECT  762000.0 2007600.0 772200.0 2021400.0 ;
      RECT  762000.0 2035200.0 772200.0 2021400.0 ;
      RECT  762000.0 2035200.0 772200.0 2049000.0 ;
      RECT  762000.0 2062800.0 772200.0 2049000.0 ;
      RECT  762000.0 2062800.0 772200.0 2076600.0 ;
      RECT  762000.0 2090400.0 772200.0 2076600.0 ;
      RECT  762000.0 2090400.0 772200.0 2104200.0 ;
      RECT  762000.0 2118000.0 772200.0 2104200.0 ;
      RECT  762000.0 2118000.0 772200.0 2131800.0 ;
      RECT  762000.0 2145600.0 772200.0 2131800.0 ;
      RECT  772200.0 379200.0 782400.0 393000.0 ;
      RECT  772200.0 406800.0 782400.0 393000.0 ;
      RECT  772200.0 406800.0 782400.0 420600.0 ;
      RECT  772200.0 434400.0 782400.0 420600.0 ;
      RECT  772200.0 434400.0 782400.0 448200.0 ;
      RECT  772200.0 462000.0 782400.0 448200.0 ;
      RECT  772200.0 462000.0 782400.0 475800.0 ;
      RECT  772200.0 489600.0 782400.0 475800.0 ;
      RECT  772200.0 489600.0 782400.0 503400.0 ;
      RECT  772200.0 517200.0 782400.0 503400.0 ;
      RECT  772200.0 517200.0 782400.0 531000.0 ;
      RECT  772200.0 544800.0 782400.0 531000.0 ;
      RECT  772200.0 544800.0 782400.0 558600.0 ;
      RECT  772200.0 572400.0 782400.0 558600.0 ;
      RECT  772200.0 572400.0 782400.0 586200.0 ;
      RECT  772200.0 600000.0 782400.0 586200.0 ;
      RECT  772200.0 600000.0 782400.0 613800.0 ;
      RECT  772200.0 627600.0 782400.0 613800.0 ;
      RECT  772200.0 627600.0 782400.0 641400.0 ;
      RECT  772200.0 655200.0 782400.0 641400.0 ;
      RECT  772200.0 655200.0 782400.0 669000.0 ;
      RECT  772200.0 682800.0 782400.0 669000.0 ;
      RECT  772200.0 682800.0 782400.0 696600.0 ;
      RECT  772200.0 710400.0 782400.0 696600.0 ;
      RECT  772200.0 710400.0 782400.0 724200.0 ;
      RECT  772200.0 738000.0 782400.0 724200.0 ;
      RECT  772200.0 738000.0 782400.0 751800.0 ;
      RECT  772200.0 765600.0 782400.0 751800.0 ;
      RECT  772200.0 765600.0 782400.0 779400.0 ;
      RECT  772200.0 793200.0 782400.0 779400.0 ;
      RECT  772200.0 793200.0 782400.0 807000.0 ;
      RECT  772200.0 820800.0 782400.0 807000.0 ;
      RECT  772200.0 820800.0 782400.0 834600.0 ;
      RECT  772200.0 848400.0 782400.0 834600.0 ;
      RECT  772200.0 848400.0 782400.0 862200.0 ;
      RECT  772200.0 876000.0 782400.0 862200.0 ;
      RECT  772200.0 876000.0 782400.0 889800.0 ;
      RECT  772200.0 903600.0 782400.0 889800.0 ;
      RECT  772200.0 903600.0 782400.0 917400.0 ;
      RECT  772200.0 931200.0 782400.0 917400.0 ;
      RECT  772200.0 931200.0 782400.0 945000.0 ;
      RECT  772200.0 958800.0 782400.0 945000.0 ;
      RECT  772200.0 958800.0 782400.0 972600.0 ;
      RECT  772200.0 986400.0 782400.0 972600.0 ;
      RECT  772200.0 986400.0 782400.0 1000200.0 ;
      RECT  772200.0 1014000.0 782400.0 1000200.0 ;
      RECT  772200.0 1014000.0 782400.0 1027800.0 ;
      RECT  772200.0 1041600.0 782400.0 1027800.0 ;
      RECT  772200.0 1041600.0 782400.0 1055400.0 ;
      RECT  772200.0 1069200.0 782400.0 1055400.0 ;
      RECT  772200.0 1069200.0 782400.0 1083000.0 ;
      RECT  772200.0 1096800.0 782400.0 1083000.0 ;
      RECT  772200.0 1096800.0 782400.0 1110600.0 ;
      RECT  772200.0 1124400.0 782400.0 1110600.0 ;
      RECT  772200.0 1124400.0 782400.0 1138200.0 ;
      RECT  772200.0 1152000.0 782400.0 1138200.0 ;
      RECT  772200.0 1152000.0 782400.0 1165800.0 ;
      RECT  772200.0 1179600.0 782400.0 1165800.0 ;
      RECT  772200.0 1179600.0 782400.0 1193400.0 ;
      RECT  772200.0 1207200.0 782400.0 1193400.0 ;
      RECT  772200.0 1207200.0 782400.0 1221000.0 ;
      RECT  772200.0 1234800.0 782400.0 1221000.0 ;
      RECT  772200.0 1234800.0 782400.0 1248600.0 ;
      RECT  772200.0 1262400.0 782400.0 1248600.0 ;
      RECT  772200.0 1262400.0 782400.0 1276200.0 ;
      RECT  772200.0 1290000.0 782400.0 1276200.0 ;
      RECT  772200.0 1290000.0 782400.0 1303800.0 ;
      RECT  772200.0 1317600.0 782400.0 1303800.0 ;
      RECT  772200.0 1317600.0 782400.0 1331400.0 ;
      RECT  772200.0 1345200.0 782400.0 1331400.0 ;
      RECT  772200.0 1345200.0 782400.0 1359000.0 ;
      RECT  772200.0 1372800.0 782400.0 1359000.0 ;
      RECT  772200.0 1372800.0 782400.0 1386600.0 ;
      RECT  772200.0 1400400.0 782400.0 1386600.0 ;
      RECT  772200.0 1400400.0 782400.0 1414200.0 ;
      RECT  772200.0 1428000.0 782400.0 1414200.0 ;
      RECT  772200.0 1428000.0 782400.0 1441800.0 ;
      RECT  772200.0 1455600.0 782400.0 1441800.0 ;
      RECT  772200.0 1455600.0 782400.0 1469400.0 ;
      RECT  772200.0 1483200.0 782400.0 1469400.0 ;
      RECT  772200.0 1483200.0 782400.0 1497000.0 ;
      RECT  772200.0 1510800.0 782400.0 1497000.0 ;
      RECT  772200.0 1510800.0 782400.0 1524600.0 ;
      RECT  772200.0 1538400.0 782400.0 1524600.0 ;
      RECT  772200.0 1538400.0 782400.0 1552200.0 ;
      RECT  772200.0 1566000.0 782400.0 1552200.0 ;
      RECT  772200.0 1566000.0 782400.0 1579800.0 ;
      RECT  772200.0 1593600.0 782400.0 1579800.0 ;
      RECT  772200.0 1593600.0 782400.0 1607400.0 ;
      RECT  772200.0 1621200.0 782400.0 1607400.0 ;
      RECT  772200.0 1621200.0 782400.0 1635000.0 ;
      RECT  772200.0 1648800.0 782400.0 1635000.0 ;
      RECT  772200.0 1648800.0 782400.0 1662600.0 ;
      RECT  772200.0 1676400.0 782400.0 1662600.0 ;
      RECT  772200.0 1676400.0 782400.0 1690200.0 ;
      RECT  772200.0 1704000.0 782400.0 1690200.0 ;
      RECT  772200.0 1704000.0 782400.0 1717800.0 ;
      RECT  772200.0 1731600.0 782400.0 1717800.0 ;
      RECT  772200.0 1731600.0 782400.0 1745400.0 ;
      RECT  772200.0 1759200.0 782400.0 1745400.0 ;
      RECT  772200.0 1759200.0 782400.0 1773000.0 ;
      RECT  772200.0 1786800.0 782400.0 1773000.0 ;
      RECT  772200.0 1786800.0 782400.0 1800600.0 ;
      RECT  772200.0 1814400.0 782400.0 1800600.0 ;
      RECT  772200.0 1814400.0 782400.0 1828200.0 ;
      RECT  772200.0 1842000.0 782400.0 1828200.0 ;
      RECT  772200.0 1842000.0 782400.0 1855800.0 ;
      RECT  772200.0 1869600.0 782400.0 1855800.0 ;
      RECT  772200.0 1869600.0 782400.0 1883400.0 ;
      RECT  772200.0 1897200.0 782400.0 1883400.0 ;
      RECT  772200.0 1897200.0 782400.0 1911000.0 ;
      RECT  772200.0 1924800.0 782400.0 1911000.0 ;
      RECT  772200.0 1924800.0 782400.0 1938600.0 ;
      RECT  772200.0 1952400.0 782400.0 1938600.0 ;
      RECT  772200.0 1952400.0 782400.0 1966200.0 ;
      RECT  772200.0 1980000.0 782400.0 1966200.0 ;
      RECT  772200.0 1980000.0 782400.0 1993800.0 ;
      RECT  772200.0 2007600.0 782400.0 1993800.0 ;
      RECT  772200.0 2007600.0 782400.0 2021400.0 ;
      RECT  772200.0 2035200.0 782400.0 2021400.0 ;
      RECT  772200.0 2035200.0 782400.0 2049000.0 ;
      RECT  772200.0 2062800.0 782400.0 2049000.0 ;
      RECT  772200.0 2062800.0 782400.0 2076600.0 ;
      RECT  772200.0 2090400.0 782400.0 2076600.0 ;
      RECT  772200.0 2090400.0 782400.0 2104200.0 ;
      RECT  772200.0 2118000.0 782400.0 2104200.0 ;
      RECT  772200.0 2118000.0 782400.0 2131800.0 ;
      RECT  772200.0 2145600.0 782400.0 2131800.0 ;
      RECT  782400.0 379200.0 792600.0 393000.0 ;
      RECT  782400.0 406800.0 792600.0 393000.0 ;
      RECT  782400.0 406800.0 792600.0 420600.0 ;
      RECT  782400.0 434400.0 792600.0 420600.0 ;
      RECT  782400.0 434400.0 792600.0 448200.0 ;
      RECT  782400.0 462000.0 792600.0 448200.0 ;
      RECT  782400.0 462000.0 792600.0 475800.0 ;
      RECT  782400.0 489600.0 792600.0 475800.0 ;
      RECT  782400.0 489600.0 792600.0 503400.0 ;
      RECT  782400.0 517200.0 792600.0 503400.0 ;
      RECT  782400.0 517200.0 792600.0 531000.0 ;
      RECT  782400.0 544800.0 792600.0 531000.0 ;
      RECT  782400.0 544800.0 792600.0 558600.0 ;
      RECT  782400.0 572400.0 792600.0 558600.0 ;
      RECT  782400.0 572400.0 792600.0 586200.0 ;
      RECT  782400.0 600000.0 792600.0 586200.0 ;
      RECT  782400.0 600000.0 792600.0 613800.0 ;
      RECT  782400.0 627600.0 792600.0 613800.0 ;
      RECT  782400.0 627600.0 792600.0 641400.0 ;
      RECT  782400.0 655200.0 792600.0 641400.0 ;
      RECT  782400.0 655200.0 792600.0 669000.0 ;
      RECT  782400.0 682800.0 792600.0 669000.0 ;
      RECT  782400.0 682800.0 792600.0 696600.0 ;
      RECT  782400.0 710400.0 792600.0 696600.0 ;
      RECT  782400.0 710400.0 792600.0 724200.0 ;
      RECT  782400.0 738000.0 792600.0 724200.0 ;
      RECT  782400.0 738000.0 792600.0 751800.0 ;
      RECT  782400.0 765600.0 792600.0 751800.0 ;
      RECT  782400.0 765600.0 792600.0 779400.0 ;
      RECT  782400.0 793200.0 792600.0 779400.0 ;
      RECT  782400.0 793200.0 792600.0 807000.0 ;
      RECT  782400.0 820800.0 792600.0 807000.0 ;
      RECT  782400.0 820800.0 792600.0 834600.0 ;
      RECT  782400.0 848400.0 792600.0 834600.0 ;
      RECT  782400.0 848400.0 792600.0 862200.0 ;
      RECT  782400.0 876000.0 792600.0 862200.0 ;
      RECT  782400.0 876000.0 792600.0 889800.0 ;
      RECT  782400.0 903600.0 792600.0 889800.0 ;
      RECT  782400.0 903600.0 792600.0 917400.0 ;
      RECT  782400.0 931200.0 792600.0 917400.0 ;
      RECT  782400.0 931200.0 792600.0 945000.0 ;
      RECT  782400.0 958800.0 792600.0 945000.0 ;
      RECT  782400.0 958800.0 792600.0 972600.0 ;
      RECT  782400.0 986400.0 792600.0 972600.0 ;
      RECT  782400.0 986400.0 792600.0 1000200.0 ;
      RECT  782400.0 1014000.0 792600.0 1000200.0 ;
      RECT  782400.0 1014000.0 792600.0 1027800.0 ;
      RECT  782400.0 1041600.0 792600.0 1027800.0 ;
      RECT  782400.0 1041600.0 792600.0 1055400.0 ;
      RECT  782400.0 1069200.0 792600.0 1055400.0 ;
      RECT  782400.0 1069200.0 792600.0 1083000.0 ;
      RECT  782400.0 1096800.0 792600.0 1083000.0 ;
      RECT  782400.0 1096800.0 792600.0 1110600.0 ;
      RECT  782400.0 1124400.0 792600.0 1110600.0 ;
      RECT  782400.0 1124400.0 792600.0 1138200.0 ;
      RECT  782400.0 1152000.0 792600.0 1138200.0 ;
      RECT  782400.0 1152000.0 792600.0 1165800.0 ;
      RECT  782400.0 1179600.0 792600.0 1165800.0 ;
      RECT  782400.0 1179600.0 792600.0 1193400.0 ;
      RECT  782400.0 1207200.0 792600.0 1193400.0 ;
      RECT  782400.0 1207200.0 792600.0 1221000.0 ;
      RECT  782400.0 1234800.0 792600.0 1221000.0 ;
      RECT  782400.0 1234800.0 792600.0 1248600.0 ;
      RECT  782400.0 1262400.0 792600.0 1248600.0 ;
      RECT  782400.0 1262400.0 792600.0 1276200.0 ;
      RECT  782400.0 1290000.0 792600.0 1276200.0 ;
      RECT  782400.0 1290000.0 792600.0 1303800.0 ;
      RECT  782400.0 1317600.0 792600.0 1303800.0 ;
      RECT  782400.0 1317600.0 792600.0 1331400.0 ;
      RECT  782400.0 1345200.0 792600.0 1331400.0 ;
      RECT  782400.0 1345200.0 792600.0 1359000.0 ;
      RECT  782400.0 1372800.0 792600.0 1359000.0 ;
      RECT  782400.0 1372800.0 792600.0 1386600.0 ;
      RECT  782400.0 1400400.0 792600.0 1386600.0 ;
      RECT  782400.0 1400400.0 792600.0 1414200.0 ;
      RECT  782400.0 1428000.0 792600.0 1414200.0 ;
      RECT  782400.0 1428000.0 792600.0 1441800.0 ;
      RECT  782400.0 1455600.0 792600.0 1441800.0 ;
      RECT  782400.0 1455600.0 792600.0 1469400.0 ;
      RECT  782400.0 1483200.0 792600.0 1469400.0 ;
      RECT  782400.0 1483200.0 792600.0 1497000.0 ;
      RECT  782400.0 1510800.0 792600.0 1497000.0 ;
      RECT  782400.0 1510800.0 792600.0 1524600.0 ;
      RECT  782400.0 1538400.0 792600.0 1524600.0 ;
      RECT  782400.0 1538400.0 792600.0 1552200.0 ;
      RECT  782400.0 1566000.0 792600.0 1552200.0 ;
      RECT  782400.0 1566000.0 792600.0 1579800.0 ;
      RECT  782400.0 1593600.0 792600.0 1579800.0 ;
      RECT  782400.0 1593600.0 792600.0 1607400.0 ;
      RECT  782400.0 1621200.0 792600.0 1607400.0 ;
      RECT  782400.0 1621200.0 792600.0 1635000.0 ;
      RECT  782400.0 1648800.0 792600.0 1635000.0 ;
      RECT  782400.0 1648800.0 792600.0 1662600.0 ;
      RECT  782400.0 1676400.0 792600.0 1662600.0 ;
      RECT  782400.0 1676400.0 792600.0 1690200.0 ;
      RECT  782400.0 1704000.0 792600.0 1690200.0 ;
      RECT  782400.0 1704000.0 792600.0 1717800.0 ;
      RECT  782400.0 1731600.0 792600.0 1717800.0 ;
      RECT  782400.0 1731600.0 792600.0 1745400.0 ;
      RECT  782400.0 1759200.0 792600.0 1745400.0 ;
      RECT  782400.0 1759200.0 792600.0 1773000.0 ;
      RECT  782400.0 1786800.0 792600.0 1773000.0 ;
      RECT  782400.0 1786800.0 792600.0 1800600.0 ;
      RECT  782400.0 1814400.0 792600.0 1800600.0 ;
      RECT  782400.0 1814400.0 792600.0 1828200.0 ;
      RECT  782400.0 1842000.0 792600.0 1828200.0 ;
      RECT  782400.0 1842000.0 792600.0 1855800.0 ;
      RECT  782400.0 1869600.0 792600.0 1855800.0 ;
      RECT  782400.0 1869600.0 792600.0 1883400.0 ;
      RECT  782400.0 1897200.0 792600.0 1883400.0 ;
      RECT  782400.0 1897200.0 792600.0 1911000.0 ;
      RECT  782400.0 1924800.0 792600.0 1911000.0 ;
      RECT  782400.0 1924800.0 792600.0 1938600.0 ;
      RECT  782400.0 1952400.0 792600.0 1938600.0 ;
      RECT  782400.0 1952400.0 792600.0 1966200.0 ;
      RECT  782400.0 1980000.0 792600.0 1966200.0 ;
      RECT  782400.0 1980000.0 792600.0 1993800.0 ;
      RECT  782400.0 2007600.0 792600.0 1993800.0 ;
      RECT  782400.0 2007600.0 792600.0 2021400.0 ;
      RECT  782400.0 2035200.0 792600.0 2021400.0 ;
      RECT  782400.0 2035200.0 792600.0 2049000.0 ;
      RECT  782400.0 2062800.0 792600.0 2049000.0 ;
      RECT  782400.0 2062800.0 792600.0 2076600.0 ;
      RECT  782400.0 2090400.0 792600.0 2076600.0 ;
      RECT  782400.0 2090400.0 792600.0 2104200.0 ;
      RECT  782400.0 2118000.0 792600.0 2104200.0 ;
      RECT  782400.0 2118000.0 792600.0 2131800.0 ;
      RECT  782400.0 2145600.0 792600.0 2131800.0 ;
      RECT  792600.0 379200.0 802800.0 393000.0 ;
      RECT  792600.0 406800.0 802800.0 393000.0 ;
      RECT  792600.0 406800.0 802800.0 420600.0 ;
      RECT  792600.0 434400.0 802800.0 420600.0 ;
      RECT  792600.0 434400.0 802800.0 448200.0 ;
      RECT  792600.0 462000.0 802800.0 448200.0 ;
      RECT  792600.0 462000.0 802800.0 475800.0 ;
      RECT  792600.0 489600.0 802800.0 475800.0 ;
      RECT  792600.0 489600.0 802800.0 503400.0 ;
      RECT  792600.0 517200.0 802800.0 503400.0 ;
      RECT  792600.0 517200.0 802800.0 531000.0 ;
      RECT  792600.0 544800.0 802800.0 531000.0 ;
      RECT  792600.0 544800.0 802800.0 558600.0 ;
      RECT  792600.0 572400.0 802800.0 558600.0 ;
      RECT  792600.0 572400.0 802800.0 586200.0 ;
      RECT  792600.0 600000.0 802800.0 586200.0 ;
      RECT  792600.0 600000.0 802800.0 613800.0 ;
      RECT  792600.0 627600.0 802800.0 613800.0 ;
      RECT  792600.0 627600.0 802800.0 641400.0 ;
      RECT  792600.0 655200.0 802800.0 641400.0 ;
      RECT  792600.0 655200.0 802800.0 669000.0 ;
      RECT  792600.0 682800.0 802800.0 669000.0 ;
      RECT  792600.0 682800.0 802800.0 696600.0 ;
      RECT  792600.0 710400.0 802800.0 696600.0 ;
      RECT  792600.0 710400.0 802800.0 724200.0 ;
      RECT  792600.0 738000.0 802800.0 724200.0 ;
      RECT  792600.0 738000.0 802800.0 751800.0 ;
      RECT  792600.0 765600.0 802800.0 751800.0 ;
      RECT  792600.0 765600.0 802800.0 779400.0 ;
      RECT  792600.0 793200.0 802800.0 779400.0 ;
      RECT  792600.0 793200.0 802800.0 807000.0 ;
      RECT  792600.0 820800.0 802800.0 807000.0 ;
      RECT  792600.0 820800.0 802800.0 834600.0 ;
      RECT  792600.0 848400.0 802800.0 834600.0 ;
      RECT  792600.0 848400.0 802800.0 862200.0 ;
      RECT  792600.0 876000.0 802800.0 862200.0 ;
      RECT  792600.0 876000.0 802800.0 889800.0 ;
      RECT  792600.0 903600.0 802800.0 889800.0 ;
      RECT  792600.0 903600.0 802800.0 917400.0 ;
      RECT  792600.0 931200.0 802800.0 917400.0 ;
      RECT  792600.0 931200.0 802800.0 945000.0 ;
      RECT  792600.0 958800.0 802800.0 945000.0 ;
      RECT  792600.0 958800.0 802800.0 972600.0 ;
      RECT  792600.0 986400.0 802800.0 972600.0 ;
      RECT  792600.0 986400.0 802800.0 1000200.0 ;
      RECT  792600.0 1014000.0 802800.0 1000200.0 ;
      RECT  792600.0 1014000.0 802800.0 1027800.0 ;
      RECT  792600.0 1041600.0 802800.0 1027800.0 ;
      RECT  792600.0 1041600.0 802800.0 1055400.0 ;
      RECT  792600.0 1069200.0 802800.0 1055400.0 ;
      RECT  792600.0 1069200.0 802800.0 1083000.0 ;
      RECT  792600.0 1096800.0 802800.0 1083000.0 ;
      RECT  792600.0 1096800.0 802800.0 1110600.0 ;
      RECT  792600.0 1124400.0 802800.0 1110600.0 ;
      RECT  792600.0 1124400.0 802800.0 1138200.0 ;
      RECT  792600.0 1152000.0 802800.0 1138200.0 ;
      RECT  792600.0 1152000.0 802800.0 1165800.0 ;
      RECT  792600.0 1179600.0 802800.0 1165800.0 ;
      RECT  792600.0 1179600.0 802800.0 1193400.0 ;
      RECT  792600.0 1207200.0 802800.0 1193400.0 ;
      RECT  792600.0 1207200.0 802800.0 1221000.0 ;
      RECT  792600.0 1234800.0 802800.0 1221000.0 ;
      RECT  792600.0 1234800.0 802800.0 1248600.0 ;
      RECT  792600.0 1262400.0 802800.0 1248600.0 ;
      RECT  792600.0 1262400.0 802800.0 1276200.0 ;
      RECT  792600.0 1290000.0 802800.0 1276200.0 ;
      RECT  792600.0 1290000.0 802800.0 1303800.0 ;
      RECT  792600.0 1317600.0 802800.0 1303800.0 ;
      RECT  792600.0 1317600.0 802800.0 1331400.0 ;
      RECT  792600.0 1345200.0 802800.0 1331400.0 ;
      RECT  792600.0 1345200.0 802800.0 1359000.0 ;
      RECT  792600.0 1372800.0 802800.0 1359000.0 ;
      RECT  792600.0 1372800.0 802800.0 1386600.0 ;
      RECT  792600.0 1400400.0 802800.0 1386600.0 ;
      RECT  792600.0 1400400.0 802800.0 1414200.0 ;
      RECT  792600.0 1428000.0 802800.0 1414200.0 ;
      RECT  792600.0 1428000.0 802800.0 1441800.0 ;
      RECT  792600.0 1455600.0 802800.0 1441800.0 ;
      RECT  792600.0 1455600.0 802800.0 1469400.0 ;
      RECT  792600.0 1483200.0 802800.0 1469400.0 ;
      RECT  792600.0 1483200.0 802800.0 1497000.0 ;
      RECT  792600.0 1510800.0 802800.0 1497000.0 ;
      RECT  792600.0 1510800.0 802800.0 1524600.0 ;
      RECT  792600.0 1538400.0 802800.0 1524600.0 ;
      RECT  792600.0 1538400.0 802800.0 1552200.0 ;
      RECT  792600.0 1566000.0 802800.0 1552200.0 ;
      RECT  792600.0 1566000.0 802800.0 1579800.0 ;
      RECT  792600.0 1593600.0 802800.0 1579800.0 ;
      RECT  792600.0 1593600.0 802800.0 1607400.0 ;
      RECT  792600.0 1621200.0 802800.0 1607400.0 ;
      RECT  792600.0 1621200.0 802800.0 1635000.0 ;
      RECT  792600.0 1648800.0 802800.0 1635000.0 ;
      RECT  792600.0 1648800.0 802800.0 1662600.0 ;
      RECT  792600.0 1676400.0 802800.0 1662600.0 ;
      RECT  792600.0 1676400.0 802800.0 1690200.0 ;
      RECT  792600.0 1704000.0 802800.0 1690200.0 ;
      RECT  792600.0 1704000.0 802800.0 1717800.0 ;
      RECT  792600.0 1731600.0 802800.0 1717800.0 ;
      RECT  792600.0 1731600.0 802800.0 1745400.0 ;
      RECT  792600.0 1759200.0 802800.0 1745400.0 ;
      RECT  792600.0 1759200.0 802800.0 1773000.0 ;
      RECT  792600.0 1786800.0 802800.0 1773000.0 ;
      RECT  792600.0 1786800.0 802800.0 1800600.0 ;
      RECT  792600.0 1814400.0 802800.0 1800600.0 ;
      RECT  792600.0 1814400.0 802800.0 1828200.0 ;
      RECT  792600.0 1842000.0 802800.0 1828200.0 ;
      RECT  792600.0 1842000.0 802800.0 1855800.0 ;
      RECT  792600.0 1869600.0 802800.0 1855800.0 ;
      RECT  792600.0 1869600.0 802800.0 1883400.0 ;
      RECT  792600.0 1897200.0 802800.0 1883400.0 ;
      RECT  792600.0 1897200.0 802800.0 1911000.0 ;
      RECT  792600.0 1924800.0 802800.0 1911000.0 ;
      RECT  792600.0 1924800.0 802800.0 1938600.0 ;
      RECT  792600.0 1952400.0 802800.0 1938600.0 ;
      RECT  792600.0 1952400.0 802800.0 1966200.0 ;
      RECT  792600.0 1980000.0 802800.0 1966200.0 ;
      RECT  792600.0 1980000.0 802800.0 1993800.0 ;
      RECT  792600.0 2007600.0 802800.0 1993800.0 ;
      RECT  792600.0 2007600.0 802800.0 2021400.0 ;
      RECT  792600.0 2035200.0 802800.0 2021400.0 ;
      RECT  792600.0 2035200.0 802800.0 2049000.0 ;
      RECT  792600.0 2062800.0 802800.0 2049000.0 ;
      RECT  792600.0 2062800.0 802800.0 2076600.0 ;
      RECT  792600.0 2090400.0 802800.0 2076600.0 ;
      RECT  792600.0 2090400.0 802800.0 2104200.0 ;
      RECT  792600.0 2118000.0 802800.0 2104200.0 ;
      RECT  792600.0 2118000.0 802800.0 2131800.0 ;
      RECT  792600.0 2145600.0 802800.0 2131800.0 ;
      RECT  802800.0 379200.0 813000.0 393000.0 ;
      RECT  802800.0 406800.0 813000.0 393000.0 ;
      RECT  802800.0 406800.0 813000.0 420600.0 ;
      RECT  802800.0 434400.0 813000.0 420600.0 ;
      RECT  802800.0 434400.0 813000.0 448200.0 ;
      RECT  802800.0 462000.0 813000.0 448200.0 ;
      RECT  802800.0 462000.0 813000.0 475800.0 ;
      RECT  802800.0 489600.0 813000.0 475800.0 ;
      RECT  802800.0 489600.0 813000.0 503400.0 ;
      RECT  802800.0 517200.0 813000.0 503400.0 ;
      RECT  802800.0 517200.0 813000.0 531000.0 ;
      RECT  802800.0 544800.0 813000.0 531000.0 ;
      RECT  802800.0 544800.0 813000.0 558600.0 ;
      RECT  802800.0 572400.0 813000.0 558600.0 ;
      RECT  802800.0 572400.0 813000.0 586200.0 ;
      RECT  802800.0 600000.0 813000.0 586200.0 ;
      RECT  802800.0 600000.0 813000.0 613800.0 ;
      RECT  802800.0 627600.0 813000.0 613800.0 ;
      RECT  802800.0 627600.0 813000.0 641400.0 ;
      RECT  802800.0 655200.0 813000.0 641400.0 ;
      RECT  802800.0 655200.0 813000.0 669000.0 ;
      RECT  802800.0 682800.0 813000.0 669000.0 ;
      RECT  802800.0 682800.0 813000.0 696600.0 ;
      RECT  802800.0 710400.0 813000.0 696600.0 ;
      RECT  802800.0 710400.0 813000.0 724200.0 ;
      RECT  802800.0 738000.0 813000.0 724200.0 ;
      RECT  802800.0 738000.0 813000.0 751800.0 ;
      RECT  802800.0 765600.0 813000.0 751800.0 ;
      RECT  802800.0 765600.0 813000.0 779400.0 ;
      RECT  802800.0 793200.0 813000.0 779400.0 ;
      RECT  802800.0 793200.0 813000.0 807000.0 ;
      RECT  802800.0 820800.0 813000.0 807000.0 ;
      RECT  802800.0 820800.0 813000.0 834600.0 ;
      RECT  802800.0 848400.0 813000.0 834600.0 ;
      RECT  802800.0 848400.0 813000.0 862200.0 ;
      RECT  802800.0 876000.0 813000.0 862200.0 ;
      RECT  802800.0 876000.0 813000.0 889800.0 ;
      RECT  802800.0 903600.0 813000.0 889800.0 ;
      RECT  802800.0 903600.0 813000.0 917400.0 ;
      RECT  802800.0 931200.0 813000.0 917400.0 ;
      RECT  802800.0 931200.0 813000.0 945000.0 ;
      RECT  802800.0 958800.0 813000.0 945000.0 ;
      RECT  802800.0 958800.0 813000.0 972600.0 ;
      RECT  802800.0 986400.0 813000.0 972600.0 ;
      RECT  802800.0 986400.0 813000.0 1000200.0 ;
      RECT  802800.0 1014000.0 813000.0 1000200.0 ;
      RECT  802800.0 1014000.0 813000.0 1027800.0 ;
      RECT  802800.0 1041600.0 813000.0 1027800.0 ;
      RECT  802800.0 1041600.0 813000.0 1055400.0 ;
      RECT  802800.0 1069200.0 813000.0 1055400.0 ;
      RECT  802800.0 1069200.0 813000.0 1083000.0 ;
      RECT  802800.0 1096800.0 813000.0 1083000.0 ;
      RECT  802800.0 1096800.0 813000.0 1110600.0 ;
      RECT  802800.0 1124400.0 813000.0 1110600.0 ;
      RECT  802800.0 1124400.0 813000.0 1138200.0 ;
      RECT  802800.0 1152000.0 813000.0 1138200.0 ;
      RECT  802800.0 1152000.0 813000.0 1165800.0 ;
      RECT  802800.0 1179600.0 813000.0 1165800.0 ;
      RECT  802800.0 1179600.0 813000.0 1193400.0 ;
      RECT  802800.0 1207200.0 813000.0 1193400.0 ;
      RECT  802800.0 1207200.0 813000.0 1221000.0 ;
      RECT  802800.0 1234800.0 813000.0 1221000.0 ;
      RECT  802800.0 1234800.0 813000.0 1248600.0 ;
      RECT  802800.0 1262400.0 813000.0 1248600.0 ;
      RECT  802800.0 1262400.0 813000.0 1276200.0 ;
      RECT  802800.0 1290000.0 813000.0 1276200.0 ;
      RECT  802800.0 1290000.0 813000.0 1303800.0 ;
      RECT  802800.0 1317600.0 813000.0 1303800.0 ;
      RECT  802800.0 1317600.0 813000.0 1331400.0 ;
      RECT  802800.0 1345200.0 813000.0 1331400.0 ;
      RECT  802800.0 1345200.0 813000.0 1359000.0 ;
      RECT  802800.0 1372800.0 813000.0 1359000.0 ;
      RECT  802800.0 1372800.0 813000.0 1386600.0 ;
      RECT  802800.0 1400400.0 813000.0 1386600.0 ;
      RECT  802800.0 1400400.0 813000.0 1414200.0 ;
      RECT  802800.0 1428000.0 813000.0 1414200.0 ;
      RECT  802800.0 1428000.0 813000.0 1441800.0 ;
      RECT  802800.0 1455600.0 813000.0 1441800.0 ;
      RECT  802800.0 1455600.0 813000.0 1469400.0 ;
      RECT  802800.0 1483200.0 813000.0 1469400.0 ;
      RECT  802800.0 1483200.0 813000.0 1497000.0 ;
      RECT  802800.0 1510800.0 813000.0 1497000.0 ;
      RECT  802800.0 1510800.0 813000.0 1524600.0 ;
      RECT  802800.0 1538400.0 813000.0 1524600.0 ;
      RECT  802800.0 1538400.0 813000.0 1552200.0 ;
      RECT  802800.0 1566000.0 813000.0 1552200.0 ;
      RECT  802800.0 1566000.0 813000.0 1579800.0 ;
      RECT  802800.0 1593600.0 813000.0 1579800.0 ;
      RECT  802800.0 1593600.0 813000.0 1607400.0 ;
      RECT  802800.0 1621200.0 813000.0 1607400.0 ;
      RECT  802800.0 1621200.0 813000.0 1635000.0 ;
      RECT  802800.0 1648800.0 813000.0 1635000.0 ;
      RECT  802800.0 1648800.0 813000.0 1662600.0 ;
      RECT  802800.0 1676400.0 813000.0 1662600.0 ;
      RECT  802800.0 1676400.0 813000.0 1690200.0 ;
      RECT  802800.0 1704000.0 813000.0 1690200.0 ;
      RECT  802800.0 1704000.0 813000.0 1717800.0 ;
      RECT  802800.0 1731600.0 813000.0 1717800.0 ;
      RECT  802800.0 1731600.0 813000.0 1745400.0 ;
      RECT  802800.0 1759200.0 813000.0 1745400.0 ;
      RECT  802800.0 1759200.0 813000.0 1773000.0 ;
      RECT  802800.0 1786800.0 813000.0 1773000.0 ;
      RECT  802800.0 1786800.0 813000.0 1800600.0 ;
      RECT  802800.0 1814400.0 813000.0 1800600.0 ;
      RECT  802800.0 1814400.0 813000.0 1828200.0 ;
      RECT  802800.0 1842000.0 813000.0 1828200.0 ;
      RECT  802800.0 1842000.0 813000.0 1855800.0 ;
      RECT  802800.0 1869600.0 813000.0 1855800.0 ;
      RECT  802800.0 1869600.0 813000.0 1883400.0 ;
      RECT  802800.0 1897200.0 813000.0 1883400.0 ;
      RECT  802800.0 1897200.0 813000.0 1911000.0 ;
      RECT  802800.0 1924800.0 813000.0 1911000.0 ;
      RECT  802800.0 1924800.0 813000.0 1938600.0 ;
      RECT  802800.0 1952400.0 813000.0 1938600.0 ;
      RECT  802800.0 1952400.0 813000.0 1966200.0 ;
      RECT  802800.0 1980000.0 813000.0 1966200.0 ;
      RECT  802800.0 1980000.0 813000.0 1993800.0 ;
      RECT  802800.0 2007600.0 813000.0 1993800.0 ;
      RECT  802800.0 2007600.0 813000.0 2021400.0 ;
      RECT  802800.0 2035200.0 813000.0 2021400.0 ;
      RECT  802800.0 2035200.0 813000.0 2049000.0 ;
      RECT  802800.0 2062800.0 813000.0 2049000.0 ;
      RECT  802800.0 2062800.0 813000.0 2076600.0 ;
      RECT  802800.0 2090400.0 813000.0 2076600.0 ;
      RECT  802800.0 2090400.0 813000.0 2104200.0 ;
      RECT  802800.0 2118000.0 813000.0 2104200.0 ;
      RECT  802800.0 2118000.0 813000.0 2131800.0 ;
      RECT  802800.0 2145600.0 813000.0 2131800.0 ;
      RECT  813000.0 379200.0 823200.0 393000.0 ;
      RECT  813000.0 406800.0 823200.0 393000.0 ;
      RECT  813000.0 406800.0 823200.0 420600.0 ;
      RECT  813000.0 434400.0 823200.0 420600.0 ;
      RECT  813000.0 434400.0 823200.0 448200.0 ;
      RECT  813000.0 462000.0 823200.0 448200.0 ;
      RECT  813000.0 462000.0 823200.0 475800.0 ;
      RECT  813000.0 489600.0 823200.0 475800.0 ;
      RECT  813000.0 489600.0 823200.0 503400.0 ;
      RECT  813000.0 517200.0 823200.0 503400.0 ;
      RECT  813000.0 517200.0 823200.0 531000.0 ;
      RECT  813000.0 544800.0 823200.0 531000.0 ;
      RECT  813000.0 544800.0 823200.0 558600.0 ;
      RECT  813000.0 572400.0 823200.0 558600.0 ;
      RECT  813000.0 572400.0 823200.0 586200.0 ;
      RECT  813000.0 600000.0 823200.0 586200.0 ;
      RECT  813000.0 600000.0 823200.0 613800.0 ;
      RECT  813000.0 627600.0 823200.0 613800.0 ;
      RECT  813000.0 627600.0 823200.0 641400.0 ;
      RECT  813000.0 655200.0 823200.0 641400.0 ;
      RECT  813000.0 655200.0 823200.0 669000.0 ;
      RECT  813000.0 682800.0 823200.0 669000.0 ;
      RECT  813000.0 682800.0 823200.0 696600.0 ;
      RECT  813000.0 710400.0 823200.0 696600.0 ;
      RECT  813000.0 710400.0 823200.0 724200.0 ;
      RECT  813000.0 738000.0 823200.0 724200.0 ;
      RECT  813000.0 738000.0 823200.0 751800.0 ;
      RECT  813000.0 765600.0 823200.0 751800.0 ;
      RECT  813000.0 765600.0 823200.0 779400.0 ;
      RECT  813000.0 793200.0 823200.0 779400.0 ;
      RECT  813000.0 793200.0 823200.0 807000.0 ;
      RECT  813000.0 820800.0 823200.0 807000.0 ;
      RECT  813000.0 820800.0 823200.0 834600.0 ;
      RECT  813000.0 848400.0 823200.0 834600.0 ;
      RECT  813000.0 848400.0 823200.0 862200.0 ;
      RECT  813000.0 876000.0 823200.0 862200.0 ;
      RECT  813000.0 876000.0 823200.0 889800.0 ;
      RECT  813000.0 903600.0 823200.0 889800.0 ;
      RECT  813000.0 903600.0 823200.0 917400.0 ;
      RECT  813000.0 931200.0 823200.0 917400.0 ;
      RECT  813000.0 931200.0 823200.0 945000.0 ;
      RECT  813000.0 958800.0 823200.0 945000.0 ;
      RECT  813000.0 958800.0 823200.0 972600.0 ;
      RECT  813000.0 986400.0 823200.0 972600.0 ;
      RECT  813000.0 986400.0 823200.0 1000200.0 ;
      RECT  813000.0 1014000.0 823200.0 1000200.0 ;
      RECT  813000.0 1014000.0 823200.0 1027800.0 ;
      RECT  813000.0 1041600.0 823200.0 1027800.0 ;
      RECT  813000.0 1041600.0 823200.0 1055400.0 ;
      RECT  813000.0 1069200.0 823200.0 1055400.0 ;
      RECT  813000.0 1069200.0 823200.0 1083000.0 ;
      RECT  813000.0 1096800.0 823200.0 1083000.0 ;
      RECT  813000.0 1096800.0 823200.0 1110600.0 ;
      RECT  813000.0 1124400.0 823200.0 1110600.0 ;
      RECT  813000.0 1124400.0 823200.0 1138200.0 ;
      RECT  813000.0 1152000.0 823200.0 1138200.0 ;
      RECT  813000.0 1152000.0 823200.0 1165800.0 ;
      RECT  813000.0 1179600.0 823200.0 1165800.0 ;
      RECT  813000.0 1179600.0 823200.0 1193400.0 ;
      RECT  813000.0 1207200.0 823200.0 1193400.0 ;
      RECT  813000.0 1207200.0 823200.0 1221000.0 ;
      RECT  813000.0 1234800.0 823200.0 1221000.0 ;
      RECT  813000.0 1234800.0 823200.0 1248600.0 ;
      RECT  813000.0 1262400.0 823200.0 1248600.0 ;
      RECT  813000.0 1262400.0 823200.0 1276200.0 ;
      RECT  813000.0 1290000.0 823200.0 1276200.0 ;
      RECT  813000.0 1290000.0 823200.0 1303800.0 ;
      RECT  813000.0 1317600.0 823200.0 1303800.0 ;
      RECT  813000.0 1317600.0 823200.0 1331400.0 ;
      RECT  813000.0 1345200.0 823200.0 1331400.0 ;
      RECT  813000.0 1345200.0 823200.0 1359000.0 ;
      RECT  813000.0 1372800.0 823200.0 1359000.0 ;
      RECT  813000.0 1372800.0 823200.0 1386600.0 ;
      RECT  813000.0 1400400.0 823200.0 1386600.0 ;
      RECT  813000.0 1400400.0 823200.0 1414200.0 ;
      RECT  813000.0 1428000.0 823200.0 1414200.0 ;
      RECT  813000.0 1428000.0 823200.0 1441800.0 ;
      RECT  813000.0 1455600.0 823200.0 1441800.0 ;
      RECT  813000.0 1455600.0 823200.0 1469400.0 ;
      RECT  813000.0 1483200.0 823200.0 1469400.0 ;
      RECT  813000.0 1483200.0 823200.0 1497000.0 ;
      RECT  813000.0 1510800.0 823200.0 1497000.0 ;
      RECT  813000.0 1510800.0 823200.0 1524600.0 ;
      RECT  813000.0 1538400.0 823200.0 1524600.0 ;
      RECT  813000.0 1538400.0 823200.0 1552200.0 ;
      RECT  813000.0 1566000.0 823200.0 1552200.0 ;
      RECT  813000.0 1566000.0 823200.0 1579800.0 ;
      RECT  813000.0 1593600.0 823200.0 1579800.0 ;
      RECT  813000.0 1593600.0 823200.0 1607400.0 ;
      RECT  813000.0 1621200.0 823200.0 1607400.0 ;
      RECT  813000.0 1621200.0 823200.0 1635000.0 ;
      RECT  813000.0 1648800.0 823200.0 1635000.0 ;
      RECT  813000.0 1648800.0 823200.0 1662600.0 ;
      RECT  813000.0 1676400.0 823200.0 1662600.0 ;
      RECT  813000.0 1676400.0 823200.0 1690200.0 ;
      RECT  813000.0 1704000.0 823200.0 1690200.0 ;
      RECT  813000.0 1704000.0 823200.0 1717800.0 ;
      RECT  813000.0 1731600.0 823200.0 1717800.0 ;
      RECT  813000.0 1731600.0 823200.0 1745400.0 ;
      RECT  813000.0 1759200.0 823200.0 1745400.0 ;
      RECT  813000.0 1759200.0 823200.0 1773000.0 ;
      RECT  813000.0 1786800.0 823200.0 1773000.0 ;
      RECT  813000.0 1786800.0 823200.0 1800600.0 ;
      RECT  813000.0 1814400.0 823200.0 1800600.0 ;
      RECT  813000.0 1814400.0 823200.0 1828200.0 ;
      RECT  813000.0 1842000.0 823200.0 1828200.0 ;
      RECT  813000.0 1842000.0 823200.0 1855800.0 ;
      RECT  813000.0 1869600.0 823200.0 1855800.0 ;
      RECT  813000.0 1869600.0 823200.0 1883400.0 ;
      RECT  813000.0 1897200.0 823200.0 1883400.0 ;
      RECT  813000.0 1897200.0 823200.0 1911000.0 ;
      RECT  813000.0 1924800.0 823200.0 1911000.0 ;
      RECT  813000.0 1924800.0 823200.0 1938600.0 ;
      RECT  813000.0 1952400.0 823200.0 1938600.0 ;
      RECT  813000.0 1952400.0 823200.0 1966200.0 ;
      RECT  813000.0 1980000.0 823200.0 1966200.0 ;
      RECT  813000.0 1980000.0 823200.0 1993800.0 ;
      RECT  813000.0 2007600.0 823200.0 1993800.0 ;
      RECT  813000.0 2007600.0 823200.0 2021400.0 ;
      RECT  813000.0 2035200.0 823200.0 2021400.0 ;
      RECT  813000.0 2035200.0 823200.0 2049000.0 ;
      RECT  813000.0 2062800.0 823200.0 2049000.0 ;
      RECT  813000.0 2062800.0 823200.0 2076600.0 ;
      RECT  813000.0 2090400.0 823200.0 2076600.0 ;
      RECT  813000.0 2090400.0 823200.0 2104200.0 ;
      RECT  813000.0 2118000.0 823200.0 2104200.0 ;
      RECT  813000.0 2118000.0 823200.0 2131800.0 ;
      RECT  813000.0 2145600.0 823200.0 2131800.0 ;
      RECT  823200.0 379200.0 833400.0 393000.0 ;
      RECT  823200.0 406800.0 833400.0 393000.0 ;
      RECT  823200.0 406800.0 833400.0 420600.0 ;
      RECT  823200.0 434400.0 833400.0 420600.0 ;
      RECT  823200.0 434400.0 833400.0 448200.0 ;
      RECT  823200.0 462000.0 833400.0 448200.0 ;
      RECT  823200.0 462000.0 833400.0 475800.0 ;
      RECT  823200.0 489600.0 833400.0 475800.0 ;
      RECT  823200.0 489600.0 833400.0 503400.0 ;
      RECT  823200.0 517200.0 833400.0 503400.0 ;
      RECT  823200.0 517200.0 833400.0 531000.0 ;
      RECT  823200.0 544800.0 833400.0 531000.0 ;
      RECT  823200.0 544800.0 833400.0 558600.0 ;
      RECT  823200.0 572400.0 833400.0 558600.0 ;
      RECT  823200.0 572400.0 833400.0 586200.0 ;
      RECT  823200.0 600000.0 833400.0 586200.0 ;
      RECT  823200.0 600000.0 833400.0 613800.0 ;
      RECT  823200.0 627600.0 833400.0 613800.0 ;
      RECT  823200.0 627600.0 833400.0 641400.0 ;
      RECT  823200.0 655200.0 833400.0 641400.0 ;
      RECT  823200.0 655200.0 833400.0 669000.0 ;
      RECT  823200.0 682800.0 833400.0 669000.0 ;
      RECT  823200.0 682800.0 833400.0 696600.0 ;
      RECT  823200.0 710400.0 833400.0 696600.0 ;
      RECT  823200.0 710400.0 833400.0 724200.0 ;
      RECT  823200.0 738000.0 833400.0 724200.0 ;
      RECT  823200.0 738000.0 833400.0 751800.0 ;
      RECT  823200.0 765600.0 833400.0 751800.0 ;
      RECT  823200.0 765600.0 833400.0 779400.0 ;
      RECT  823200.0 793200.0 833400.0 779400.0 ;
      RECT  823200.0 793200.0 833400.0 807000.0 ;
      RECT  823200.0 820800.0 833400.0 807000.0 ;
      RECT  823200.0 820800.0 833400.0 834600.0 ;
      RECT  823200.0 848400.0 833400.0 834600.0 ;
      RECT  823200.0 848400.0 833400.0 862200.0 ;
      RECT  823200.0 876000.0 833400.0 862200.0 ;
      RECT  823200.0 876000.0 833400.0 889800.0 ;
      RECT  823200.0 903600.0 833400.0 889800.0 ;
      RECT  823200.0 903600.0 833400.0 917400.0 ;
      RECT  823200.0 931200.0 833400.0 917400.0 ;
      RECT  823200.0 931200.0 833400.0 945000.0 ;
      RECT  823200.0 958800.0 833400.0 945000.0 ;
      RECT  823200.0 958800.0 833400.0 972600.0 ;
      RECT  823200.0 986400.0 833400.0 972600.0 ;
      RECT  823200.0 986400.0 833400.0 1000200.0 ;
      RECT  823200.0 1014000.0 833400.0 1000200.0 ;
      RECT  823200.0 1014000.0 833400.0 1027800.0 ;
      RECT  823200.0 1041600.0 833400.0 1027800.0 ;
      RECT  823200.0 1041600.0 833400.0 1055400.0 ;
      RECT  823200.0 1069200.0 833400.0 1055400.0 ;
      RECT  823200.0 1069200.0 833400.0 1083000.0 ;
      RECT  823200.0 1096800.0 833400.0 1083000.0 ;
      RECT  823200.0 1096800.0 833400.0 1110600.0 ;
      RECT  823200.0 1124400.0 833400.0 1110600.0 ;
      RECT  823200.0 1124400.0 833400.0 1138200.0 ;
      RECT  823200.0 1152000.0 833400.0 1138200.0 ;
      RECT  823200.0 1152000.0 833400.0 1165800.0 ;
      RECT  823200.0 1179600.0 833400.0 1165800.0 ;
      RECT  823200.0 1179600.0 833400.0 1193400.0 ;
      RECT  823200.0 1207200.0 833400.0 1193400.0 ;
      RECT  823200.0 1207200.0 833400.0 1221000.0 ;
      RECT  823200.0 1234800.0 833400.0 1221000.0 ;
      RECT  823200.0 1234800.0 833400.0 1248600.0 ;
      RECT  823200.0 1262400.0 833400.0 1248600.0 ;
      RECT  823200.0 1262400.0 833400.0 1276200.0 ;
      RECT  823200.0 1290000.0 833400.0 1276200.0 ;
      RECT  823200.0 1290000.0 833400.0 1303800.0 ;
      RECT  823200.0 1317600.0 833400.0 1303800.0 ;
      RECT  823200.0 1317600.0 833400.0 1331400.0 ;
      RECT  823200.0 1345200.0 833400.0 1331400.0 ;
      RECT  823200.0 1345200.0 833400.0 1359000.0 ;
      RECT  823200.0 1372800.0 833400.0 1359000.0 ;
      RECT  823200.0 1372800.0 833400.0 1386600.0 ;
      RECT  823200.0 1400400.0 833400.0 1386600.0 ;
      RECT  823200.0 1400400.0 833400.0 1414200.0 ;
      RECT  823200.0 1428000.0 833400.0 1414200.0 ;
      RECT  823200.0 1428000.0 833400.0 1441800.0 ;
      RECT  823200.0 1455600.0 833400.0 1441800.0 ;
      RECT  823200.0 1455600.0 833400.0 1469400.0 ;
      RECT  823200.0 1483200.0 833400.0 1469400.0 ;
      RECT  823200.0 1483200.0 833400.0 1497000.0 ;
      RECT  823200.0 1510800.0 833400.0 1497000.0 ;
      RECT  823200.0 1510800.0 833400.0 1524600.0 ;
      RECT  823200.0 1538400.0 833400.0 1524600.0 ;
      RECT  823200.0 1538400.0 833400.0 1552200.0 ;
      RECT  823200.0 1566000.0 833400.0 1552200.0 ;
      RECT  823200.0 1566000.0 833400.0 1579800.0 ;
      RECT  823200.0 1593600.0 833400.0 1579800.0 ;
      RECT  823200.0 1593600.0 833400.0 1607400.0 ;
      RECT  823200.0 1621200.0 833400.0 1607400.0 ;
      RECT  823200.0 1621200.0 833400.0 1635000.0 ;
      RECT  823200.0 1648800.0 833400.0 1635000.0 ;
      RECT  823200.0 1648800.0 833400.0 1662600.0 ;
      RECT  823200.0 1676400.0 833400.0 1662600.0 ;
      RECT  823200.0 1676400.0 833400.0 1690200.0 ;
      RECT  823200.0 1704000.0 833400.0 1690200.0 ;
      RECT  823200.0 1704000.0 833400.0 1717800.0 ;
      RECT  823200.0 1731600.0 833400.0 1717800.0 ;
      RECT  823200.0 1731600.0 833400.0 1745400.0 ;
      RECT  823200.0 1759200.0 833400.0 1745400.0 ;
      RECT  823200.0 1759200.0 833400.0 1773000.0 ;
      RECT  823200.0 1786800.0 833400.0 1773000.0 ;
      RECT  823200.0 1786800.0 833400.0 1800600.0 ;
      RECT  823200.0 1814400.0 833400.0 1800600.0 ;
      RECT  823200.0 1814400.0 833400.0 1828200.0 ;
      RECT  823200.0 1842000.0 833400.0 1828200.0 ;
      RECT  823200.0 1842000.0 833400.0 1855800.0 ;
      RECT  823200.0 1869600.0 833400.0 1855800.0 ;
      RECT  823200.0 1869600.0 833400.0 1883400.0 ;
      RECT  823200.0 1897200.0 833400.0 1883400.0 ;
      RECT  823200.0 1897200.0 833400.0 1911000.0 ;
      RECT  823200.0 1924800.0 833400.0 1911000.0 ;
      RECT  823200.0 1924800.0 833400.0 1938600.0 ;
      RECT  823200.0 1952400.0 833400.0 1938600.0 ;
      RECT  823200.0 1952400.0 833400.0 1966200.0 ;
      RECT  823200.0 1980000.0 833400.0 1966200.0 ;
      RECT  823200.0 1980000.0 833400.0 1993800.0 ;
      RECT  823200.0 2007600.0 833400.0 1993800.0 ;
      RECT  823200.0 2007600.0 833400.0 2021400.0 ;
      RECT  823200.0 2035200.0 833400.0 2021400.0 ;
      RECT  823200.0 2035200.0 833400.0 2049000.0 ;
      RECT  823200.0 2062800.0 833400.0 2049000.0 ;
      RECT  823200.0 2062800.0 833400.0 2076600.0 ;
      RECT  823200.0 2090400.0 833400.0 2076600.0 ;
      RECT  823200.0 2090400.0 833400.0 2104200.0 ;
      RECT  823200.0 2118000.0 833400.0 2104200.0 ;
      RECT  823200.0 2118000.0 833400.0 2131800.0 ;
      RECT  823200.0 2145600.0 833400.0 2131800.0 ;
      RECT  833400.0 379200.0 843600.0 393000.0 ;
      RECT  833400.0 406800.0 843600.0 393000.0 ;
      RECT  833400.0 406800.0 843600.0 420600.0 ;
      RECT  833400.0 434400.0 843600.0 420600.0 ;
      RECT  833400.0 434400.0 843600.0 448200.0 ;
      RECT  833400.0 462000.0 843600.0 448200.0 ;
      RECT  833400.0 462000.0 843600.0 475800.0 ;
      RECT  833400.0 489600.0 843600.0 475800.0 ;
      RECT  833400.0 489600.0 843600.0 503400.0 ;
      RECT  833400.0 517200.0 843600.0 503400.0 ;
      RECT  833400.0 517200.0 843600.0 531000.0 ;
      RECT  833400.0 544800.0 843600.0 531000.0 ;
      RECT  833400.0 544800.0 843600.0 558600.0 ;
      RECT  833400.0 572400.0 843600.0 558600.0 ;
      RECT  833400.0 572400.0 843600.0 586200.0 ;
      RECT  833400.0 600000.0 843600.0 586200.0 ;
      RECT  833400.0 600000.0 843600.0 613800.0 ;
      RECT  833400.0 627600.0 843600.0 613800.0 ;
      RECT  833400.0 627600.0 843600.0 641400.0 ;
      RECT  833400.0 655200.0 843600.0 641400.0 ;
      RECT  833400.0 655200.0 843600.0 669000.0 ;
      RECT  833400.0 682800.0 843600.0 669000.0 ;
      RECT  833400.0 682800.0 843600.0 696600.0 ;
      RECT  833400.0 710400.0 843600.0 696600.0 ;
      RECT  833400.0 710400.0 843600.0 724200.0 ;
      RECT  833400.0 738000.0 843600.0 724200.0 ;
      RECT  833400.0 738000.0 843600.0 751800.0 ;
      RECT  833400.0 765600.0 843600.0 751800.0 ;
      RECT  833400.0 765600.0 843600.0 779400.0 ;
      RECT  833400.0 793200.0 843600.0 779400.0 ;
      RECT  833400.0 793200.0 843600.0 807000.0 ;
      RECT  833400.0 820800.0 843600.0 807000.0 ;
      RECT  833400.0 820800.0 843600.0 834600.0 ;
      RECT  833400.0 848400.0 843600.0 834600.0 ;
      RECT  833400.0 848400.0 843600.0 862200.0 ;
      RECT  833400.0 876000.0 843600.0 862200.0 ;
      RECT  833400.0 876000.0 843600.0 889800.0 ;
      RECT  833400.0 903600.0 843600.0 889800.0 ;
      RECT  833400.0 903600.0 843600.0 917400.0 ;
      RECT  833400.0 931200.0 843600.0 917400.0 ;
      RECT  833400.0 931200.0 843600.0 945000.0 ;
      RECT  833400.0 958800.0 843600.0 945000.0 ;
      RECT  833400.0 958800.0 843600.0 972600.0 ;
      RECT  833400.0 986400.0 843600.0 972600.0 ;
      RECT  833400.0 986400.0 843600.0 1000200.0 ;
      RECT  833400.0 1014000.0 843600.0 1000200.0 ;
      RECT  833400.0 1014000.0 843600.0 1027800.0 ;
      RECT  833400.0 1041600.0 843600.0 1027800.0 ;
      RECT  833400.0 1041600.0 843600.0 1055400.0 ;
      RECT  833400.0 1069200.0 843600.0 1055400.0 ;
      RECT  833400.0 1069200.0 843600.0 1083000.0 ;
      RECT  833400.0 1096800.0 843600.0 1083000.0 ;
      RECT  833400.0 1096800.0 843600.0 1110600.0 ;
      RECT  833400.0 1124400.0 843600.0 1110600.0 ;
      RECT  833400.0 1124400.0 843600.0 1138200.0 ;
      RECT  833400.0 1152000.0 843600.0 1138200.0 ;
      RECT  833400.0 1152000.0 843600.0 1165800.0 ;
      RECT  833400.0 1179600.0 843600.0 1165800.0 ;
      RECT  833400.0 1179600.0 843600.0 1193400.0 ;
      RECT  833400.0 1207200.0 843600.0 1193400.0 ;
      RECT  833400.0 1207200.0 843600.0 1221000.0 ;
      RECT  833400.0 1234800.0 843600.0 1221000.0 ;
      RECT  833400.0 1234800.0 843600.0 1248600.0 ;
      RECT  833400.0 1262400.0 843600.0 1248600.0 ;
      RECT  833400.0 1262400.0 843600.0 1276200.0 ;
      RECT  833400.0 1290000.0 843600.0 1276200.0 ;
      RECT  833400.0 1290000.0 843600.0 1303800.0 ;
      RECT  833400.0 1317600.0 843600.0 1303800.0 ;
      RECT  833400.0 1317600.0 843600.0 1331400.0 ;
      RECT  833400.0 1345200.0 843600.0 1331400.0 ;
      RECT  833400.0 1345200.0 843600.0 1359000.0 ;
      RECT  833400.0 1372800.0 843600.0 1359000.0 ;
      RECT  833400.0 1372800.0 843600.0 1386600.0 ;
      RECT  833400.0 1400400.0 843600.0 1386600.0 ;
      RECT  833400.0 1400400.0 843600.0 1414200.0 ;
      RECT  833400.0 1428000.0 843600.0 1414200.0 ;
      RECT  833400.0 1428000.0 843600.0 1441800.0 ;
      RECT  833400.0 1455600.0 843600.0 1441800.0 ;
      RECT  833400.0 1455600.0 843600.0 1469400.0 ;
      RECT  833400.0 1483200.0 843600.0 1469400.0 ;
      RECT  833400.0 1483200.0 843600.0 1497000.0 ;
      RECT  833400.0 1510800.0 843600.0 1497000.0 ;
      RECT  833400.0 1510800.0 843600.0 1524600.0 ;
      RECT  833400.0 1538400.0 843600.0 1524600.0 ;
      RECT  833400.0 1538400.0 843600.0 1552200.0 ;
      RECT  833400.0 1566000.0 843600.0 1552200.0 ;
      RECT  833400.0 1566000.0 843600.0 1579800.0 ;
      RECT  833400.0 1593600.0 843600.0 1579800.0 ;
      RECT  833400.0 1593600.0 843600.0 1607400.0 ;
      RECT  833400.0 1621200.0 843600.0 1607400.0 ;
      RECT  833400.0 1621200.0 843600.0 1635000.0 ;
      RECT  833400.0 1648800.0 843600.0 1635000.0 ;
      RECT  833400.0 1648800.0 843600.0 1662600.0 ;
      RECT  833400.0 1676400.0 843600.0 1662600.0 ;
      RECT  833400.0 1676400.0 843600.0 1690200.0 ;
      RECT  833400.0 1704000.0 843600.0 1690200.0 ;
      RECT  833400.0 1704000.0 843600.0 1717800.0 ;
      RECT  833400.0 1731600.0 843600.0 1717800.0 ;
      RECT  833400.0 1731600.0 843600.0 1745400.0 ;
      RECT  833400.0 1759200.0 843600.0 1745400.0 ;
      RECT  833400.0 1759200.0 843600.0 1773000.0 ;
      RECT  833400.0 1786800.0 843600.0 1773000.0 ;
      RECT  833400.0 1786800.0 843600.0 1800600.0 ;
      RECT  833400.0 1814400.0 843600.0 1800600.0 ;
      RECT  833400.0 1814400.0 843600.0 1828200.0 ;
      RECT  833400.0 1842000.0 843600.0 1828200.0 ;
      RECT  833400.0 1842000.0 843600.0 1855800.0 ;
      RECT  833400.0 1869600.0 843600.0 1855800.0 ;
      RECT  833400.0 1869600.0 843600.0 1883400.0 ;
      RECT  833400.0 1897200.0 843600.0 1883400.0 ;
      RECT  833400.0 1897200.0 843600.0 1911000.0 ;
      RECT  833400.0 1924800.0 843600.0 1911000.0 ;
      RECT  833400.0 1924800.0 843600.0 1938600.0 ;
      RECT  833400.0 1952400.0 843600.0 1938600.0 ;
      RECT  833400.0 1952400.0 843600.0 1966200.0 ;
      RECT  833400.0 1980000.0 843600.0 1966200.0 ;
      RECT  833400.0 1980000.0 843600.0 1993800.0 ;
      RECT  833400.0 2007600.0 843600.0 1993800.0 ;
      RECT  833400.0 2007600.0 843600.0 2021400.0 ;
      RECT  833400.0 2035200.0 843600.0 2021400.0 ;
      RECT  833400.0 2035200.0 843600.0 2049000.0 ;
      RECT  833400.0 2062800.0 843600.0 2049000.0 ;
      RECT  833400.0 2062800.0 843600.0 2076600.0 ;
      RECT  833400.0 2090400.0 843600.0 2076600.0 ;
      RECT  833400.0 2090400.0 843600.0 2104200.0 ;
      RECT  833400.0 2118000.0 843600.0 2104200.0 ;
      RECT  833400.0 2118000.0 843600.0 2131800.0 ;
      RECT  833400.0 2145600.0 843600.0 2131800.0 ;
      RECT  843600.0 379200.0 853800.0 393000.0 ;
      RECT  843600.0 406800.0 853800.0 393000.0 ;
      RECT  843600.0 406800.0 853800.0 420600.0 ;
      RECT  843600.0 434400.0 853800.0 420600.0 ;
      RECT  843600.0 434400.0 853800.0 448200.0 ;
      RECT  843600.0 462000.0 853800.0 448200.0 ;
      RECT  843600.0 462000.0 853800.0 475800.0 ;
      RECT  843600.0 489600.0 853800.0 475800.0 ;
      RECT  843600.0 489600.0 853800.0 503400.0 ;
      RECT  843600.0 517200.0 853800.0 503400.0 ;
      RECT  843600.0 517200.0 853800.0 531000.0 ;
      RECT  843600.0 544800.0 853800.0 531000.0 ;
      RECT  843600.0 544800.0 853800.0 558600.0 ;
      RECT  843600.0 572400.0 853800.0 558600.0 ;
      RECT  843600.0 572400.0 853800.0 586200.0 ;
      RECT  843600.0 600000.0 853800.0 586200.0 ;
      RECT  843600.0 600000.0 853800.0 613800.0 ;
      RECT  843600.0 627600.0 853800.0 613800.0 ;
      RECT  843600.0 627600.0 853800.0 641400.0 ;
      RECT  843600.0 655200.0 853800.0 641400.0 ;
      RECT  843600.0 655200.0 853800.0 669000.0 ;
      RECT  843600.0 682800.0 853800.0 669000.0 ;
      RECT  843600.0 682800.0 853800.0 696600.0 ;
      RECT  843600.0 710400.0 853800.0 696600.0 ;
      RECT  843600.0 710400.0 853800.0 724200.0 ;
      RECT  843600.0 738000.0 853800.0 724200.0 ;
      RECT  843600.0 738000.0 853800.0 751800.0 ;
      RECT  843600.0 765600.0 853800.0 751800.0 ;
      RECT  843600.0 765600.0 853800.0 779400.0 ;
      RECT  843600.0 793200.0 853800.0 779400.0 ;
      RECT  843600.0 793200.0 853800.0 807000.0 ;
      RECT  843600.0 820800.0 853800.0 807000.0 ;
      RECT  843600.0 820800.0 853800.0 834600.0 ;
      RECT  843600.0 848400.0 853800.0 834600.0 ;
      RECT  843600.0 848400.0 853800.0 862200.0 ;
      RECT  843600.0 876000.0 853800.0 862200.0 ;
      RECT  843600.0 876000.0 853800.0 889800.0 ;
      RECT  843600.0 903600.0 853800.0 889800.0 ;
      RECT  843600.0 903600.0 853800.0 917400.0 ;
      RECT  843600.0 931200.0 853800.0 917400.0 ;
      RECT  843600.0 931200.0 853800.0 945000.0 ;
      RECT  843600.0 958800.0 853800.0 945000.0 ;
      RECT  843600.0 958800.0 853800.0 972600.0 ;
      RECT  843600.0 986400.0 853800.0 972600.0 ;
      RECT  843600.0 986400.0 853800.0 1000200.0 ;
      RECT  843600.0 1014000.0 853800.0 1000200.0 ;
      RECT  843600.0 1014000.0 853800.0 1027800.0 ;
      RECT  843600.0 1041600.0 853800.0 1027800.0 ;
      RECT  843600.0 1041600.0 853800.0 1055400.0 ;
      RECT  843600.0 1069200.0 853800.0 1055400.0 ;
      RECT  843600.0 1069200.0 853800.0 1083000.0 ;
      RECT  843600.0 1096800.0 853800.0 1083000.0 ;
      RECT  843600.0 1096800.0 853800.0 1110600.0 ;
      RECT  843600.0 1124400.0 853800.0 1110600.0 ;
      RECT  843600.0 1124400.0 853800.0 1138200.0 ;
      RECT  843600.0 1152000.0 853800.0 1138200.0 ;
      RECT  843600.0 1152000.0 853800.0 1165800.0 ;
      RECT  843600.0 1179600.0 853800.0 1165800.0 ;
      RECT  843600.0 1179600.0 853800.0 1193400.0 ;
      RECT  843600.0 1207200.0 853800.0 1193400.0 ;
      RECT  843600.0 1207200.0 853800.0 1221000.0 ;
      RECT  843600.0 1234800.0 853800.0 1221000.0 ;
      RECT  843600.0 1234800.0 853800.0 1248600.0 ;
      RECT  843600.0 1262400.0 853800.0 1248600.0 ;
      RECT  843600.0 1262400.0 853800.0 1276200.0 ;
      RECT  843600.0 1290000.0 853800.0 1276200.0 ;
      RECT  843600.0 1290000.0 853800.0 1303800.0 ;
      RECT  843600.0 1317600.0 853800.0 1303800.0 ;
      RECT  843600.0 1317600.0 853800.0 1331400.0 ;
      RECT  843600.0 1345200.0 853800.0 1331400.0 ;
      RECT  843600.0 1345200.0 853800.0 1359000.0 ;
      RECT  843600.0 1372800.0 853800.0 1359000.0 ;
      RECT  843600.0 1372800.0 853800.0 1386600.0 ;
      RECT  843600.0 1400400.0 853800.0 1386600.0 ;
      RECT  843600.0 1400400.0 853800.0 1414200.0 ;
      RECT  843600.0 1428000.0 853800.0 1414200.0 ;
      RECT  843600.0 1428000.0 853800.0 1441800.0 ;
      RECT  843600.0 1455600.0 853800.0 1441800.0 ;
      RECT  843600.0 1455600.0 853800.0 1469400.0 ;
      RECT  843600.0 1483200.0 853800.0 1469400.0 ;
      RECT  843600.0 1483200.0 853800.0 1497000.0 ;
      RECT  843600.0 1510800.0 853800.0 1497000.0 ;
      RECT  843600.0 1510800.0 853800.0 1524600.0 ;
      RECT  843600.0 1538400.0 853800.0 1524600.0 ;
      RECT  843600.0 1538400.0 853800.0 1552200.0 ;
      RECT  843600.0 1566000.0 853800.0 1552200.0 ;
      RECT  843600.0 1566000.0 853800.0 1579800.0 ;
      RECT  843600.0 1593600.0 853800.0 1579800.0 ;
      RECT  843600.0 1593600.0 853800.0 1607400.0 ;
      RECT  843600.0 1621200.0 853800.0 1607400.0 ;
      RECT  843600.0 1621200.0 853800.0 1635000.0 ;
      RECT  843600.0 1648800.0 853800.0 1635000.0 ;
      RECT  843600.0 1648800.0 853800.0 1662600.0 ;
      RECT  843600.0 1676400.0 853800.0 1662600.0 ;
      RECT  843600.0 1676400.0 853800.0 1690200.0 ;
      RECT  843600.0 1704000.0 853800.0 1690200.0 ;
      RECT  843600.0 1704000.0 853800.0 1717800.0 ;
      RECT  843600.0 1731600.0 853800.0 1717800.0 ;
      RECT  843600.0 1731600.0 853800.0 1745400.0 ;
      RECT  843600.0 1759200.0 853800.0 1745400.0 ;
      RECT  843600.0 1759200.0 853800.0 1773000.0 ;
      RECT  843600.0 1786800.0 853800.0 1773000.0 ;
      RECT  843600.0 1786800.0 853800.0 1800600.0 ;
      RECT  843600.0 1814400.0 853800.0 1800600.0 ;
      RECT  843600.0 1814400.0 853800.0 1828200.0 ;
      RECT  843600.0 1842000.0 853800.0 1828200.0 ;
      RECT  843600.0 1842000.0 853800.0 1855800.0 ;
      RECT  843600.0 1869600.0 853800.0 1855800.0 ;
      RECT  843600.0 1869600.0 853800.0 1883400.0 ;
      RECT  843600.0 1897200.0 853800.0 1883400.0 ;
      RECT  843600.0 1897200.0 853800.0 1911000.0 ;
      RECT  843600.0 1924800.0 853800.0 1911000.0 ;
      RECT  843600.0 1924800.0 853800.0 1938600.0 ;
      RECT  843600.0 1952400.0 853800.0 1938600.0 ;
      RECT  843600.0 1952400.0 853800.0 1966200.0 ;
      RECT  843600.0 1980000.0 853800.0 1966200.0 ;
      RECT  843600.0 1980000.0 853800.0 1993800.0 ;
      RECT  843600.0 2007600.0 853800.0 1993800.0 ;
      RECT  843600.0 2007600.0 853800.0 2021400.0 ;
      RECT  843600.0 2035200.0 853800.0 2021400.0 ;
      RECT  843600.0 2035200.0 853800.0 2049000.0 ;
      RECT  843600.0 2062800.0 853800.0 2049000.0 ;
      RECT  843600.0 2062800.0 853800.0 2076600.0 ;
      RECT  843600.0 2090400.0 853800.0 2076600.0 ;
      RECT  843600.0 2090400.0 853800.0 2104200.0 ;
      RECT  843600.0 2118000.0 853800.0 2104200.0 ;
      RECT  843600.0 2118000.0 853800.0 2131800.0 ;
      RECT  843600.0 2145600.0 853800.0 2131800.0 ;
      RECT  853800.0 379200.0 864000.0 393000.0 ;
      RECT  853800.0 406800.0 864000.0 393000.0 ;
      RECT  853800.0 406800.0 864000.0 420600.0 ;
      RECT  853800.0 434400.0 864000.0 420600.0 ;
      RECT  853800.0 434400.0 864000.0 448200.0 ;
      RECT  853800.0 462000.0 864000.0 448200.0 ;
      RECT  853800.0 462000.0 864000.0 475800.0 ;
      RECT  853800.0 489600.0 864000.0 475800.0 ;
      RECT  853800.0 489600.0 864000.0 503400.0 ;
      RECT  853800.0 517200.0 864000.0 503400.0 ;
      RECT  853800.0 517200.0 864000.0 531000.0 ;
      RECT  853800.0 544800.0 864000.0 531000.0 ;
      RECT  853800.0 544800.0 864000.0 558600.0 ;
      RECT  853800.0 572400.0 864000.0 558600.0 ;
      RECT  853800.0 572400.0 864000.0 586200.0 ;
      RECT  853800.0 600000.0 864000.0 586200.0 ;
      RECT  853800.0 600000.0 864000.0 613800.0 ;
      RECT  853800.0 627600.0 864000.0 613800.0 ;
      RECT  853800.0 627600.0 864000.0 641400.0 ;
      RECT  853800.0 655200.0 864000.0 641400.0 ;
      RECT  853800.0 655200.0 864000.0 669000.0 ;
      RECT  853800.0 682800.0 864000.0 669000.0 ;
      RECT  853800.0 682800.0 864000.0 696600.0 ;
      RECT  853800.0 710400.0 864000.0 696600.0 ;
      RECT  853800.0 710400.0 864000.0 724200.0 ;
      RECT  853800.0 738000.0 864000.0 724200.0 ;
      RECT  853800.0 738000.0 864000.0 751800.0 ;
      RECT  853800.0 765600.0 864000.0 751800.0 ;
      RECT  853800.0 765600.0 864000.0 779400.0 ;
      RECT  853800.0 793200.0 864000.0 779400.0 ;
      RECT  853800.0 793200.0 864000.0 807000.0 ;
      RECT  853800.0 820800.0 864000.0 807000.0 ;
      RECT  853800.0 820800.0 864000.0 834600.0 ;
      RECT  853800.0 848400.0 864000.0 834600.0 ;
      RECT  853800.0 848400.0 864000.0 862200.0 ;
      RECT  853800.0 876000.0 864000.0 862200.0 ;
      RECT  853800.0 876000.0 864000.0 889800.0 ;
      RECT  853800.0 903600.0 864000.0 889800.0 ;
      RECT  853800.0 903600.0 864000.0 917400.0 ;
      RECT  853800.0 931200.0 864000.0 917400.0 ;
      RECT  853800.0 931200.0 864000.0 945000.0 ;
      RECT  853800.0 958800.0 864000.0 945000.0 ;
      RECT  853800.0 958800.0 864000.0 972600.0 ;
      RECT  853800.0 986400.0 864000.0 972600.0 ;
      RECT  853800.0 986400.0 864000.0 1000200.0 ;
      RECT  853800.0 1014000.0 864000.0 1000200.0 ;
      RECT  853800.0 1014000.0 864000.0 1027800.0 ;
      RECT  853800.0 1041600.0 864000.0 1027800.0 ;
      RECT  853800.0 1041600.0 864000.0 1055400.0 ;
      RECT  853800.0 1069200.0 864000.0 1055400.0 ;
      RECT  853800.0 1069200.0 864000.0 1083000.0 ;
      RECT  853800.0 1096800.0 864000.0 1083000.0 ;
      RECT  853800.0 1096800.0 864000.0 1110600.0 ;
      RECT  853800.0 1124400.0 864000.0 1110600.0 ;
      RECT  853800.0 1124400.0 864000.0 1138200.0 ;
      RECT  853800.0 1152000.0 864000.0 1138200.0 ;
      RECT  853800.0 1152000.0 864000.0 1165800.0 ;
      RECT  853800.0 1179600.0 864000.0 1165800.0 ;
      RECT  853800.0 1179600.0 864000.0 1193400.0 ;
      RECT  853800.0 1207200.0 864000.0 1193400.0 ;
      RECT  853800.0 1207200.0 864000.0 1221000.0 ;
      RECT  853800.0 1234800.0 864000.0 1221000.0 ;
      RECT  853800.0 1234800.0 864000.0 1248600.0 ;
      RECT  853800.0 1262400.0 864000.0 1248600.0 ;
      RECT  853800.0 1262400.0 864000.0 1276200.0 ;
      RECT  853800.0 1290000.0 864000.0 1276200.0 ;
      RECT  853800.0 1290000.0 864000.0 1303800.0 ;
      RECT  853800.0 1317600.0 864000.0 1303800.0 ;
      RECT  853800.0 1317600.0 864000.0 1331400.0 ;
      RECT  853800.0 1345200.0 864000.0 1331400.0 ;
      RECT  853800.0 1345200.0 864000.0 1359000.0 ;
      RECT  853800.0 1372800.0 864000.0 1359000.0 ;
      RECT  853800.0 1372800.0 864000.0 1386600.0 ;
      RECT  853800.0 1400400.0 864000.0 1386600.0 ;
      RECT  853800.0 1400400.0 864000.0 1414200.0 ;
      RECT  853800.0 1428000.0 864000.0 1414200.0 ;
      RECT  853800.0 1428000.0 864000.0 1441800.0 ;
      RECT  853800.0 1455600.0 864000.0 1441800.0 ;
      RECT  853800.0 1455600.0 864000.0 1469400.0 ;
      RECT  853800.0 1483200.0 864000.0 1469400.0 ;
      RECT  853800.0 1483200.0 864000.0 1497000.0 ;
      RECT  853800.0 1510800.0 864000.0 1497000.0 ;
      RECT  853800.0 1510800.0 864000.0 1524600.0 ;
      RECT  853800.0 1538400.0 864000.0 1524600.0 ;
      RECT  853800.0 1538400.0 864000.0 1552200.0 ;
      RECT  853800.0 1566000.0 864000.0 1552200.0 ;
      RECT  853800.0 1566000.0 864000.0 1579800.0 ;
      RECT  853800.0 1593600.0 864000.0 1579800.0 ;
      RECT  853800.0 1593600.0 864000.0 1607400.0 ;
      RECT  853800.0 1621200.0 864000.0 1607400.0 ;
      RECT  853800.0 1621200.0 864000.0 1635000.0 ;
      RECT  853800.0 1648800.0 864000.0 1635000.0 ;
      RECT  853800.0 1648800.0 864000.0 1662600.0 ;
      RECT  853800.0 1676400.0 864000.0 1662600.0 ;
      RECT  853800.0 1676400.0 864000.0 1690200.0 ;
      RECT  853800.0 1704000.0 864000.0 1690200.0 ;
      RECT  853800.0 1704000.0 864000.0 1717800.0 ;
      RECT  853800.0 1731600.0 864000.0 1717800.0 ;
      RECT  853800.0 1731600.0 864000.0 1745400.0 ;
      RECT  853800.0 1759200.0 864000.0 1745400.0 ;
      RECT  853800.0 1759200.0 864000.0 1773000.0 ;
      RECT  853800.0 1786800.0 864000.0 1773000.0 ;
      RECT  853800.0 1786800.0 864000.0 1800600.0 ;
      RECT  853800.0 1814400.0 864000.0 1800600.0 ;
      RECT  853800.0 1814400.0 864000.0 1828200.0 ;
      RECT  853800.0 1842000.0 864000.0 1828200.0 ;
      RECT  853800.0 1842000.0 864000.0 1855800.0 ;
      RECT  853800.0 1869600.0 864000.0 1855800.0 ;
      RECT  853800.0 1869600.0 864000.0 1883400.0 ;
      RECT  853800.0 1897200.0 864000.0 1883400.0 ;
      RECT  853800.0 1897200.0 864000.0 1911000.0 ;
      RECT  853800.0 1924800.0 864000.0 1911000.0 ;
      RECT  853800.0 1924800.0 864000.0 1938600.0 ;
      RECT  853800.0 1952400.0 864000.0 1938600.0 ;
      RECT  853800.0 1952400.0 864000.0 1966200.0 ;
      RECT  853800.0 1980000.0 864000.0 1966200.0 ;
      RECT  853800.0 1980000.0 864000.0 1993800.0 ;
      RECT  853800.0 2007600.0 864000.0 1993800.0 ;
      RECT  853800.0 2007600.0 864000.0 2021400.0 ;
      RECT  853800.0 2035200.0 864000.0 2021400.0 ;
      RECT  853800.0 2035200.0 864000.0 2049000.0 ;
      RECT  853800.0 2062800.0 864000.0 2049000.0 ;
      RECT  853800.0 2062800.0 864000.0 2076600.0 ;
      RECT  853800.0 2090400.0 864000.0 2076600.0 ;
      RECT  853800.0 2090400.0 864000.0 2104200.0 ;
      RECT  853800.0 2118000.0 864000.0 2104200.0 ;
      RECT  853800.0 2118000.0 864000.0 2131800.0 ;
      RECT  853800.0 2145600.0 864000.0 2131800.0 ;
      RECT  864000.0 379200.0 874200.0 393000.0 ;
      RECT  864000.0 406800.0 874200.0 393000.0 ;
      RECT  864000.0 406800.0 874200.0 420600.0 ;
      RECT  864000.0 434400.0 874200.0 420600.0 ;
      RECT  864000.0 434400.0 874200.0 448200.0 ;
      RECT  864000.0 462000.0 874200.0 448200.0 ;
      RECT  864000.0 462000.0 874200.0 475800.0 ;
      RECT  864000.0 489600.0 874200.0 475800.0 ;
      RECT  864000.0 489600.0 874200.0 503400.0 ;
      RECT  864000.0 517200.0 874200.0 503400.0 ;
      RECT  864000.0 517200.0 874200.0 531000.0 ;
      RECT  864000.0 544800.0 874200.0 531000.0 ;
      RECT  864000.0 544800.0 874200.0 558600.0 ;
      RECT  864000.0 572400.0 874200.0 558600.0 ;
      RECT  864000.0 572400.0 874200.0 586200.0 ;
      RECT  864000.0 600000.0 874200.0 586200.0 ;
      RECT  864000.0 600000.0 874200.0 613800.0 ;
      RECT  864000.0 627600.0 874200.0 613800.0 ;
      RECT  864000.0 627600.0 874200.0 641400.0 ;
      RECT  864000.0 655200.0 874200.0 641400.0 ;
      RECT  864000.0 655200.0 874200.0 669000.0 ;
      RECT  864000.0 682800.0 874200.0 669000.0 ;
      RECT  864000.0 682800.0 874200.0 696600.0 ;
      RECT  864000.0 710400.0 874200.0 696600.0 ;
      RECT  864000.0 710400.0 874200.0 724200.0 ;
      RECT  864000.0 738000.0 874200.0 724200.0 ;
      RECT  864000.0 738000.0 874200.0 751800.0 ;
      RECT  864000.0 765600.0 874200.0 751800.0 ;
      RECT  864000.0 765600.0 874200.0 779400.0 ;
      RECT  864000.0 793200.0 874200.0 779400.0 ;
      RECT  864000.0 793200.0 874200.0 807000.0 ;
      RECT  864000.0 820800.0 874200.0 807000.0 ;
      RECT  864000.0 820800.0 874200.0 834600.0 ;
      RECT  864000.0 848400.0 874200.0 834600.0 ;
      RECT  864000.0 848400.0 874200.0 862200.0 ;
      RECT  864000.0 876000.0 874200.0 862200.0 ;
      RECT  864000.0 876000.0 874200.0 889800.0 ;
      RECT  864000.0 903600.0 874200.0 889800.0 ;
      RECT  864000.0 903600.0 874200.0 917400.0 ;
      RECT  864000.0 931200.0 874200.0 917400.0 ;
      RECT  864000.0 931200.0 874200.0 945000.0 ;
      RECT  864000.0 958800.0 874200.0 945000.0 ;
      RECT  864000.0 958800.0 874200.0 972600.0 ;
      RECT  864000.0 986400.0 874200.0 972600.0 ;
      RECT  864000.0 986400.0 874200.0 1000200.0 ;
      RECT  864000.0 1014000.0 874200.0 1000200.0 ;
      RECT  864000.0 1014000.0 874200.0 1027800.0 ;
      RECT  864000.0 1041600.0 874200.0 1027800.0 ;
      RECT  864000.0 1041600.0 874200.0 1055400.0 ;
      RECT  864000.0 1069200.0 874200.0 1055400.0 ;
      RECT  864000.0 1069200.0 874200.0 1083000.0 ;
      RECT  864000.0 1096800.0 874200.0 1083000.0 ;
      RECT  864000.0 1096800.0 874200.0 1110600.0 ;
      RECT  864000.0 1124400.0 874200.0 1110600.0 ;
      RECT  864000.0 1124400.0 874200.0 1138200.0 ;
      RECT  864000.0 1152000.0 874200.0 1138200.0 ;
      RECT  864000.0 1152000.0 874200.0 1165800.0 ;
      RECT  864000.0 1179600.0 874200.0 1165800.0 ;
      RECT  864000.0 1179600.0 874200.0 1193400.0 ;
      RECT  864000.0 1207200.0 874200.0 1193400.0 ;
      RECT  864000.0 1207200.0 874200.0 1221000.0 ;
      RECT  864000.0 1234800.0 874200.0 1221000.0 ;
      RECT  864000.0 1234800.0 874200.0 1248600.0 ;
      RECT  864000.0 1262400.0 874200.0 1248600.0 ;
      RECT  864000.0 1262400.0 874200.0 1276200.0 ;
      RECT  864000.0 1290000.0 874200.0 1276200.0 ;
      RECT  864000.0 1290000.0 874200.0 1303800.0 ;
      RECT  864000.0 1317600.0 874200.0 1303800.0 ;
      RECT  864000.0 1317600.0 874200.0 1331400.0 ;
      RECT  864000.0 1345200.0 874200.0 1331400.0 ;
      RECT  864000.0 1345200.0 874200.0 1359000.0 ;
      RECT  864000.0 1372800.0 874200.0 1359000.0 ;
      RECT  864000.0 1372800.0 874200.0 1386600.0 ;
      RECT  864000.0 1400400.0 874200.0 1386600.0 ;
      RECT  864000.0 1400400.0 874200.0 1414200.0 ;
      RECT  864000.0 1428000.0 874200.0 1414200.0 ;
      RECT  864000.0 1428000.0 874200.0 1441800.0 ;
      RECT  864000.0 1455600.0 874200.0 1441800.0 ;
      RECT  864000.0 1455600.0 874200.0 1469400.0 ;
      RECT  864000.0 1483200.0 874200.0 1469400.0 ;
      RECT  864000.0 1483200.0 874200.0 1497000.0 ;
      RECT  864000.0 1510800.0 874200.0 1497000.0 ;
      RECT  864000.0 1510800.0 874200.0 1524600.0 ;
      RECT  864000.0 1538400.0 874200.0 1524600.0 ;
      RECT  864000.0 1538400.0 874200.0 1552200.0 ;
      RECT  864000.0 1566000.0 874200.0 1552200.0 ;
      RECT  864000.0 1566000.0 874200.0 1579800.0 ;
      RECT  864000.0 1593600.0 874200.0 1579800.0 ;
      RECT  864000.0 1593600.0 874200.0 1607400.0 ;
      RECT  864000.0 1621200.0 874200.0 1607400.0 ;
      RECT  864000.0 1621200.0 874200.0 1635000.0 ;
      RECT  864000.0 1648800.0 874200.0 1635000.0 ;
      RECT  864000.0 1648800.0 874200.0 1662600.0 ;
      RECT  864000.0 1676400.0 874200.0 1662600.0 ;
      RECT  864000.0 1676400.0 874200.0 1690200.0 ;
      RECT  864000.0 1704000.0 874200.0 1690200.0 ;
      RECT  864000.0 1704000.0 874200.0 1717800.0 ;
      RECT  864000.0 1731600.0 874200.0 1717800.0 ;
      RECT  864000.0 1731600.0 874200.0 1745400.0 ;
      RECT  864000.0 1759200.0 874200.0 1745400.0 ;
      RECT  864000.0 1759200.0 874200.0 1773000.0 ;
      RECT  864000.0 1786800.0 874200.0 1773000.0 ;
      RECT  864000.0 1786800.0 874200.0 1800600.0 ;
      RECT  864000.0 1814400.0 874200.0 1800600.0 ;
      RECT  864000.0 1814400.0 874200.0 1828200.0 ;
      RECT  864000.0 1842000.0 874200.0 1828200.0 ;
      RECT  864000.0 1842000.0 874200.0 1855800.0 ;
      RECT  864000.0 1869600.0 874200.0 1855800.0 ;
      RECT  864000.0 1869600.0 874200.0 1883400.0 ;
      RECT  864000.0 1897200.0 874200.0 1883400.0 ;
      RECT  864000.0 1897200.0 874200.0 1911000.0 ;
      RECT  864000.0 1924800.0 874200.0 1911000.0 ;
      RECT  864000.0 1924800.0 874200.0 1938600.0 ;
      RECT  864000.0 1952400.0 874200.0 1938600.0 ;
      RECT  864000.0 1952400.0 874200.0 1966200.0 ;
      RECT  864000.0 1980000.0 874200.0 1966200.0 ;
      RECT  864000.0 1980000.0 874200.0 1993800.0 ;
      RECT  864000.0 2007600.0 874200.0 1993800.0 ;
      RECT  864000.0 2007600.0 874200.0 2021400.0 ;
      RECT  864000.0 2035200.0 874200.0 2021400.0 ;
      RECT  864000.0 2035200.0 874200.0 2049000.0 ;
      RECT  864000.0 2062800.0 874200.0 2049000.0 ;
      RECT  864000.0 2062800.0 874200.0 2076600.0 ;
      RECT  864000.0 2090400.0 874200.0 2076600.0 ;
      RECT  864000.0 2090400.0 874200.0 2104200.0 ;
      RECT  864000.0 2118000.0 874200.0 2104200.0 ;
      RECT  864000.0 2118000.0 874200.0 2131800.0 ;
      RECT  864000.0 2145600.0 874200.0 2131800.0 ;
      RECT  874200.0 379200.0 884400.0 393000.0 ;
      RECT  874200.0 406800.0 884400.0 393000.0 ;
      RECT  874200.0 406800.0 884400.0 420600.0 ;
      RECT  874200.0 434400.0 884400.0 420600.0 ;
      RECT  874200.0 434400.0 884400.0 448200.0 ;
      RECT  874200.0 462000.0 884400.0 448200.0 ;
      RECT  874200.0 462000.0 884400.0 475800.0 ;
      RECT  874200.0 489600.0 884400.0 475800.0 ;
      RECT  874200.0 489600.0 884400.0 503400.0 ;
      RECT  874200.0 517200.0 884400.0 503400.0 ;
      RECT  874200.0 517200.0 884400.0 531000.0 ;
      RECT  874200.0 544800.0 884400.0 531000.0 ;
      RECT  874200.0 544800.0 884400.0 558600.0 ;
      RECT  874200.0 572400.0 884400.0 558600.0 ;
      RECT  874200.0 572400.0 884400.0 586200.0 ;
      RECT  874200.0 600000.0 884400.0 586200.0 ;
      RECT  874200.0 600000.0 884400.0 613800.0 ;
      RECT  874200.0 627600.0 884400.0 613800.0 ;
      RECT  874200.0 627600.0 884400.0 641400.0 ;
      RECT  874200.0 655200.0 884400.0 641400.0 ;
      RECT  874200.0 655200.0 884400.0 669000.0 ;
      RECT  874200.0 682800.0 884400.0 669000.0 ;
      RECT  874200.0 682800.0 884400.0 696600.0 ;
      RECT  874200.0 710400.0 884400.0 696600.0 ;
      RECT  874200.0 710400.0 884400.0 724200.0 ;
      RECT  874200.0 738000.0 884400.0 724200.0 ;
      RECT  874200.0 738000.0 884400.0 751800.0 ;
      RECT  874200.0 765600.0 884400.0 751800.0 ;
      RECT  874200.0 765600.0 884400.0 779400.0 ;
      RECT  874200.0 793200.0 884400.0 779400.0 ;
      RECT  874200.0 793200.0 884400.0 807000.0 ;
      RECT  874200.0 820800.0 884400.0 807000.0 ;
      RECT  874200.0 820800.0 884400.0 834600.0 ;
      RECT  874200.0 848400.0 884400.0 834600.0 ;
      RECT  874200.0 848400.0 884400.0 862200.0 ;
      RECT  874200.0 876000.0 884400.0 862200.0 ;
      RECT  874200.0 876000.0 884400.0 889800.0 ;
      RECT  874200.0 903600.0 884400.0 889800.0 ;
      RECT  874200.0 903600.0 884400.0 917400.0 ;
      RECT  874200.0 931200.0 884400.0 917400.0 ;
      RECT  874200.0 931200.0 884400.0 945000.0 ;
      RECT  874200.0 958800.0 884400.0 945000.0 ;
      RECT  874200.0 958800.0 884400.0 972600.0 ;
      RECT  874200.0 986400.0 884400.0 972600.0 ;
      RECT  874200.0 986400.0 884400.0 1000200.0 ;
      RECT  874200.0 1014000.0 884400.0 1000200.0 ;
      RECT  874200.0 1014000.0 884400.0 1027800.0 ;
      RECT  874200.0 1041600.0 884400.0 1027800.0 ;
      RECT  874200.0 1041600.0 884400.0 1055400.0 ;
      RECT  874200.0 1069200.0 884400.0 1055400.0 ;
      RECT  874200.0 1069200.0 884400.0 1083000.0 ;
      RECT  874200.0 1096800.0 884400.0 1083000.0 ;
      RECT  874200.0 1096800.0 884400.0 1110600.0 ;
      RECT  874200.0 1124400.0 884400.0 1110600.0 ;
      RECT  874200.0 1124400.0 884400.0 1138200.0 ;
      RECT  874200.0 1152000.0 884400.0 1138200.0 ;
      RECT  874200.0 1152000.0 884400.0 1165800.0 ;
      RECT  874200.0 1179600.0 884400.0 1165800.0 ;
      RECT  874200.0 1179600.0 884400.0 1193400.0 ;
      RECT  874200.0 1207200.0 884400.0 1193400.0 ;
      RECT  874200.0 1207200.0 884400.0 1221000.0 ;
      RECT  874200.0 1234800.0 884400.0 1221000.0 ;
      RECT  874200.0 1234800.0 884400.0 1248600.0 ;
      RECT  874200.0 1262400.0 884400.0 1248600.0 ;
      RECT  874200.0 1262400.0 884400.0 1276200.0 ;
      RECT  874200.0 1290000.0 884400.0 1276200.0 ;
      RECT  874200.0 1290000.0 884400.0 1303800.0 ;
      RECT  874200.0 1317600.0 884400.0 1303800.0 ;
      RECT  874200.0 1317600.0 884400.0 1331400.0 ;
      RECT  874200.0 1345200.0 884400.0 1331400.0 ;
      RECT  874200.0 1345200.0 884400.0 1359000.0 ;
      RECT  874200.0 1372800.0 884400.0 1359000.0 ;
      RECT  874200.0 1372800.0 884400.0 1386600.0 ;
      RECT  874200.0 1400400.0 884400.0 1386600.0 ;
      RECT  874200.0 1400400.0 884400.0 1414200.0 ;
      RECT  874200.0 1428000.0 884400.0 1414200.0 ;
      RECT  874200.0 1428000.0 884400.0 1441800.0 ;
      RECT  874200.0 1455600.0 884400.0 1441800.0 ;
      RECT  874200.0 1455600.0 884400.0 1469400.0 ;
      RECT  874200.0 1483200.0 884400.0 1469400.0 ;
      RECT  874200.0 1483200.0 884400.0 1497000.0 ;
      RECT  874200.0 1510800.0 884400.0 1497000.0 ;
      RECT  874200.0 1510800.0 884400.0 1524600.0 ;
      RECT  874200.0 1538400.0 884400.0 1524600.0 ;
      RECT  874200.0 1538400.0 884400.0 1552200.0 ;
      RECT  874200.0 1566000.0 884400.0 1552200.0 ;
      RECT  874200.0 1566000.0 884400.0 1579800.0 ;
      RECT  874200.0 1593600.0 884400.0 1579800.0 ;
      RECT  874200.0 1593600.0 884400.0 1607400.0 ;
      RECT  874200.0 1621200.0 884400.0 1607400.0 ;
      RECT  874200.0 1621200.0 884400.0 1635000.0 ;
      RECT  874200.0 1648800.0 884400.0 1635000.0 ;
      RECT  874200.0 1648800.0 884400.0 1662600.0 ;
      RECT  874200.0 1676400.0 884400.0 1662600.0 ;
      RECT  874200.0 1676400.0 884400.0 1690200.0 ;
      RECT  874200.0 1704000.0 884400.0 1690200.0 ;
      RECT  874200.0 1704000.0 884400.0 1717800.0 ;
      RECT  874200.0 1731600.0 884400.0 1717800.0 ;
      RECT  874200.0 1731600.0 884400.0 1745400.0 ;
      RECT  874200.0 1759200.0 884400.0 1745400.0 ;
      RECT  874200.0 1759200.0 884400.0 1773000.0 ;
      RECT  874200.0 1786800.0 884400.0 1773000.0 ;
      RECT  874200.0 1786800.0 884400.0 1800600.0 ;
      RECT  874200.0 1814400.0 884400.0 1800600.0 ;
      RECT  874200.0 1814400.0 884400.0 1828200.0 ;
      RECT  874200.0 1842000.0 884400.0 1828200.0 ;
      RECT  874200.0 1842000.0 884400.0 1855800.0 ;
      RECT  874200.0 1869600.0 884400.0 1855800.0 ;
      RECT  874200.0 1869600.0 884400.0 1883400.0 ;
      RECT  874200.0 1897200.0 884400.0 1883400.0 ;
      RECT  874200.0 1897200.0 884400.0 1911000.0 ;
      RECT  874200.0 1924800.0 884400.0 1911000.0 ;
      RECT  874200.0 1924800.0 884400.0 1938600.0 ;
      RECT  874200.0 1952400.0 884400.0 1938600.0 ;
      RECT  874200.0 1952400.0 884400.0 1966200.0 ;
      RECT  874200.0 1980000.0 884400.0 1966200.0 ;
      RECT  874200.0 1980000.0 884400.0 1993800.0 ;
      RECT  874200.0 2007600.0 884400.0 1993800.0 ;
      RECT  874200.0 2007600.0 884400.0 2021400.0 ;
      RECT  874200.0 2035200.0 884400.0 2021400.0 ;
      RECT  874200.0 2035200.0 884400.0 2049000.0 ;
      RECT  874200.0 2062800.0 884400.0 2049000.0 ;
      RECT  874200.0 2062800.0 884400.0 2076600.0 ;
      RECT  874200.0 2090400.0 884400.0 2076600.0 ;
      RECT  874200.0 2090400.0 884400.0 2104200.0 ;
      RECT  874200.0 2118000.0 884400.0 2104200.0 ;
      RECT  874200.0 2118000.0 884400.0 2131800.0 ;
      RECT  874200.0 2145600.0 884400.0 2131800.0 ;
      RECT  884400.0 379200.0 894600.0 393000.0 ;
      RECT  884400.0 406800.0 894600.0 393000.0 ;
      RECT  884400.0 406800.0 894600.0 420600.0 ;
      RECT  884400.0 434400.0 894600.0 420600.0 ;
      RECT  884400.0 434400.0 894600.0 448200.0 ;
      RECT  884400.0 462000.0 894600.0 448200.0 ;
      RECT  884400.0 462000.0 894600.0 475800.0 ;
      RECT  884400.0 489600.0 894600.0 475800.0 ;
      RECT  884400.0 489600.0 894600.0 503400.0 ;
      RECT  884400.0 517200.0 894600.0 503400.0 ;
      RECT  884400.0 517200.0 894600.0 531000.0 ;
      RECT  884400.0 544800.0 894600.0 531000.0 ;
      RECT  884400.0 544800.0 894600.0 558600.0 ;
      RECT  884400.0 572400.0 894600.0 558600.0 ;
      RECT  884400.0 572400.0 894600.0 586200.0 ;
      RECT  884400.0 600000.0 894600.0 586200.0 ;
      RECT  884400.0 600000.0 894600.0 613800.0 ;
      RECT  884400.0 627600.0 894600.0 613800.0 ;
      RECT  884400.0 627600.0 894600.0 641400.0 ;
      RECT  884400.0 655200.0 894600.0 641400.0 ;
      RECT  884400.0 655200.0 894600.0 669000.0 ;
      RECT  884400.0 682800.0 894600.0 669000.0 ;
      RECT  884400.0 682800.0 894600.0 696600.0 ;
      RECT  884400.0 710400.0 894600.0 696600.0 ;
      RECT  884400.0 710400.0 894600.0 724200.0 ;
      RECT  884400.0 738000.0 894600.0 724200.0 ;
      RECT  884400.0 738000.0 894600.0 751800.0 ;
      RECT  884400.0 765600.0 894600.0 751800.0 ;
      RECT  884400.0 765600.0 894600.0 779400.0 ;
      RECT  884400.0 793200.0 894600.0 779400.0 ;
      RECT  884400.0 793200.0 894600.0 807000.0 ;
      RECT  884400.0 820800.0 894600.0 807000.0 ;
      RECT  884400.0 820800.0 894600.0 834600.0 ;
      RECT  884400.0 848400.0 894600.0 834600.0 ;
      RECT  884400.0 848400.0 894600.0 862200.0 ;
      RECT  884400.0 876000.0 894600.0 862200.0 ;
      RECT  884400.0 876000.0 894600.0 889800.0 ;
      RECT  884400.0 903600.0 894600.0 889800.0 ;
      RECT  884400.0 903600.0 894600.0 917400.0 ;
      RECT  884400.0 931200.0 894600.0 917400.0 ;
      RECT  884400.0 931200.0 894600.0 945000.0 ;
      RECT  884400.0 958800.0 894600.0 945000.0 ;
      RECT  884400.0 958800.0 894600.0 972600.0 ;
      RECT  884400.0 986400.0 894600.0 972600.0 ;
      RECT  884400.0 986400.0 894600.0 1000200.0 ;
      RECT  884400.0 1014000.0 894600.0 1000200.0 ;
      RECT  884400.0 1014000.0 894600.0 1027800.0 ;
      RECT  884400.0 1041600.0 894600.0 1027800.0 ;
      RECT  884400.0 1041600.0 894600.0 1055400.0 ;
      RECT  884400.0 1069200.0 894600.0 1055400.0 ;
      RECT  884400.0 1069200.0 894600.0 1083000.0 ;
      RECT  884400.0 1096800.0 894600.0 1083000.0 ;
      RECT  884400.0 1096800.0 894600.0 1110600.0 ;
      RECT  884400.0 1124400.0 894600.0 1110600.0 ;
      RECT  884400.0 1124400.0 894600.0 1138200.0 ;
      RECT  884400.0 1152000.0 894600.0 1138200.0 ;
      RECT  884400.0 1152000.0 894600.0 1165800.0 ;
      RECT  884400.0 1179600.0 894600.0 1165800.0 ;
      RECT  884400.0 1179600.0 894600.0 1193400.0 ;
      RECT  884400.0 1207200.0 894600.0 1193400.0 ;
      RECT  884400.0 1207200.0 894600.0 1221000.0 ;
      RECT  884400.0 1234800.0 894600.0 1221000.0 ;
      RECT  884400.0 1234800.0 894600.0 1248600.0 ;
      RECT  884400.0 1262400.0 894600.0 1248600.0 ;
      RECT  884400.0 1262400.0 894600.0 1276200.0 ;
      RECT  884400.0 1290000.0 894600.0 1276200.0 ;
      RECT  884400.0 1290000.0 894600.0 1303800.0 ;
      RECT  884400.0 1317600.0 894600.0 1303800.0 ;
      RECT  884400.0 1317600.0 894600.0 1331400.0 ;
      RECT  884400.0 1345200.0 894600.0 1331400.0 ;
      RECT  884400.0 1345200.0 894600.0 1359000.0 ;
      RECT  884400.0 1372800.0 894600.0 1359000.0 ;
      RECT  884400.0 1372800.0 894600.0 1386600.0 ;
      RECT  884400.0 1400400.0 894600.0 1386600.0 ;
      RECT  884400.0 1400400.0 894600.0 1414200.0 ;
      RECT  884400.0 1428000.0 894600.0 1414200.0 ;
      RECT  884400.0 1428000.0 894600.0 1441800.0 ;
      RECT  884400.0 1455600.0 894600.0 1441800.0 ;
      RECT  884400.0 1455600.0 894600.0 1469400.0 ;
      RECT  884400.0 1483200.0 894600.0 1469400.0 ;
      RECT  884400.0 1483200.0 894600.0 1497000.0 ;
      RECT  884400.0 1510800.0 894600.0 1497000.0 ;
      RECT  884400.0 1510800.0 894600.0 1524600.0 ;
      RECT  884400.0 1538400.0 894600.0 1524600.0 ;
      RECT  884400.0 1538400.0 894600.0 1552200.0 ;
      RECT  884400.0 1566000.0 894600.0 1552200.0 ;
      RECT  884400.0 1566000.0 894600.0 1579800.0 ;
      RECT  884400.0 1593600.0 894600.0 1579800.0 ;
      RECT  884400.0 1593600.0 894600.0 1607400.0 ;
      RECT  884400.0 1621200.0 894600.0 1607400.0 ;
      RECT  884400.0 1621200.0 894600.0 1635000.0 ;
      RECT  884400.0 1648800.0 894600.0 1635000.0 ;
      RECT  884400.0 1648800.0 894600.0 1662600.0 ;
      RECT  884400.0 1676400.0 894600.0 1662600.0 ;
      RECT  884400.0 1676400.0 894600.0 1690200.0 ;
      RECT  884400.0 1704000.0 894600.0 1690200.0 ;
      RECT  884400.0 1704000.0 894600.0 1717800.0 ;
      RECT  884400.0 1731600.0 894600.0 1717800.0 ;
      RECT  884400.0 1731600.0 894600.0 1745400.0 ;
      RECT  884400.0 1759200.0 894600.0 1745400.0 ;
      RECT  884400.0 1759200.0 894600.0 1773000.0 ;
      RECT  884400.0 1786800.0 894600.0 1773000.0 ;
      RECT  884400.0 1786800.0 894600.0 1800600.0 ;
      RECT  884400.0 1814400.0 894600.0 1800600.0 ;
      RECT  884400.0 1814400.0 894600.0 1828200.0 ;
      RECT  884400.0 1842000.0 894600.0 1828200.0 ;
      RECT  884400.0 1842000.0 894600.0 1855800.0 ;
      RECT  884400.0 1869600.0 894600.0 1855800.0 ;
      RECT  884400.0 1869600.0 894600.0 1883400.0 ;
      RECT  884400.0 1897200.0 894600.0 1883400.0 ;
      RECT  884400.0 1897200.0 894600.0 1911000.0 ;
      RECT  884400.0 1924800.0 894600.0 1911000.0 ;
      RECT  884400.0 1924800.0 894600.0 1938600.0 ;
      RECT  884400.0 1952400.0 894600.0 1938600.0 ;
      RECT  884400.0 1952400.0 894600.0 1966200.0 ;
      RECT  884400.0 1980000.0 894600.0 1966200.0 ;
      RECT  884400.0 1980000.0 894600.0 1993800.0 ;
      RECT  884400.0 2007600.0 894600.0 1993800.0 ;
      RECT  884400.0 2007600.0 894600.0 2021400.0 ;
      RECT  884400.0 2035200.0 894600.0 2021400.0 ;
      RECT  884400.0 2035200.0 894600.0 2049000.0 ;
      RECT  884400.0 2062800.0 894600.0 2049000.0 ;
      RECT  884400.0 2062800.0 894600.0 2076600.0 ;
      RECT  884400.0 2090400.0 894600.0 2076600.0 ;
      RECT  884400.0 2090400.0 894600.0 2104200.0 ;
      RECT  884400.0 2118000.0 894600.0 2104200.0 ;
      RECT  884400.0 2118000.0 894600.0 2131800.0 ;
      RECT  884400.0 2145600.0 894600.0 2131800.0 ;
      RECT  894600.0 379200.0 904800.0 393000.0 ;
      RECT  894600.0 406800.0 904800.0 393000.0 ;
      RECT  894600.0 406800.0 904800.0 420600.0 ;
      RECT  894600.0 434400.0 904800.0 420600.0 ;
      RECT  894600.0 434400.0 904800.0 448200.0 ;
      RECT  894600.0 462000.0 904800.0 448200.0 ;
      RECT  894600.0 462000.0 904800.0 475800.0 ;
      RECT  894600.0 489600.0 904800.0 475800.0 ;
      RECT  894600.0 489600.0 904800.0 503400.0 ;
      RECT  894600.0 517200.0 904800.0 503400.0 ;
      RECT  894600.0 517200.0 904800.0 531000.0 ;
      RECT  894600.0 544800.0 904800.0 531000.0 ;
      RECT  894600.0 544800.0 904800.0 558600.0 ;
      RECT  894600.0 572400.0 904800.0 558600.0 ;
      RECT  894600.0 572400.0 904800.0 586200.0 ;
      RECT  894600.0 600000.0 904800.0 586200.0 ;
      RECT  894600.0 600000.0 904800.0 613800.0 ;
      RECT  894600.0 627600.0 904800.0 613800.0 ;
      RECT  894600.0 627600.0 904800.0 641400.0 ;
      RECT  894600.0 655200.0 904800.0 641400.0 ;
      RECT  894600.0 655200.0 904800.0 669000.0 ;
      RECT  894600.0 682800.0 904800.0 669000.0 ;
      RECT  894600.0 682800.0 904800.0 696600.0 ;
      RECT  894600.0 710400.0 904800.0 696600.0 ;
      RECT  894600.0 710400.0 904800.0 724200.0 ;
      RECT  894600.0 738000.0 904800.0 724200.0 ;
      RECT  894600.0 738000.0 904800.0 751800.0 ;
      RECT  894600.0 765600.0 904800.0 751800.0 ;
      RECT  894600.0 765600.0 904800.0 779400.0 ;
      RECT  894600.0 793200.0 904800.0 779400.0 ;
      RECT  894600.0 793200.0 904800.0 807000.0 ;
      RECT  894600.0 820800.0 904800.0 807000.0 ;
      RECT  894600.0 820800.0 904800.0 834600.0 ;
      RECT  894600.0 848400.0 904800.0 834600.0 ;
      RECT  894600.0 848400.0 904800.0 862200.0 ;
      RECT  894600.0 876000.0 904800.0 862200.0 ;
      RECT  894600.0 876000.0 904800.0 889800.0 ;
      RECT  894600.0 903600.0 904800.0 889800.0 ;
      RECT  894600.0 903600.0 904800.0 917400.0 ;
      RECT  894600.0 931200.0 904800.0 917400.0 ;
      RECT  894600.0 931200.0 904800.0 945000.0 ;
      RECT  894600.0 958800.0 904800.0 945000.0 ;
      RECT  894600.0 958800.0 904800.0 972600.0 ;
      RECT  894600.0 986400.0 904800.0 972600.0 ;
      RECT  894600.0 986400.0 904800.0 1000200.0 ;
      RECT  894600.0 1014000.0 904800.0 1000200.0 ;
      RECT  894600.0 1014000.0 904800.0 1027800.0 ;
      RECT  894600.0 1041600.0 904800.0 1027800.0 ;
      RECT  894600.0 1041600.0 904800.0 1055400.0 ;
      RECT  894600.0 1069200.0 904800.0 1055400.0 ;
      RECT  894600.0 1069200.0 904800.0 1083000.0 ;
      RECT  894600.0 1096800.0 904800.0 1083000.0 ;
      RECT  894600.0 1096800.0 904800.0 1110600.0 ;
      RECT  894600.0 1124400.0 904800.0 1110600.0 ;
      RECT  894600.0 1124400.0 904800.0 1138200.0 ;
      RECT  894600.0 1152000.0 904800.0 1138200.0 ;
      RECT  894600.0 1152000.0 904800.0 1165800.0 ;
      RECT  894600.0 1179600.0 904800.0 1165800.0 ;
      RECT  894600.0 1179600.0 904800.0 1193400.0 ;
      RECT  894600.0 1207200.0 904800.0 1193400.0 ;
      RECT  894600.0 1207200.0 904800.0 1221000.0 ;
      RECT  894600.0 1234800.0 904800.0 1221000.0 ;
      RECT  894600.0 1234800.0 904800.0 1248600.0 ;
      RECT  894600.0 1262400.0 904800.0 1248600.0 ;
      RECT  894600.0 1262400.0 904800.0 1276200.0 ;
      RECT  894600.0 1290000.0 904800.0 1276200.0 ;
      RECT  894600.0 1290000.0 904800.0 1303800.0 ;
      RECT  894600.0 1317600.0 904800.0 1303800.0 ;
      RECT  894600.0 1317600.0 904800.0 1331400.0 ;
      RECT  894600.0 1345200.0 904800.0 1331400.0 ;
      RECT  894600.0 1345200.0 904800.0 1359000.0 ;
      RECT  894600.0 1372800.0 904800.0 1359000.0 ;
      RECT  894600.0 1372800.0 904800.0 1386600.0 ;
      RECT  894600.0 1400400.0 904800.0 1386600.0 ;
      RECT  894600.0 1400400.0 904800.0 1414200.0 ;
      RECT  894600.0 1428000.0 904800.0 1414200.0 ;
      RECT  894600.0 1428000.0 904800.0 1441800.0 ;
      RECT  894600.0 1455600.0 904800.0 1441800.0 ;
      RECT  894600.0 1455600.0 904800.0 1469400.0 ;
      RECT  894600.0 1483200.0 904800.0 1469400.0 ;
      RECT  894600.0 1483200.0 904800.0 1497000.0 ;
      RECT  894600.0 1510800.0 904800.0 1497000.0 ;
      RECT  894600.0 1510800.0 904800.0 1524600.0 ;
      RECT  894600.0 1538400.0 904800.0 1524600.0 ;
      RECT  894600.0 1538400.0 904800.0 1552200.0 ;
      RECT  894600.0 1566000.0 904800.0 1552200.0 ;
      RECT  894600.0 1566000.0 904800.0 1579800.0 ;
      RECT  894600.0 1593600.0 904800.0 1579800.0 ;
      RECT  894600.0 1593600.0 904800.0 1607400.0 ;
      RECT  894600.0 1621200.0 904800.0 1607400.0 ;
      RECT  894600.0 1621200.0 904800.0 1635000.0 ;
      RECT  894600.0 1648800.0 904800.0 1635000.0 ;
      RECT  894600.0 1648800.0 904800.0 1662600.0 ;
      RECT  894600.0 1676400.0 904800.0 1662600.0 ;
      RECT  894600.0 1676400.0 904800.0 1690200.0 ;
      RECT  894600.0 1704000.0 904800.0 1690200.0 ;
      RECT  894600.0 1704000.0 904800.0 1717800.0 ;
      RECT  894600.0 1731600.0 904800.0 1717800.0 ;
      RECT  894600.0 1731600.0 904800.0 1745400.0 ;
      RECT  894600.0 1759200.0 904800.0 1745400.0 ;
      RECT  894600.0 1759200.0 904800.0 1773000.0 ;
      RECT  894600.0 1786800.0 904800.0 1773000.0 ;
      RECT  894600.0 1786800.0 904800.0 1800600.0 ;
      RECT  894600.0 1814400.0 904800.0 1800600.0 ;
      RECT  894600.0 1814400.0 904800.0 1828200.0 ;
      RECT  894600.0 1842000.0 904800.0 1828200.0 ;
      RECT  894600.0 1842000.0 904800.0 1855800.0 ;
      RECT  894600.0 1869600.0 904800.0 1855800.0 ;
      RECT  894600.0 1869600.0 904800.0 1883400.0 ;
      RECT  894600.0 1897200.0 904800.0 1883400.0 ;
      RECT  894600.0 1897200.0 904800.0 1911000.0 ;
      RECT  894600.0 1924800.0 904800.0 1911000.0 ;
      RECT  894600.0 1924800.0 904800.0 1938600.0 ;
      RECT  894600.0 1952400.0 904800.0 1938600.0 ;
      RECT  894600.0 1952400.0 904800.0 1966200.0 ;
      RECT  894600.0 1980000.0 904800.0 1966200.0 ;
      RECT  894600.0 1980000.0 904800.0 1993800.0 ;
      RECT  894600.0 2007600.0 904800.0 1993800.0 ;
      RECT  894600.0 2007600.0 904800.0 2021400.0 ;
      RECT  894600.0 2035200.0 904800.0 2021400.0 ;
      RECT  894600.0 2035200.0 904800.0 2049000.0 ;
      RECT  894600.0 2062800.0 904800.0 2049000.0 ;
      RECT  894600.0 2062800.0 904800.0 2076600.0 ;
      RECT  894600.0 2090400.0 904800.0 2076600.0 ;
      RECT  894600.0 2090400.0 904800.0 2104200.0 ;
      RECT  894600.0 2118000.0 904800.0 2104200.0 ;
      RECT  894600.0 2118000.0 904800.0 2131800.0 ;
      RECT  894600.0 2145600.0 904800.0 2131800.0 ;
      RECT  904800.0 379200.0 915000.0 393000.0 ;
      RECT  904800.0 406800.0 915000.0 393000.0 ;
      RECT  904800.0 406800.0 915000.0 420600.0 ;
      RECT  904800.0 434400.0 915000.0 420600.0 ;
      RECT  904800.0 434400.0 915000.0 448200.0 ;
      RECT  904800.0 462000.0 915000.0 448200.0 ;
      RECT  904800.0 462000.0 915000.0 475800.0 ;
      RECT  904800.0 489600.0 915000.0 475800.0 ;
      RECT  904800.0 489600.0 915000.0 503400.0 ;
      RECT  904800.0 517200.0 915000.0 503400.0 ;
      RECT  904800.0 517200.0 915000.0 531000.0 ;
      RECT  904800.0 544800.0 915000.0 531000.0 ;
      RECT  904800.0 544800.0 915000.0 558600.0 ;
      RECT  904800.0 572400.0 915000.0 558600.0 ;
      RECT  904800.0 572400.0 915000.0 586200.0 ;
      RECT  904800.0 600000.0 915000.0 586200.0 ;
      RECT  904800.0 600000.0 915000.0 613800.0 ;
      RECT  904800.0 627600.0 915000.0 613800.0 ;
      RECT  904800.0 627600.0 915000.0 641400.0 ;
      RECT  904800.0 655200.0 915000.0 641400.0 ;
      RECT  904800.0 655200.0 915000.0 669000.0 ;
      RECT  904800.0 682800.0 915000.0 669000.0 ;
      RECT  904800.0 682800.0 915000.0 696600.0 ;
      RECT  904800.0 710400.0 915000.0 696600.0 ;
      RECT  904800.0 710400.0 915000.0 724200.0 ;
      RECT  904800.0 738000.0 915000.0 724200.0 ;
      RECT  904800.0 738000.0 915000.0 751800.0 ;
      RECT  904800.0 765600.0 915000.0 751800.0 ;
      RECT  904800.0 765600.0 915000.0 779400.0 ;
      RECT  904800.0 793200.0 915000.0 779400.0 ;
      RECT  904800.0 793200.0 915000.0 807000.0 ;
      RECT  904800.0 820800.0 915000.0 807000.0 ;
      RECT  904800.0 820800.0 915000.0 834600.0 ;
      RECT  904800.0 848400.0 915000.0 834600.0 ;
      RECT  904800.0 848400.0 915000.0 862200.0 ;
      RECT  904800.0 876000.0 915000.0 862200.0 ;
      RECT  904800.0 876000.0 915000.0 889800.0 ;
      RECT  904800.0 903600.0 915000.0 889800.0 ;
      RECT  904800.0 903600.0 915000.0 917400.0 ;
      RECT  904800.0 931200.0 915000.0 917400.0 ;
      RECT  904800.0 931200.0 915000.0 945000.0 ;
      RECT  904800.0 958800.0 915000.0 945000.0 ;
      RECT  904800.0 958800.0 915000.0 972600.0 ;
      RECT  904800.0 986400.0 915000.0 972600.0 ;
      RECT  904800.0 986400.0 915000.0 1000200.0 ;
      RECT  904800.0 1014000.0 915000.0 1000200.0 ;
      RECT  904800.0 1014000.0 915000.0 1027800.0 ;
      RECT  904800.0 1041600.0 915000.0 1027800.0 ;
      RECT  904800.0 1041600.0 915000.0 1055400.0 ;
      RECT  904800.0 1069200.0 915000.0 1055400.0 ;
      RECT  904800.0 1069200.0 915000.0 1083000.0 ;
      RECT  904800.0 1096800.0 915000.0 1083000.0 ;
      RECT  904800.0 1096800.0 915000.0 1110600.0 ;
      RECT  904800.0 1124400.0 915000.0 1110600.0 ;
      RECT  904800.0 1124400.0 915000.0 1138200.0 ;
      RECT  904800.0 1152000.0 915000.0 1138200.0 ;
      RECT  904800.0 1152000.0 915000.0 1165800.0 ;
      RECT  904800.0 1179600.0 915000.0 1165800.0 ;
      RECT  904800.0 1179600.0 915000.0 1193400.0 ;
      RECT  904800.0 1207200.0 915000.0 1193400.0 ;
      RECT  904800.0 1207200.0 915000.0 1221000.0 ;
      RECT  904800.0 1234800.0 915000.0 1221000.0 ;
      RECT  904800.0 1234800.0 915000.0 1248600.0 ;
      RECT  904800.0 1262400.0 915000.0 1248600.0 ;
      RECT  904800.0 1262400.0 915000.0 1276200.0 ;
      RECT  904800.0 1290000.0 915000.0 1276200.0 ;
      RECT  904800.0 1290000.0 915000.0 1303800.0 ;
      RECT  904800.0 1317600.0 915000.0 1303800.0 ;
      RECT  904800.0 1317600.0 915000.0 1331400.0 ;
      RECT  904800.0 1345200.0 915000.0 1331400.0 ;
      RECT  904800.0 1345200.0 915000.0 1359000.0 ;
      RECT  904800.0 1372800.0 915000.0 1359000.0 ;
      RECT  904800.0 1372800.0 915000.0 1386600.0 ;
      RECT  904800.0 1400400.0 915000.0 1386600.0 ;
      RECT  904800.0 1400400.0 915000.0 1414200.0 ;
      RECT  904800.0 1428000.0 915000.0 1414200.0 ;
      RECT  904800.0 1428000.0 915000.0 1441800.0 ;
      RECT  904800.0 1455600.0 915000.0 1441800.0 ;
      RECT  904800.0 1455600.0 915000.0 1469400.0 ;
      RECT  904800.0 1483200.0 915000.0 1469400.0 ;
      RECT  904800.0 1483200.0 915000.0 1497000.0 ;
      RECT  904800.0 1510800.0 915000.0 1497000.0 ;
      RECT  904800.0 1510800.0 915000.0 1524600.0 ;
      RECT  904800.0 1538400.0 915000.0 1524600.0 ;
      RECT  904800.0 1538400.0 915000.0 1552200.0 ;
      RECT  904800.0 1566000.0 915000.0 1552200.0 ;
      RECT  904800.0 1566000.0 915000.0 1579800.0 ;
      RECT  904800.0 1593600.0 915000.0 1579800.0 ;
      RECT  904800.0 1593600.0 915000.0 1607400.0 ;
      RECT  904800.0 1621200.0 915000.0 1607400.0 ;
      RECT  904800.0 1621200.0 915000.0 1635000.0 ;
      RECT  904800.0 1648800.0 915000.0 1635000.0 ;
      RECT  904800.0 1648800.0 915000.0 1662600.0 ;
      RECT  904800.0 1676400.0 915000.0 1662600.0 ;
      RECT  904800.0 1676400.0 915000.0 1690200.0 ;
      RECT  904800.0 1704000.0 915000.0 1690200.0 ;
      RECT  904800.0 1704000.0 915000.0 1717800.0 ;
      RECT  904800.0 1731600.0 915000.0 1717800.0 ;
      RECT  904800.0 1731600.0 915000.0 1745400.0 ;
      RECT  904800.0 1759200.0 915000.0 1745400.0 ;
      RECT  904800.0 1759200.0 915000.0 1773000.0 ;
      RECT  904800.0 1786800.0 915000.0 1773000.0 ;
      RECT  904800.0 1786800.0 915000.0 1800600.0 ;
      RECT  904800.0 1814400.0 915000.0 1800600.0 ;
      RECT  904800.0 1814400.0 915000.0 1828200.0 ;
      RECT  904800.0 1842000.0 915000.0 1828200.0 ;
      RECT  904800.0 1842000.0 915000.0 1855800.0 ;
      RECT  904800.0 1869600.0 915000.0 1855800.0 ;
      RECT  904800.0 1869600.0 915000.0 1883400.0 ;
      RECT  904800.0 1897200.0 915000.0 1883400.0 ;
      RECT  904800.0 1897200.0 915000.0 1911000.0 ;
      RECT  904800.0 1924800.0 915000.0 1911000.0 ;
      RECT  904800.0 1924800.0 915000.0 1938600.0 ;
      RECT  904800.0 1952400.0 915000.0 1938600.0 ;
      RECT  904800.0 1952400.0 915000.0 1966200.0 ;
      RECT  904800.0 1980000.0 915000.0 1966200.0 ;
      RECT  904800.0 1980000.0 915000.0 1993800.0 ;
      RECT  904800.0 2007600.0 915000.0 1993800.0 ;
      RECT  904800.0 2007600.0 915000.0 2021400.0 ;
      RECT  904800.0 2035200.0 915000.0 2021400.0 ;
      RECT  904800.0 2035200.0 915000.0 2049000.0 ;
      RECT  904800.0 2062800.0 915000.0 2049000.0 ;
      RECT  904800.0 2062800.0 915000.0 2076600.0 ;
      RECT  904800.0 2090400.0 915000.0 2076600.0 ;
      RECT  904800.0 2090400.0 915000.0 2104200.0 ;
      RECT  904800.0 2118000.0 915000.0 2104200.0 ;
      RECT  904800.0 2118000.0 915000.0 2131800.0 ;
      RECT  904800.0 2145600.0 915000.0 2131800.0 ;
      RECT  915000.0 379200.0 925200.0 393000.0 ;
      RECT  915000.0 406800.0 925200.0 393000.0 ;
      RECT  915000.0 406800.0 925200.0 420600.0 ;
      RECT  915000.0 434400.0 925200.0 420600.0 ;
      RECT  915000.0 434400.0 925200.0 448200.0 ;
      RECT  915000.0 462000.0 925200.0 448200.0 ;
      RECT  915000.0 462000.0 925200.0 475800.0 ;
      RECT  915000.0 489600.0 925200.0 475800.0 ;
      RECT  915000.0 489600.0 925200.0 503400.0 ;
      RECT  915000.0 517200.0 925200.0 503400.0 ;
      RECT  915000.0 517200.0 925200.0 531000.0 ;
      RECT  915000.0 544800.0 925200.0 531000.0 ;
      RECT  915000.0 544800.0 925200.0 558600.0 ;
      RECT  915000.0 572400.0 925200.0 558600.0 ;
      RECT  915000.0 572400.0 925200.0 586200.0 ;
      RECT  915000.0 600000.0 925200.0 586200.0 ;
      RECT  915000.0 600000.0 925200.0 613800.0 ;
      RECT  915000.0 627600.0 925200.0 613800.0 ;
      RECT  915000.0 627600.0 925200.0 641400.0 ;
      RECT  915000.0 655200.0 925200.0 641400.0 ;
      RECT  915000.0 655200.0 925200.0 669000.0 ;
      RECT  915000.0 682800.0 925200.0 669000.0 ;
      RECT  915000.0 682800.0 925200.0 696600.0 ;
      RECT  915000.0 710400.0 925200.0 696600.0 ;
      RECT  915000.0 710400.0 925200.0 724200.0 ;
      RECT  915000.0 738000.0 925200.0 724200.0 ;
      RECT  915000.0 738000.0 925200.0 751800.0 ;
      RECT  915000.0 765600.0 925200.0 751800.0 ;
      RECT  915000.0 765600.0 925200.0 779400.0 ;
      RECT  915000.0 793200.0 925200.0 779400.0 ;
      RECT  915000.0 793200.0 925200.0 807000.0 ;
      RECT  915000.0 820800.0 925200.0 807000.0 ;
      RECT  915000.0 820800.0 925200.0 834600.0 ;
      RECT  915000.0 848400.0 925200.0 834600.0 ;
      RECT  915000.0 848400.0 925200.0 862200.0 ;
      RECT  915000.0 876000.0 925200.0 862200.0 ;
      RECT  915000.0 876000.0 925200.0 889800.0 ;
      RECT  915000.0 903600.0 925200.0 889800.0 ;
      RECT  915000.0 903600.0 925200.0 917400.0 ;
      RECT  915000.0 931200.0 925200.0 917400.0 ;
      RECT  915000.0 931200.0 925200.0 945000.0 ;
      RECT  915000.0 958800.0 925200.0 945000.0 ;
      RECT  915000.0 958800.0 925200.0 972600.0 ;
      RECT  915000.0 986400.0 925200.0 972600.0 ;
      RECT  915000.0 986400.0 925200.0 1000200.0 ;
      RECT  915000.0 1014000.0 925200.0 1000200.0 ;
      RECT  915000.0 1014000.0 925200.0 1027800.0 ;
      RECT  915000.0 1041600.0 925200.0 1027800.0 ;
      RECT  915000.0 1041600.0 925200.0 1055400.0 ;
      RECT  915000.0 1069200.0 925200.0 1055400.0 ;
      RECT  915000.0 1069200.0 925200.0 1083000.0 ;
      RECT  915000.0 1096800.0 925200.0 1083000.0 ;
      RECT  915000.0 1096800.0 925200.0 1110600.0 ;
      RECT  915000.0 1124400.0 925200.0 1110600.0 ;
      RECT  915000.0 1124400.0 925200.0 1138200.0 ;
      RECT  915000.0 1152000.0 925200.0 1138200.0 ;
      RECT  915000.0 1152000.0 925200.0 1165800.0 ;
      RECT  915000.0 1179600.0 925200.0 1165800.0 ;
      RECT  915000.0 1179600.0 925200.0 1193400.0 ;
      RECT  915000.0 1207200.0 925200.0 1193400.0 ;
      RECT  915000.0 1207200.0 925200.0 1221000.0 ;
      RECT  915000.0 1234800.0 925200.0 1221000.0 ;
      RECT  915000.0 1234800.0 925200.0 1248600.0 ;
      RECT  915000.0 1262400.0 925200.0 1248600.0 ;
      RECT  915000.0 1262400.0 925200.0 1276200.0 ;
      RECT  915000.0 1290000.0 925200.0 1276200.0 ;
      RECT  915000.0 1290000.0 925200.0 1303800.0 ;
      RECT  915000.0 1317600.0 925200.0 1303800.0 ;
      RECT  915000.0 1317600.0 925200.0 1331400.0 ;
      RECT  915000.0 1345200.0 925200.0 1331400.0 ;
      RECT  915000.0 1345200.0 925200.0 1359000.0 ;
      RECT  915000.0 1372800.0 925200.0 1359000.0 ;
      RECT  915000.0 1372800.0 925200.0 1386600.0 ;
      RECT  915000.0 1400400.0 925200.0 1386600.0 ;
      RECT  915000.0 1400400.0 925200.0 1414200.0 ;
      RECT  915000.0 1428000.0 925200.0 1414200.0 ;
      RECT  915000.0 1428000.0 925200.0 1441800.0 ;
      RECT  915000.0 1455600.0 925200.0 1441800.0 ;
      RECT  915000.0 1455600.0 925200.0 1469400.0 ;
      RECT  915000.0 1483200.0 925200.0 1469400.0 ;
      RECT  915000.0 1483200.0 925200.0 1497000.0 ;
      RECT  915000.0 1510800.0 925200.0 1497000.0 ;
      RECT  915000.0 1510800.0 925200.0 1524600.0 ;
      RECT  915000.0 1538400.0 925200.0 1524600.0 ;
      RECT  915000.0 1538400.0 925200.0 1552200.0 ;
      RECT  915000.0 1566000.0 925200.0 1552200.0 ;
      RECT  915000.0 1566000.0 925200.0 1579800.0 ;
      RECT  915000.0 1593600.0 925200.0 1579800.0 ;
      RECT  915000.0 1593600.0 925200.0 1607400.0 ;
      RECT  915000.0 1621200.0 925200.0 1607400.0 ;
      RECT  915000.0 1621200.0 925200.0 1635000.0 ;
      RECT  915000.0 1648800.0 925200.0 1635000.0 ;
      RECT  915000.0 1648800.0 925200.0 1662600.0 ;
      RECT  915000.0 1676400.0 925200.0 1662600.0 ;
      RECT  915000.0 1676400.0 925200.0 1690200.0 ;
      RECT  915000.0 1704000.0 925200.0 1690200.0 ;
      RECT  915000.0 1704000.0 925200.0 1717800.0 ;
      RECT  915000.0 1731600.0 925200.0 1717800.0 ;
      RECT  915000.0 1731600.0 925200.0 1745400.0 ;
      RECT  915000.0 1759200.0 925200.0 1745400.0 ;
      RECT  915000.0 1759200.0 925200.0 1773000.0 ;
      RECT  915000.0 1786800.0 925200.0 1773000.0 ;
      RECT  915000.0 1786800.0 925200.0 1800600.0 ;
      RECT  915000.0 1814400.0 925200.0 1800600.0 ;
      RECT  915000.0 1814400.0 925200.0 1828200.0 ;
      RECT  915000.0 1842000.0 925200.0 1828200.0 ;
      RECT  915000.0 1842000.0 925200.0 1855800.0 ;
      RECT  915000.0 1869600.0 925200.0 1855800.0 ;
      RECT  915000.0 1869600.0 925200.0 1883400.0 ;
      RECT  915000.0 1897200.0 925200.0 1883400.0 ;
      RECT  915000.0 1897200.0 925200.0 1911000.0 ;
      RECT  915000.0 1924800.0 925200.0 1911000.0 ;
      RECT  915000.0 1924800.0 925200.0 1938600.0 ;
      RECT  915000.0 1952400.0 925200.0 1938600.0 ;
      RECT  915000.0 1952400.0 925200.0 1966200.0 ;
      RECT  915000.0 1980000.0 925200.0 1966200.0 ;
      RECT  915000.0 1980000.0 925200.0 1993800.0 ;
      RECT  915000.0 2007600.0 925200.0 1993800.0 ;
      RECT  915000.0 2007600.0 925200.0 2021400.0 ;
      RECT  915000.0 2035200.0 925200.0 2021400.0 ;
      RECT  915000.0 2035200.0 925200.0 2049000.0 ;
      RECT  915000.0 2062800.0 925200.0 2049000.0 ;
      RECT  915000.0 2062800.0 925200.0 2076600.0 ;
      RECT  915000.0 2090400.0 925200.0 2076600.0 ;
      RECT  915000.0 2090400.0 925200.0 2104200.0 ;
      RECT  915000.0 2118000.0 925200.0 2104200.0 ;
      RECT  915000.0 2118000.0 925200.0 2131800.0 ;
      RECT  915000.0 2145600.0 925200.0 2131800.0 ;
      RECT  925200.0 379200.0 935400.0 393000.0 ;
      RECT  925200.0 406800.0 935400.0 393000.0 ;
      RECT  925200.0 406800.0 935400.0 420600.0 ;
      RECT  925200.0 434400.0 935400.0 420600.0 ;
      RECT  925200.0 434400.0 935400.0 448200.0 ;
      RECT  925200.0 462000.0 935400.0 448200.0 ;
      RECT  925200.0 462000.0 935400.0 475800.0 ;
      RECT  925200.0 489600.0 935400.0 475800.0 ;
      RECT  925200.0 489600.0 935400.0 503400.0 ;
      RECT  925200.0 517200.0 935400.0 503400.0 ;
      RECT  925200.0 517200.0 935400.0 531000.0 ;
      RECT  925200.0 544800.0 935400.0 531000.0 ;
      RECT  925200.0 544800.0 935400.0 558600.0 ;
      RECT  925200.0 572400.0 935400.0 558600.0 ;
      RECT  925200.0 572400.0 935400.0 586200.0 ;
      RECT  925200.0 600000.0 935400.0 586200.0 ;
      RECT  925200.0 600000.0 935400.0 613800.0 ;
      RECT  925200.0 627600.0 935400.0 613800.0 ;
      RECT  925200.0 627600.0 935400.0 641400.0 ;
      RECT  925200.0 655200.0 935400.0 641400.0 ;
      RECT  925200.0 655200.0 935400.0 669000.0 ;
      RECT  925200.0 682800.0 935400.0 669000.0 ;
      RECT  925200.0 682800.0 935400.0 696600.0 ;
      RECT  925200.0 710400.0 935400.0 696600.0 ;
      RECT  925200.0 710400.0 935400.0 724200.0 ;
      RECT  925200.0 738000.0 935400.0 724200.0 ;
      RECT  925200.0 738000.0 935400.0 751800.0 ;
      RECT  925200.0 765600.0 935400.0 751800.0 ;
      RECT  925200.0 765600.0 935400.0 779400.0 ;
      RECT  925200.0 793200.0 935400.0 779400.0 ;
      RECT  925200.0 793200.0 935400.0 807000.0 ;
      RECT  925200.0 820800.0 935400.0 807000.0 ;
      RECT  925200.0 820800.0 935400.0 834600.0 ;
      RECT  925200.0 848400.0 935400.0 834600.0 ;
      RECT  925200.0 848400.0 935400.0 862200.0 ;
      RECT  925200.0 876000.0 935400.0 862200.0 ;
      RECT  925200.0 876000.0 935400.0 889800.0 ;
      RECT  925200.0 903600.0 935400.0 889800.0 ;
      RECT  925200.0 903600.0 935400.0 917400.0 ;
      RECT  925200.0 931200.0 935400.0 917400.0 ;
      RECT  925200.0 931200.0 935400.0 945000.0 ;
      RECT  925200.0 958800.0 935400.0 945000.0 ;
      RECT  925200.0 958800.0 935400.0 972600.0 ;
      RECT  925200.0 986400.0 935400.0 972600.0 ;
      RECT  925200.0 986400.0 935400.0 1000200.0 ;
      RECT  925200.0 1014000.0 935400.0 1000200.0 ;
      RECT  925200.0 1014000.0 935400.0 1027800.0 ;
      RECT  925200.0 1041600.0 935400.0 1027800.0 ;
      RECT  925200.0 1041600.0 935400.0 1055400.0 ;
      RECT  925200.0 1069200.0 935400.0 1055400.0 ;
      RECT  925200.0 1069200.0 935400.0 1083000.0 ;
      RECT  925200.0 1096800.0 935400.0 1083000.0 ;
      RECT  925200.0 1096800.0 935400.0 1110600.0 ;
      RECT  925200.0 1124400.0 935400.0 1110600.0 ;
      RECT  925200.0 1124400.0 935400.0 1138200.0 ;
      RECT  925200.0 1152000.0 935400.0 1138200.0 ;
      RECT  925200.0 1152000.0 935400.0 1165800.0 ;
      RECT  925200.0 1179600.0 935400.0 1165800.0 ;
      RECT  925200.0 1179600.0 935400.0 1193400.0 ;
      RECT  925200.0 1207200.0 935400.0 1193400.0 ;
      RECT  925200.0 1207200.0 935400.0 1221000.0 ;
      RECT  925200.0 1234800.0 935400.0 1221000.0 ;
      RECT  925200.0 1234800.0 935400.0 1248600.0 ;
      RECT  925200.0 1262400.0 935400.0 1248600.0 ;
      RECT  925200.0 1262400.0 935400.0 1276200.0 ;
      RECT  925200.0 1290000.0 935400.0 1276200.0 ;
      RECT  925200.0 1290000.0 935400.0 1303800.0 ;
      RECT  925200.0 1317600.0 935400.0 1303800.0 ;
      RECT  925200.0 1317600.0 935400.0 1331400.0 ;
      RECT  925200.0 1345200.0 935400.0 1331400.0 ;
      RECT  925200.0 1345200.0 935400.0 1359000.0 ;
      RECT  925200.0 1372800.0 935400.0 1359000.0 ;
      RECT  925200.0 1372800.0 935400.0 1386600.0 ;
      RECT  925200.0 1400400.0 935400.0 1386600.0 ;
      RECT  925200.0 1400400.0 935400.0 1414200.0 ;
      RECT  925200.0 1428000.0 935400.0 1414200.0 ;
      RECT  925200.0 1428000.0 935400.0 1441800.0 ;
      RECT  925200.0 1455600.0 935400.0 1441800.0 ;
      RECT  925200.0 1455600.0 935400.0 1469400.0 ;
      RECT  925200.0 1483200.0 935400.0 1469400.0 ;
      RECT  925200.0 1483200.0 935400.0 1497000.0 ;
      RECT  925200.0 1510800.0 935400.0 1497000.0 ;
      RECT  925200.0 1510800.0 935400.0 1524600.0 ;
      RECT  925200.0 1538400.0 935400.0 1524600.0 ;
      RECT  925200.0 1538400.0 935400.0 1552200.0 ;
      RECT  925200.0 1566000.0 935400.0 1552200.0 ;
      RECT  925200.0 1566000.0 935400.0 1579800.0 ;
      RECT  925200.0 1593600.0 935400.0 1579800.0 ;
      RECT  925200.0 1593600.0 935400.0 1607400.0 ;
      RECT  925200.0 1621200.0 935400.0 1607400.0 ;
      RECT  925200.0 1621200.0 935400.0 1635000.0 ;
      RECT  925200.0 1648800.0 935400.0 1635000.0 ;
      RECT  925200.0 1648800.0 935400.0 1662600.0 ;
      RECT  925200.0 1676400.0 935400.0 1662600.0 ;
      RECT  925200.0 1676400.0 935400.0 1690200.0 ;
      RECT  925200.0 1704000.0 935400.0 1690200.0 ;
      RECT  925200.0 1704000.0 935400.0 1717800.0 ;
      RECT  925200.0 1731600.0 935400.0 1717800.0 ;
      RECT  925200.0 1731600.0 935400.0 1745400.0 ;
      RECT  925200.0 1759200.0 935400.0 1745400.0 ;
      RECT  925200.0 1759200.0 935400.0 1773000.0 ;
      RECT  925200.0 1786800.0 935400.0 1773000.0 ;
      RECT  925200.0 1786800.0 935400.0 1800600.0 ;
      RECT  925200.0 1814400.0 935400.0 1800600.0 ;
      RECT  925200.0 1814400.0 935400.0 1828200.0 ;
      RECT  925200.0 1842000.0 935400.0 1828200.0 ;
      RECT  925200.0 1842000.0 935400.0 1855800.0 ;
      RECT  925200.0 1869600.0 935400.0 1855800.0 ;
      RECT  925200.0 1869600.0 935400.0 1883400.0 ;
      RECT  925200.0 1897200.0 935400.0 1883400.0 ;
      RECT  925200.0 1897200.0 935400.0 1911000.0 ;
      RECT  925200.0 1924800.0 935400.0 1911000.0 ;
      RECT  925200.0 1924800.0 935400.0 1938600.0 ;
      RECT  925200.0 1952400.0 935400.0 1938600.0 ;
      RECT  925200.0 1952400.0 935400.0 1966200.0 ;
      RECT  925200.0 1980000.0 935400.0 1966200.0 ;
      RECT  925200.0 1980000.0 935400.0 1993800.0 ;
      RECT  925200.0 2007600.0 935400.0 1993800.0 ;
      RECT  925200.0 2007600.0 935400.0 2021400.0 ;
      RECT  925200.0 2035200.0 935400.0 2021400.0 ;
      RECT  925200.0 2035200.0 935400.0 2049000.0 ;
      RECT  925200.0 2062800.0 935400.0 2049000.0 ;
      RECT  925200.0 2062800.0 935400.0 2076600.0 ;
      RECT  925200.0 2090400.0 935400.0 2076600.0 ;
      RECT  925200.0 2090400.0 935400.0 2104200.0 ;
      RECT  925200.0 2118000.0 935400.0 2104200.0 ;
      RECT  925200.0 2118000.0 935400.0 2131800.0 ;
      RECT  925200.0 2145600.0 935400.0 2131800.0 ;
      RECT  935400.0 379200.0 945600.0 393000.0 ;
      RECT  935400.0 406800.0 945600.0 393000.0 ;
      RECT  935400.0 406800.0 945600.0 420600.0 ;
      RECT  935400.0 434400.0 945600.0 420600.0 ;
      RECT  935400.0 434400.0 945600.0 448200.0 ;
      RECT  935400.0 462000.0 945600.0 448200.0 ;
      RECT  935400.0 462000.0 945600.0 475800.0 ;
      RECT  935400.0 489600.0 945600.0 475800.0 ;
      RECT  935400.0 489600.0 945600.0 503400.0 ;
      RECT  935400.0 517200.0 945600.0 503400.0 ;
      RECT  935400.0 517200.0 945600.0 531000.0 ;
      RECT  935400.0 544800.0 945600.0 531000.0 ;
      RECT  935400.0 544800.0 945600.0 558600.0 ;
      RECT  935400.0 572400.0 945600.0 558600.0 ;
      RECT  935400.0 572400.0 945600.0 586200.0 ;
      RECT  935400.0 600000.0 945600.0 586200.0 ;
      RECT  935400.0 600000.0 945600.0 613800.0 ;
      RECT  935400.0 627600.0 945600.0 613800.0 ;
      RECT  935400.0 627600.0 945600.0 641400.0 ;
      RECT  935400.0 655200.0 945600.0 641400.0 ;
      RECT  935400.0 655200.0 945600.0 669000.0 ;
      RECT  935400.0 682800.0 945600.0 669000.0 ;
      RECT  935400.0 682800.0 945600.0 696600.0 ;
      RECT  935400.0 710400.0 945600.0 696600.0 ;
      RECT  935400.0 710400.0 945600.0 724200.0 ;
      RECT  935400.0 738000.0 945600.0 724200.0 ;
      RECT  935400.0 738000.0 945600.0 751800.0 ;
      RECT  935400.0 765600.0 945600.0 751800.0 ;
      RECT  935400.0 765600.0 945600.0 779400.0 ;
      RECT  935400.0 793200.0 945600.0 779400.0 ;
      RECT  935400.0 793200.0 945600.0 807000.0 ;
      RECT  935400.0 820800.0 945600.0 807000.0 ;
      RECT  935400.0 820800.0 945600.0 834600.0 ;
      RECT  935400.0 848400.0 945600.0 834600.0 ;
      RECT  935400.0 848400.0 945600.0 862200.0 ;
      RECT  935400.0 876000.0 945600.0 862200.0 ;
      RECT  935400.0 876000.0 945600.0 889800.0 ;
      RECT  935400.0 903600.0 945600.0 889800.0 ;
      RECT  935400.0 903600.0 945600.0 917400.0 ;
      RECT  935400.0 931200.0 945600.0 917400.0 ;
      RECT  935400.0 931200.0 945600.0 945000.0 ;
      RECT  935400.0 958800.0 945600.0 945000.0 ;
      RECT  935400.0 958800.0 945600.0 972600.0 ;
      RECT  935400.0 986400.0 945600.0 972600.0 ;
      RECT  935400.0 986400.0 945600.0 1000200.0 ;
      RECT  935400.0 1014000.0 945600.0 1000200.0 ;
      RECT  935400.0 1014000.0 945600.0 1027800.0 ;
      RECT  935400.0 1041600.0 945600.0 1027800.0 ;
      RECT  935400.0 1041600.0 945600.0 1055400.0 ;
      RECT  935400.0 1069200.0 945600.0 1055400.0 ;
      RECT  935400.0 1069200.0 945600.0 1083000.0 ;
      RECT  935400.0 1096800.0 945600.0 1083000.0 ;
      RECT  935400.0 1096800.0 945600.0 1110600.0 ;
      RECT  935400.0 1124400.0 945600.0 1110600.0 ;
      RECT  935400.0 1124400.0 945600.0 1138200.0 ;
      RECT  935400.0 1152000.0 945600.0 1138200.0 ;
      RECT  935400.0 1152000.0 945600.0 1165800.0 ;
      RECT  935400.0 1179600.0 945600.0 1165800.0 ;
      RECT  935400.0 1179600.0 945600.0 1193400.0 ;
      RECT  935400.0 1207200.0 945600.0 1193400.0 ;
      RECT  935400.0 1207200.0 945600.0 1221000.0 ;
      RECT  935400.0 1234800.0 945600.0 1221000.0 ;
      RECT  935400.0 1234800.0 945600.0 1248600.0 ;
      RECT  935400.0 1262400.0 945600.0 1248600.0 ;
      RECT  935400.0 1262400.0 945600.0 1276200.0 ;
      RECT  935400.0 1290000.0 945600.0 1276200.0 ;
      RECT  935400.0 1290000.0 945600.0 1303800.0 ;
      RECT  935400.0 1317600.0 945600.0 1303800.0 ;
      RECT  935400.0 1317600.0 945600.0 1331400.0 ;
      RECT  935400.0 1345200.0 945600.0 1331400.0 ;
      RECT  935400.0 1345200.0 945600.0 1359000.0 ;
      RECT  935400.0 1372800.0 945600.0 1359000.0 ;
      RECT  935400.0 1372800.0 945600.0 1386600.0 ;
      RECT  935400.0 1400400.0 945600.0 1386600.0 ;
      RECT  935400.0 1400400.0 945600.0 1414200.0 ;
      RECT  935400.0 1428000.0 945600.0 1414200.0 ;
      RECT  935400.0 1428000.0 945600.0 1441800.0 ;
      RECT  935400.0 1455600.0 945600.0 1441800.0 ;
      RECT  935400.0 1455600.0 945600.0 1469400.0 ;
      RECT  935400.0 1483200.0 945600.0 1469400.0 ;
      RECT  935400.0 1483200.0 945600.0 1497000.0 ;
      RECT  935400.0 1510800.0 945600.0 1497000.0 ;
      RECT  935400.0 1510800.0 945600.0 1524600.0 ;
      RECT  935400.0 1538400.0 945600.0 1524600.0 ;
      RECT  935400.0 1538400.0 945600.0 1552200.0 ;
      RECT  935400.0 1566000.0 945600.0 1552200.0 ;
      RECT  935400.0 1566000.0 945600.0 1579800.0 ;
      RECT  935400.0 1593600.0 945600.0 1579800.0 ;
      RECT  935400.0 1593600.0 945600.0 1607400.0 ;
      RECT  935400.0 1621200.0 945600.0 1607400.0 ;
      RECT  935400.0 1621200.0 945600.0 1635000.0 ;
      RECT  935400.0 1648800.0 945600.0 1635000.0 ;
      RECT  935400.0 1648800.0 945600.0 1662600.0 ;
      RECT  935400.0 1676400.0 945600.0 1662600.0 ;
      RECT  935400.0 1676400.0 945600.0 1690200.0 ;
      RECT  935400.0 1704000.0 945600.0 1690200.0 ;
      RECT  935400.0 1704000.0 945600.0 1717800.0 ;
      RECT  935400.0 1731600.0 945600.0 1717800.0 ;
      RECT  935400.0 1731600.0 945600.0 1745400.0 ;
      RECT  935400.0 1759200.0 945600.0 1745400.0 ;
      RECT  935400.0 1759200.0 945600.0 1773000.0 ;
      RECT  935400.0 1786800.0 945600.0 1773000.0 ;
      RECT  935400.0 1786800.0 945600.0 1800600.0 ;
      RECT  935400.0 1814400.0 945600.0 1800600.0 ;
      RECT  935400.0 1814400.0 945600.0 1828200.0 ;
      RECT  935400.0 1842000.0 945600.0 1828200.0 ;
      RECT  935400.0 1842000.0 945600.0 1855800.0 ;
      RECT  935400.0 1869600.0 945600.0 1855800.0 ;
      RECT  935400.0 1869600.0 945600.0 1883400.0 ;
      RECT  935400.0 1897200.0 945600.0 1883400.0 ;
      RECT  935400.0 1897200.0 945600.0 1911000.0 ;
      RECT  935400.0 1924800.0 945600.0 1911000.0 ;
      RECT  935400.0 1924800.0 945600.0 1938600.0 ;
      RECT  935400.0 1952400.0 945600.0 1938600.0 ;
      RECT  935400.0 1952400.0 945600.0 1966200.0 ;
      RECT  935400.0 1980000.0 945600.0 1966200.0 ;
      RECT  935400.0 1980000.0 945600.0 1993800.0 ;
      RECT  935400.0 2007600.0 945600.0 1993800.0 ;
      RECT  935400.0 2007600.0 945600.0 2021400.0 ;
      RECT  935400.0 2035200.0 945600.0 2021400.0 ;
      RECT  935400.0 2035200.0 945600.0 2049000.0 ;
      RECT  935400.0 2062800.0 945600.0 2049000.0 ;
      RECT  935400.0 2062800.0 945600.0 2076600.0 ;
      RECT  935400.0 2090400.0 945600.0 2076600.0 ;
      RECT  935400.0 2090400.0 945600.0 2104200.0 ;
      RECT  935400.0 2118000.0 945600.0 2104200.0 ;
      RECT  935400.0 2118000.0 945600.0 2131800.0 ;
      RECT  935400.0 2145600.0 945600.0 2131800.0 ;
      RECT  945600.0 379200.0 955800.0 393000.0 ;
      RECT  945600.0 406800.0 955800.0 393000.0 ;
      RECT  945600.0 406800.0 955800.0 420600.0 ;
      RECT  945600.0 434400.0 955800.0 420600.0 ;
      RECT  945600.0 434400.0 955800.0 448200.0 ;
      RECT  945600.0 462000.0 955800.0 448200.0 ;
      RECT  945600.0 462000.0 955800.0 475800.0 ;
      RECT  945600.0 489600.0 955800.0 475800.0 ;
      RECT  945600.0 489600.0 955800.0 503400.0 ;
      RECT  945600.0 517200.0 955800.0 503400.0 ;
      RECT  945600.0 517200.0 955800.0 531000.0 ;
      RECT  945600.0 544800.0 955800.0 531000.0 ;
      RECT  945600.0 544800.0 955800.0 558600.0 ;
      RECT  945600.0 572400.0 955800.0 558600.0 ;
      RECT  945600.0 572400.0 955800.0 586200.0 ;
      RECT  945600.0 600000.0 955800.0 586200.0 ;
      RECT  945600.0 600000.0 955800.0 613800.0 ;
      RECT  945600.0 627600.0 955800.0 613800.0 ;
      RECT  945600.0 627600.0 955800.0 641400.0 ;
      RECT  945600.0 655200.0 955800.0 641400.0 ;
      RECT  945600.0 655200.0 955800.0 669000.0 ;
      RECT  945600.0 682800.0 955800.0 669000.0 ;
      RECT  945600.0 682800.0 955800.0 696600.0 ;
      RECT  945600.0 710400.0 955800.0 696600.0 ;
      RECT  945600.0 710400.0 955800.0 724200.0 ;
      RECT  945600.0 738000.0 955800.0 724200.0 ;
      RECT  945600.0 738000.0 955800.0 751800.0 ;
      RECT  945600.0 765600.0 955800.0 751800.0 ;
      RECT  945600.0 765600.0 955800.0 779400.0 ;
      RECT  945600.0 793200.0 955800.0 779400.0 ;
      RECT  945600.0 793200.0 955800.0 807000.0 ;
      RECT  945600.0 820800.0 955800.0 807000.0 ;
      RECT  945600.0 820800.0 955800.0 834600.0 ;
      RECT  945600.0 848400.0 955800.0 834600.0 ;
      RECT  945600.0 848400.0 955800.0 862200.0 ;
      RECT  945600.0 876000.0 955800.0 862200.0 ;
      RECT  945600.0 876000.0 955800.0 889800.0 ;
      RECT  945600.0 903600.0 955800.0 889800.0 ;
      RECT  945600.0 903600.0 955800.0 917400.0 ;
      RECT  945600.0 931200.0 955800.0 917400.0 ;
      RECT  945600.0 931200.0 955800.0 945000.0 ;
      RECT  945600.0 958800.0 955800.0 945000.0 ;
      RECT  945600.0 958800.0 955800.0 972600.0 ;
      RECT  945600.0 986400.0 955800.0 972600.0 ;
      RECT  945600.0 986400.0 955800.0 1000200.0 ;
      RECT  945600.0 1014000.0 955800.0 1000200.0 ;
      RECT  945600.0 1014000.0 955800.0 1027800.0 ;
      RECT  945600.0 1041600.0 955800.0 1027800.0 ;
      RECT  945600.0 1041600.0 955800.0 1055400.0 ;
      RECT  945600.0 1069200.0 955800.0 1055400.0 ;
      RECT  945600.0 1069200.0 955800.0 1083000.0 ;
      RECT  945600.0 1096800.0 955800.0 1083000.0 ;
      RECT  945600.0 1096800.0 955800.0 1110600.0 ;
      RECT  945600.0 1124400.0 955800.0 1110600.0 ;
      RECT  945600.0 1124400.0 955800.0 1138200.0 ;
      RECT  945600.0 1152000.0 955800.0 1138200.0 ;
      RECT  945600.0 1152000.0 955800.0 1165800.0 ;
      RECT  945600.0 1179600.0 955800.0 1165800.0 ;
      RECT  945600.0 1179600.0 955800.0 1193400.0 ;
      RECT  945600.0 1207200.0 955800.0 1193400.0 ;
      RECT  945600.0 1207200.0 955800.0 1221000.0 ;
      RECT  945600.0 1234800.0 955800.0 1221000.0 ;
      RECT  945600.0 1234800.0 955800.0 1248600.0 ;
      RECT  945600.0 1262400.0 955800.0 1248600.0 ;
      RECT  945600.0 1262400.0 955800.0 1276200.0 ;
      RECT  945600.0 1290000.0 955800.0 1276200.0 ;
      RECT  945600.0 1290000.0 955800.0 1303800.0 ;
      RECT  945600.0 1317600.0 955800.0 1303800.0 ;
      RECT  945600.0 1317600.0 955800.0 1331400.0 ;
      RECT  945600.0 1345200.0 955800.0 1331400.0 ;
      RECT  945600.0 1345200.0 955800.0 1359000.0 ;
      RECT  945600.0 1372800.0 955800.0 1359000.0 ;
      RECT  945600.0 1372800.0 955800.0 1386600.0 ;
      RECT  945600.0 1400400.0 955800.0 1386600.0 ;
      RECT  945600.0 1400400.0 955800.0 1414200.0 ;
      RECT  945600.0 1428000.0 955800.0 1414200.0 ;
      RECT  945600.0 1428000.0 955800.0 1441800.0 ;
      RECT  945600.0 1455600.0 955800.0 1441800.0 ;
      RECT  945600.0 1455600.0 955800.0 1469400.0 ;
      RECT  945600.0 1483200.0 955800.0 1469400.0 ;
      RECT  945600.0 1483200.0 955800.0 1497000.0 ;
      RECT  945600.0 1510800.0 955800.0 1497000.0 ;
      RECT  945600.0 1510800.0 955800.0 1524600.0 ;
      RECT  945600.0 1538400.0 955800.0 1524600.0 ;
      RECT  945600.0 1538400.0 955800.0 1552200.0 ;
      RECT  945600.0 1566000.0 955800.0 1552200.0 ;
      RECT  945600.0 1566000.0 955800.0 1579800.0 ;
      RECT  945600.0 1593600.0 955800.0 1579800.0 ;
      RECT  945600.0 1593600.0 955800.0 1607400.0 ;
      RECT  945600.0 1621200.0 955800.0 1607400.0 ;
      RECT  945600.0 1621200.0 955800.0 1635000.0 ;
      RECT  945600.0 1648800.0 955800.0 1635000.0 ;
      RECT  945600.0 1648800.0 955800.0 1662600.0 ;
      RECT  945600.0 1676400.0 955800.0 1662600.0 ;
      RECT  945600.0 1676400.0 955800.0 1690200.0 ;
      RECT  945600.0 1704000.0 955800.0 1690200.0 ;
      RECT  945600.0 1704000.0 955800.0 1717800.0 ;
      RECT  945600.0 1731600.0 955800.0 1717800.0 ;
      RECT  945600.0 1731600.0 955800.0 1745400.0 ;
      RECT  945600.0 1759200.0 955800.0 1745400.0 ;
      RECT  945600.0 1759200.0 955800.0 1773000.0 ;
      RECT  945600.0 1786800.0 955800.0 1773000.0 ;
      RECT  945600.0 1786800.0 955800.0 1800600.0 ;
      RECT  945600.0 1814400.0 955800.0 1800600.0 ;
      RECT  945600.0 1814400.0 955800.0 1828200.0 ;
      RECT  945600.0 1842000.0 955800.0 1828200.0 ;
      RECT  945600.0 1842000.0 955800.0 1855800.0 ;
      RECT  945600.0 1869600.0 955800.0 1855800.0 ;
      RECT  945600.0 1869600.0 955800.0 1883400.0 ;
      RECT  945600.0 1897200.0 955800.0 1883400.0 ;
      RECT  945600.0 1897200.0 955800.0 1911000.0 ;
      RECT  945600.0 1924800.0 955800.0 1911000.0 ;
      RECT  945600.0 1924800.0 955800.0 1938600.0 ;
      RECT  945600.0 1952400.0 955800.0 1938600.0 ;
      RECT  945600.0 1952400.0 955800.0 1966200.0 ;
      RECT  945600.0 1980000.0 955800.0 1966200.0 ;
      RECT  945600.0 1980000.0 955800.0 1993800.0 ;
      RECT  945600.0 2007600.0 955800.0 1993800.0 ;
      RECT  945600.0 2007600.0 955800.0 2021400.0 ;
      RECT  945600.0 2035200.0 955800.0 2021400.0 ;
      RECT  945600.0 2035200.0 955800.0 2049000.0 ;
      RECT  945600.0 2062800.0 955800.0 2049000.0 ;
      RECT  945600.0 2062800.0 955800.0 2076600.0 ;
      RECT  945600.0 2090400.0 955800.0 2076600.0 ;
      RECT  945600.0 2090400.0 955800.0 2104200.0 ;
      RECT  945600.0 2118000.0 955800.0 2104200.0 ;
      RECT  945600.0 2118000.0 955800.0 2131800.0 ;
      RECT  945600.0 2145600.0 955800.0 2131800.0 ;
      RECT  955800.0 379200.0 966000.0 393000.0 ;
      RECT  955800.0 406800.0 966000.0 393000.0 ;
      RECT  955800.0 406800.0 966000.0 420600.0 ;
      RECT  955800.0 434400.0 966000.0 420600.0 ;
      RECT  955800.0 434400.0 966000.0 448200.0 ;
      RECT  955800.0 462000.0 966000.0 448200.0 ;
      RECT  955800.0 462000.0 966000.0 475800.0 ;
      RECT  955800.0 489600.0 966000.0 475800.0 ;
      RECT  955800.0 489600.0 966000.0 503400.0 ;
      RECT  955800.0 517200.0 966000.0 503400.0 ;
      RECT  955800.0 517200.0 966000.0 531000.0 ;
      RECT  955800.0 544800.0 966000.0 531000.0 ;
      RECT  955800.0 544800.0 966000.0 558600.0 ;
      RECT  955800.0 572400.0 966000.0 558600.0 ;
      RECT  955800.0 572400.0 966000.0 586200.0 ;
      RECT  955800.0 600000.0 966000.0 586200.0 ;
      RECT  955800.0 600000.0 966000.0 613800.0 ;
      RECT  955800.0 627600.0 966000.0 613800.0 ;
      RECT  955800.0 627600.0 966000.0 641400.0 ;
      RECT  955800.0 655200.0 966000.0 641400.0 ;
      RECT  955800.0 655200.0 966000.0 669000.0 ;
      RECT  955800.0 682800.0 966000.0 669000.0 ;
      RECT  955800.0 682800.0 966000.0 696600.0 ;
      RECT  955800.0 710400.0 966000.0 696600.0 ;
      RECT  955800.0 710400.0 966000.0 724200.0 ;
      RECT  955800.0 738000.0 966000.0 724200.0 ;
      RECT  955800.0 738000.0 966000.0 751800.0 ;
      RECT  955800.0 765600.0 966000.0 751800.0 ;
      RECT  955800.0 765600.0 966000.0 779400.0 ;
      RECT  955800.0 793200.0 966000.0 779400.0 ;
      RECT  955800.0 793200.0 966000.0 807000.0 ;
      RECT  955800.0 820800.0 966000.0 807000.0 ;
      RECT  955800.0 820800.0 966000.0 834600.0 ;
      RECT  955800.0 848400.0 966000.0 834600.0 ;
      RECT  955800.0 848400.0 966000.0 862200.0 ;
      RECT  955800.0 876000.0 966000.0 862200.0 ;
      RECT  955800.0 876000.0 966000.0 889800.0 ;
      RECT  955800.0 903600.0 966000.0 889800.0 ;
      RECT  955800.0 903600.0 966000.0 917400.0 ;
      RECT  955800.0 931200.0 966000.0 917400.0 ;
      RECT  955800.0 931200.0 966000.0 945000.0 ;
      RECT  955800.0 958800.0 966000.0 945000.0 ;
      RECT  955800.0 958800.0 966000.0 972600.0 ;
      RECT  955800.0 986400.0 966000.0 972600.0 ;
      RECT  955800.0 986400.0 966000.0 1000200.0 ;
      RECT  955800.0 1014000.0 966000.0 1000200.0 ;
      RECT  955800.0 1014000.0 966000.0 1027800.0 ;
      RECT  955800.0 1041600.0 966000.0 1027800.0 ;
      RECT  955800.0 1041600.0 966000.0 1055400.0 ;
      RECT  955800.0 1069200.0 966000.0 1055400.0 ;
      RECT  955800.0 1069200.0 966000.0 1083000.0 ;
      RECT  955800.0 1096800.0 966000.0 1083000.0 ;
      RECT  955800.0 1096800.0 966000.0 1110600.0 ;
      RECT  955800.0 1124400.0 966000.0 1110600.0 ;
      RECT  955800.0 1124400.0 966000.0 1138200.0 ;
      RECT  955800.0 1152000.0 966000.0 1138200.0 ;
      RECT  955800.0 1152000.0 966000.0 1165800.0 ;
      RECT  955800.0 1179600.0 966000.0 1165800.0 ;
      RECT  955800.0 1179600.0 966000.0 1193400.0 ;
      RECT  955800.0 1207200.0 966000.0 1193400.0 ;
      RECT  955800.0 1207200.0 966000.0 1221000.0 ;
      RECT  955800.0 1234800.0 966000.0 1221000.0 ;
      RECT  955800.0 1234800.0 966000.0 1248600.0 ;
      RECT  955800.0 1262400.0 966000.0 1248600.0 ;
      RECT  955800.0 1262400.0 966000.0 1276200.0 ;
      RECT  955800.0 1290000.0 966000.0 1276200.0 ;
      RECT  955800.0 1290000.0 966000.0 1303800.0 ;
      RECT  955800.0 1317600.0 966000.0 1303800.0 ;
      RECT  955800.0 1317600.0 966000.0 1331400.0 ;
      RECT  955800.0 1345200.0 966000.0 1331400.0 ;
      RECT  955800.0 1345200.0 966000.0 1359000.0 ;
      RECT  955800.0 1372800.0 966000.0 1359000.0 ;
      RECT  955800.0 1372800.0 966000.0 1386600.0 ;
      RECT  955800.0 1400400.0 966000.0 1386600.0 ;
      RECT  955800.0 1400400.0 966000.0 1414200.0 ;
      RECT  955800.0 1428000.0 966000.0 1414200.0 ;
      RECT  955800.0 1428000.0 966000.0 1441800.0 ;
      RECT  955800.0 1455600.0 966000.0 1441800.0 ;
      RECT  955800.0 1455600.0 966000.0 1469400.0 ;
      RECT  955800.0 1483200.0 966000.0 1469400.0 ;
      RECT  955800.0 1483200.0 966000.0 1497000.0 ;
      RECT  955800.0 1510800.0 966000.0 1497000.0 ;
      RECT  955800.0 1510800.0 966000.0 1524600.0 ;
      RECT  955800.0 1538400.0 966000.0 1524600.0 ;
      RECT  955800.0 1538400.0 966000.0 1552200.0 ;
      RECT  955800.0 1566000.0 966000.0 1552200.0 ;
      RECT  955800.0 1566000.0 966000.0 1579800.0 ;
      RECT  955800.0 1593600.0 966000.0 1579800.0 ;
      RECT  955800.0 1593600.0 966000.0 1607400.0 ;
      RECT  955800.0 1621200.0 966000.0 1607400.0 ;
      RECT  955800.0 1621200.0 966000.0 1635000.0 ;
      RECT  955800.0 1648800.0 966000.0 1635000.0 ;
      RECT  955800.0 1648800.0 966000.0 1662600.0 ;
      RECT  955800.0 1676400.0 966000.0 1662600.0 ;
      RECT  955800.0 1676400.0 966000.0 1690200.0 ;
      RECT  955800.0 1704000.0 966000.0 1690200.0 ;
      RECT  955800.0 1704000.0 966000.0 1717800.0 ;
      RECT  955800.0 1731600.0 966000.0 1717800.0 ;
      RECT  955800.0 1731600.0 966000.0 1745400.0 ;
      RECT  955800.0 1759200.0 966000.0 1745400.0 ;
      RECT  955800.0 1759200.0 966000.0 1773000.0 ;
      RECT  955800.0 1786800.0 966000.0 1773000.0 ;
      RECT  955800.0 1786800.0 966000.0 1800600.0 ;
      RECT  955800.0 1814400.0 966000.0 1800600.0 ;
      RECT  955800.0 1814400.0 966000.0 1828200.0 ;
      RECT  955800.0 1842000.0 966000.0 1828200.0 ;
      RECT  955800.0 1842000.0 966000.0 1855800.0 ;
      RECT  955800.0 1869600.0 966000.0 1855800.0 ;
      RECT  955800.0 1869600.0 966000.0 1883400.0 ;
      RECT  955800.0 1897200.0 966000.0 1883400.0 ;
      RECT  955800.0 1897200.0 966000.0 1911000.0 ;
      RECT  955800.0 1924800.0 966000.0 1911000.0 ;
      RECT  955800.0 1924800.0 966000.0 1938600.0 ;
      RECT  955800.0 1952400.0 966000.0 1938600.0 ;
      RECT  955800.0 1952400.0 966000.0 1966200.0 ;
      RECT  955800.0 1980000.0 966000.0 1966200.0 ;
      RECT  955800.0 1980000.0 966000.0 1993800.0 ;
      RECT  955800.0 2007600.0 966000.0 1993800.0 ;
      RECT  955800.0 2007600.0 966000.0 2021400.0 ;
      RECT  955800.0 2035200.0 966000.0 2021400.0 ;
      RECT  955800.0 2035200.0 966000.0 2049000.0 ;
      RECT  955800.0 2062800.0 966000.0 2049000.0 ;
      RECT  955800.0 2062800.0 966000.0 2076600.0 ;
      RECT  955800.0 2090400.0 966000.0 2076600.0 ;
      RECT  955800.0 2090400.0 966000.0 2104200.0 ;
      RECT  955800.0 2118000.0 966000.0 2104200.0 ;
      RECT  955800.0 2118000.0 966000.0 2131800.0 ;
      RECT  955800.0 2145600.0 966000.0 2131800.0 ;
      RECT  966000.0 379200.0 976200.0 393000.0 ;
      RECT  966000.0 406800.0 976200.0 393000.0 ;
      RECT  966000.0 406800.0 976200.0 420600.0 ;
      RECT  966000.0 434400.0 976200.0 420600.0 ;
      RECT  966000.0 434400.0 976200.0 448200.0 ;
      RECT  966000.0 462000.0 976200.0 448200.0 ;
      RECT  966000.0 462000.0 976200.0 475800.0 ;
      RECT  966000.0 489600.0 976200.0 475800.0 ;
      RECT  966000.0 489600.0 976200.0 503400.0 ;
      RECT  966000.0 517200.0 976200.0 503400.0 ;
      RECT  966000.0 517200.0 976200.0 531000.0 ;
      RECT  966000.0 544800.0 976200.0 531000.0 ;
      RECT  966000.0 544800.0 976200.0 558600.0 ;
      RECT  966000.0 572400.0 976200.0 558600.0 ;
      RECT  966000.0 572400.0 976200.0 586200.0 ;
      RECT  966000.0 600000.0 976200.0 586200.0 ;
      RECT  966000.0 600000.0 976200.0 613800.0 ;
      RECT  966000.0 627600.0 976200.0 613800.0 ;
      RECT  966000.0 627600.0 976200.0 641400.0 ;
      RECT  966000.0 655200.0 976200.0 641400.0 ;
      RECT  966000.0 655200.0 976200.0 669000.0 ;
      RECT  966000.0 682800.0 976200.0 669000.0 ;
      RECT  966000.0 682800.0 976200.0 696600.0 ;
      RECT  966000.0 710400.0 976200.0 696600.0 ;
      RECT  966000.0 710400.0 976200.0 724200.0 ;
      RECT  966000.0 738000.0 976200.0 724200.0 ;
      RECT  966000.0 738000.0 976200.0 751800.0 ;
      RECT  966000.0 765600.0 976200.0 751800.0 ;
      RECT  966000.0 765600.0 976200.0 779400.0 ;
      RECT  966000.0 793200.0 976200.0 779400.0 ;
      RECT  966000.0 793200.0 976200.0 807000.0 ;
      RECT  966000.0 820800.0 976200.0 807000.0 ;
      RECT  966000.0 820800.0 976200.0 834600.0 ;
      RECT  966000.0 848400.0 976200.0 834600.0 ;
      RECT  966000.0 848400.0 976200.0 862200.0 ;
      RECT  966000.0 876000.0 976200.0 862200.0 ;
      RECT  966000.0 876000.0 976200.0 889800.0 ;
      RECT  966000.0 903600.0 976200.0 889800.0 ;
      RECT  966000.0 903600.0 976200.0 917400.0 ;
      RECT  966000.0 931200.0 976200.0 917400.0 ;
      RECT  966000.0 931200.0 976200.0 945000.0 ;
      RECT  966000.0 958800.0 976200.0 945000.0 ;
      RECT  966000.0 958800.0 976200.0 972600.0 ;
      RECT  966000.0 986400.0 976200.0 972600.0 ;
      RECT  966000.0 986400.0 976200.0 1000200.0 ;
      RECT  966000.0 1014000.0 976200.0 1000200.0 ;
      RECT  966000.0 1014000.0 976200.0 1027800.0 ;
      RECT  966000.0 1041600.0 976200.0 1027800.0 ;
      RECT  966000.0 1041600.0 976200.0 1055400.0 ;
      RECT  966000.0 1069200.0 976200.0 1055400.0 ;
      RECT  966000.0 1069200.0 976200.0 1083000.0 ;
      RECT  966000.0 1096800.0 976200.0 1083000.0 ;
      RECT  966000.0 1096800.0 976200.0 1110600.0 ;
      RECT  966000.0 1124400.0 976200.0 1110600.0 ;
      RECT  966000.0 1124400.0 976200.0 1138200.0 ;
      RECT  966000.0 1152000.0 976200.0 1138200.0 ;
      RECT  966000.0 1152000.0 976200.0 1165800.0 ;
      RECT  966000.0 1179600.0 976200.0 1165800.0 ;
      RECT  966000.0 1179600.0 976200.0 1193400.0 ;
      RECT  966000.0 1207200.0 976200.0 1193400.0 ;
      RECT  966000.0 1207200.0 976200.0 1221000.0 ;
      RECT  966000.0 1234800.0 976200.0 1221000.0 ;
      RECT  966000.0 1234800.0 976200.0 1248600.0 ;
      RECT  966000.0 1262400.0 976200.0 1248600.0 ;
      RECT  966000.0 1262400.0 976200.0 1276200.0 ;
      RECT  966000.0 1290000.0 976200.0 1276200.0 ;
      RECT  966000.0 1290000.0 976200.0 1303800.0 ;
      RECT  966000.0 1317600.0 976200.0 1303800.0 ;
      RECT  966000.0 1317600.0 976200.0 1331400.0 ;
      RECT  966000.0 1345200.0 976200.0 1331400.0 ;
      RECT  966000.0 1345200.0 976200.0 1359000.0 ;
      RECT  966000.0 1372800.0 976200.0 1359000.0 ;
      RECT  966000.0 1372800.0 976200.0 1386600.0 ;
      RECT  966000.0 1400400.0 976200.0 1386600.0 ;
      RECT  966000.0 1400400.0 976200.0 1414200.0 ;
      RECT  966000.0 1428000.0 976200.0 1414200.0 ;
      RECT  966000.0 1428000.0 976200.0 1441800.0 ;
      RECT  966000.0 1455600.0 976200.0 1441800.0 ;
      RECT  966000.0 1455600.0 976200.0 1469400.0 ;
      RECT  966000.0 1483200.0 976200.0 1469400.0 ;
      RECT  966000.0 1483200.0 976200.0 1497000.0 ;
      RECT  966000.0 1510800.0 976200.0 1497000.0 ;
      RECT  966000.0 1510800.0 976200.0 1524600.0 ;
      RECT  966000.0 1538400.0 976200.0 1524600.0 ;
      RECT  966000.0 1538400.0 976200.0 1552200.0 ;
      RECT  966000.0 1566000.0 976200.0 1552200.0 ;
      RECT  966000.0 1566000.0 976200.0 1579800.0 ;
      RECT  966000.0 1593600.0 976200.0 1579800.0 ;
      RECT  966000.0 1593600.0 976200.0 1607400.0 ;
      RECT  966000.0 1621200.0 976200.0 1607400.0 ;
      RECT  966000.0 1621200.0 976200.0 1635000.0 ;
      RECT  966000.0 1648800.0 976200.0 1635000.0 ;
      RECT  966000.0 1648800.0 976200.0 1662600.0 ;
      RECT  966000.0 1676400.0 976200.0 1662600.0 ;
      RECT  966000.0 1676400.0 976200.0 1690200.0 ;
      RECT  966000.0 1704000.0 976200.0 1690200.0 ;
      RECT  966000.0 1704000.0 976200.0 1717800.0 ;
      RECT  966000.0 1731600.0 976200.0 1717800.0 ;
      RECT  966000.0 1731600.0 976200.0 1745400.0 ;
      RECT  966000.0 1759200.0 976200.0 1745400.0 ;
      RECT  966000.0 1759200.0 976200.0 1773000.0 ;
      RECT  966000.0 1786800.0 976200.0 1773000.0 ;
      RECT  966000.0 1786800.0 976200.0 1800600.0 ;
      RECT  966000.0 1814400.0 976200.0 1800600.0 ;
      RECT  966000.0 1814400.0 976200.0 1828200.0 ;
      RECT  966000.0 1842000.0 976200.0 1828200.0 ;
      RECT  966000.0 1842000.0 976200.0 1855800.0 ;
      RECT  966000.0 1869600.0 976200.0 1855800.0 ;
      RECT  966000.0 1869600.0 976200.0 1883400.0 ;
      RECT  966000.0 1897200.0 976200.0 1883400.0 ;
      RECT  966000.0 1897200.0 976200.0 1911000.0 ;
      RECT  966000.0 1924800.0 976200.0 1911000.0 ;
      RECT  966000.0 1924800.0 976200.0 1938600.0 ;
      RECT  966000.0 1952400.0 976200.0 1938600.0 ;
      RECT  966000.0 1952400.0 976200.0 1966200.0 ;
      RECT  966000.0 1980000.0 976200.0 1966200.0 ;
      RECT  966000.0 1980000.0 976200.0 1993800.0 ;
      RECT  966000.0 2007600.0 976200.0 1993800.0 ;
      RECT  966000.0 2007600.0 976200.0 2021400.0 ;
      RECT  966000.0 2035200.0 976200.0 2021400.0 ;
      RECT  966000.0 2035200.0 976200.0 2049000.0 ;
      RECT  966000.0 2062800.0 976200.0 2049000.0 ;
      RECT  966000.0 2062800.0 976200.0 2076600.0 ;
      RECT  966000.0 2090400.0 976200.0 2076600.0 ;
      RECT  966000.0 2090400.0 976200.0 2104200.0 ;
      RECT  966000.0 2118000.0 976200.0 2104200.0 ;
      RECT  966000.0 2118000.0 976200.0 2131800.0 ;
      RECT  966000.0 2145600.0 976200.0 2131800.0 ;
      RECT  976200.0 379200.0 986400.0 393000.0 ;
      RECT  976200.0 406800.0 986400.0 393000.0 ;
      RECT  976200.0 406800.0 986400.0 420600.0 ;
      RECT  976200.0 434400.0 986400.0 420600.0 ;
      RECT  976200.0 434400.0 986400.0 448200.0 ;
      RECT  976200.0 462000.0 986400.0 448200.0 ;
      RECT  976200.0 462000.0 986400.0 475800.0 ;
      RECT  976200.0 489600.0 986400.0 475800.0 ;
      RECT  976200.0 489600.0 986400.0 503400.0 ;
      RECT  976200.0 517200.0 986400.0 503400.0 ;
      RECT  976200.0 517200.0 986400.0 531000.0 ;
      RECT  976200.0 544800.0 986400.0 531000.0 ;
      RECT  976200.0 544800.0 986400.0 558600.0 ;
      RECT  976200.0 572400.0 986400.0 558600.0 ;
      RECT  976200.0 572400.0 986400.0 586200.0 ;
      RECT  976200.0 600000.0 986400.0 586200.0 ;
      RECT  976200.0 600000.0 986400.0 613800.0 ;
      RECT  976200.0 627600.0 986400.0 613800.0 ;
      RECT  976200.0 627600.0 986400.0 641400.0 ;
      RECT  976200.0 655200.0 986400.0 641400.0 ;
      RECT  976200.0 655200.0 986400.0 669000.0 ;
      RECT  976200.0 682800.0 986400.0 669000.0 ;
      RECT  976200.0 682800.0 986400.0 696600.0 ;
      RECT  976200.0 710400.0 986400.0 696600.0 ;
      RECT  976200.0 710400.0 986400.0 724200.0 ;
      RECT  976200.0 738000.0 986400.0 724200.0 ;
      RECT  976200.0 738000.0 986400.0 751800.0 ;
      RECT  976200.0 765600.0 986400.0 751800.0 ;
      RECT  976200.0 765600.0 986400.0 779400.0 ;
      RECT  976200.0 793200.0 986400.0 779400.0 ;
      RECT  976200.0 793200.0 986400.0 807000.0 ;
      RECT  976200.0 820800.0 986400.0 807000.0 ;
      RECT  976200.0 820800.0 986400.0 834600.0 ;
      RECT  976200.0 848400.0 986400.0 834600.0 ;
      RECT  976200.0 848400.0 986400.0 862200.0 ;
      RECT  976200.0 876000.0 986400.0 862200.0 ;
      RECT  976200.0 876000.0 986400.0 889800.0 ;
      RECT  976200.0 903600.0 986400.0 889800.0 ;
      RECT  976200.0 903600.0 986400.0 917400.0 ;
      RECT  976200.0 931200.0 986400.0 917400.0 ;
      RECT  976200.0 931200.0 986400.0 945000.0 ;
      RECT  976200.0 958800.0 986400.0 945000.0 ;
      RECT  976200.0 958800.0 986400.0 972600.0 ;
      RECT  976200.0 986400.0 986400.0 972600.0 ;
      RECT  976200.0 986400.0 986400.0 1000200.0 ;
      RECT  976200.0 1014000.0 986400.0 1000200.0 ;
      RECT  976200.0 1014000.0 986400.0 1027800.0 ;
      RECT  976200.0 1041600.0 986400.0 1027800.0 ;
      RECT  976200.0 1041600.0 986400.0 1055400.0 ;
      RECT  976200.0 1069200.0 986400.0 1055400.0 ;
      RECT  976200.0 1069200.0 986400.0 1083000.0 ;
      RECT  976200.0 1096800.0 986400.0 1083000.0 ;
      RECT  976200.0 1096800.0 986400.0 1110600.0 ;
      RECT  976200.0 1124400.0 986400.0 1110600.0 ;
      RECT  976200.0 1124400.0 986400.0 1138200.0 ;
      RECT  976200.0 1152000.0 986400.0 1138200.0 ;
      RECT  976200.0 1152000.0 986400.0 1165800.0 ;
      RECT  976200.0 1179600.0 986400.0 1165800.0 ;
      RECT  976200.0 1179600.0 986400.0 1193400.0 ;
      RECT  976200.0 1207200.0 986400.0 1193400.0 ;
      RECT  976200.0 1207200.0 986400.0 1221000.0 ;
      RECT  976200.0 1234800.0 986400.0 1221000.0 ;
      RECT  976200.0 1234800.0 986400.0 1248600.0 ;
      RECT  976200.0 1262400.0 986400.0 1248600.0 ;
      RECT  976200.0 1262400.0 986400.0 1276200.0 ;
      RECT  976200.0 1290000.0 986400.0 1276200.0 ;
      RECT  976200.0 1290000.0 986400.0 1303800.0 ;
      RECT  976200.0 1317600.0 986400.0 1303800.0 ;
      RECT  976200.0 1317600.0 986400.0 1331400.0 ;
      RECT  976200.0 1345200.0 986400.0 1331400.0 ;
      RECT  976200.0 1345200.0 986400.0 1359000.0 ;
      RECT  976200.0 1372800.0 986400.0 1359000.0 ;
      RECT  976200.0 1372800.0 986400.0 1386600.0 ;
      RECT  976200.0 1400400.0 986400.0 1386600.0 ;
      RECT  976200.0 1400400.0 986400.0 1414200.0 ;
      RECT  976200.0 1428000.0 986400.0 1414200.0 ;
      RECT  976200.0 1428000.0 986400.0 1441800.0 ;
      RECT  976200.0 1455600.0 986400.0 1441800.0 ;
      RECT  976200.0 1455600.0 986400.0 1469400.0 ;
      RECT  976200.0 1483200.0 986400.0 1469400.0 ;
      RECT  976200.0 1483200.0 986400.0 1497000.0 ;
      RECT  976200.0 1510800.0 986400.0 1497000.0 ;
      RECT  976200.0 1510800.0 986400.0 1524600.0 ;
      RECT  976200.0 1538400.0 986400.0 1524600.0 ;
      RECT  976200.0 1538400.0 986400.0 1552200.0 ;
      RECT  976200.0 1566000.0 986400.0 1552200.0 ;
      RECT  976200.0 1566000.0 986400.0 1579800.0 ;
      RECT  976200.0 1593600.0 986400.0 1579800.0 ;
      RECT  976200.0 1593600.0 986400.0 1607400.0 ;
      RECT  976200.0 1621200.0 986400.0 1607400.0 ;
      RECT  976200.0 1621200.0 986400.0 1635000.0 ;
      RECT  976200.0 1648800.0 986400.0 1635000.0 ;
      RECT  976200.0 1648800.0 986400.0 1662600.0 ;
      RECT  976200.0 1676400.0 986400.0 1662600.0 ;
      RECT  976200.0 1676400.0 986400.0 1690200.0 ;
      RECT  976200.0 1704000.0 986400.0 1690200.0 ;
      RECT  976200.0 1704000.0 986400.0 1717800.0 ;
      RECT  976200.0 1731600.0 986400.0 1717800.0 ;
      RECT  976200.0 1731600.0 986400.0 1745400.0 ;
      RECT  976200.0 1759200.0 986400.0 1745400.0 ;
      RECT  976200.0 1759200.0 986400.0 1773000.0 ;
      RECT  976200.0 1786800.0 986400.0 1773000.0 ;
      RECT  976200.0 1786800.0 986400.0 1800600.0 ;
      RECT  976200.0 1814400.0 986400.0 1800600.0 ;
      RECT  976200.0 1814400.0 986400.0 1828200.0 ;
      RECT  976200.0 1842000.0 986400.0 1828200.0 ;
      RECT  976200.0 1842000.0 986400.0 1855800.0 ;
      RECT  976200.0 1869600.0 986400.0 1855800.0 ;
      RECT  976200.0 1869600.0 986400.0 1883400.0 ;
      RECT  976200.0 1897200.0 986400.0 1883400.0 ;
      RECT  976200.0 1897200.0 986400.0 1911000.0 ;
      RECT  976200.0 1924800.0 986400.0 1911000.0 ;
      RECT  976200.0 1924800.0 986400.0 1938600.0 ;
      RECT  976200.0 1952400.0 986400.0 1938600.0 ;
      RECT  976200.0 1952400.0 986400.0 1966200.0 ;
      RECT  976200.0 1980000.0 986400.0 1966200.0 ;
      RECT  976200.0 1980000.0 986400.0 1993800.0 ;
      RECT  976200.0 2007600.0 986400.0 1993800.0 ;
      RECT  976200.0 2007600.0 986400.0 2021400.0 ;
      RECT  976200.0 2035200.0 986400.0 2021400.0 ;
      RECT  976200.0 2035200.0 986400.0 2049000.0 ;
      RECT  976200.0 2062800.0 986400.0 2049000.0 ;
      RECT  976200.0 2062800.0 986400.0 2076600.0 ;
      RECT  976200.0 2090400.0 986400.0 2076600.0 ;
      RECT  976200.0 2090400.0 986400.0 2104200.0 ;
      RECT  976200.0 2118000.0 986400.0 2104200.0 ;
      RECT  976200.0 2118000.0 986400.0 2131800.0 ;
      RECT  976200.0 2145600.0 986400.0 2131800.0 ;
      RECT  986400.0 379200.0 996600.0 393000.0 ;
      RECT  986400.0 406800.0 996600.0 393000.0 ;
      RECT  986400.0 406800.0 996600.0 420600.0 ;
      RECT  986400.0 434400.0 996600.0 420600.0 ;
      RECT  986400.0 434400.0 996600.0 448200.0 ;
      RECT  986400.0 462000.0 996600.0 448200.0 ;
      RECT  986400.0 462000.0 996600.0 475800.0 ;
      RECT  986400.0 489600.0 996600.0 475800.0 ;
      RECT  986400.0 489600.0 996600.0 503400.0 ;
      RECT  986400.0 517200.0 996600.0 503400.0 ;
      RECT  986400.0 517200.0 996600.0 531000.0 ;
      RECT  986400.0 544800.0 996600.0 531000.0 ;
      RECT  986400.0 544800.0 996600.0 558600.0 ;
      RECT  986400.0 572400.0 996600.0 558600.0 ;
      RECT  986400.0 572400.0 996600.0 586200.0 ;
      RECT  986400.0 600000.0 996600.0 586200.0 ;
      RECT  986400.0 600000.0 996600.0 613800.0 ;
      RECT  986400.0 627600.0 996600.0 613800.0 ;
      RECT  986400.0 627600.0 996600.0 641400.0 ;
      RECT  986400.0 655200.0 996600.0 641400.0 ;
      RECT  986400.0 655200.0 996600.0 669000.0 ;
      RECT  986400.0 682800.0 996600.0 669000.0 ;
      RECT  986400.0 682800.0 996600.0 696600.0 ;
      RECT  986400.0 710400.0 996600.0 696600.0 ;
      RECT  986400.0 710400.0 996600.0 724200.0 ;
      RECT  986400.0 738000.0 996600.0 724200.0 ;
      RECT  986400.0 738000.0 996600.0 751800.0 ;
      RECT  986400.0 765600.0 996600.0 751800.0 ;
      RECT  986400.0 765600.0 996600.0 779400.0 ;
      RECT  986400.0 793200.0 996600.0 779400.0 ;
      RECT  986400.0 793200.0 996600.0 807000.0 ;
      RECT  986400.0 820800.0 996600.0 807000.0 ;
      RECT  986400.0 820800.0 996600.0 834600.0 ;
      RECT  986400.0 848400.0 996600.0 834600.0 ;
      RECT  986400.0 848400.0 996600.0 862200.0 ;
      RECT  986400.0 876000.0 996600.0 862200.0 ;
      RECT  986400.0 876000.0 996600.0 889800.0 ;
      RECT  986400.0 903600.0 996600.0 889800.0 ;
      RECT  986400.0 903600.0 996600.0 917400.0 ;
      RECT  986400.0 931200.0 996600.0 917400.0 ;
      RECT  986400.0 931200.0 996600.0 945000.0 ;
      RECT  986400.0 958800.0 996600.0 945000.0 ;
      RECT  986400.0 958800.0 996600.0 972600.0 ;
      RECT  986400.0 986400.0 996600.0 972600.0 ;
      RECT  986400.0 986400.0 996600.0 1000200.0 ;
      RECT  986400.0 1014000.0 996600.0 1000200.0 ;
      RECT  986400.0 1014000.0 996600.0 1027800.0 ;
      RECT  986400.0 1041600.0 996600.0 1027800.0 ;
      RECT  986400.0 1041600.0 996600.0 1055400.0 ;
      RECT  986400.0 1069200.0 996600.0 1055400.0 ;
      RECT  986400.0 1069200.0 996600.0 1083000.0 ;
      RECT  986400.0 1096800.0 996600.0 1083000.0 ;
      RECT  986400.0 1096800.0 996600.0 1110600.0 ;
      RECT  986400.0 1124400.0 996600.0 1110600.0 ;
      RECT  986400.0 1124400.0 996600.0 1138200.0 ;
      RECT  986400.0 1152000.0 996600.0 1138200.0 ;
      RECT  986400.0 1152000.0 996600.0 1165800.0 ;
      RECT  986400.0 1179600.0 996600.0 1165800.0 ;
      RECT  986400.0 1179600.0 996600.0 1193400.0 ;
      RECT  986400.0 1207200.0 996600.0 1193400.0 ;
      RECT  986400.0 1207200.0 996600.0 1221000.0 ;
      RECT  986400.0 1234800.0 996600.0 1221000.0 ;
      RECT  986400.0 1234800.0 996600.0 1248600.0 ;
      RECT  986400.0 1262400.0 996600.0 1248600.0 ;
      RECT  986400.0 1262400.0 996600.0 1276200.0 ;
      RECT  986400.0 1290000.0 996600.0 1276200.0 ;
      RECT  986400.0 1290000.0 996600.0 1303800.0 ;
      RECT  986400.0 1317600.0 996600.0 1303800.0 ;
      RECT  986400.0 1317600.0 996600.0 1331400.0 ;
      RECT  986400.0 1345200.0 996600.0 1331400.0 ;
      RECT  986400.0 1345200.0 996600.0 1359000.0 ;
      RECT  986400.0 1372800.0 996600.0 1359000.0 ;
      RECT  986400.0 1372800.0 996600.0 1386600.0 ;
      RECT  986400.0 1400400.0 996600.0 1386600.0 ;
      RECT  986400.0 1400400.0 996600.0 1414200.0 ;
      RECT  986400.0 1428000.0 996600.0 1414200.0 ;
      RECT  986400.0 1428000.0 996600.0 1441800.0 ;
      RECT  986400.0 1455600.0 996600.0 1441800.0 ;
      RECT  986400.0 1455600.0 996600.0 1469400.0 ;
      RECT  986400.0 1483200.0 996600.0 1469400.0 ;
      RECT  986400.0 1483200.0 996600.0 1497000.0 ;
      RECT  986400.0 1510800.0 996600.0 1497000.0 ;
      RECT  986400.0 1510800.0 996600.0 1524600.0 ;
      RECT  986400.0 1538400.0 996600.0 1524600.0 ;
      RECT  986400.0 1538400.0 996600.0 1552200.0 ;
      RECT  986400.0 1566000.0 996600.0 1552200.0 ;
      RECT  986400.0 1566000.0 996600.0 1579800.0 ;
      RECT  986400.0 1593600.0 996600.0 1579800.0 ;
      RECT  986400.0 1593600.0 996600.0 1607400.0 ;
      RECT  986400.0 1621200.0 996600.0 1607400.0 ;
      RECT  986400.0 1621200.0 996600.0 1635000.0 ;
      RECT  986400.0 1648800.0 996600.0 1635000.0 ;
      RECT  986400.0 1648800.0 996600.0 1662600.0 ;
      RECT  986400.0 1676400.0 996600.0 1662600.0 ;
      RECT  986400.0 1676400.0 996600.0 1690200.0 ;
      RECT  986400.0 1704000.0 996600.0 1690200.0 ;
      RECT  986400.0 1704000.0 996600.0 1717800.0 ;
      RECT  986400.0 1731600.0 996600.0 1717800.0 ;
      RECT  986400.0 1731600.0 996600.0 1745400.0 ;
      RECT  986400.0 1759200.0 996600.0 1745400.0 ;
      RECT  986400.0 1759200.0 996600.0 1773000.0 ;
      RECT  986400.0 1786800.0 996600.0 1773000.0 ;
      RECT  986400.0 1786800.0 996600.0 1800600.0 ;
      RECT  986400.0 1814400.0 996600.0 1800600.0 ;
      RECT  986400.0 1814400.0 996600.0 1828200.0 ;
      RECT  986400.0 1842000.0 996600.0 1828200.0 ;
      RECT  986400.0 1842000.0 996600.0 1855800.0 ;
      RECT  986400.0 1869600.0 996600.0 1855800.0 ;
      RECT  986400.0 1869600.0 996600.0 1883400.0 ;
      RECT  986400.0 1897200.0 996600.0 1883400.0 ;
      RECT  986400.0 1897200.0 996600.0 1911000.0 ;
      RECT  986400.0 1924800.0 996600.0 1911000.0 ;
      RECT  986400.0 1924800.0 996600.0 1938600.0 ;
      RECT  986400.0 1952400.0 996600.0 1938600.0 ;
      RECT  986400.0 1952400.0 996600.0 1966200.0 ;
      RECT  986400.0 1980000.0 996600.0 1966200.0 ;
      RECT  986400.0 1980000.0 996600.0 1993800.0 ;
      RECT  986400.0 2007600.0 996600.0 1993800.0 ;
      RECT  986400.0 2007600.0 996600.0 2021400.0 ;
      RECT  986400.0 2035200.0 996600.0 2021400.0 ;
      RECT  986400.0 2035200.0 996600.0 2049000.0 ;
      RECT  986400.0 2062800.0 996600.0 2049000.0 ;
      RECT  986400.0 2062800.0 996600.0 2076600.0 ;
      RECT  986400.0 2090400.0 996600.0 2076600.0 ;
      RECT  986400.0 2090400.0 996600.0 2104200.0 ;
      RECT  986400.0 2118000.0 996600.0 2104200.0 ;
      RECT  986400.0 2118000.0 996600.0 2131800.0 ;
      RECT  986400.0 2145600.0 996600.0 2131800.0 ;
      RECT  996600.0 379200.0 1006800.0 393000.0 ;
      RECT  996600.0 406800.0 1006800.0 393000.0 ;
      RECT  996600.0 406800.0 1006800.0 420600.0 ;
      RECT  996600.0 434400.0 1006800.0 420600.0 ;
      RECT  996600.0 434400.0 1006800.0 448200.0 ;
      RECT  996600.0 462000.0 1006800.0 448200.0 ;
      RECT  996600.0 462000.0 1006800.0 475800.0 ;
      RECT  996600.0 489600.0 1006800.0 475800.0 ;
      RECT  996600.0 489600.0 1006800.0 503400.0 ;
      RECT  996600.0 517200.0 1006800.0 503400.0 ;
      RECT  996600.0 517200.0 1006800.0 531000.0 ;
      RECT  996600.0 544800.0 1006800.0 531000.0 ;
      RECT  996600.0 544800.0 1006800.0 558600.0 ;
      RECT  996600.0 572400.0 1006800.0 558600.0 ;
      RECT  996600.0 572400.0 1006800.0 586200.0 ;
      RECT  996600.0 600000.0 1006800.0 586200.0 ;
      RECT  996600.0 600000.0 1006800.0 613800.0 ;
      RECT  996600.0 627600.0 1006800.0 613800.0 ;
      RECT  996600.0 627600.0 1006800.0 641400.0 ;
      RECT  996600.0 655200.0 1006800.0 641400.0 ;
      RECT  996600.0 655200.0 1006800.0 669000.0 ;
      RECT  996600.0 682800.0 1006800.0 669000.0 ;
      RECT  996600.0 682800.0 1006800.0 696600.0 ;
      RECT  996600.0 710400.0 1006800.0 696600.0 ;
      RECT  996600.0 710400.0 1006800.0 724200.0 ;
      RECT  996600.0 738000.0 1006800.0 724200.0 ;
      RECT  996600.0 738000.0 1006800.0 751800.0 ;
      RECT  996600.0 765600.0 1006800.0 751800.0 ;
      RECT  996600.0 765600.0 1006800.0 779400.0 ;
      RECT  996600.0 793200.0 1006800.0 779400.0 ;
      RECT  996600.0 793200.0 1006800.0 807000.0 ;
      RECT  996600.0 820800.0 1006800.0 807000.0 ;
      RECT  996600.0 820800.0 1006800.0 834600.0 ;
      RECT  996600.0 848400.0 1006800.0 834600.0 ;
      RECT  996600.0 848400.0 1006800.0 862200.0 ;
      RECT  996600.0 876000.0 1006800.0 862200.0 ;
      RECT  996600.0 876000.0 1006800.0 889800.0 ;
      RECT  996600.0 903600.0 1006800.0 889800.0 ;
      RECT  996600.0 903600.0 1006800.0 917400.0 ;
      RECT  996600.0 931200.0 1006800.0 917400.0 ;
      RECT  996600.0 931200.0 1006800.0 945000.0 ;
      RECT  996600.0 958800.0 1006800.0 945000.0 ;
      RECT  996600.0 958800.0 1006800.0 972600.0 ;
      RECT  996600.0 986400.0 1006800.0 972600.0 ;
      RECT  996600.0 986400.0 1006800.0 1000200.0 ;
      RECT  996600.0 1014000.0 1006800.0 1000200.0 ;
      RECT  996600.0 1014000.0 1006800.0 1027800.0 ;
      RECT  996600.0 1041600.0 1006800.0 1027800.0 ;
      RECT  996600.0 1041600.0 1006800.0 1055400.0 ;
      RECT  996600.0 1069200.0 1006800.0 1055400.0 ;
      RECT  996600.0 1069200.0 1006800.0 1083000.0 ;
      RECT  996600.0 1096800.0 1006800.0 1083000.0 ;
      RECT  996600.0 1096800.0 1006800.0 1110600.0 ;
      RECT  996600.0 1124400.0 1006800.0 1110600.0 ;
      RECT  996600.0 1124400.0 1006800.0 1138200.0 ;
      RECT  996600.0 1152000.0 1006800.0 1138200.0 ;
      RECT  996600.0 1152000.0 1006800.0 1165800.0 ;
      RECT  996600.0 1179600.0 1006800.0 1165800.0 ;
      RECT  996600.0 1179600.0 1006800.0 1193400.0 ;
      RECT  996600.0 1207200.0 1006800.0 1193400.0 ;
      RECT  996600.0 1207200.0 1006800.0 1221000.0 ;
      RECT  996600.0 1234800.0 1006800.0 1221000.0 ;
      RECT  996600.0 1234800.0 1006800.0 1248600.0 ;
      RECT  996600.0 1262400.0 1006800.0 1248600.0 ;
      RECT  996600.0 1262400.0 1006800.0 1276200.0 ;
      RECT  996600.0 1290000.0 1006800.0 1276200.0 ;
      RECT  996600.0 1290000.0 1006800.0 1303800.0 ;
      RECT  996600.0 1317600.0 1006800.0 1303800.0 ;
      RECT  996600.0 1317600.0 1006800.0 1331400.0 ;
      RECT  996600.0 1345200.0 1006800.0 1331400.0 ;
      RECT  996600.0 1345200.0 1006800.0 1359000.0 ;
      RECT  996600.0 1372800.0 1006800.0 1359000.0 ;
      RECT  996600.0 1372800.0 1006800.0 1386600.0 ;
      RECT  996600.0 1400400.0 1006800.0 1386600.0 ;
      RECT  996600.0 1400400.0 1006800.0 1414200.0 ;
      RECT  996600.0 1428000.0 1006800.0 1414200.0 ;
      RECT  996600.0 1428000.0 1006800.0 1441800.0 ;
      RECT  996600.0 1455600.0 1006800.0 1441800.0 ;
      RECT  996600.0 1455600.0 1006800.0 1469400.0 ;
      RECT  996600.0 1483200.0 1006800.0 1469400.0 ;
      RECT  996600.0 1483200.0 1006800.0 1497000.0 ;
      RECT  996600.0 1510800.0 1006800.0 1497000.0 ;
      RECT  996600.0 1510800.0 1006800.0 1524600.0 ;
      RECT  996600.0 1538400.0 1006800.0 1524600.0 ;
      RECT  996600.0 1538400.0 1006800.0 1552200.0 ;
      RECT  996600.0 1566000.0 1006800.0 1552200.0 ;
      RECT  996600.0 1566000.0 1006800.0 1579800.0 ;
      RECT  996600.0 1593600.0 1006800.0 1579800.0 ;
      RECT  996600.0 1593600.0 1006800.0 1607400.0 ;
      RECT  996600.0 1621200.0 1006800.0 1607400.0 ;
      RECT  996600.0 1621200.0 1006800.0 1635000.0 ;
      RECT  996600.0 1648800.0 1006800.0 1635000.0 ;
      RECT  996600.0 1648800.0 1006800.0 1662600.0 ;
      RECT  996600.0 1676400.0 1006800.0 1662600.0 ;
      RECT  996600.0 1676400.0 1006800.0 1690200.0 ;
      RECT  996600.0 1704000.0 1006800.0 1690200.0 ;
      RECT  996600.0 1704000.0 1006800.0 1717800.0 ;
      RECT  996600.0 1731600.0 1006800.0 1717800.0 ;
      RECT  996600.0 1731600.0 1006800.0 1745400.0 ;
      RECT  996600.0 1759200.0 1006800.0 1745400.0 ;
      RECT  996600.0 1759200.0 1006800.0 1773000.0 ;
      RECT  996600.0 1786800.0 1006800.0 1773000.0 ;
      RECT  996600.0 1786800.0 1006800.0 1800600.0 ;
      RECT  996600.0 1814400.0 1006800.0 1800600.0 ;
      RECT  996600.0 1814400.0 1006800.0 1828200.0 ;
      RECT  996600.0 1842000.0 1006800.0 1828200.0 ;
      RECT  996600.0 1842000.0 1006800.0 1855800.0 ;
      RECT  996600.0 1869600.0 1006800.0 1855800.0 ;
      RECT  996600.0 1869600.0 1006800.0 1883400.0 ;
      RECT  996600.0 1897200.0 1006800.0 1883400.0 ;
      RECT  996600.0 1897200.0 1006800.0 1911000.0 ;
      RECT  996600.0 1924800.0 1006800.0 1911000.0 ;
      RECT  996600.0 1924800.0 1006800.0 1938600.0 ;
      RECT  996600.0 1952400.0 1006800.0 1938600.0 ;
      RECT  996600.0 1952400.0 1006800.0 1966200.0 ;
      RECT  996600.0 1980000.0 1006800.0 1966200.0 ;
      RECT  996600.0 1980000.0 1006800.0 1993800.0 ;
      RECT  996600.0 2007600.0 1006800.0 1993800.0 ;
      RECT  996600.0 2007600.0 1006800.0 2021400.0 ;
      RECT  996600.0 2035200.0 1006800.0 2021400.0 ;
      RECT  996600.0 2035200.0 1006800.0 2049000.0 ;
      RECT  996600.0 2062800.0 1006800.0 2049000.0 ;
      RECT  996600.0 2062800.0 1006800.0 2076600.0 ;
      RECT  996600.0 2090400.0 1006800.0 2076600.0 ;
      RECT  996600.0 2090400.0 1006800.0 2104200.0 ;
      RECT  996600.0 2118000.0 1006800.0 2104200.0 ;
      RECT  996600.0 2118000.0 1006800.0 2131800.0 ;
      RECT  996600.0 2145600.0 1006800.0 2131800.0 ;
      RECT  1006800.0 379200.0 1017000.0 393000.0 ;
      RECT  1006800.0 406800.0 1017000.0 393000.0 ;
      RECT  1006800.0 406800.0 1017000.0 420600.0 ;
      RECT  1006800.0 434400.0 1017000.0 420600.0 ;
      RECT  1006800.0 434400.0 1017000.0 448200.0 ;
      RECT  1006800.0 462000.0 1017000.0 448200.0 ;
      RECT  1006800.0 462000.0 1017000.0 475800.0 ;
      RECT  1006800.0 489600.0 1017000.0 475800.0 ;
      RECT  1006800.0 489600.0 1017000.0 503400.0 ;
      RECT  1006800.0 517200.0 1017000.0 503400.0 ;
      RECT  1006800.0 517200.0 1017000.0 531000.0 ;
      RECT  1006800.0 544800.0 1017000.0 531000.0 ;
      RECT  1006800.0 544800.0 1017000.0 558600.0 ;
      RECT  1006800.0 572400.0 1017000.0 558600.0 ;
      RECT  1006800.0 572400.0 1017000.0 586200.0 ;
      RECT  1006800.0 600000.0 1017000.0 586200.0 ;
      RECT  1006800.0 600000.0 1017000.0 613800.0 ;
      RECT  1006800.0 627600.0 1017000.0 613800.0 ;
      RECT  1006800.0 627600.0 1017000.0 641400.0 ;
      RECT  1006800.0 655200.0 1017000.0 641400.0 ;
      RECT  1006800.0 655200.0 1017000.0 669000.0 ;
      RECT  1006800.0 682800.0 1017000.0 669000.0 ;
      RECT  1006800.0 682800.0 1017000.0 696600.0 ;
      RECT  1006800.0 710400.0 1017000.0 696600.0 ;
      RECT  1006800.0 710400.0 1017000.0 724200.0 ;
      RECT  1006800.0 738000.0 1017000.0 724200.0 ;
      RECT  1006800.0 738000.0 1017000.0 751800.0 ;
      RECT  1006800.0 765600.0 1017000.0 751800.0 ;
      RECT  1006800.0 765600.0 1017000.0 779400.0 ;
      RECT  1006800.0 793200.0 1017000.0 779400.0 ;
      RECT  1006800.0 793200.0 1017000.0 807000.0 ;
      RECT  1006800.0 820800.0 1017000.0 807000.0 ;
      RECT  1006800.0 820800.0 1017000.0 834600.0 ;
      RECT  1006800.0 848400.0 1017000.0 834600.0 ;
      RECT  1006800.0 848400.0 1017000.0 862200.0 ;
      RECT  1006800.0 876000.0 1017000.0 862200.0 ;
      RECT  1006800.0 876000.0 1017000.0 889800.0 ;
      RECT  1006800.0 903600.0 1017000.0 889800.0 ;
      RECT  1006800.0 903600.0 1017000.0 917400.0 ;
      RECT  1006800.0 931200.0 1017000.0 917400.0 ;
      RECT  1006800.0 931200.0 1017000.0 945000.0 ;
      RECT  1006800.0 958800.0 1017000.0 945000.0 ;
      RECT  1006800.0 958800.0 1017000.0 972600.0 ;
      RECT  1006800.0 986400.0 1017000.0 972600.0 ;
      RECT  1006800.0 986400.0 1017000.0 1000200.0 ;
      RECT  1006800.0 1014000.0 1017000.0 1000200.0 ;
      RECT  1006800.0 1014000.0 1017000.0 1027800.0 ;
      RECT  1006800.0 1041600.0 1017000.0 1027800.0 ;
      RECT  1006800.0 1041600.0 1017000.0 1055400.0 ;
      RECT  1006800.0 1069200.0 1017000.0 1055400.0 ;
      RECT  1006800.0 1069200.0 1017000.0 1083000.0 ;
      RECT  1006800.0 1096800.0 1017000.0 1083000.0 ;
      RECT  1006800.0 1096800.0 1017000.0 1110600.0 ;
      RECT  1006800.0 1124400.0 1017000.0 1110600.0 ;
      RECT  1006800.0 1124400.0 1017000.0 1138200.0 ;
      RECT  1006800.0 1152000.0 1017000.0 1138200.0 ;
      RECT  1006800.0 1152000.0 1017000.0 1165800.0 ;
      RECT  1006800.0 1179600.0 1017000.0 1165800.0 ;
      RECT  1006800.0 1179600.0 1017000.0 1193400.0 ;
      RECT  1006800.0 1207200.0 1017000.0 1193400.0 ;
      RECT  1006800.0 1207200.0 1017000.0 1221000.0 ;
      RECT  1006800.0 1234800.0 1017000.0 1221000.0 ;
      RECT  1006800.0 1234800.0 1017000.0 1248600.0 ;
      RECT  1006800.0 1262400.0 1017000.0 1248600.0 ;
      RECT  1006800.0 1262400.0 1017000.0 1276200.0 ;
      RECT  1006800.0 1290000.0 1017000.0 1276200.0 ;
      RECT  1006800.0 1290000.0 1017000.0 1303800.0 ;
      RECT  1006800.0 1317600.0 1017000.0 1303800.0 ;
      RECT  1006800.0 1317600.0 1017000.0 1331400.0 ;
      RECT  1006800.0 1345200.0 1017000.0 1331400.0 ;
      RECT  1006800.0 1345200.0 1017000.0 1359000.0 ;
      RECT  1006800.0 1372800.0 1017000.0 1359000.0 ;
      RECT  1006800.0 1372800.0 1017000.0 1386600.0 ;
      RECT  1006800.0 1400400.0 1017000.0 1386600.0 ;
      RECT  1006800.0 1400400.0 1017000.0 1414200.0 ;
      RECT  1006800.0 1428000.0 1017000.0 1414200.0 ;
      RECT  1006800.0 1428000.0 1017000.0 1441800.0 ;
      RECT  1006800.0 1455600.0 1017000.0 1441800.0 ;
      RECT  1006800.0 1455600.0 1017000.0 1469400.0 ;
      RECT  1006800.0 1483200.0 1017000.0 1469400.0 ;
      RECT  1006800.0 1483200.0 1017000.0 1497000.0 ;
      RECT  1006800.0 1510800.0 1017000.0 1497000.0 ;
      RECT  1006800.0 1510800.0 1017000.0 1524600.0 ;
      RECT  1006800.0 1538400.0 1017000.0 1524600.0 ;
      RECT  1006800.0 1538400.0 1017000.0 1552200.0 ;
      RECT  1006800.0 1566000.0 1017000.0 1552200.0 ;
      RECT  1006800.0 1566000.0 1017000.0 1579800.0 ;
      RECT  1006800.0 1593600.0 1017000.0 1579800.0 ;
      RECT  1006800.0 1593600.0 1017000.0 1607400.0 ;
      RECT  1006800.0 1621200.0 1017000.0 1607400.0 ;
      RECT  1006800.0 1621200.0 1017000.0 1635000.0 ;
      RECT  1006800.0 1648800.0 1017000.0 1635000.0 ;
      RECT  1006800.0 1648800.0 1017000.0 1662600.0 ;
      RECT  1006800.0 1676400.0 1017000.0 1662600.0 ;
      RECT  1006800.0 1676400.0 1017000.0 1690200.0 ;
      RECT  1006800.0 1704000.0 1017000.0 1690200.0 ;
      RECT  1006800.0 1704000.0 1017000.0 1717800.0 ;
      RECT  1006800.0 1731600.0 1017000.0 1717800.0 ;
      RECT  1006800.0 1731600.0 1017000.0 1745400.0 ;
      RECT  1006800.0 1759200.0 1017000.0 1745400.0 ;
      RECT  1006800.0 1759200.0 1017000.0 1773000.0 ;
      RECT  1006800.0 1786800.0 1017000.0 1773000.0 ;
      RECT  1006800.0 1786800.0 1017000.0 1800600.0 ;
      RECT  1006800.0 1814400.0 1017000.0 1800600.0 ;
      RECT  1006800.0 1814400.0 1017000.0 1828200.0 ;
      RECT  1006800.0 1842000.0 1017000.0 1828200.0 ;
      RECT  1006800.0 1842000.0 1017000.0 1855800.0 ;
      RECT  1006800.0 1869600.0 1017000.0 1855800.0 ;
      RECT  1006800.0 1869600.0 1017000.0 1883400.0 ;
      RECT  1006800.0 1897200.0 1017000.0 1883400.0 ;
      RECT  1006800.0 1897200.0 1017000.0 1911000.0 ;
      RECT  1006800.0 1924800.0 1017000.0 1911000.0 ;
      RECT  1006800.0 1924800.0 1017000.0 1938600.0 ;
      RECT  1006800.0 1952400.0 1017000.0 1938600.0 ;
      RECT  1006800.0 1952400.0 1017000.0 1966200.0 ;
      RECT  1006800.0 1980000.0 1017000.0 1966200.0 ;
      RECT  1006800.0 1980000.0 1017000.0 1993800.0 ;
      RECT  1006800.0 2007600.0 1017000.0 1993800.0 ;
      RECT  1006800.0 2007600.0 1017000.0 2021400.0 ;
      RECT  1006800.0 2035200.0 1017000.0 2021400.0 ;
      RECT  1006800.0 2035200.0 1017000.0 2049000.0 ;
      RECT  1006800.0 2062800.0 1017000.0 2049000.0 ;
      RECT  1006800.0 2062800.0 1017000.0 2076600.0 ;
      RECT  1006800.0 2090400.0 1017000.0 2076600.0 ;
      RECT  1006800.0 2090400.0 1017000.0 2104200.0 ;
      RECT  1006800.0 2118000.0 1017000.0 2104200.0 ;
      RECT  1006800.0 2118000.0 1017000.0 2131800.0 ;
      RECT  1006800.0 2145600.0 1017000.0 2131800.0 ;
      RECT  1017000.0 379200.0 1027200.0 393000.0 ;
      RECT  1017000.0 406800.0 1027200.0 393000.0 ;
      RECT  1017000.0 406800.0 1027200.0 420600.0 ;
      RECT  1017000.0 434400.0 1027200.0 420600.0 ;
      RECT  1017000.0 434400.0 1027200.0 448200.0 ;
      RECT  1017000.0 462000.0 1027200.0 448200.0 ;
      RECT  1017000.0 462000.0 1027200.0 475800.0 ;
      RECT  1017000.0 489600.0 1027200.0 475800.0 ;
      RECT  1017000.0 489600.0 1027200.0 503400.0 ;
      RECT  1017000.0 517200.0 1027200.0 503400.0 ;
      RECT  1017000.0 517200.0 1027200.0 531000.0 ;
      RECT  1017000.0 544800.0 1027200.0 531000.0 ;
      RECT  1017000.0 544800.0 1027200.0 558600.0 ;
      RECT  1017000.0 572400.0 1027200.0 558600.0 ;
      RECT  1017000.0 572400.0 1027200.0 586200.0 ;
      RECT  1017000.0 600000.0 1027200.0 586200.0 ;
      RECT  1017000.0 600000.0 1027200.0 613800.0 ;
      RECT  1017000.0 627600.0 1027200.0 613800.0 ;
      RECT  1017000.0 627600.0 1027200.0 641400.0 ;
      RECT  1017000.0 655200.0 1027200.0 641400.0 ;
      RECT  1017000.0 655200.0 1027200.0 669000.0 ;
      RECT  1017000.0 682800.0 1027200.0 669000.0 ;
      RECT  1017000.0 682800.0 1027200.0 696600.0 ;
      RECT  1017000.0 710400.0 1027200.0 696600.0 ;
      RECT  1017000.0 710400.0 1027200.0 724200.0 ;
      RECT  1017000.0 738000.0 1027200.0 724200.0 ;
      RECT  1017000.0 738000.0 1027200.0 751800.0 ;
      RECT  1017000.0 765600.0 1027200.0 751800.0 ;
      RECT  1017000.0 765600.0 1027200.0 779400.0 ;
      RECT  1017000.0 793200.0 1027200.0 779400.0 ;
      RECT  1017000.0 793200.0 1027200.0 807000.0 ;
      RECT  1017000.0 820800.0 1027200.0 807000.0 ;
      RECT  1017000.0 820800.0 1027200.0 834600.0 ;
      RECT  1017000.0 848400.0 1027200.0 834600.0 ;
      RECT  1017000.0 848400.0 1027200.0 862200.0 ;
      RECT  1017000.0 876000.0 1027200.0 862200.0 ;
      RECT  1017000.0 876000.0 1027200.0 889800.0 ;
      RECT  1017000.0 903600.0 1027200.0 889800.0 ;
      RECT  1017000.0 903600.0 1027200.0 917400.0 ;
      RECT  1017000.0 931200.0 1027200.0 917400.0 ;
      RECT  1017000.0 931200.0 1027200.0 945000.0 ;
      RECT  1017000.0 958800.0 1027200.0 945000.0 ;
      RECT  1017000.0 958800.0 1027200.0 972600.0 ;
      RECT  1017000.0 986400.0 1027200.0 972600.0 ;
      RECT  1017000.0 986400.0 1027200.0 1000200.0 ;
      RECT  1017000.0 1014000.0 1027200.0 1000200.0 ;
      RECT  1017000.0 1014000.0 1027200.0 1027800.0 ;
      RECT  1017000.0 1041600.0 1027200.0 1027800.0 ;
      RECT  1017000.0 1041600.0 1027200.0 1055400.0 ;
      RECT  1017000.0 1069200.0 1027200.0 1055400.0 ;
      RECT  1017000.0 1069200.0 1027200.0 1083000.0 ;
      RECT  1017000.0 1096800.0 1027200.0 1083000.0 ;
      RECT  1017000.0 1096800.0 1027200.0 1110600.0 ;
      RECT  1017000.0 1124400.0 1027200.0 1110600.0 ;
      RECT  1017000.0 1124400.0 1027200.0 1138200.0 ;
      RECT  1017000.0 1152000.0 1027200.0 1138200.0 ;
      RECT  1017000.0 1152000.0 1027200.0 1165800.0 ;
      RECT  1017000.0 1179600.0 1027200.0 1165800.0 ;
      RECT  1017000.0 1179600.0 1027200.0 1193400.0 ;
      RECT  1017000.0 1207200.0 1027200.0 1193400.0 ;
      RECT  1017000.0 1207200.0 1027200.0 1221000.0 ;
      RECT  1017000.0 1234800.0 1027200.0 1221000.0 ;
      RECT  1017000.0 1234800.0 1027200.0 1248600.0 ;
      RECT  1017000.0 1262400.0 1027200.0 1248600.0 ;
      RECT  1017000.0 1262400.0 1027200.0 1276200.0 ;
      RECT  1017000.0 1290000.0 1027200.0 1276200.0 ;
      RECT  1017000.0 1290000.0 1027200.0 1303800.0 ;
      RECT  1017000.0 1317600.0 1027200.0 1303800.0 ;
      RECT  1017000.0 1317600.0 1027200.0 1331400.0 ;
      RECT  1017000.0 1345200.0 1027200.0 1331400.0 ;
      RECT  1017000.0 1345200.0 1027200.0 1359000.0 ;
      RECT  1017000.0 1372800.0 1027200.0 1359000.0 ;
      RECT  1017000.0 1372800.0 1027200.0 1386600.0 ;
      RECT  1017000.0 1400400.0 1027200.0 1386600.0 ;
      RECT  1017000.0 1400400.0 1027200.0 1414200.0 ;
      RECT  1017000.0 1428000.0 1027200.0 1414200.0 ;
      RECT  1017000.0 1428000.0 1027200.0 1441800.0 ;
      RECT  1017000.0 1455600.0 1027200.0 1441800.0 ;
      RECT  1017000.0 1455600.0 1027200.0 1469400.0 ;
      RECT  1017000.0 1483200.0 1027200.0 1469400.0 ;
      RECT  1017000.0 1483200.0 1027200.0 1497000.0 ;
      RECT  1017000.0 1510800.0 1027200.0 1497000.0 ;
      RECT  1017000.0 1510800.0 1027200.0 1524600.0 ;
      RECT  1017000.0 1538400.0 1027200.0 1524600.0 ;
      RECT  1017000.0 1538400.0 1027200.0 1552200.0 ;
      RECT  1017000.0 1566000.0 1027200.0 1552200.0 ;
      RECT  1017000.0 1566000.0 1027200.0 1579800.0 ;
      RECT  1017000.0 1593600.0 1027200.0 1579800.0 ;
      RECT  1017000.0 1593600.0 1027200.0 1607400.0 ;
      RECT  1017000.0 1621200.0 1027200.0 1607400.0 ;
      RECT  1017000.0 1621200.0 1027200.0 1635000.0 ;
      RECT  1017000.0 1648800.0 1027200.0 1635000.0 ;
      RECT  1017000.0 1648800.0 1027200.0 1662600.0 ;
      RECT  1017000.0 1676400.0 1027200.0 1662600.0 ;
      RECT  1017000.0 1676400.0 1027200.0 1690200.0 ;
      RECT  1017000.0 1704000.0 1027200.0 1690200.0 ;
      RECT  1017000.0 1704000.0 1027200.0 1717800.0 ;
      RECT  1017000.0 1731600.0 1027200.0 1717800.0 ;
      RECT  1017000.0 1731600.0 1027200.0 1745400.0 ;
      RECT  1017000.0 1759200.0 1027200.0 1745400.0 ;
      RECT  1017000.0 1759200.0 1027200.0 1773000.0 ;
      RECT  1017000.0 1786800.0 1027200.0 1773000.0 ;
      RECT  1017000.0 1786800.0 1027200.0 1800600.0 ;
      RECT  1017000.0 1814400.0 1027200.0 1800600.0 ;
      RECT  1017000.0 1814400.0 1027200.0 1828200.0 ;
      RECT  1017000.0 1842000.0 1027200.0 1828200.0 ;
      RECT  1017000.0 1842000.0 1027200.0 1855800.0 ;
      RECT  1017000.0 1869600.0 1027200.0 1855800.0 ;
      RECT  1017000.0 1869600.0 1027200.0 1883400.0 ;
      RECT  1017000.0 1897200.0 1027200.0 1883400.0 ;
      RECT  1017000.0 1897200.0 1027200.0 1911000.0 ;
      RECT  1017000.0 1924800.0 1027200.0 1911000.0 ;
      RECT  1017000.0 1924800.0 1027200.0 1938600.0 ;
      RECT  1017000.0 1952400.0 1027200.0 1938600.0 ;
      RECT  1017000.0 1952400.0 1027200.0 1966200.0 ;
      RECT  1017000.0 1980000.0 1027200.0 1966200.0 ;
      RECT  1017000.0 1980000.0 1027200.0 1993800.0 ;
      RECT  1017000.0 2007600.0 1027200.0 1993800.0 ;
      RECT  1017000.0 2007600.0 1027200.0 2021400.0 ;
      RECT  1017000.0 2035200.0 1027200.0 2021400.0 ;
      RECT  1017000.0 2035200.0 1027200.0 2049000.0 ;
      RECT  1017000.0 2062800.0 1027200.0 2049000.0 ;
      RECT  1017000.0 2062800.0 1027200.0 2076600.0 ;
      RECT  1017000.0 2090400.0 1027200.0 2076600.0 ;
      RECT  1017000.0 2090400.0 1027200.0 2104200.0 ;
      RECT  1017000.0 2118000.0 1027200.0 2104200.0 ;
      RECT  1017000.0 2118000.0 1027200.0 2131800.0 ;
      RECT  1017000.0 2145600.0 1027200.0 2131800.0 ;
      RECT  1027200.0 379200.0 1037400.0 393000.0 ;
      RECT  1027200.0 406800.0 1037400.0 393000.0 ;
      RECT  1027200.0 406800.0 1037400.0 420600.0 ;
      RECT  1027200.0 434400.0 1037400.0 420600.0 ;
      RECT  1027200.0 434400.0 1037400.0 448200.0 ;
      RECT  1027200.0 462000.0 1037400.0 448200.0 ;
      RECT  1027200.0 462000.0 1037400.0 475800.0 ;
      RECT  1027200.0 489600.0 1037400.0 475800.0 ;
      RECT  1027200.0 489600.0 1037400.0 503400.0 ;
      RECT  1027200.0 517200.0 1037400.0 503400.0 ;
      RECT  1027200.0 517200.0 1037400.0 531000.0 ;
      RECT  1027200.0 544800.0 1037400.0 531000.0 ;
      RECT  1027200.0 544800.0 1037400.0 558600.0 ;
      RECT  1027200.0 572400.0 1037400.0 558600.0 ;
      RECT  1027200.0 572400.0 1037400.0 586200.0 ;
      RECT  1027200.0 600000.0 1037400.0 586200.0 ;
      RECT  1027200.0 600000.0 1037400.0 613800.0 ;
      RECT  1027200.0 627600.0 1037400.0 613800.0 ;
      RECT  1027200.0 627600.0 1037400.0 641400.0 ;
      RECT  1027200.0 655200.0 1037400.0 641400.0 ;
      RECT  1027200.0 655200.0 1037400.0 669000.0 ;
      RECT  1027200.0 682800.0 1037400.0 669000.0 ;
      RECT  1027200.0 682800.0 1037400.0 696600.0 ;
      RECT  1027200.0 710400.0 1037400.0 696600.0 ;
      RECT  1027200.0 710400.0 1037400.0 724200.0 ;
      RECT  1027200.0 738000.0 1037400.0 724200.0 ;
      RECT  1027200.0 738000.0 1037400.0 751800.0 ;
      RECT  1027200.0 765600.0 1037400.0 751800.0 ;
      RECT  1027200.0 765600.0 1037400.0 779400.0 ;
      RECT  1027200.0 793200.0 1037400.0 779400.0 ;
      RECT  1027200.0 793200.0 1037400.0 807000.0 ;
      RECT  1027200.0 820800.0 1037400.0 807000.0 ;
      RECT  1027200.0 820800.0 1037400.0 834600.0 ;
      RECT  1027200.0 848400.0 1037400.0 834600.0 ;
      RECT  1027200.0 848400.0 1037400.0 862200.0 ;
      RECT  1027200.0 876000.0 1037400.0 862200.0 ;
      RECT  1027200.0 876000.0 1037400.0 889800.0 ;
      RECT  1027200.0 903600.0 1037400.0 889800.0 ;
      RECT  1027200.0 903600.0 1037400.0 917400.0 ;
      RECT  1027200.0 931200.0 1037400.0 917400.0 ;
      RECT  1027200.0 931200.0 1037400.0 945000.0 ;
      RECT  1027200.0 958800.0 1037400.0 945000.0 ;
      RECT  1027200.0 958800.0 1037400.0 972600.0 ;
      RECT  1027200.0 986400.0 1037400.0 972600.0 ;
      RECT  1027200.0 986400.0 1037400.0 1000200.0 ;
      RECT  1027200.0 1014000.0 1037400.0 1000200.0 ;
      RECT  1027200.0 1014000.0 1037400.0 1027800.0 ;
      RECT  1027200.0 1041600.0 1037400.0 1027800.0 ;
      RECT  1027200.0 1041600.0 1037400.0 1055400.0 ;
      RECT  1027200.0 1069200.0 1037400.0 1055400.0 ;
      RECT  1027200.0 1069200.0 1037400.0 1083000.0 ;
      RECT  1027200.0 1096800.0 1037400.0 1083000.0 ;
      RECT  1027200.0 1096800.0 1037400.0 1110600.0 ;
      RECT  1027200.0 1124400.0 1037400.0 1110600.0 ;
      RECT  1027200.0 1124400.0 1037400.0 1138200.0 ;
      RECT  1027200.0 1152000.0 1037400.0 1138200.0 ;
      RECT  1027200.0 1152000.0 1037400.0 1165800.0 ;
      RECT  1027200.0 1179600.0 1037400.0 1165800.0 ;
      RECT  1027200.0 1179600.0 1037400.0 1193400.0 ;
      RECT  1027200.0 1207200.0 1037400.0 1193400.0 ;
      RECT  1027200.0 1207200.0 1037400.0 1221000.0 ;
      RECT  1027200.0 1234800.0 1037400.0 1221000.0 ;
      RECT  1027200.0 1234800.0 1037400.0 1248600.0 ;
      RECT  1027200.0 1262400.0 1037400.0 1248600.0 ;
      RECT  1027200.0 1262400.0 1037400.0 1276200.0 ;
      RECT  1027200.0 1290000.0 1037400.0 1276200.0 ;
      RECT  1027200.0 1290000.0 1037400.0 1303800.0 ;
      RECT  1027200.0 1317600.0 1037400.0 1303800.0 ;
      RECT  1027200.0 1317600.0 1037400.0 1331400.0 ;
      RECT  1027200.0 1345200.0 1037400.0 1331400.0 ;
      RECT  1027200.0 1345200.0 1037400.0 1359000.0 ;
      RECT  1027200.0 1372800.0 1037400.0 1359000.0 ;
      RECT  1027200.0 1372800.0 1037400.0 1386600.0 ;
      RECT  1027200.0 1400400.0 1037400.0 1386600.0 ;
      RECT  1027200.0 1400400.0 1037400.0 1414200.0 ;
      RECT  1027200.0 1428000.0 1037400.0 1414200.0 ;
      RECT  1027200.0 1428000.0 1037400.0 1441800.0 ;
      RECT  1027200.0 1455600.0 1037400.0 1441800.0 ;
      RECT  1027200.0 1455600.0 1037400.0 1469400.0 ;
      RECT  1027200.0 1483200.0 1037400.0 1469400.0 ;
      RECT  1027200.0 1483200.0 1037400.0 1497000.0 ;
      RECT  1027200.0 1510800.0 1037400.0 1497000.0 ;
      RECT  1027200.0 1510800.0 1037400.0 1524600.0 ;
      RECT  1027200.0 1538400.0 1037400.0 1524600.0 ;
      RECT  1027200.0 1538400.0 1037400.0 1552200.0 ;
      RECT  1027200.0 1566000.0 1037400.0 1552200.0 ;
      RECT  1027200.0 1566000.0 1037400.0 1579800.0 ;
      RECT  1027200.0 1593600.0 1037400.0 1579800.0 ;
      RECT  1027200.0 1593600.0 1037400.0 1607400.0 ;
      RECT  1027200.0 1621200.0 1037400.0 1607400.0 ;
      RECT  1027200.0 1621200.0 1037400.0 1635000.0 ;
      RECT  1027200.0 1648800.0 1037400.0 1635000.0 ;
      RECT  1027200.0 1648800.0 1037400.0 1662600.0 ;
      RECT  1027200.0 1676400.0 1037400.0 1662600.0 ;
      RECT  1027200.0 1676400.0 1037400.0 1690200.0 ;
      RECT  1027200.0 1704000.0 1037400.0 1690200.0 ;
      RECT  1027200.0 1704000.0 1037400.0 1717800.0 ;
      RECT  1027200.0 1731600.0 1037400.0 1717800.0 ;
      RECT  1027200.0 1731600.0 1037400.0 1745400.0 ;
      RECT  1027200.0 1759200.0 1037400.0 1745400.0 ;
      RECT  1027200.0 1759200.0 1037400.0 1773000.0 ;
      RECT  1027200.0 1786800.0 1037400.0 1773000.0 ;
      RECT  1027200.0 1786800.0 1037400.0 1800600.0 ;
      RECT  1027200.0 1814400.0 1037400.0 1800600.0 ;
      RECT  1027200.0 1814400.0 1037400.0 1828200.0 ;
      RECT  1027200.0 1842000.0 1037400.0 1828200.0 ;
      RECT  1027200.0 1842000.0 1037400.0 1855800.0 ;
      RECT  1027200.0 1869600.0 1037400.0 1855800.0 ;
      RECT  1027200.0 1869600.0 1037400.0 1883400.0 ;
      RECT  1027200.0 1897200.0 1037400.0 1883400.0 ;
      RECT  1027200.0 1897200.0 1037400.0 1911000.0 ;
      RECT  1027200.0 1924800.0 1037400.0 1911000.0 ;
      RECT  1027200.0 1924800.0 1037400.0 1938600.0 ;
      RECT  1027200.0 1952400.0 1037400.0 1938600.0 ;
      RECT  1027200.0 1952400.0 1037400.0 1966200.0 ;
      RECT  1027200.0 1980000.0 1037400.0 1966200.0 ;
      RECT  1027200.0 1980000.0 1037400.0 1993800.0 ;
      RECT  1027200.0 2007600.0 1037400.0 1993800.0 ;
      RECT  1027200.0 2007600.0 1037400.0 2021400.0 ;
      RECT  1027200.0 2035200.0 1037400.0 2021400.0 ;
      RECT  1027200.0 2035200.0 1037400.0 2049000.0 ;
      RECT  1027200.0 2062800.0 1037400.0 2049000.0 ;
      RECT  1027200.0 2062800.0 1037400.0 2076600.0 ;
      RECT  1027200.0 2090400.0 1037400.0 2076600.0 ;
      RECT  1027200.0 2090400.0 1037400.0 2104200.0 ;
      RECT  1027200.0 2118000.0 1037400.0 2104200.0 ;
      RECT  1027200.0 2118000.0 1037400.0 2131800.0 ;
      RECT  1027200.0 2145600.0 1037400.0 2131800.0 ;
      RECT  1037400.0 379200.0 1047600.0 393000.0 ;
      RECT  1037400.0 406800.0 1047600.0 393000.0 ;
      RECT  1037400.0 406800.0 1047600.0 420600.0 ;
      RECT  1037400.0 434400.0 1047600.0 420600.0 ;
      RECT  1037400.0 434400.0 1047600.0 448200.0 ;
      RECT  1037400.0 462000.0 1047600.0 448200.0 ;
      RECT  1037400.0 462000.0 1047600.0 475800.0 ;
      RECT  1037400.0 489600.0 1047600.0 475800.0 ;
      RECT  1037400.0 489600.0 1047600.0 503400.0 ;
      RECT  1037400.0 517200.0 1047600.0 503400.0 ;
      RECT  1037400.0 517200.0 1047600.0 531000.0 ;
      RECT  1037400.0 544800.0 1047600.0 531000.0 ;
      RECT  1037400.0 544800.0 1047600.0 558600.0 ;
      RECT  1037400.0 572400.0 1047600.0 558600.0 ;
      RECT  1037400.0 572400.0 1047600.0 586200.0 ;
      RECT  1037400.0 600000.0 1047600.0 586200.0 ;
      RECT  1037400.0 600000.0 1047600.0 613800.0 ;
      RECT  1037400.0 627600.0 1047600.0 613800.0 ;
      RECT  1037400.0 627600.0 1047600.0 641400.0 ;
      RECT  1037400.0 655200.0 1047600.0 641400.0 ;
      RECT  1037400.0 655200.0 1047600.0 669000.0 ;
      RECT  1037400.0 682800.0 1047600.0 669000.0 ;
      RECT  1037400.0 682800.0 1047600.0 696600.0 ;
      RECT  1037400.0 710400.0 1047600.0 696600.0 ;
      RECT  1037400.0 710400.0 1047600.0 724200.0 ;
      RECT  1037400.0 738000.0 1047600.0 724200.0 ;
      RECT  1037400.0 738000.0 1047600.0 751800.0 ;
      RECT  1037400.0 765600.0 1047600.0 751800.0 ;
      RECT  1037400.0 765600.0 1047600.0 779400.0 ;
      RECT  1037400.0 793200.0 1047600.0 779400.0 ;
      RECT  1037400.0 793200.0 1047600.0 807000.0 ;
      RECT  1037400.0 820800.0 1047600.0 807000.0 ;
      RECT  1037400.0 820800.0 1047600.0 834600.0 ;
      RECT  1037400.0 848400.0 1047600.0 834600.0 ;
      RECT  1037400.0 848400.0 1047600.0 862200.0 ;
      RECT  1037400.0 876000.0 1047600.0 862200.0 ;
      RECT  1037400.0 876000.0 1047600.0 889800.0 ;
      RECT  1037400.0 903600.0 1047600.0 889800.0 ;
      RECT  1037400.0 903600.0 1047600.0 917400.0 ;
      RECT  1037400.0 931200.0 1047600.0 917400.0 ;
      RECT  1037400.0 931200.0 1047600.0 945000.0 ;
      RECT  1037400.0 958800.0 1047600.0 945000.0 ;
      RECT  1037400.0 958800.0 1047600.0 972600.0 ;
      RECT  1037400.0 986400.0 1047600.0 972600.0 ;
      RECT  1037400.0 986400.0 1047600.0 1000200.0 ;
      RECT  1037400.0 1014000.0 1047600.0 1000200.0 ;
      RECT  1037400.0 1014000.0 1047600.0 1027800.0 ;
      RECT  1037400.0 1041600.0 1047600.0 1027800.0 ;
      RECT  1037400.0 1041600.0 1047600.0 1055400.0 ;
      RECT  1037400.0 1069200.0 1047600.0 1055400.0 ;
      RECT  1037400.0 1069200.0 1047600.0 1083000.0 ;
      RECT  1037400.0 1096800.0 1047600.0 1083000.0 ;
      RECT  1037400.0 1096800.0 1047600.0 1110600.0 ;
      RECT  1037400.0 1124400.0 1047600.0 1110600.0 ;
      RECT  1037400.0 1124400.0 1047600.0 1138200.0 ;
      RECT  1037400.0 1152000.0 1047600.0 1138200.0 ;
      RECT  1037400.0 1152000.0 1047600.0 1165800.0 ;
      RECT  1037400.0 1179600.0 1047600.0 1165800.0 ;
      RECT  1037400.0 1179600.0 1047600.0 1193400.0 ;
      RECT  1037400.0 1207200.0 1047600.0 1193400.0 ;
      RECT  1037400.0 1207200.0 1047600.0 1221000.0 ;
      RECT  1037400.0 1234800.0 1047600.0 1221000.0 ;
      RECT  1037400.0 1234800.0 1047600.0 1248600.0 ;
      RECT  1037400.0 1262400.0 1047600.0 1248600.0 ;
      RECT  1037400.0 1262400.0 1047600.0 1276200.0 ;
      RECT  1037400.0 1290000.0 1047600.0 1276200.0 ;
      RECT  1037400.0 1290000.0 1047600.0 1303800.0 ;
      RECT  1037400.0 1317600.0 1047600.0 1303800.0 ;
      RECT  1037400.0 1317600.0 1047600.0 1331400.0 ;
      RECT  1037400.0 1345200.0 1047600.0 1331400.0 ;
      RECT  1037400.0 1345200.0 1047600.0 1359000.0 ;
      RECT  1037400.0 1372800.0 1047600.0 1359000.0 ;
      RECT  1037400.0 1372800.0 1047600.0 1386600.0 ;
      RECT  1037400.0 1400400.0 1047600.0 1386600.0 ;
      RECT  1037400.0 1400400.0 1047600.0 1414200.0 ;
      RECT  1037400.0 1428000.0 1047600.0 1414200.0 ;
      RECT  1037400.0 1428000.0 1047600.0 1441800.0 ;
      RECT  1037400.0 1455600.0 1047600.0 1441800.0 ;
      RECT  1037400.0 1455600.0 1047600.0 1469400.0 ;
      RECT  1037400.0 1483200.0 1047600.0 1469400.0 ;
      RECT  1037400.0 1483200.0 1047600.0 1497000.0 ;
      RECT  1037400.0 1510800.0 1047600.0 1497000.0 ;
      RECT  1037400.0 1510800.0 1047600.0 1524600.0 ;
      RECT  1037400.0 1538400.0 1047600.0 1524600.0 ;
      RECT  1037400.0 1538400.0 1047600.0 1552200.0 ;
      RECT  1037400.0 1566000.0 1047600.0 1552200.0 ;
      RECT  1037400.0 1566000.0 1047600.0 1579800.0 ;
      RECT  1037400.0 1593600.0 1047600.0 1579800.0 ;
      RECT  1037400.0 1593600.0 1047600.0 1607400.0 ;
      RECT  1037400.0 1621200.0 1047600.0 1607400.0 ;
      RECT  1037400.0 1621200.0 1047600.0 1635000.0 ;
      RECT  1037400.0 1648800.0 1047600.0 1635000.0 ;
      RECT  1037400.0 1648800.0 1047600.0 1662600.0 ;
      RECT  1037400.0 1676400.0 1047600.0 1662600.0 ;
      RECT  1037400.0 1676400.0 1047600.0 1690200.0 ;
      RECT  1037400.0 1704000.0 1047600.0 1690200.0 ;
      RECT  1037400.0 1704000.0 1047600.0 1717800.0 ;
      RECT  1037400.0 1731600.0 1047600.0 1717800.0 ;
      RECT  1037400.0 1731600.0 1047600.0 1745400.0 ;
      RECT  1037400.0 1759200.0 1047600.0 1745400.0 ;
      RECT  1037400.0 1759200.0 1047600.0 1773000.0 ;
      RECT  1037400.0 1786800.0 1047600.0 1773000.0 ;
      RECT  1037400.0 1786800.0 1047600.0 1800600.0 ;
      RECT  1037400.0 1814400.0 1047600.0 1800600.0 ;
      RECT  1037400.0 1814400.0 1047600.0 1828200.0 ;
      RECT  1037400.0 1842000.0 1047600.0 1828200.0 ;
      RECT  1037400.0 1842000.0 1047600.0 1855800.0 ;
      RECT  1037400.0 1869600.0 1047600.0 1855800.0 ;
      RECT  1037400.0 1869600.0 1047600.0 1883400.0 ;
      RECT  1037400.0 1897200.0 1047600.0 1883400.0 ;
      RECT  1037400.0 1897200.0 1047600.0 1911000.0 ;
      RECT  1037400.0 1924800.0 1047600.0 1911000.0 ;
      RECT  1037400.0 1924800.0 1047600.0 1938600.0 ;
      RECT  1037400.0 1952400.0 1047600.0 1938600.0 ;
      RECT  1037400.0 1952400.0 1047600.0 1966200.0 ;
      RECT  1037400.0 1980000.0 1047600.0 1966200.0 ;
      RECT  1037400.0 1980000.0 1047600.0 1993800.0 ;
      RECT  1037400.0 2007600.0 1047600.0 1993800.0 ;
      RECT  1037400.0 2007600.0 1047600.0 2021400.0 ;
      RECT  1037400.0 2035200.0 1047600.0 2021400.0 ;
      RECT  1037400.0 2035200.0 1047600.0 2049000.0 ;
      RECT  1037400.0 2062800.0 1047600.0 2049000.0 ;
      RECT  1037400.0 2062800.0 1047600.0 2076600.0 ;
      RECT  1037400.0 2090400.0 1047600.0 2076600.0 ;
      RECT  1037400.0 2090400.0 1047600.0 2104200.0 ;
      RECT  1037400.0 2118000.0 1047600.0 2104200.0 ;
      RECT  1037400.0 2118000.0 1047600.0 2131800.0 ;
      RECT  1037400.0 2145600.0 1047600.0 2131800.0 ;
      RECT  1047600.0 379200.0 1057800.0 393000.0 ;
      RECT  1047600.0 406800.0 1057800.0 393000.0 ;
      RECT  1047600.0 406800.0 1057800.0 420600.0 ;
      RECT  1047600.0 434400.0 1057800.0 420600.0 ;
      RECT  1047600.0 434400.0 1057800.0 448200.0 ;
      RECT  1047600.0 462000.0 1057800.0 448200.0 ;
      RECT  1047600.0 462000.0 1057800.0 475800.0 ;
      RECT  1047600.0 489600.0 1057800.0 475800.0 ;
      RECT  1047600.0 489600.0 1057800.0 503400.0 ;
      RECT  1047600.0 517200.0 1057800.0 503400.0 ;
      RECT  1047600.0 517200.0 1057800.0 531000.0 ;
      RECT  1047600.0 544800.0 1057800.0 531000.0 ;
      RECT  1047600.0 544800.0 1057800.0 558600.0 ;
      RECT  1047600.0 572400.0 1057800.0 558600.0 ;
      RECT  1047600.0 572400.0 1057800.0 586200.0 ;
      RECT  1047600.0 600000.0 1057800.0 586200.0 ;
      RECT  1047600.0 600000.0 1057800.0 613800.0 ;
      RECT  1047600.0 627600.0 1057800.0 613800.0 ;
      RECT  1047600.0 627600.0 1057800.0 641400.0 ;
      RECT  1047600.0 655200.0 1057800.0 641400.0 ;
      RECT  1047600.0 655200.0 1057800.0 669000.0 ;
      RECT  1047600.0 682800.0 1057800.0 669000.0 ;
      RECT  1047600.0 682800.0 1057800.0 696600.0 ;
      RECT  1047600.0 710400.0 1057800.0 696600.0 ;
      RECT  1047600.0 710400.0 1057800.0 724200.0 ;
      RECT  1047600.0 738000.0 1057800.0 724200.0 ;
      RECT  1047600.0 738000.0 1057800.0 751800.0 ;
      RECT  1047600.0 765600.0 1057800.0 751800.0 ;
      RECT  1047600.0 765600.0 1057800.0 779400.0 ;
      RECT  1047600.0 793200.0 1057800.0 779400.0 ;
      RECT  1047600.0 793200.0 1057800.0 807000.0 ;
      RECT  1047600.0 820800.0 1057800.0 807000.0 ;
      RECT  1047600.0 820800.0 1057800.0 834600.0 ;
      RECT  1047600.0 848400.0 1057800.0 834600.0 ;
      RECT  1047600.0 848400.0 1057800.0 862200.0 ;
      RECT  1047600.0 876000.0 1057800.0 862200.0 ;
      RECT  1047600.0 876000.0 1057800.0 889800.0 ;
      RECT  1047600.0 903600.0 1057800.0 889800.0 ;
      RECT  1047600.0 903600.0 1057800.0 917400.0 ;
      RECT  1047600.0 931200.0 1057800.0 917400.0 ;
      RECT  1047600.0 931200.0 1057800.0 945000.0 ;
      RECT  1047600.0 958800.0 1057800.0 945000.0 ;
      RECT  1047600.0 958800.0 1057800.0 972600.0 ;
      RECT  1047600.0 986400.0 1057800.0 972600.0 ;
      RECT  1047600.0 986400.0 1057800.0 1000200.0 ;
      RECT  1047600.0 1014000.0 1057800.0 1000200.0 ;
      RECT  1047600.0 1014000.0 1057800.0 1027800.0 ;
      RECT  1047600.0 1041600.0 1057800.0 1027800.0 ;
      RECT  1047600.0 1041600.0 1057800.0 1055400.0 ;
      RECT  1047600.0 1069200.0 1057800.0 1055400.0 ;
      RECT  1047600.0 1069200.0 1057800.0 1083000.0 ;
      RECT  1047600.0 1096800.0 1057800.0 1083000.0 ;
      RECT  1047600.0 1096800.0 1057800.0 1110600.0 ;
      RECT  1047600.0 1124400.0 1057800.0 1110600.0 ;
      RECT  1047600.0 1124400.0 1057800.0 1138200.0 ;
      RECT  1047600.0 1152000.0 1057800.0 1138200.0 ;
      RECT  1047600.0 1152000.0 1057800.0 1165800.0 ;
      RECT  1047600.0 1179600.0 1057800.0 1165800.0 ;
      RECT  1047600.0 1179600.0 1057800.0 1193400.0 ;
      RECT  1047600.0 1207200.0 1057800.0 1193400.0 ;
      RECT  1047600.0 1207200.0 1057800.0 1221000.0 ;
      RECT  1047600.0 1234800.0 1057800.0 1221000.0 ;
      RECT  1047600.0 1234800.0 1057800.0 1248600.0 ;
      RECT  1047600.0 1262400.0 1057800.0 1248600.0 ;
      RECT  1047600.0 1262400.0 1057800.0 1276200.0 ;
      RECT  1047600.0 1290000.0 1057800.0 1276200.0 ;
      RECT  1047600.0 1290000.0 1057800.0 1303800.0 ;
      RECT  1047600.0 1317600.0 1057800.0 1303800.0 ;
      RECT  1047600.0 1317600.0 1057800.0 1331400.0 ;
      RECT  1047600.0 1345200.0 1057800.0 1331400.0 ;
      RECT  1047600.0 1345200.0 1057800.0 1359000.0 ;
      RECT  1047600.0 1372800.0 1057800.0 1359000.0 ;
      RECT  1047600.0 1372800.0 1057800.0 1386600.0 ;
      RECT  1047600.0 1400400.0 1057800.0 1386600.0 ;
      RECT  1047600.0 1400400.0 1057800.0 1414200.0 ;
      RECT  1047600.0 1428000.0 1057800.0 1414200.0 ;
      RECT  1047600.0 1428000.0 1057800.0 1441800.0 ;
      RECT  1047600.0 1455600.0 1057800.0 1441800.0 ;
      RECT  1047600.0 1455600.0 1057800.0 1469400.0 ;
      RECT  1047600.0 1483200.0 1057800.0 1469400.0 ;
      RECT  1047600.0 1483200.0 1057800.0 1497000.0 ;
      RECT  1047600.0 1510800.0 1057800.0 1497000.0 ;
      RECT  1047600.0 1510800.0 1057800.0 1524600.0 ;
      RECT  1047600.0 1538400.0 1057800.0 1524600.0 ;
      RECT  1047600.0 1538400.0 1057800.0 1552200.0 ;
      RECT  1047600.0 1566000.0 1057800.0 1552200.0 ;
      RECT  1047600.0 1566000.0 1057800.0 1579800.0 ;
      RECT  1047600.0 1593600.0 1057800.0 1579800.0 ;
      RECT  1047600.0 1593600.0 1057800.0 1607400.0 ;
      RECT  1047600.0 1621200.0 1057800.0 1607400.0 ;
      RECT  1047600.0 1621200.0 1057800.0 1635000.0 ;
      RECT  1047600.0 1648800.0 1057800.0 1635000.0 ;
      RECT  1047600.0 1648800.0 1057800.0 1662600.0 ;
      RECT  1047600.0 1676400.0 1057800.0 1662600.0 ;
      RECT  1047600.0 1676400.0 1057800.0 1690200.0 ;
      RECT  1047600.0 1704000.0 1057800.0 1690200.0 ;
      RECT  1047600.0 1704000.0 1057800.0 1717800.0 ;
      RECT  1047600.0 1731600.0 1057800.0 1717800.0 ;
      RECT  1047600.0 1731600.0 1057800.0 1745400.0 ;
      RECT  1047600.0 1759200.0 1057800.0 1745400.0 ;
      RECT  1047600.0 1759200.0 1057800.0 1773000.0 ;
      RECT  1047600.0 1786800.0 1057800.0 1773000.0 ;
      RECT  1047600.0 1786800.0 1057800.0 1800600.0 ;
      RECT  1047600.0 1814400.0 1057800.0 1800600.0 ;
      RECT  1047600.0 1814400.0 1057800.0 1828200.0 ;
      RECT  1047600.0 1842000.0 1057800.0 1828200.0 ;
      RECT  1047600.0 1842000.0 1057800.0 1855800.0 ;
      RECT  1047600.0 1869600.0 1057800.0 1855800.0 ;
      RECT  1047600.0 1869600.0 1057800.0 1883400.0 ;
      RECT  1047600.0 1897200.0 1057800.0 1883400.0 ;
      RECT  1047600.0 1897200.0 1057800.0 1911000.0 ;
      RECT  1047600.0 1924800.0 1057800.0 1911000.0 ;
      RECT  1047600.0 1924800.0 1057800.0 1938600.0 ;
      RECT  1047600.0 1952400.0 1057800.0 1938600.0 ;
      RECT  1047600.0 1952400.0 1057800.0 1966200.0 ;
      RECT  1047600.0 1980000.0 1057800.0 1966200.0 ;
      RECT  1047600.0 1980000.0 1057800.0 1993800.0 ;
      RECT  1047600.0 2007600.0 1057800.0 1993800.0 ;
      RECT  1047600.0 2007600.0 1057800.0 2021400.0 ;
      RECT  1047600.0 2035200.0 1057800.0 2021400.0 ;
      RECT  1047600.0 2035200.0 1057800.0 2049000.0 ;
      RECT  1047600.0 2062800.0 1057800.0 2049000.0 ;
      RECT  1047600.0 2062800.0 1057800.0 2076600.0 ;
      RECT  1047600.0 2090400.0 1057800.0 2076600.0 ;
      RECT  1047600.0 2090400.0 1057800.0 2104200.0 ;
      RECT  1047600.0 2118000.0 1057800.0 2104200.0 ;
      RECT  1047600.0 2118000.0 1057800.0 2131800.0 ;
      RECT  1047600.0 2145600.0 1057800.0 2131800.0 ;
      RECT  1057800.0 379200.0 1068000.0 393000.0 ;
      RECT  1057800.0 406800.0 1068000.0 393000.0 ;
      RECT  1057800.0 406800.0 1068000.0 420600.0 ;
      RECT  1057800.0 434400.0 1068000.0 420600.0 ;
      RECT  1057800.0 434400.0 1068000.0 448200.0 ;
      RECT  1057800.0 462000.0 1068000.0 448200.0 ;
      RECT  1057800.0 462000.0 1068000.0 475800.0 ;
      RECT  1057800.0 489600.0 1068000.0 475800.0 ;
      RECT  1057800.0 489600.0 1068000.0 503400.0 ;
      RECT  1057800.0 517200.0 1068000.0 503400.0 ;
      RECT  1057800.0 517200.0 1068000.0 531000.0 ;
      RECT  1057800.0 544800.0 1068000.0 531000.0 ;
      RECT  1057800.0 544800.0 1068000.0 558600.0 ;
      RECT  1057800.0 572400.0 1068000.0 558600.0 ;
      RECT  1057800.0 572400.0 1068000.0 586200.0 ;
      RECT  1057800.0 600000.0 1068000.0 586200.0 ;
      RECT  1057800.0 600000.0 1068000.0 613800.0 ;
      RECT  1057800.0 627600.0 1068000.0 613800.0 ;
      RECT  1057800.0 627600.0 1068000.0 641400.0 ;
      RECT  1057800.0 655200.0 1068000.0 641400.0 ;
      RECT  1057800.0 655200.0 1068000.0 669000.0 ;
      RECT  1057800.0 682800.0 1068000.0 669000.0 ;
      RECT  1057800.0 682800.0 1068000.0 696600.0 ;
      RECT  1057800.0 710400.0 1068000.0 696600.0 ;
      RECT  1057800.0 710400.0 1068000.0 724200.0 ;
      RECT  1057800.0 738000.0 1068000.0 724200.0 ;
      RECT  1057800.0 738000.0 1068000.0 751800.0 ;
      RECT  1057800.0 765600.0 1068000.0 751800.0 ;
      RECT  1057800.0 765600.0 1068000.0 779400.0 ;
      RECT  1057800.0 793200.0 1068000.0 779400.0 ;
      RECT  1057800.0 793200.0 1068000.0 807000.0 ;
      RECT  1057800.0 820800.0 1068000.0 807000.0 ;
      RECT  1057800.0 820800.0 1068000.0 834600.0 ;
      RECT  1057800.0 848400.0 1068000.0 834600.0 ;
      RECT  1057800.0 848400.0 1068000.0 862200.0 ;
      RECT  1057800.0 876000.0 1068000.0 862200.0 ;
      RECT  1057800.0 876000.0 1068000.0 889800.0 ;
      RECT  1057800.0 903600.0 1068000.0 889800.0 ;
      RECT  1057800.0 903600.0 1068000.0 917400.0 ;
      RECT  1057800.0 931200.0 1068000.0 917400.0 ;
      RECT  1057800.0 931200.0 1068000.0 945000.0 ;
      RECT  1057800.0 958800.0 1068000.0 945000.0 ;
      RECT  1057800.0 958800.0 1068000.0 972600.0 ;
      RECT  1057800.0 986400.0 1068000.0 972600.0 ;
      RECT  1057800.0 986400.0 1068000.0 1000200.0 ;
      RECT  1057800.0 1014000.0 1068000.0 1000200.0 ;
      RECT  1057800.0 1014000.0 1068000.0 1027800.0 ;
      RECT  1057800.0 1041600.0 1068000.0 1027800.0 ;
      RECT  1057800.0 1041600.0 1068000.0 1055400.0 ;
      RECT  1057800.0 1069200.0 1068000.0 1055400.0 ;
      RECT  1057800.0 1069200.0 1068000.0 1083000.0 ;
      RECT  1057800.0 1096800.0 1068000.0 1083000.0 ;
      RECT  1057800.0 1096800.0 1068000.0 1110600.0 ;
      RECT  1057800.0 1124400.0 1068000.0 1110600.0 ;
      RECT  1057800.0 1124400.0 1068000.0 1138200.0 ;
      RECT  1057800.0 1152000.0 1068000.0 1138200.0 ;
      RECT  1057800.0 1152000.0 1068000.0 1165800.0 ;
      RECT  1057800.0 1179600.0 1068000.0 1165800.0 ;
      RECT  1057800.0 1179600.0 1068000.0 1193400.0 ;
      RECT  1057800.0 1207200.0 1068000.0 1193400.0 ;
      RECT  1057800.0 1207200.0 1068000.0 1221000.0 ;
      RECT  1057800.0 1234800.0 1068000.0 1221000.0 ;
      RECT  1057800.0 1234800.0 1068000.0 1248600.0 ;
      RECT  1057800.0 1262400.0 1068000.0 1248600.0 ;
      RECT  1057800.0 1262400.0 1068000.0 1276200.0 ;
      RECT  1057800.0 1290000.0 1068000.0 1276200.0 ;
      RECT  1057800.0 1290000.0 1068000.0 1303800.0 ;
      RECT  1057800.0 1317600.0 1068000.0 1303800.0 ;
      RECT  1057800.0 1317600.0 1068000.0 1331400.0 ;
      RECT  1057800.0 1345200.0 1068000.0 1331400.0 ;
      RECT  1057800.0 1345200.0 1068000.0 1359000.0 ;
      RECT  1057800.0 1372800.0 1068000.0 1359000.0 ;
      RECT  1057800.0 1372800.0 1068000.0 1386600.0 ;
      RECT  1057800.0 1400400.0 1068000.0 1386600.0 ;
      RECT  1057800.0 1400400.0 1068000.0 1414200.0 ;
      RECT  1057800.0 1428000.0 1068000.0 1414200.0 ;
      RECT  1057800.0 1428000.0 1068000.0 1441800.0 ;
      RECT  1057800.0 1455600.0 1068000.0 1441800.0 ;
      RECT  1057800.0 1455600.0 1068000.0 1469400.0 ;
      RECT  1057800.0 1483200.0 1068000.0 1469400.0 ;
      RECT  1057800.0 1483200.0 1068000.0 1497000.0 ;
      RECT  1057800.0 1510800.0 1068000.0 1497000.0 ;
      RECT  1057800.0 1510800.0 1068000.0 1524600.0 ;
      RECT  1057800.0 1538400.0 1068000.0 1524600.0 ;
      RECT  1057800.0 1538400.0 1068000.0 1552200.0 ;
      RECT  1057800.0 1566000.0 1068000.0 1552200.0 ;
      RECT  1057800.0 1566000.0 1068000.0 1579800.0 ;
      RECT  1057800.0 1593600.0 1068000.0 1579800.0 ;
      RECT  1057800.0 1593600.0 1068000.0 1607400.0 ;
      RECT  1057800.0 1621200.0 1068000.0 1607400.0 ;
      RECT  1057800.0 1621200.0 1068000.0 1635000.0 ;
      RECT  1057800.0 1648800.0 1068000.0 1635000.0 ;
      RECT  1057800.0 1648800.0 1068000.0 1662600.0 ;
      RECT  1057800.0 1676400.0 1068000.0 1662600.0 ;
      RECT  1057800.0 1676400.0 1068000.0 1690200.0 ;
      RECT  1057800.0 1704000.0 1068000.0 1690200.0 ;
      RECT  1057800.0 1704000.0 1068000.0 1717800.0 ;
      RECT  1057800.0 1731600.0 1068000.0 1717800.0 ;
      RECT  1057800.0 1731600.0 1068000.0 1745400.0 ;
      RECT  1057800.0 1759200.0 1068000.0 1745400.0 ;
      RECT  1057800.0 1759200.0 1068000.0 1773000.0 ;
      RECT  1057800.0 1786800.0 1068000.0 1773000.0 ;
      RECT  1057800.0 1786800.0 1068000.0 1800600.0 ;
      RECT  1057800.0 1814400.0 1068000.0 1800600.0 ;
      RECT  1057800.0 1814400.0 1068000.0 1828200.0 ;
      RECT  1057800.0 1842000.0 1068000.0 1828200.0 ;
      RECT  1057800.0 1842000.0 1068000.0 1855800.0 ;
      RECT  1057800.0 1869600.0 1068000.0 1855800.0 ;
      RECT  1057800.0 1869600.0 1068000.0 1883400.0 ;
      RECT  1057800.0 1897200.0 1068000.0 1883400.0 ;
      RECT  1057800.0 1897200.0 1068000.0 1911000.0 ;
      RECT  1057800.0 1924800.0 1068000.0 1911000.0 ;
      RECT  1057800.0 1924800.0 1068000.0 1938600.0 ;
      RECT  1057800.0 1952400.0 1068000.0 1938600.0 ;
      RECT  1057800.0 1952400.0 1068000.0 1966200.0 ;
      RECT  1057800.0 1980000.0 1068000.0 1966200.0 ;
      RECT  1057800.0 1980000.0 1068000.0 1993800.0 ;
      RECT  1057800.0 2007600.0 1068000.0 1993800.0 ;
      RECT  1057800.0 2007600.0 1068000.0 2021400.0 ;
      RECT  1057800.0 2035200.0 1068000.0 2021400.0 ;
      RECT  1057800.0 2035200.0 1068000.0 2049000.0 ;
      RECT  1057800.0 2062800.0 1068000.0 2049000.0 ;
      RECT  1057800.0 2062800.0 1068000.0 2076600.0 ;
      RECT  1057800.0 2090400.0 1068000.0 2076600.0 ;
      RECT  1057800.0 2090400.0 1068000.0 2104200.0 ;
      RECT  1057800.0 2118000.0 1068000.0 2104200.0 ;
      RECT  1057800.0 2118000.0 1068000.0 2131800.0 ;
      RECT  1057800.0 2145600.0 1068000.0 2131800.0 ;
      RECT  1068000.0 379200.0 1078200.0 393000.0 ;
      RECT  1068000.0 406800.0 1078200.0 393000.0 ;
      RECT  1068000.0 406800.0 1078200.0 420600.0 ;
      RECT  1068000.0 434400.0 1078200.0 420600.0 ;
      RECT  1068000.0 434400.0 1078200.0 448200.0 ;
      RECT  1068000.0 462000.0 1078200.0 448200.0 ;
      RECT  1068000.0 462000.0 1078200.0 475800.0 ;
      RECT  1068000.0 489600.0 1078200.0 475800.0 ;
      RECT  1068000.0 489600.0 1078200.0 503400.0 ;
      RECT  1068000.0 517200.0 1078200.0 503400.0 ;
      RECT  1068000.0 517200.0 1078200.0 531000.0 ;
      RECT  1068000.0 544800.0 1078200.0 531000.0 ;
      RECT  1068000.0 544800.0 1078200.0 558600.0 ;
      RECT  1068000.0 572400.0 1078200.0 558600.0 ;
      RECT  1068000.0 572400.0 1078200.0 586200.0 ;
      RECT  1068000.0 600000.0 1078200.0 586200.0 ;
      RECT  1068000.0 600000.0 1078200.0 613800.0 ;
      RECT  1068000.0 627600.0 1078200.0 613800.0 ;
      RECT  1068000.0 627600.0 1078200.0 641400.0 ;
      RECT  1068000.0 655200.0 1078200.0 641400.0 ;
      RECT  1068000.0 655200.0 1078200.0 669000.0 ;
      RECT  1068000.0 682800.0 1078200.0 669000.0 ;
      RECT  1068000.0 682800.0 1078200.0 696600.0 ;
      RECT  1068000.0 710400.0 1078200.0 696600.0 ;
      RECT  1068000.0 710400.0 1078200.0 724200.0 ;
      RECT  1068000.0 738000.0 1078200.0 724200.0 ;
      RECT  1068000.0 738000.0 1078200.0 751800.0 ;
      RECT  1068000.0 765600.0 1078200.0 751800.0 ;
      RECT  1068000.0 765600.0 1078200.0 779400.0 ;
      RECT  1068000.0 793200.0 1078200.0 779400.0 ;
      RECT  1068000.0 793200.0 1078200.0 807000.0 ;
      RECT  1068000.0 820800.0 1078200.0 807000.0 ;
      RECT  1068000.0 820800.0 1078200.0 834600.0 ;
      RECT  1068000.0 848400.0 1078200.0 834600.0 ;
      RECT  1068000.0 848400.0 1078200.0 862200.0 ;
      RECT  1068000.0 876000.0 1078200.0 862200.0 ;
      RECT  1068000.0 876000.0 1078200.0 889800.0 ;
      RECT  1068000.0 903600.0 1078200.0 889800.0 ;
      RECT  1068000.0 903600.0 1078200.0 917400.0 ;
      RECT  1068000.0 931200.0 1078200.0 917400.0 ;
      RECT  1068000.0 931200.0 1078200.0 945000.0 ;
      RECT  1068000.0 958800.0 1078200.0 945000.0 ;
      RECT  1068000.0 958800.0 1078200.0 972600.0 ;
      RECT  1068000.0 986400.0 1078200.0 972600.0 ;
      RECT  1068000.0 986400.0 1078200.0 1000200.0 ;
      RECT  1068000.0 1014000.0 1078200.0 1000200.0 ;
      RECT  1068000.0 1014000.0 1078200.0 1027800.0 ;
      RECT  1068000.0 1041600.0 1078200.0 1027800.0 ;
      RECT  1068000.0 1041600.0 1078200.0 1055400.0 ;
      RECT  1068000.0 1069200.0 1078200.0 1055400.0 ;
      RECT  1068000.0 1069200.0 1078200.0 1083000.0 ;
      RECT  1068000.0 1096800.0 1078200.0 1083000.0 ;
      RECT  1068000.0 1096800.0 1078200.0 1110600.0 ;
      RECT  1068000.0 1124400.0 1078200.0 1110600.0 ;
      RECT  1068000.0 1124400.0 1078200.0 1138200.0 ;
      RECT  1068000.0 1152000.0 1078200.0 1138200.0 ;
      RECT  1068000.0 1152000.0 1078200.0 1165800.0 ;
      RECT  1068000.0 1179600.0 1078200.0 1165800.0 ;
      RECT  1068000.0 1179600.0 1078200.0 1193400.0 ;
      RECT  1068000.0 1207200.0 1078200.0 1193400.0 ;
      RECT  1068000.0 1207200.0 1078200.0 1221000.0 ;
      RECT  1068000.0 1234800.0 1078200.0 1221000.0 ;
      RECT  1068000.0 1234800.0 1078200.0 1248600.0 ;
      RECT  1068000.0 1262400.0 1078200.0 1248600.0 ;
      RECT  1068000.0 1262400.0 1078200.0 1276200.0 ;
      RECT  1068000.0 1290000.0 1078200.0 1276200.0 ;
      RECT  1068000.0 1290000.0 1078200.0 1303800.0 ;
      RECT  1068000.0 1317600.0 1078200.0 1303800.0 ;
      RECT  1068000.0 1317600.0 1078200.0 1331400.0 ;
      RECT  1068000.0 1345200.0 1078200.0 1331400.0 ;
      RECT  1068000.0 1345200.0 1078200.0 1359000.0 ;
      RECT  1068000.0 1372800.0 1078200.0 1359000.0 ;
      RECT  1068000.0 1372800.0 1078200.0 1386600.0 ;
      RECT  1068000.0 1400400.0 1078200.0 1386600.0 ;
      RECT  1068000.0 1400400.0 1078200.0 1414200.0 ;
      RECT  1068000.0 1428000.0 1078200.0 1414200.0 ;
      RECT  1068000.0 1428000.0 1078200.0 1441800.0 ;
      RECT  1068000.0 1455600.0 1078200.0 1441800.0 ;
      RECT  1068000.0 1455600.0 1078200.0 1469400.0 ;
      RECT  1068000.0 1483200.0 1078200.0 1469400.0 ;
      RECT  1068000.0 1483200.0 1078200.0 1497000.0 ;
      RECT  1068000.0 1510800.0 1078200.0 1497000.0 ;
      RECT  1068000.0 1510800.0 1078200.0 1524600.0 ;
      RECT  1068000.0 1538400.0 1078200.0 1524600.0 ;
      RECT  1068000.0 1538400.0 1078200.0 1552200.0 ;
      RECT  1068000.0 1566000.0 1078200.0 1552200.0 ;
      RECT  1068000.0 1566000.0 1078200.0 1579800.0 ;
      RECT  1068000.0 1593600.0 1078200.0 1579800.0 ;
      RECT  1068000.0 1593600.0 1078200.0 1607400.0 ;
      RECT  1068000.0 1621200.0 1078200.0 1607400.0 ;
      RECT  1068000.0 1621200.0 1078200.0 1635000.0 ;
      RECT  1068000.0 1648800.0 1078200.0 1635000.0 ;
      RECT  1068000.0 1648800.0 1078200.0 1662600.0 ;
      RECT  1068000.0 1676400.0 1078200.0 1662600.0 ;
      RECT  1068000.0 1676400.0 1078200.0 1690200.0 ;
      RECT  1068000.0 1704000.0 1078200.0 1690200.0 ;
      RECT  1068000.0 1704000.0 1078200.0 1717800.0 ;
      RECT  1068000.0 1731600.0 1078200.0 1717800.0 ;
      RECT  1068000.0 1731600.0 1078200.0 1745400.0 ;
      RECT  1068000.0 1759200.0 1078200.0 1745400.0 ;
      RECT  1068000.0 1759200.0 1078200.0 1773000.0 ;
      RECT  1068000.0 1786800.0 1078200.0 1773000.0 ;
      RECT  1068000.0 1786800.0 1078200.0 1800600.0 ;
      RECT  1068000.0 1814400.0 1078200.0 1800600.0 ;
      RECT  1068000.0 1814400.0 1078200.0 1828200.0 ;
      RECT  1068000.0 1842000.0 1078200.0 1828200.0 ;
      RECT  1068000.0 1842000.0 1078200.0 1855800.0 ;
      RECT  1068000.0 1869600.0 1078200.0 1855800.0 ;
      RECT  1068000.0 1869600.0 1078200.0 1883400.0 ;
      RECT  1068000.0 1897200.0 1078200.0 1883400.0 ;
      RECT  1068000.0 1897200.0 1078200.0 1911000.0 ;
      RECT  1068000.0 1924800.0 1078200.0 1911000.0 ;
      RECT  1068000.0 1924800.0 1078200.0 1938600.0 ;
      RECT  1068000.0 1952400.0 1078200.0 1938600.0 ;
      RECT  1068000.0 1952400.0 1078200.0 1966200.0 ;
      RECT  1068000.0 1980000.0 1078200.0 1966200.0 ;
      RECT  1068000.0 1980000.0 1078200.0 1993800.0 ;
      RECT  1068000.0 2007600.0 1078200.0 1993800.0 ;
      RECT  1068000.0 2007600.0 1078200.0 2021400.0 ;
      RECT  1068000.0 2035200.0 1078200.0 2021400.0 ;
      RECT  1068000.0 2035200.0 1078200.0 2049000.0 ;
      RECT  1068000.0 2062800.0 1078200.0 2049000.0 ;
      RECT  1068000.0 2062800.0 1078200.0 2076600.0 ;
      RECT  1068000.0 2090400.0 1078200.0 2076600.0 ;
      RECT  1068000.0 2090400.0 1078200.0 2104200.0 ;
      RECT  1068000.0 2118000.0 1078200.0 2104200.0 ;
      RECT  1068000.0 2118000.0 1078200.0 2131800.0 ;
      RECT  1068000.0 2145600.0 1078200.0 2131800.0 ;
      RECT  1078200.0 379200.0 1088400.0 393000.0 ;
      RECT  1078200.0 406800.0 1088400.0 393000.0 ;
      RECT  1078200.0 406800.0 1088400.0 420600.0 ;
      RECT  1078200.0 434400.0 1088400.0 420600.0 ;
      RECT  1078200.0 434400.0 1088400.0 448200.0 ;
      RECT  1078200.0 462000.0 1088400.0 448200.0 ;
      RECT  1078200.0 462000.0 1088400.0 475800.0 ;
      RECT  1078200.0 489600.0 1088400.0 475800.0 ;
      RECT  1078200.0 489600.0 1088400.0 503400.0 ;
      RECT  1078200.0 517200.0 1088400.0 503400.0 ;
      RECT  1078200.0 517200.0 1088400.0 531000.0 ;
      RECT  1078200.0 544800.0 1088400.0 531000.0 ;
      RECT  1078200.0 544800.0 1088400.0 558600.0 ;
      RECT  1078200.0 572400.0 1088400.0 558600.0 ;
      RECT  1078200.0 572400.0 1088400.0 586200.0 ;
      RECT  1078200.0 600000.0 1088400.0 586200.0 ;
      RECT  1078200.0 600000.0 1088400.0 613800.0 ;
      RECT  1078200.0 627600.0 1088400.0 613800.0 ;
      RECT  1078200.0 627600.0 1088400.0 641400.0 ;
      RECT  1078200.0 655200.0 1088400.0 641400.0 ;
      RECT  1078200.0 655200.0 1088400.0 669000.0 ;
      RECT  1078200.0 682800.0 1088400.0 669000.0 ;
      RECT  1078200.0 682800.0 1088400.0 696600.0 ;
      RECT  1078200.0 710400.0 1088400.0 696600.0 ;
      RECT  1078200.0 710400.0 1088400.0 724200.0 ;
      RECT  1078200.0 738000.0 1088400.0 724200.0 ;
      RECT  1078200.0 738000.0 1088400.0 751800.0 ;
      RECT  1078200.0 765600.0 1088400.0 751800.0 ;
      RECT  1078200.0 765600.0 1088400.0 779400.0 ;
      RECT  1078200.0 793200.0 1088400.0 779400.0 ;
      RECT  1078200.0 793200.0 1088400.0 807000.0 ;
      RECT  1078200.0 820800.0 1088400.0 807000.0 ;
      RECT  1078200.0 820800.0 1088400.0 834600.0 ;
      RECT  1078200.0 848400.0 1088400.0 834600.0 ;
      RECT  1078200.0 848400.0 1088400.0 862200.0 ;
      RECT  1078200.0 876000.0 1088400.0 862200.0 ;
      RECT  1078200.0 876000.0 1088400.0 889800.0 ;
      RECT  1078200.0 903600.0 1088400.0 889800.0 ;
      RECT  1078200.0 903600.0 1088400.0 917400.0 ;
      RECT  1078200.0 931200.0 1088400.0 917400.0 ;
      RECT  1078200.0 931200.0 1088400.0 945000.0 ;
      RECT  1078200.0 958800.0 1088400.0 945000.0 ;
      RECT  1078200.0 958800.0 1088400.0 972600.0 ;
      RECT  1078200.0 986400.0 1088400.0 972600.0 ;
      RECT  1078200.0 986400.0 1088400.0 1000200.0 ;
      RECT  1078200.0 1014000.0 1088400.0 1000200.0 ;
      RECT  1078200.0 1014000.0 1088400.0 1027800.0 ;
      RECT  1078200.0 1041600.0 1088400.0 1027800.0 ;
      RECT  1078200.0 1041600.0 1088400.0 1055400.0 ;
      RECT  1078200.0 1069200.0 1088400.0 1055400.0 ;
      RECT  1078200.0 1069200.0 1088400.0 1083000.0 ;
      RECT  1078200.0 1096800.0 1088400.0 1083000.0 ;
      RECT  1078200.0 1096800.0 1088400.0 1110600.0 ;
      RECT  1078200.0 1124400.0 1088400.0 1110600.0 ;
      RECT  1078200.0 1124400.0 1088400.0 1138200.0 ;
      RECT  1078200.0 1152000.0 1088400.0 1138200.0 ;
      RECT  1078200.0 1152000.0 1088400.0 1165800.0 ;
      RECT  1078200.0 1179600.0 1088400.0 1165800.0 ;
      RECT  1078200.0 1179600.0 1088400.0 1193400.0 ;
      RECT  1078200.0 1207200.0 1088400.0 1193400.0 ;
      RECT  1078200.0 1207200.0 1088400.0 1221000.0 ;
      RECT  1078200.0 1234800.0 1088400.0 1221000.0 ;
      RECT  1078200.0 1234800.0 1088400.0 1248600.0 ;
      RECT  1078200.0 1262400.0 1088400.0 1248600.0 ;
      RECT  1078200.0 1262400.0 1088400.0 1276200.0 ;
      RECT  1078200.0 1290000.0 1088400.0 1276200.0 ;
      RECT  1078200.0 1290000.0 1088400.0 1303800.0 ;
      RECT  1078200.0 1317600.0 1088400.0 1303800.0 ;
      RECT  1078200.0 1317600.0 1088400.0 1331400.0 ;
      RECT  1078200.0 1345200.0 1088400.0 1331400.0 ;
      RECT  1078200.0 1345200.0 1088400.0 1359000.0 ;
      RECT  1078200.0 1372800.0 1088400.0 1359000.0 ;
      RECT  1078200.0 1372800.0 1088400.0 1386600.0 ;
      RECT  1078200.0 1400400.0 1088400.0 1386600.0 ;
      RECT  1078200.0 1400400.0 1088400.0 1414200.0 ;
      RECT  1078200.0 1428000.0 1088400.0 1414200.0 ;
      RECT  1078200.0 1428000.0 1088400.0 1441800.0 ;
      RECT  1078200.0 1455600.0 1088400.0 1441800.0 ;
      RECT  1078200.0 1455600.0 1088400.0 1469400.0 ;
      RECT  1078200.0 1483200.0 1088400.0 1469400.0 ;
      RECT  1078200.0 1483200.0 1088400.0 1497000.0 ;
      RECT  1078200.0 1510800.0 1088400.0 1497000.0 ;
      RECT  1078200.0 1510800.0 1088400.0 1524600.0 ;
      RECT  1078200.0 1538400.0 1088400.0 1524600.0 ;
      RECT  1078200.0 1538400.0 1088400.0 1552200.0 ;
      RECT  1078200.0 1566000.0 1088400.0 1552200.0 ;
      RECT  1078200.0 1566000.0 1088400.0 1579800.0 ;
      RECT  1078200.0 1593600.0 1088400.0 1579800.0 ;
      RECT  1078200.0 1593600.0 1088400.0 1607400.0 ;
      RECT  1078200.0 1621200.0 1088400.0 1607400.0 ;
      RECT  1078200.0 1621200.0 1088400.0 1635000.0 ;
      RECT  1078200.0 1648800.0 1088400.0 1635000.0 ;
      RECT  1078200.0 1648800.0 1088400.0 1662600.0 ;
      RECT  1078200.0 1676400.0 1088400.0 1662600.0 ;
      RECT  1078200.0 1676400.0 1088400.0 1690200.0 ;
      RECT  1078200.0 1704000.0 1088400.0 1690200.0 ;
      RECT  1078200.0 1704000.0 1088400.0 1717800.0 ;
      RECT  1078200.0 1731600.0 1088400.0 1717800.0 ;
      RECT  1078200.0 1731600.0 1088400.0 1745400.0 ;
      RECT  1078200.0 1759200.0 1088400.0 1745400.0 ;
      RECT  1078200.0 1759200.0 1088400.0 1773000.0 ;
      RECT  1078200.0 1786800.0 1088400.0 1773000.0 ;
      RECT  1078200.0 1786800.0 1088400.0 1800600.0 ;
      RECT  1078200.0 1814400.0 1088400.0 1800600.0 ;
      RECT  1078200.0 1814400.0 1088400.0 1828200.0 ;
      RECT  1078200.0 1842000.0 1088400.0 1828200.0 ;
      RECT  1078200.0 1842000.0 1088400.0 1855800.0 ;
      RECT  1078200.0 1869600.0 1088400.0 1855800.0 ;
      RECT  1078200.0 1869600.0 1088400.0 1883400.0 ;
      RECT  1078200.0 1897200.0 1088400.0 1883400.0 ;
      RECT  1078200.0 1897200.0 1088400.0 1911000.0 ;
      RECT  1078200.0 1924800.0 1088400.0 1911000.0 ;
      RECT  1078200.0 1924800.0 1088400.0 1938600.0 ;
      RECT  1078200.0 1952400.0 1088400.0 1938600.0 ;
      RECT  1078200.0 1952400.0 1088400.0 1966200.0 ;
      RECT  1078200.0 1980000.0 1088400.0 1966200.0 ;
      RECT  1078200.0 1980000.0 1088400.0 1993800.0 ;
      RECT  1078200.0 2007600.0 1088400.0 1993800.0 ;
      RECT  1078200.0 2007600.0 1088400.0 2021400.0 ;
      RECT  1078200.0 2035200.0 1088400.0 2021400.0 ;
      RECT  1078200.0 2035200.0 1088400.0 2049000.0 ;
      RECT  1078200.0 2062800.0 1088400.0 2049000.0 ;
      RECT  1078200.0 2062800.0 1088400.0 2076600.0 ;
      RECT  1078200.0 2090400.0 1088400.0 2076600.0 ;
      RECT  1078200.0 2090400.0 1088400.0 2104200.0 ;
      RECT  1078200.0 2118000.0 1088400.0 2104200.0 ;
      RECT  1078200.0 2118000.0 1088400.0 2131800.0 ;
      RECT  1078200.0 2145600.0 1088400.0 2131800.0 ;
      RECT  1088400.0 379200.0 1098600.0 393000.0 ;
      RECT  1088400.0 406800.0 1098600.0 393000.0 ;
      RECT  1088400.0 406800.0 1098600.0 420600.0 ;
      RECT  1088400.0 434400.0 1098600.0 420600.0 ;
      RECT  1088400.0 434400.0 1098600.0 448200.0 ;
      RECT  1088400.0 462000.0 1098600.0 448200.0 ;
      RECT  1088400.0 462000.0 1098600.0 475800.0 ;
      RECT  1088400.0 489600.0 1098600.0 475800.0 ;
      RECT  1088400.0 489600.0 1098600.0 503400.0 ;
      RECT  1088400.0 517200.0 1098600.0 503400.0 ;
      RECT  1088400.0 517200.0 1098600.0 531000.0 ;
      RECT  1088400.0 544800.0 1098600.0 531000.0 ;
      RECT  1088400.0 544800.0 1098600.0 558600.0 ;
      RECT  1088400.0 572400.0 1098600.0 558600.0 ;
      RECT  1088400.0 572400.0 1098600.0 586200.0 ;
      RECT  1088400.0 600000.0 1098600.0 586200.0 ;
      RECT  1088400.0 600000.0 1098600.0 613800.0 ;
      RECT  1088400.0 627600.0 1098600.0 613800.0 ;
      RECT  1088400.0 627600.0 1098600.0 641400.0 ;
      RECT  1088400.0 655200.0 1098600.0 641400.0 ;
      RECT  1088400.0 655200.0 1098600.0 669000.0 ;
      RECT  1088400.0 682800.0 1098600.0 669000.0 ;
      RECT  1088400.0 682800.0 1098600.0 696600.0 ;
      RECT  1088400.0 710400.0 1098600.0 696600.0 ;
      RECT  1088400.0 710400.0 1098600.0 724200.0 ;
      RECT  1088400.0 738000.0 1098600.0 724200.0 ;
      RECT  1088400.0 738000.0 1098600.0 751800.0 ;
      RECT  1088400.0 765600.0 1098600.0 751800.0 ;
      RECT  1088400.0 765600.0 1098600.0 779400.0 ;
      RECT  1088400.0 793200.0 1098600.0 779400.0 ;
      RECT  1088400.0 793200.0 1098600.0 807000.0 ;
      RECT  1088400.0 820800.0 1098600.0 807000.0 ;
      RECT  1088400.0 820800.0 1098600.0 834600.0 ;
      RECT  1088400.0 848400.0 1098600.0 834600.0 ;
      RECT  1088400.0 848400.0 1098600.0 862200.0 ;
      RECT  1088400.0 876000.0 1098600.0 862200.0 ;
      RECT  1088400.0 876000.0 1098600.0 889800.0 ;
      RECT  1088400.0 903600.0 1098600.0 889800.0 ;
      RECT  1088400.0 903600.0 1098600.0 917400.0 ;
      RECT  1088400.0 931200.0 1098600.0 917400.0 ;
      RECT  1088400.0 931200.0 1098600.0 945000.0 ;
      RECT  1088400.0 958800.0 1098600.0 945000.0 ;
      RECT  1088400.0 958800.0 1098600.0 972600.0 ;
      RECT  1088400.0 986400.0 1098600.0 972600.0 ;
      RECT  1088400.0 986400.0 1098600.0 1000200.0 ;
      RECT  1088400.0 1014000.0 1098600.0 1000200.0 ;
      RECT  1088400.0 1014000.0 1098600.0 1027800.0 ;
      RECT  1088400.0 1041600.0 1098600.0 1027800.0 ;
      RECT  1088400.0 1041600.0 1098600.0 1055400.0 ;
      RECT  1088400.0 1069200.0 1098600.0 1055400.0 ;
      RECT  1088400.0 1069200.0 1098600.0 1083000.0 ;
      RECT  1088400.0 1096800.0 1098600.0 1083000.0 ;
      RECT  1088400.0 1096800.0 1098600.0 1110600.0 ;
      RECT  1088400.0 1124400.0 1098600.0 1110600.0 ;
      RECT  1088400.0 1124400.0 1098600.0 1138200.0 ;
      RECT  1088400.0 1152000.0 1098600.0 1138200.0 ;
      RECT  1088400.0 1152000.0 1098600.0 1165800.0 ;
      RECT  1088400.0 1179600.0 1098600.0 1165800.0 ;
      RECT  1088400.0 1179600.0 1098600.0 1193400.0 ;
      RECT  1088400.0 1207200.0 1098600.0 1193400.0 ;
      RECT  1088400.0 1207200.0 1098600.0 1221000.0 ;
      RECT  1088400.0 1234800.0 1098600.0 1221000.0 ;
      RECT  1088400.0 1234800.0 1098600.0 1248600.0 ;
      RECT  1088400.0 1262400.0 1098600.0 1248600.0 ;
      RECT  1088400.0 1262400.0 1098600.0 1276200.0 ;
      RECT  1088400.0 1290000.0 1098600.0 1276200.0 ;
      RECT  1088400.0 1290000.0 1098600.0 1303800.0 ;
      RECT  1088400.0 1317600.0 1098600.0 1303800.0 ;
      RECT  1088400.0 1317600.0 1098600.0 1331400.0 ;
      RECT  1088400.0 1345200.0 1098600.0 1331400.0 ;
      RECT  1088400.0 1345200.0 1098600.0 1359000.0 ;
      RECT  1088400.0 1372800.0 1098600.0 1359000.0 ;
      RECT  1088400.0 1372800.0 1098600.0 1386600.0 ;
      RECT  1088400.0 1400400.0 1098600.0 1386600.0 ;
      RECT  1088400.0 1400400.0 1098600.0 1414200.0 ;
      RECT  1088400.0 1428000.0 1098600.0 1414200.0 ;
      RECT  1088400.0 1428000.0 1098600.0 1441800.0 ;
      RECT  1088400.0 1455600.0 1098600.0 1441800.0 ;
      RECT  1088400.0 1455600.0 1098600.0 1469400.0 ;
      RECT  1088400.0 1483200.0 1098600.0 1469400.0 ;
      RECT  1088400.0 1483200.0 1098600.0 1497000.0 ;
      RECT  1088400.0 1510800.0 1098600.0 1497000.0 ;
      RECT  1088400.0 1510800.0 1098600.0 1524600.0 ;
      RECT  1088400.0 1538400.0 1098600.0 1524600.0 ;
      RECT  1088400.0 1538400.0 1098600.0 1552200.0 ;
      RECT  1088400.0 1566000.0 1098600.0 1552200.0 ;
      RECT  1088400.0 1566000.0 1098600.0 1579800.0 ;
      RECT  1088400.0 1593600.0 1098600.0 1579800.0 ;
      RECT  1088400.0 1593600.0 1098600.0 1607400.0 ;
      RECT  1088400.0 1621200.0 1098600.0 1607400.0 ;
      RECT  1088400.0 1621200.0 1098600.0 1635000.0 ;
      RECT  1088400.0 1648800.0 1098600.0 1635000.0 ;
      RECT  1088400.0 1648800.0 1098600.0 1662600.0 ;
      RECT  1088400.0 1676400.0 1098600.0 1662600.0 ;
      RECT  1088400.0 1676400.0 1098600.0 1690200.0 ;
      RECT  1088400.0 1704000.0 1098600.0 1690200.0 ;
      RECT  1088400.0 1704000.0 1098600.0 1717800.0 ;
      RECT  1088400.0 1731600.0 1098600.0 1717800.0 ;
      RECT  1088400.0 1731600.0 1098600.0 1745400.0 ;
      RECT  1088400.0 1759200.0 1098600.0 1745400.0 ;
      RECT  1088400.0 1759200.0 1098600.0 1773000.0 ;
      RECT  1088400.0 1786800.0 1098600.0 1773000.0 ;
      RECT  1088400.0 1786800.0 1098600.0 1800600.0 ;
      RECT  1088400.0 1814400.0 1098600.0 1800600.0 ;
      RECT  1088400.0 1814400.0 1098600.0 1828200.0 ;
      RECT  1088400.0 1842000.0 1098600.0 1828200.0 ;
      RECT  1088400.0 1842000.0 1098600.0 1855800.0 ;
      RECT  1088400.0 1869600.0 1098600.0 1855800.0 ;
      RECT  1088400.0 1869600.0 1098600.0 1883400.0 ;
      RECT  1088400.0 1897200.0 1098600.0 1883400.0 ;
      RECT  1088400.0 1897200.0 1098600.0 1911000.0 ;
      RECT  1088400.0 1924800.0 1098600.0 1911000.0 ;
      RECT  1088400.0 1924800.0 1098600.0 1938600.0 ;
      RECT  1088400.0 1952400.0 1098600.0 1938600.0 ;
      RECT  1088400.0 1952400.0 1098600.0 1966200.0 ;
      RECT  1088400.0 1980000.0 1098600.0 1966200.0 ;
      RECT  1088400.0 1980000.0 1098600.0 1993800.0 ;
      RECT  1088400.0 2007600.0 1098600.0 1993800.0 ;
      RECT  1088400.0 2007600.0 1098600.0 2021400.0 ;
      RECT  1088400.0 2035200.0 1098600.0 2021400.0 ;
      RECT  1088400.0 2035200.0 1098600.0 2049000.0 ;
      RECT  1088400.0 2062800.0 1098600.0 2049000.0 ;
      RECT  1088400.0 2062800.0 1098600.0 2076600.0 ;
      RECT  1088400.0 2090400.0 1098600.0 2076600.0 ;
      RECT  1088400.0 2090400.0 1098600.0 2104200.0 ;
      RECT  1088400.0 2118000.0 1098600.0 2104200.0 ;
      RECT  1088400.0 2118000.0 1098600.0 2131800.0 ;
      RECT  1088400.0 2145600.0 1098600.0 2131800.0 ;
      RECT  1098600.0 379200.0 1108800.0 393000.0 ;
      RECT  1098600.0 406800.0 1108800.0 393000.0 ;
      RECT  1098600.0 406800.0 1108800.0 420600.0 ;
      RECT  1098600.0 434400.0 1108800.0 420600.0 ;
      RECT  1098600.0 434400.0 1108800.0 448200.0 ;
      RECT  1098600.0 462000.0 1108800.0 448200.0 ;
      RECT  1098600.0 462000.0 1108800.0 475800.0 ;
      RECT  1098600.0 489600.0 1108800.0 475800.0 ;
      RECT  1098600.0 489600.0 1108800.0 503400.0 ;
      RECT  1098600.0 517200.0 1108800.0 503400.0 ;
      RECT  1098600.0 517200.0 1108800.0 531000.0 ;
      RECT  1098600.0 544800.0 1108800.0 531000.0 ;
      RECT  1098600.0 544800.0 1108800.0 558600.0 ;
      RECT  1098600.0 572400.0 1108800.0 558600.0 ;
      RECT  1098600.0 572400.0 1108800.0 586200.0 ;
      RECT  1098600.0 600000.0 1108800.0 586200.0 ;
      RECT  1098600.0 600000.0 1108800.0 613800.0 ;
      RECT  1098600.0 627600.0 1108800.0 613800.0 ;
      RECT  1098600.0 627600.0 1108800.0 641400.0 ;
      RECT  1098600.0 655200.0 1108800.0 641400.0 ;
      RECT  1098600.0 655200.0 1108800.0 669000.0 ;
      RECT  1098600.0 682800.0 1108800.0 669000.0 ;
      RECT  1098600.0 682800.0 1108800.0 696600.0 ;
      RECT  1098600.0 710400.0 1108800.0 696600.0 ;
      RECT  1098600.0 710400.0 1108800.0 724200.0 ;
      RECT  1098600.0 738000.0 1108800.0 724200.0 ;
      RECT  1098600.0 738000.0 1108800.0 751800.0 ;
      RECT  1098600.0 765600.0 1108800.0 751800.0 ;
      RECT  1098600.0 765600.0 1108800.0 779400.0 ;
      RECT  1098600.0 793200.0 1108800.0 779400.0 ;
      RECT  1098600.0 793200.0 1108800.0 807000.0 ;
      RECT  1098600.0 820800.0 1108800.0 807000.0 ;
      RECT  1098600.0 820800.0 1108800.0 834600.0 ;
      RECT  1098600.0 848400.0 1108800.0 834600.0 ;
      RECT  1098600.0 848400.0 1108800.0 862200.0 ;
      RECT  1098600.0 876000.0 1108800.0 862200.0 ;
      RECT  1098600.0 876000.0 1108800.0 889800.0 ;
      RECT  1098600.0 903600.0 1108800.0 889800.0 ;
      RECT  1098600.0 903600.0 1108800.0 917400.0 ;
      RECT  1098600.0 931200.0 1108800.0 917400.0 ;
      RECT  1098600.0 931200.0 1108800.0 945000.0 ;
      RECT  1098600.0 958800.0 1108800.0 945000.0 ;
      RECT  1098600.0 958800.0 1108800.0 972600.0 ;
      RECT  1098600.0 986400.0 1108800.0 972600.0 ;
      RECT  1098600.0 986400.0 1108800.0 1000200.0 ;
      RECT  1098600.0 1014000.0 1108800.0 1000200.0 ;
      RECT  1098600.0 1014000.0 1108800.0 1027800.0 ;
      RECT  1098600.0 1041600.0 1108800.0 1027800.0 ;
      RECT  1098600.0 1041600.0 1108800.0 1055400.0 ;
      RECT  1098600.0 1069200.0 1108800.0 1055400.0 ;
      RECT  1098600.0 1069200.0 1108800.0 1083000.0 ;
      RECT  1098600.0 1096800.0 1108800.0 1083000.0 ;
      RECT  1098600.0 1096800.0 1108800.0 1110600.0 ;
      RECT  1098600.0 1124400.0 1108800.0 1110600.0 ;
      RECT  1098600.0 1124400.0 1108800.0 1138200.0 ;
      RECT  1098600.0 1152000.0 1108800.0 1138200.0 ;
      RECT  1098600.0 1152000.0 1108800.0 1165800.0 ;
      RECT  1098600.0 1179600.0 1108800.0 1165800.0 ;
      RECT  1098600.0 1179600.0 1108800.0 1193400.0 ;
      RECT  1098600.0 1207200.0 1108800.0 1193400.0 ;
      RECT  1098600.0 1207200.0 1108800.0 1221000.0 ;
      RECT  1098600.0 1234800.0 1108800.0 1221000.0 ;
      RECT  1098600.0 1234800.0 1108800.0 1248600.0 ;
      RECT  1098600.0 1262400.0 1108800.0 1248600.0 ;
      RECT  1098600.0 1262400.0 1108800.0 1276200.0 ;
      RECT  1098600.0 1290000.0 1108800.0 1276200.0 ;
      RECT  1098600.0 1290000.0 1108800.0 1303800.0 ;
      RECT  1098600.0 1317600.0 1108800.0 1303800.0 ;
      RECT  1098600.0 1317600.0 1108800.0 1331400.0 ;
      RECT  1098600.0 1345200.0 1108800.0 1331400.0 ;
      RECT  1098600.0 1345200.0 1108800.0 1359000.0 ;
      RECT  1098600.0 1372800.0 1108800.0 1359000.0 ;
      RECT  1098600.0 1372800.0 1108800.0 1386600.0 ;
      RECT  1098600.0 1400400.0 1108800.0 1386600.0 ;
      RECT  1098600.0 1400400.0 1108800.0 1414200.0 ;
      RECT  1098600.0 1428000.0 1108800.0 1414200.0 ;
      RECT  1098600.0 1428000.0 1108800.0 1441800.0 ;
      RECT  1098600.0 1455600.0 1108800.0 1441800.0 ;
      RECT  1098600.0 1455600.0 1108800.0 1469400.0 ;
      RECT  1098600.0 1483200.0 1108800.0 1469400.0 ;
      RECT  1098600.0 1483200.0 1108800.0 1497000.0 ;
      RECT  1098600.0 1510800.0 1108800.0 1497000.0 ;
      RECT  1098600.0 1510800.0 1108800.0 1524600.0 ;
      RECT  1098600.0 1538400.0 1108800.0 1524600.0 ;
      RECT  1098600.0 1538400.0 1108800.0 1552200.0 ;
      RECT  1098600.0 1566000.0 1108800.0 1552200.0 ;
      RECT  1098600.0 1566000.0 1108800.0 1579800.0 ;
      RECT  1098600.0 1593600.0 1108800.0 1579800.0 ;
      RECT  1098600.0 1593600.0 1108800.0 1607400.0 ;
      RECT  1098600.0 1621200.0 1108800.0 1607400.0 ;
      RECT  1098600.0 1621200.0 1108800.0 1635000.0 ;
      RECT  1098600.0 1648800.0 1108800.0 1635000.0 ;
      RECT  1098600.0 1648800.0 1108800.0 1662600.0 ;
      RECT  1098600.0 1676400.0 1108800.0 1662600.0 ;
      RECT  1098600.0 1676400.0 1108800.0 1690200.0 ;
      RECT  1098600.0 1704000.0 1108800.0 1690200.0 ;
      RECT  1098600.0 1704000.0 1108800.0 1717800.0 ;
      RECT  1098600.0 1731600.0 1108800.0 1717800.0 ;
      RECT  1098600.0 1731600.0 1108800.0 1745400.0 ;
      RECT  1098600.0 1759200.0 1108800.0 1745400.0 ;
      RECT  1098600.0 1759200.0 1108800.0 1773000.0 ;
      RECT  1098600.0 1786800.0 1108800.0 1773000.0 ;
      RECT  1098600.0 1786800.0 1108800.0 1800600.0 ;
      RECT  1098600.0 1814400.0 1108800.0 1800600.0 ;
      RECT  1098600.0 1814400.0 1108800.0 1828200.0 ;
      RECT  1098600.0 1842000.0 1108800.0 1828200.0 ;
      RECT  1098600.0 1842000.0 1108800.0 1855800.0 ;
      RECT  1098600.0 1869600.0 1108800.0 1855800.0 ;
      RECT  1098600.0 1869600.0 1108800.0 1883400.0 ;
      RECT  1098600.0 1897200.0 1108800.0 1883400.0 ;
      RECT  1098600.0 1897200.0 1108800.0 1911000.0 ;
      RECT  1098600.0 1924800.0 1108800.0 1911000.0 ;
      RECT  1098600.0 1924800.0 1108800.0 1938600.0 ;
      RECT  1098600.0 1952400.0 1108800.0 1938600.0 ;
      RECT  1098600.0 1952400.0 1108800.0 1966200.0 ;
      RECT  1098600.0 1980000.0 1108800.0 1966200.0 ;
      RECT  1098600.0 1980000.0 1108800.0 1993800.0 ;
      RECT  1098600.0 2007600.0 1108800.0 1993800.0 ;
      RECT  1098600.0 2007600.0 1108800.0 2021400.0 ;
      RECT  1098600.0 2035200.0 1108800.0 2021400.0 ;
      RECT  1098600.0 2035200.0 1108800.0 2049000.0 ;
      RECT  1098600.0 2062800.0 1108800.0 2049000.0 ;
      RECT  1098600.0 2062800.0 1108800.0 2076600.0 ;
      RECT  1098600.0 2090400.0 1108800.0 2076600.0 ;
      RECT  1098600.0 2090400.0 1108800.0 2104200.0 ;
      RECT  1098600.0 2118000.0 1108800.0 2104200.0 ;
      RECT  1098600.0 2118000.0 1108800.0 2131800.0 ;
      RECT  1098600.0 2145600.0 1108800.0 2131800.0 ;
      RECT  1108800.0 379200.0 1119000.0 393000.0 ;
      RECT  1108800.0 406800.0 1119000.0 393000.0 ;
      RECT  1108800.0 406800.0 1119000.0 420600.0 ;
      RECT  1108800.0 434400.0 1119000.0 420600.0 ;
      RECT  1108800.0 434400.0 1119000.0 448200.0 ;
      RECT  1108800.0 462000.0 1119000.0 448200.0 ;
      RECT  1108800.0 462000.0 1119000.0 475800.0 ;
      RECT  1108800.0 489600.0 1119000.0 475800.0 ;
      RECT  1108800.0 489600.0 1119000.0 503400.0 ;
      RECT  1108800.0 517200.0 1119000.0 503400.0 ;
      RECT  1108800.0 517200.0 1119000.0 531000.0 ;
      RECT  1108800.0 544800.0 1119000.0 531000.0 ;
      RECT  1108800.0 544800.0 1119000.0 558600.0 ;
      RECT  1108800.0 572400.0 1119000.0 558600.0 ;
      RECT  1108800.0 572400.0 1119000.0 586200.0 ;
      RECT  1108800.0 600000.0 1119000.0 586200.0 ;
      RECT  1108800.0 600000.0 1119000.0 613800.0 ;
      RECT  1108800.0 627600.0 1119000.0 613800.0 ;
      RECT  1108800.0 627600.0 1119000.0 641400.0 ;
      RECT  1108800.0 655200.0 1119000.0 641400.0 ;
      RECT  1108800.0 655200.0 1119000.0 669000.0 ;
      RECT  1108800.0 682800.0 1119000.0 669000.0 ;
      RECT  1108800.0 682800.0 1119000.0 696600.0 ;
      RECT  1108800.0 710400.0 1119000.0 696600.0 ;
      RECT  1108800.0 710400.0 1119000.0 724200.0 ;
      RECT  1108800.0 738000.0 1119000.0 724200.0 ;
      RECT  1108800.0 738000.0 1119000.0 751800.0 ;
      RECT  1108800.0 765600.0 1119000.0 751800.0 ;
      RECT  1108800.0 765600.0 1119000.0 779400.0 ;
      RECT  1108800.0 793200.0 1119000.0 779400.0 ;
      RECT  1108800.0 793200.0 1119000.0 807000.0 ;
      RECT  1108800.0 820800.0 1119000.0 807000.0 ;
      RECT  1108800.0 820800.0 1119000.0 834600.0 ;
      RECT  1108800.0 848400.0 1119000.0 834600.0 ;
      RECT  1108800.0 848400.0 1119000.0 862200.0 ;
      RECT  1108800.0 876000.0 1119000.0 862200.0 ;
      RECT  1108800.0 876000.0 1119000.0 889800.0 ;
      RECT  1108800.0 903600.0 1119000.0 889800.0 ;
      RECT  1108800.0 903600.0 1119000.0 917400.0 ;
      RECT  1108800.0 931200.0 1119000.0 917400.0 ;
      RECT  1108800.0 931200.0 1119000.0 945000.0 ;
      RECT  1108800.0 958800.0 1119000.0 945000.0 ;
      RECT  1108800.0 958800.0 1119000.0 972600.0 ;
      RECT  1108800.0 986400.0 1119000.0 972600.0 ;
      RECT  1108800.0 986400.0 1119000.0 1000200.0 ;
      RECT  1108800.0 1014000.0 1119000.0 1000200.0 ;
      RECT  1108800.0 1014000.0 1119000.0 1027800.0 ;
      RECT  1108800.0 1041600.0 1119000.0 1027800.0 ;
      RECT  1108800.0 1041600.0 1119000.0 1055400.0 ;
      RECT  1108800.0 1069200.0 1119000.0 1055400.0 ;
      RECT  1108800.0 1069200.0 1119000.0 1083000.0 ;
      RECT  1108800.0 1096800.0 1119000.0 1083000.0 ;
      RECT  1108800.0 1096800.0 1119000.0 1110600.0 ;
      RECT  1108800.0 1124400.0 1119000.0 1110600.0 ;
      RECT  1108800.0 1124400.0 1119000.0 1138200.0 ;
      RECT  1108800.0 1152000.0 1119000.0 1138200.0 ;
      RECT  1108800.0 1152000.0 1119000.0 1165800.0 ;
      RECT  1108800.0 1179600.0 1119000.0 1165800.0 ;
      RECT  1108800.0 1179600.0 1119000.0 1193400.0 ;
      RECT  1108800.0 1207200.0 1119000.0 1193400.0 ;
      RECT  1108800.0 1207200.0 1119000.0 1221000.0 ;
      RECT  1108800.0 1234800.0 1119000.0 1221000.0 ;
      RECT  1108800.0 1234800.0 1119000.0 1248600.0 ;
      RECT  1108800.0 1262400.0 1119000.0 1248600.0 ;
      RECT  1108800.0 1262400.0 1119000.0 1276200.0 ;
      RECT  1108800.0 1290000.0 1119000.0 1276200.0 ;
      RECT  1108800.0 1290000.0 1119000.0 1303800.0 ;
      RECT  1108800.0 1317600.0 1119000.0 1303800.0 ;
      RECT  1108800.0 1317600.0 1119000.0 1331400.0 ;
      RECT  1108800.0 1345200.0 1119000.0 1331400.0 ;
      RECT  1108800.0 1345200.0 1119000.0 1359000.0 ;
      RECT  1108800.0 1372800.0 1119000.0 1359000.0 ;
      RECT  1108800.0 1372800.0 1119000.0 1386600.0 ;
      RECT  1108800.0 1400400.0 1119000.0 1386600.0 ;
      RECT  1108800.0 1400400.0 1119000.0 1414200.0 ;
      RECT  1108800.0 1428000.0 1119000.0 1414200.0 ;
      RECT  1108800.0 1428000.0 1119000.0 1441800.0 ;
      RECT  1108800.0 1455600.0 1119000.0 1441800.0 ;
      RECT  1108800.0 1455600.0 1119000.0 1469400.0 ;
      RECT  1108800.0 1483200.0 1119000.0 1469400.0 ;
      RECT  1108800.0 1483200.0 1119000.0 1497000.0 ;
      RECT  1108800.0 1510800.0 1119000.0 1497000.0 ;
      RECT  1108800.0 1510800.0 1119000.0 1524600.0 ;
      RECT  1108800.0 1538400.0 1119000.0 1524600.0 ;
      RECT  1108800.0 1538400.0 1119000.0 1552200.0 ;
      RECT  1108800.0 1566000.0 1119000.0 1552200.0 ;
      RECT  1108800.0 1566000.0 1119000.0 1579800.0 ;
      RECT  1108800.0 1593600.0 1119000.0 1579800.0 ;
      RECT  1108800.0 1593600.0 1119000.0 1607400.0 ;
      RECT  1108800.0 1621200.0 1119000.0 1607400.0 ;
      RECT  1108800.0 1621200.0 1119000.0 1635000.0 ;
      RECT  1108800.0 1648800.0 1119000.0 1635000.0 ;
      RECT  1108800.0 1648800.0 1119000.0 1662600.0 ;
      RECT  1108800.0 1676400.0 1119000.0 1662600.0 ;
      RECT  1108800.0 1676400.0 1119000.0 1690200.0 ;
      RECT  1108800.0 1704000.0 1119000.0 1690200.0 ;
      RECT  1108800.0 1704000.0 1119000.0 1717800.0 ;
      RECT  1108800.0 1731600.0 1119000.0 1717800.0 ;
      RECT  1108800.0 1731600.0 1119000.0 1745400.0 ;
      RECT  1108800.0 1759200.0 1119000.0 1745400.0 ;
      RECT  1108800.0 1759200.0 1119000.0 1773000.0 ;
      RECT  1108800.0 1786800.0 1119000.0 1773000.0 ;
      RECT  1108800.0 1786800.0 1119000.0 1800600.0 ;
      RECT  1108800.0 1814400.0 1119000.0 1800600.0 ;
      RECT  1108800.0 1814400.0 1119000.0 1828200.0 ;
      RECT  1108800.0 1842000.0 1119000.0 1828200.0 ;
      RECT  1108800.0 1842000.0 1119000.0 1855800.0 ;
      RECT  1108800.0 1869600.0 1119000.0 1855800.0 ;
      RECT  1108800.0 1869600.0 1119000.0 1883400.0 ;
      RECT  1108800.0 1897200.0 1119000.0 1883400.0 ;
      RECT  1108800.0 1897200.0 1119000.0 1911000.0 ;
      RECT  1108800.0 1924800.0 1119000.0 1911000.0 ;
      RECT  1108800.0 1924800.0 1119000.0 1938600.0 ;
      RECT  1108800.0 1952400.0 1119000.0 1938600.0 ;
      RECT  1108800.0 1952400.0 1119000.0 1966200.0 ;
      RECT  1108800.0 1980000.0 1119000.0 1966200.0 ;
      RECT  1108800.0 1980000.0 1119000.0 1993800.0 ;
      RECT  1108800.0 2007600.0 1119000.0 1993800.0 ;
      RECT  1108800.0 2007600.0 1119000.0 2021400.0 ;
      RECT  1108800.0 2035200.0 1119000.0 2021400.0 ;
      RECT  1108800.0 2035200.0 1119000.0 2049000.0 ;
      RECT  1108800.0 2062800.0 1119000.0 2049000.0 ;
      RECT  1108800.0 2062800.0 1119000.0 2076600.0 ;
      RECT  1108800.0 2090400.0 1119000.0 2076600.0 ;
      RECT  1108800.0 2090400.0 1119000.0 2104200.0 ;
      RECT  1108800.0 2118000.0 1119000.0 2104200.0 ;
      RECT  1108800.0 2118000.0 1119000.0 2131800.0 ;
      RECT  1108800.0 2145600.0 1119000.0 2131800.0 ;
      RECT  1119000.0 379200.0 1129200.0 393000.0 ;
      RECT  1119000.0 406800.0 1129200.0 393000.0 ;
      RECT  1119000.0 406800.0 1129200.0 420600.0 ;
      RECT  1119000.0 434400.0 1129200.0 420600.0 ;
      RECT  1119000.0 434400.0 1129200.0 448200.0 ;
      RECT  1119000.0 462000.0 1129200.0 448200.0 ;
      RECT  1119000.0 462000.0 1129200.0 475800.0 ;
      RECT  1119000.0 489600.0 1129200.0 475800.0 ;
      RECT  1119000.0 489600.0 1129200.0 503400.0 ;
      RECT  1119000.0 517200.0 1129200.0 503400.0 ;
      RECT  1119000.0 517200.0 1129200.0 531000.0 ;
      RECT  1119000.0 544800.0 1129200.0 531000.0 ;
      RECT  1119000.0 544800.0 1129200.0 558600.0 ;
      RECT  1119000.0 572400.0 1129200.0 558600.0 ;
      RECT  1119000.0 572400.0 1129200.0 586200.0 ;
      RECT  1119000.0 600000.0 1129200.0 586200.0 ;
      RECT  1119000.0 600000.0 1129200.0 613800.0 ;
      RECT  1119000.0 627600.0 1129200.0 613800.0 ;
      RECT  1119000.0 627600.0 1129200.0 641400.0 ;
      RECT  1119000.0 655200.0 1129200.0 641400.0 ;
      RECT  1119000.0 655200.0 1129200.0 669000.0 ;
      RECT  1119000.0 682800.0 1129200.0 669000.0 ;
      RECT  1119000.0 682800.0 1129200.0 696600.0 ;
      RECT  1119000.0 710400.0 1129200.0 696600.0 ;
      RECT  1119000.0 710400.0 1129200.0 724200.0 ;
      RECT  1119000.0 738000.0 1129200.0 724200.0 ;
      RECT  1119000.0 738000.0 1129200.0 751800.0 ;
      RECT  1119000.0 765600.0 1129200.0 751800.0 ;
      RECT  1119000.0 765600.0 1129200.0 779400.0 ;
      RECT  1119000.0 793200.0 1129200.0 779400.0 ;
      RECT  1119000.0 793200.0 1129200.0 807000.0 ;
      RECT  1119000.0 820800.0 1129200.0 807000.0 ;
      RECT  1119000.0 820800.0 1129200.0 834600.0 ;
      RECT  1119000.0 848400.0 1129200.0 834600.0 ;
      RECT  1119000.0 848400.0 1129200.0 862200.0 ;
      RECT  1119000.0 876000.0 1129200.0 862200.0 ;
      RECT  1119000.0 876000.0 1129200.0 889800.0 ;
      RECT  1119000.0 903600.0 1129200.0 889800.0 ;
      RECT  1119000.0 903600.0 1129200.0 917400.0 ;
      RECT  1119000.0 931200.0 1129200.0 917400.0 ;
      RECT  1119000.0 931200.0 1129200.0 945000.0 ;
      RECT  1119000.0 958800.0 1129200.0 945000.0 ;
      RECT  1119000.0 958800.0 1129200.0 972600.0 ;
      RECT  1119000.0 986400.0 1129200.0 972600.0 ;
      RECT  1119000.0 986400.0 1129200.0 1000200.0 ;
      RECT  1119000.0 1014000.0 1129200.0 1000200.0 ;
      RECT  1119000.0 1014000.0 1129200.0 1027800.0 ;
      RECT  1119000.0 1041600.0 1129200.0 1027800.0 ;
      RECT  1119000.0 1041600.0 1129200.0 1055400.0 ;
      RECT  1119000.0 1069200.0 1129200.0 1055400.0 ;
      RECT  1119000.0 1069200.0 1129200.0 1083000.0 ;
      RECT  1119000.0 1096800.0 1129200.0 1083000.0 ;
      RECT  1119000.0 1096800.0 1129200.0 1110600.0 ;
      RECT  1119000.0 1124400.0 1129200.0 1110600.0 ;
      RECT  1119000.0 1124400.0 1129200.0 1138200.0 ;
      RECT  1119000.0 1152000.0 1129200.0 1138200.0 ;
      RECT  1119000.0 1152000.0 1129200.0 1165800.0 ;
      RECT  1119000.0 1179600.0 1129200.0 1165800.0 ;
      RECT  1119000.0 1179600.0 1129200.0 1193400.0 ;
      RECT  1119000.0 1207200.0 1129200.0 1193400.0 ;
      RECT  1119000.0 1207200.0 1129200.0 1221000.0 ;
      RECT  1119000.0 1234800.0 1129200.0 1221000.0 ;
      RECT  1119000.0 1234800.0 1129200.0 1248600.0 ;
      RECT  1119000.0 1262400.0 1129200.0 1248600.0 ;
      RECT  1119000.0 1262400.0 1129200.0 1276200.0 ;
      RECT  1119000.0 1290000.0 1129200.0 1276200.0 ;
      RECT  1119000.0 1290000.0 1129200.0 1303800.0 ;
      RECT  1119000.0 1317600.0 1129200.0 1303800.0 ;
      RECT  1119000.0 1317600.0 1129200.0 1331400.0 ;
      RECT  1119000.0 1345200.0 1129200.0 1331400.0 ;
      RECT  1119000.0 1345200.0 1129200.0 1359000.0 ;
      RECT  1119000.0 1372800.0 1129200.0 1359000.0 ;
      RECT  1119000.0 1372800.0 1129200.0 1386600.0 ;
      RECT  1119000.0 1400400.0 1129200.0 1386600.0 ;
      RECT  1119000.0 1400400.0 1129200.0 1414200.0 ;
      RECT  1119000.0 1428000.0 1129200.0 1414200.0 ;
      RECT  1119000.0 1428000.0 1129200.0 1441800.0 ;
      RECT  1119000.0 1455600.0 1129200.0 1441800.0 ;
      RECT  1119000.0 1455600.0 1129200.0 1469400.0 ;
      RECT  1119000.0 1483200.0 1129200.0 1469400.0 ;
      RECT  1119000.0 1483200.0 1129200.0 1497000.0 ;
      RECT  1119000.0 1510800.0 1129200.0 1497000.0 ;
      RECT  1119000.0 1510800.0 1129200.0 1524600.0 ;
      RECT  1119000.0 1538400.0 1129200.0 1524600.0 ;
      RECT  1119000.0 1538400.0 1129200.0 1552200.0 ;
      RECT  1119000.0 1566000.0 1129200.0 1552200.0 ;
      RECT  1119000.0 1566000.0 1129200.0 1579800.0 ;
      RECT  1119000.0 1593600.0 1129200.0 1579800.0 ;
      RECT  1119000.0 1593600.0 1129200.0 1607400.0 ;
      RECT  1119000.0 1621200.0 1129200.0 1607400.0 ;
      RECT  1119000.0 1621200.0 1129200.0 1635000.0 ;
      RECT  1119000.0 1648800.0 1129200.0 1635000.0 ;
      RECT  1119000.0 1648800.0 1129200.0 1662600.0 ;
      RECT  1119000.0 1676400.0 1129200.0 1662600.0 ;
      RECT  1119000.0 1676400.0 1129200.0 1690200.0 ;
      RECT  1119000.0 1704000.0 1129200.0 1690200.0 ;
      RECT  1119000.0 1704000.0 1129200.0 1717800.0 ;
      RECT  1119000.0 1731600.0 1129200.0 1717800.0 ;
      RECT  1119000.0 1731600.0 1129200.0 1745400.0 ;
      RECT  1119000.0 1759200.0 1129200.0 1745400.0 ;
      RECT  1119000.0 1759200.0 1129200.0 1773000.0 ;
      RECT  1119000.0 1786800.0 1129200.0 1773000.0 ;
      RECT  1119000.0 1786800.0 1129200.0 1800600.0 ;
      RECT  1119000.0 1814400.0 1129200.0 1800600.0 ;
      RECT  1119000.0 1814400.0 1129200.0 1828200.0 ;
      RECT  1119000.0 1842000.0 1129200.0 1828200.0 ;
      RECT  1119000.0 1842000.0 1129200.0 1855800.0 ;
      RECT  1119000.0 1869600.0 1129200.0 1855800.0 ;
      RECT  1119000.0 1869600.0 1129200.0 1883400.0 ;
      RECT  1119000.0 1897200.0 1129200.0 1883400.0 ;
      RECT  1119000.0 1897200.0 1129200.0 1911000.0 ;
      RECT  1119000.0 1924800.0 1129200.0 1911000.0 ;
      RECT  1119000.0 1924800.0 1129200.0 1938600.0 ;
      RECT  1119000.0 1952400.0 1129200.0 1938600.0 ;
      RECT  1119000.0 1952400.0 1129200.0 1966200.0 ;
      RECT  1119000.0 1980000.0 1129200.0 1966200.0 ;
      RECT  1119000.0 1980000.0 1129200.0 1993800.0 ;
      RECT  1119000.0 2007600.0 1129200.0 1993800.0 ;
      RECT  1119000.0 2007600.0 1129200.0 2021400.0 ;
      RECT  1119000.0 2035200.0 1129200.0 2021400.0 ;
      RECT  1119000.0 2035200.0 1129200.0 2049000.0 ;
      RECT  1119000.0 2062800.0 1129200.0 2049000.0 ;
      RECT  1119000.0 2062800.0 1129200.0 2076600.0 ;
      RECT  1119000.0 2090400.0 1129200.0 2076600.0 ;
      RECT  1119000.0 2090400.0 1129200.0 2104200.0 ;
      RECT  1119000.0 2118000.0 1129200.0 2104200.0 ;
      RECT  1119000.0 2118000.0 1129200.0 2131800.0 ;
      RECT  1119000.0 2145600.0 1129200.0 2131800.0 ;
      RECT  1129200.0 379200.0 1139400.0 393000.0 ;
      RECT  1129200.0 406800.0 1139400.0 393000.0 ;
      RECT  1129200.0 406800.0 1139400.0 420600.0 ;
      RECT  1129200.0 434400.0 1139400.0 420600.0 ;
      RECT  1129200.0 434400.0 1139400.0 448200.0 ;
      RECT  1129200.0 462000.0 1139400.0 448200.0 ;
      RECT  1129200.0 462000.0 1139400.0 475800.0 ;
      RECT  1129200.0 489600.0 1139400.0 475800.0 ;
      RECT  1129200.0 489600.0 1139400.0 503400.0 ;
      RECT  1129200.0 517200.0 1139400.0 503400.0 ;
      RECT  1129200.0 517200.0 1139400.0 531000.0 ;
      RECT  1129200.0 544800.0 1139400.0 531000.0 ;
      RECT  1129200.0 544800.0 1139400.0 558600.0 ;
      RECT  1129200.0 572400.0 1139400.0 558600.0 ;
      RECT  1129200.0 572400.0 1139400.0 586200.0 ;
      RECT  1129200.0 600000.0 1139400.0 586200.0 ;
      RECT  1129200.0 600000.0 1139400.0 613800.0 ;
      RECT  1129200.0 627600.0 1139400.0 613800.0 ;
      RECT  1129200.0 627600.0 1139400.0 641400.0 ;
      RECT  1129200.0 655200.0 1139400.0 641400.0 ;
      RECT  1129200.0 655200.0 1139400.0 669000.0 ;
      RECT  1129200.0 682800.0 1139400.0 669000.0 ;
      RECT  1129200.0 682800.0 1139400.0 696600.0 ;
      RECT  1129200.0 710400.0 1139400.0 696600.0 ;
      RECT  1129200.0 710400.0 1139400.0 724200.0 ;
      RECT  1129200.0 738000.0 1139400.0 724200.0 ;
      RECT  1129200.0 738000.0 1139400.0 751800.0 ;
      RECT  1129200.0 765600.0 1139400.0 751800.0 ;
      RECT  1129200.0 765600.0 1139400.0 779400.0 ;
      RECT  1129200.0 793200.0 1139400.0 779400.0 ;
      RECT  1129200.0 793200.0 1139400.0 807000.0 ;
      RECT  1129200.0 820800.0 1139400.0 807000.0 ;
      RECT  1129200.0 820800.0 1139400.0 834600.0 ;
      RECT  1129200.0 848400.0 1139400.0 834600.0 ;
      RECT  1129200.0 848400.0 1139400.0 862200.0 ;
      RECT  1129200.0 876000.0 1139400.0 862200.0 ;
      RECT  1129200.0 876000.0 1139400.0 889800.0 ;
      RECT  1129200.0 903600.0 1139400.0 889800.0 ;
      RECT  1129200.0 903600.0 1139400.0 917400.0 ;
      RECT  1129200.0 931200.0 1139400.0 917400.0 ;
      RECT  1129200.0 931200.0 1139400.0 945000.0 ;
      RECT  1129200.0 958800.0 1139400.0 945000.0 ;
      RECT  1129200.0 958800.0 1139400.0 972600.0 ;
      RECT  1129200.0 986400.0 1139400.0 972600.0 ;
      RECT  1129200.0 986400.0 1139400.0 1000200.0 ;
      RECT  1129200.0 1014000.0 1139400.0 1000200.0 ;
      RECT  1129200.0 1014000.0 1139400.0 1027800.0 ;
      RECT  1129200.0 1041600.0 1139400.0 1027800.0 ;
      RECT  1129200.0 1041600.0 1139400.0 1055400.0 ;
      RECT  1129200.0 1069200.0 1139400.0 1055400.0 ;
      RECT  1129200.0 1069200.0 1139400.0 1083000.0 ;
      RECT  1129200.0 1096800.0 1139400.0 1083000.0 ;
      RECT  1129200.0 1096800.0 1139400.0 1110600.0 ;
      RECT  1129200.0 1124400.0 1139400.0 1110600.0 ;
      RECT  1129200.0 1124400.0 1139400.0 1138200.0 ;
      RECT  1129200.0 1152000.0 1139400.0 1138200.0 ;
      RECT  1129200.0 1152000.0 1139400.0 1165800.0 ;
      RECT  1129200.0 1179600.0 1139400.0 1165800.0 ;
      RECT  1129200.0 1179600.0 1139400.0 1193400.0 ;
      RECT  1129200.0 1207200.0 1139400.0 1193400.0 ;
      RECT  1129200.0 1207200.0 1139400.0 1221000.0 ;
      RECT  1129200.0 1234800.0 1139400.0 1221000.0 ;
      RECT  1129200.0 1234800.0 1139400.0 1248600.0 ;
      RECT  1129200.0 1262400.0 1139400.0 1248600.0 ;
      RECT  1129200.0 1262400.0 1139400.0 1276200.0 ;
      RECT  1129200.0 1290000.0 1139400.0 1276200.0 ;
      RECT  1129200.0 1290000.0 1139400.0 1303800.0 ;
      RECT  1129200.0 1317600.0 1139400.0 1303800.0 ;
      RECT  1129200.0 1317600.0 1139400.0 1331400.0 ;
      RECT  1129200.0 1345200.0 1139400.0 1331400.0 ;
      RECT  1129200.0 1345200.0 1139400.0 1359000.0 ;
      RECT  1129200.0 1372800.0 1139400.0 1359000.0 ;
      RECT  1129200.0 1372800.0 1139400.0 1386600.0 ;
      RECT  1129200.0 1400400.0 1139400.0 1386600.0 ;
      RECT  1129200.0 1400400.0 1139400.0 1414200.0 ;
      RECT  1129200.0 1428000.0 1139400.0 1414200.0 ;
      RECT  1129200.0 1428000.0 1139400.0 1441800.0 ;
      RECT  1129200.0 1455600.0 1139400.0 1441800.0 ;
      RECT  1129200.0 1455600.0 1139400.0 1469400.0 ;
      RECT  1129200.0 1483200.0 1139400.0 1469400.0 ;
      RECT  1129200.0 1483200.0 1139400.0 1497000.0 ;
      RECT  1129200.0 1510800.0 1139400.0 1497000.0 ;
      RECT  1129200.0 1510800.0 1139400.0 1524600.0 ;
      RECT  1129200.0 1538400.0 1139400.0 1524600.0 ;
      RECT  1129200.0 1538400.0 1139400.0 1552200.0 ;
      RECT  1129200.0 1566000.0 1139400.0 1552200.0 ;
      RECT  1129200.0 1566000.0 1139400.0 1579800.0 ;
      RECT  1129200.0 1593600.0 1139400.0 1579800.0 ;
      RECT  1129200.0 1593600.0 1139400.0 1607400.0 ;
      RECT  1129200.0 1621200.0 1139400.0 1607400.0 ;
      RECT  1129200.0 1621200.0 1139400.0 1635000.0 ;
      RECT  1129200.0 1648800.0 1139400.0 1635000.0 ;
      RECT  1129200.0 1648800.0 1139400.0 1662600.0 ;
      RECT  1129200.0 1676400.0 1139400.0 1662600.0 ;
      RECT  1129200.0 1676400.0 1139400.0 1690200.0 ;
      RECT  1129200.0 1704000.0 1139400.0 1690200.0 ;
      RECT  1129200.0 1704000.0 1139400.0 1717800.0 ;
      RECT  1129200.0 1731600.0 1139400.0 1717800.0 ;
      RECT  1129200.0 1731600.0 1139400.0 1745400.0 ;
      RECT  1129200.0 1759200.0 1139400.0 1745400.0 ;
      RECT  1129200.0 1759200.0 1139400.0 1773000.0 ;
      RECT  1129200.0 1786800.0 1139400.0 1773000.0 ;
      RECT  1129200.0 1786800.0 1139400.0 1800600.0 ;
      RECT  1129200.0 1814400.0 1139400.0 1800600.0 ;
      RECT  1129200.0 1814400.0 1139400.0 1828200.0 ;
      RECT  1129200.0 1842000.0 1139400.0 1828200.0 ;
      RECT  1129200.0 1842000.0 1139400.0 1855800.0 ;
      RECT  1129200.0 1869600.0 1139400.0 1855800.0 ;
      RECT  1129200.0 1869600.0 1139400.0 1883400.0 ;
      RECT  1129200.0 1897200.0 1139400.0 1883400.0 ;
      RECT  1129200.0 1897200.0 1139400.0 1911000.0 ;
      RECT  1129200.0 1924800.0 1139400.0 1911000.0 ;
      RECT  1129200.0 1924800.0 1139400.0 1938600.0 ;
      RECT  1129200.0 1952400.0 1139400.0 1938600.0 ;
      RECT  1129200.0 1952400.0 1139400.0 1966200.0 ;
      RECT  1129200.0 1980000.0 1139400.0 1966200.0 ;
      RECT  1129200.0 1980000.0 1139400.0 1993800.0 ;
      RECT  1129200.0 2007600.0 1139400.0 1993800.0 ;
      RECT  1129200.0 2007600.0 1139400.0 2021400.0 ;
      RECT  1129200.0 2035200.0 1139400.0 2021400.0 ;
      RECT  1129200.0 2035200.0 1139400.0 2049000.0 ;
      RECT  1129200.0 2062800.0 1139400.0 2049000.0 ;
      RECT  1129200.0 2062800.0 1139400.0 2076600.0 ;
      RECT  1129200.0 2090400.0 1139400.0 2076600.0 ;
      RECT  1129200.0 2090400.0 1139400.0 2104200.0 ;
      RECT  1129200.0 2118000.0 1139400.0 2104200.0 ;
      RECT  1129200.0 2118000.0 1139400.0 2131800.0 ;
      RECT  1129200.0 2145600.0 1139400.0 2131800.0 ;
      RECT  1139400.0 379200.0 1149600.0 393000.0 ;
      RECT  1139400.0 406800.0 1149600.0 393000.0 ;
      RECT  1139400.0 406800.0 1149600.0 420600.0 ;
      RECT  1139400.0 434400.0 1149600.0 420600.0 ;
      RECT  1139400.0 434400.0 1149600.0 448200.0 ;
      RECT  1139400.0 462000.0 1149600.0 448200.0 ;
      RECT  1139400.0 462000.0 1149600.0 475800.0 ;
      RECT  1139400.0 489600.0 1149600.0 475800.0 ;
      RECT  1139400.0 489600.0 1149600.0 503400.0 ;
      RECT  1139400.0 517200.0 1149600.0 503400.0 ;
      RECT  1139400.0 517200.0 1149600.0 531000.0 ;
      RECT  1139400.0 544800.0 1149600.0 531000.0 ;
      RECT  1139400.0 544800.0 1149600.0 558600.0 ;
      RECT  1139400.0 572400.0 1149600.0 558600.0 ;
      RECT  1139400.0 572400.0 1149600.0 586200.0 ;
      RECT  1139400.0 600000.0 1149600.0 586200.0 ;
      RECT  1139400.0 600000.0 1149600.0 613800.0 ;
      RECT  1139400.0 627600.0 1149600.0 613800.0 ;
      RECT  1139400.0 627600.0 1149600.0 641400.0 ;
      RECT  1139400.0 655200.0 1149600.0 641400.0 ;
      RECT  1139400.0 655200.0 1149600.0 669000.0 ;
      RECT  1139400.0 682800.0 1149600.0 669000.0 ;
      RECT  1139400.0 682800.0 1149600.0 696600.0 ;
      RECT  1139400.0 710400.0 1149600.0 696600.0 ;
      RECT  1139400.0 710400.0 1149600.0 724200.0 ;
      RECT  1139400.0 738000.0 1149600.0 724200.0 ;
      RECT  1139400.0 738000.0 1149600.0 751800.0 ;
      RECT  1139400.0 765600.0 1149600.0 751800.0 ;
      RECT  1139400.0 765600.0 1149600.0 779400.0 ;
      RECT  1139400.0 793200.0 1149600.0 779400.0 ;
      RECT  1139400.0 793200.0 1149600.0 807000.0 ;
      RECT  1139400.0 820800.0 1149600.0 807000.0 ;
      RECT  1139400.0 820800.0 1149600.0 834600.0 ;
      RECT  1139400.0 848400.0 1149600.0 834600.0 ;
      RECT  1139400.0 848400.0 1149600.0 862200.0 ;
      RECT  1139400.0 876000.0 1149600.0 862200.0 ;
      RECT  1139400.0 876000.0 1149600.0 889800.0 ;
      RECT  1139400.0 903600.0 1149600.0 889800.0 ;
      RECT  1139400.0 903600.0 1149600.0 917400.0 ;
      RECT  1139400.0 931200.0 1149600.0 917400.0 ;
      RECT  1139400.0 931200.0 1149600.0 945000.0 ;
      RECT  1139400.0 958800.0 1149600.0 945000.0 ;
      RECT  1139400.0 958800.0 1149600.0 972600.0 ;
      RECT  1139400.0 986400.0 1149600.0 972600.0 ;
      RECT  1139400.0 986400.0 1149600.0 1000200.0 ;
      RECT  1139400.0 1014000.0 1149600.0 1000200.0 ;
      RECT  1139400.0 1014000.0 1149600.0 1027800.0 ;
      RECT  1139400.0 1041600.0 1149600.0 1027800.0 ;
      RECT  1139400.0 1041600.0 1149600.0 1055400.0 ;
      RECT  1139400.0 1069200.0 1149600.0 1055400.0 ;
      RECT  1139400.0 1069200.0 1149600.0 1083000.0 ;
      RECT  1139400.0 1096800.0 1149600.0 1083000.0 ;
      RECT  1139400.0 1096800.0 1149600.0 1110600.0 ;
      RECT  1139400.0 1124400.0 1149600.0 1110600.0 ;
      RECT  1139400.0 1124400.0 1149600.0 1138200.0 ;
      RECT  1139400.0 1152000.0 1149600.0 1138200.0 ;
      RECT  1139400.0 1152000.0 1149600.0 1165800.0 ;
      RECT  1139400.0 1179600.0 1149600.0 1165800.0 ;
      RECT  1139400.0 1179600.0 1149600.0 1193400.0 ;
      RECT  1139400.0 1207200.0 1149600.0 1193400.0 ;
      RECT  1139400.0 1207200.0 1149600.0 1221000.0 ;
      RECT  1139400.0 1234800.0 1149600.0 1221000.0 ;
      RECT  1139400.0 1234800.0 1149600.0 1248600.0 ;
      RECT  1139400.0 1262400.0 1149600.0 1248600.0 ;
      RECT  1139400.0 1262400.0 1149600.0 1276200.0 ;
      RECT  1139400.0 1290000.0 1149600.0 1276200.0 ;
      RECT  1139400.0 1290000.0 1149600.0 1303800.0 ;
      RECT  1139400.0 1317600.0 1149600.0 1303800.0 ;
      RECT  1139400.0 1317600.0 1149600.0 1331400.0 ;
      RECT  1139400.0 1345200.0 1149600.0 1331400.0 ;
      RECT  1139400.0 1345200.0 1149600.0 1359000.0 ;
      RECT  1139400.0 1372800.0 1149600.0 1359000.0 ;
      RECT  1139400.0 1372800.0 1149600.0 1386600.0 ;
      RECT  1139400.0 1400400.0 1149600.0 1386600.0 ;
      RECT  1139400.0 1400400.0 1149600.0 1414200.0 ;
      RECT  1139400.0 1428000.0 1149600.0 1414200.0 ;
      RECT  1139400.0 1428000.0 1149600.0 1441800.0 ;
      RECT  1139400.0 1455600.0 1149600.0 1441800.0 ;
      RECT  1139400.0 1455600.0 1149600.0 1469400.0 ;
      RECT  1139400.0 1483200.0 1149600.0 1469400.0 ;
      RECT  1139400.0 1483200.0 1149600.0 1497000.0 ;
      RECT  1139400.0 1510800.0 1149600.0 1497000.0 ;
      RECT  1139400.0 1510800.0 1149600.0 1524600.0 ;
      RECT  1139400.0 1538400.0 1149600.0 1524600.0 ;
      RECT  1139400.0 1538400.0 1149600.0 1552200.0 ;
      RECT  1139400.0 1566000.0 1149600.0 1552200.0 ;
      RECT  1139400.0 1566000.0 1149600.0 1579800.0 ;
      RECT  1139400.0 1593600.0 1149600.0 1579800.0 ;
      RECT  1139400.0 1593600.0 1149600.0 1607400.0 ;
      RECT  1139400.0 1621200.0 1149600.0 1607400.0 ;
      RECT  1139400.0 1621200.0 1149600.0 1635000.0 ;
      RECT  1139400.0 1648800.0 1149600.0 1635000.0 ;
      RECT  1139400.0 1648800.0 1149600.0 1662600.0 ;
      RECT  1139400.0 1676400.0 1149600.0 1662600.0 ;
      RECT  1139400.0 1676400.0 1149600.0 1690200.0 ;
      RECT  1139400.0 1704000.0 1149600.0 1690200.0 ;
      RECT  1139400.0 1704000.0 1149600.0 1717800.0 ;
      RECT  1139400.0 1731600.0 1149600.0 1717800.0 ;
      RECT  1139400.0 1731600.0 1149600.0 1745400.0 ;
      RECT  1139400.0 1759200.0 1149600.0 1745400.0 ;
      RECT  1139400.0 1759200.0 1149600.0 1773000.0 ;
      RECT  1139400.0 1786800.0 1149600.0 1773000.0 ;
      RECT  1139400.0 1786800.0 1149600.0 1800600.0 ;
      RECT  1139400.0 1814400.0 1149600.0 1800600.0 ;
      RECT  1139400.0 1814400.0 1149600.0 1828200.0 ;
      RECT  1139400.0 1842000.0 1149600.0 1828200.0 ;
      RECT  1139400.0 1842000.0 1149600.0 1855800.0 ;
      RECT  1139400.0 1869600.0 1149600.0 1855800.0 ;
      RECT  1139400.0 1869600.0 1149600.0 1883400.0 ;
      RECT  1139400.0 1897200.0 1149600.0 1883400.0 ;
      RECT  1139400.0 1897200.0 1149600.0 1911000.0 ;
      RECT  1139400.0 1924800.0 1149600.0 1911000.0 ;
      RECT  1139400.0 1924800.0 1149600.0 1938600.0 ;
      RECT  1139400.0 1952400.0 1149600.0 1938600.0 ;
      RECT  1139400.0 1952400.0 1149600.0 1966200.0 ;
      RECT  1139400.0 1980000.0 1149600.0 1966200.0 ;
      RECT  1139400.0 1980000.0 1149600.0 1993800.0 ;
      RECT  1139400.0 2007600.0 1149600.0 1993800.0 ;
      RECT  1139400.0 2007600.0 1149600.0 2021400.0 ;
      RECT  1139400.0 2035200.0 1149600.0 2021400.0 ;
      RECT  1139400.0 2035200.0 1149600.0 2049000.0 ;
      RECT  1139400.0 2062800.0 1149600.0 2049000.0 ;
      RECT  1139400.0 2062800.0 1149600.0 2076600.0 ;
      RECT  1139400.0 2090400.0 1149600.0 2076600.0 ;
      RECT  1139400.0 2090400.0 1149600.0 2104200.0 ;
      RECT  1139400.0 2118000.0 1149600.0 2104200.0 ;
      RECT  1139400.0 2118000.0 1149600.0 2131800.0 ;
      RECT  1139400.0 2145600.0 1149600.0 2131800.0 ;
      RECT  1149600.0 379200.0 1159800.0 393000.0 ;
      RECT  1149600.0 406800.0 1159800.0 393000.0 ;
      RECT  1149600.0 406800.0 1159800.0 420600.0 ;
      RECT  1149600.0 434400.0 1159800.0 420600.0 ;
      RECT  1149600.0 434400.0 1159800.0 448200.0 ;
      RECT  1149600.0 462000.0 1159800.0 448200.0 ;
      RECT  1149600.0 462000.0 1159800.0 475800.0 ;
      RECT  1149600.0 489600.0 1159800.0 475800.0 ;
      RECT  1149600.0 489600.0 1159800.0 503400.0 ;
      RECT  1149600.0 517200.0 1159800.0 503400.0 ;
      RECT  1149600.0 517200.0 1159800.0 531000.0 ;
      RECT  1149600.0 544800.0 1159800.0 531000.0 ;
      RECT  1149600.0 544800.0 1159800.0 558600.0 ;
      RECT  1149600.0 572400.0 1159800.0 558600.0 ;
      RECT  1149600.0 572400.0 1159800.0 586200.0 ;
      RECT  1149600.0 600000.0 1159800.0 586200.0 ;
      RECT  1149600.0 600000.0 1159800.0 613800.0 ;
      RECT  1149600.0 627600.0 1159800.0 613800.0 ;
      RECT  1149600.0 627600.0 1159800.0 641400.0 ;
      RECT  1149600.0 655200.0 1159800.0 641400.0 ;
      RECT  1149600.0 655200.0 1159800.0 669000.0 ;
      RECT  1149600.0 682800.0 1159800.0 669000.0 ;
      RECT  1149600.0 682800.0 1159800.0 696600.0 ;
      RECT  1149600.0 710400.0 1159800.0 696600.0 ;
      RECT  1149600.0 710400.0 1159800.0 724200.0 ;
      RECT  1149600.0 738000.0 1159800.0 724200.0 ;
      RECT  1149600.0 738000.0 1159800.0 751800.0 ;
      RECT  1149600.0 765600.0 1159800.0 751800.0 ;
      RECT  1149600.0 765600.0 1159800.0 779400.0 ;
      RECT  1149600.0 793200.0 1159800.0 779400.0 ;
      RECT  1149600.0 793200.0 1159800.0 807000.0 ;
      RECT  1149600.0 820800.0 1159800.0 807000.0 ;
      RECT  1149600.0 820800.0 1159800.0 834600.0 ;
      RECT  1149600.0 848400.0 1159800.0 834600.0 ;
      RECT  1149600.0 848400.0 1159800.0 862200.0 ;
      RECT  1149600.0 876000.0 1159800.0 862200.0 ;
      RECT  1149600.0 876000.0 1159800.0 889800.0 ;
      RECT  1149600.0 903600.0 1159800.0 889800.0 ;
      RECT  1149600.0 903600.0 1159800.0 917400.0 ;
      RECT  1149600.0 931200.0 1159800.0 917400.0 ;
      RECT  1149600.0 931200.0 1159800.0 945000.0 ;
      RECT  1149600.0 958800.0 1159800.0 945000.0 ;
      RECT  1149600.0 958800.0 1159800.0 972600.0 ;
      RECT  1149600.0 986400.0 1159800.0 972600.0 ;
      RECT  1149600.0 986400.0 1159800.0 1000200.0 ;
      RECT  1149600.0 1014000.0 1159800.0 1000200.0 ;
      RECT  1149600.0 1014000.0 1159800.0 1027800.0 ;
      RECT  1149600.0 1041600.0 1159800.0 1027800.0 ;
      RECT  1149600.0 1041600.0 1159800.0 1055400.0 ;
      RECT  1149600.0 1069200.0 1159800.0 1055400.0 ;
      RECT  1149600.0 1069200.0 1159800.0 1083000.0 ;
      RECT  1149600.0 1096800.0 1159800.0 1083000.0 ;
      RECT  1149600.0 1096800.0 1159800.0 1110600.0 ;
      RECT  1149600.0 1124400.0 1159800.0 1110600.0 ;
      RECT  1149600.0 1124400.0 1159800.0 1138200.0 ;
      RECT  1149600.0 1152000.0 1159800.0 1138200.0 ;
      RECT  1149600.0 1152000.0 1159800.0 1165800.0 ;
      RECT  1149600.0 1179600.0 1159800.0 1165800.0 ;
      RECT  1149600.0 1179600.0 1159800.0 1193400.0 ;
      RECT  1149600.0 1207200.0 1159800.0 1193400.0 ;
      RECT  1149600.0 1207200.0 1159800.0 1221000.0 ;
      RECT  1149600.0 1234800.0 1159800.0 1221000.0 ;
      RECT  1149600.0 1234800.0 1159800.0 1248600.0 ;
      RECT  1149600.0 1262400.0 1159800.0 1248600.0 ;
      RECT  1149600.0 1262400.0 1159800.0 1276200.0 ;
      RECT  1149600.0 1290000.0 1159800.0 1276200.0 ;
      RECT  1149600.0 1290000.0 1159800.0 1303800.0 ;
      RECT  1149600.0 1317600.0 1159800.0 1303800.0 ;
      RECT  1149600.0 1317600.0 1159800.0 1331400.0 ;
      RECT  1149600.0 1345200.0 1159800.0 1331400.0 ;
      RECT  1149600.0 1345200.0 1159800.0 1359000.0 ;
      RECT  1149600.0 1372800.0 1159800.0 1359000.0 ;
      RECT  1149600.0 1372800.0 1159800.0 1386600.0 ;
      RECT  1149600.0 1400400.0 1159800.0 1386600.0 ;
      RECT  1149600.0 1400400.0 1159800.0 1414200.0 ;
      RECT  1149600.0 1428000.0 1159800.0 1414200.0 ;
      RECT  1149600.0 1428000.0 1159800.0 1441800.0 ;
      RECT  1149600.0 1455600.0 1159800.0 1441800.0 ;
      RECT  1149600.0 1455600.0 1159800.0 1469400.0 ;
      RECT  1149600.0 1483200.0 1159800.0 1469400.0 ;
      RECT  1149600.0 1483200.0 1159800.0 1497000.0 ;
      RECT  1149600.0 1510800.0 1159800.0 1497000.0 ;
      RECT  1149600.0 1510800.0 1159800.0 1524600.0 ;
      RECT  1149600.0 1538400.0 1159800.0 1524600.0 ;
      RECT  1149600.0 1538400.0 1159800.0 1552200.0 ;
      RECT  1149600.0 1566000.0 1159800.0 1552200.0 ;
      RECT  1149600.0 1566000.0 1159800.0 1579800.0 ;
      RECT  1149600.0 1593600.0 1159800.0 1579800.0 ;
      RECT  1149600.0 1593600.0 1159800.0 1607400.0 ;
      RECT  1149600.0 1621200.0 1159800.0 1607400.0 ;
      RECT  1149600.0 1621200.0 1159800.0 1635000.0 ;
      RECT  1149600.0 1648800.0 1159800.0 1635000.0 ;
      RECT  1149600.0 1648800.0 1159800.0 1662600.0 ;
      RECT  1149600.0 1676400.0 1159800.0 1662600.0 ;
      RECT  1149600.0 1676400.0 1159800.0 1690200.0 ;
      RECT  1149600.0 1704000.0 1159800.0 1690200.0 ;
      RECT  1149600.0 1704000.0 1159800.0 1717800.0 ;
      RECT  1149600.0 1731600.0 1159800.0 1717800.0 ;
      RECT  1149600.0 1731600.0 1159800.0 1745400.0 ;
      RECT  1149600.0 1759200.0 1159800.0 1745400.0 ;
      RECT  1149600.0 1759200.0 1159800.0 1773000.0 ;
      RECT  1149600.0 1786800.0 1159800.0 1773000.0 ;
      RECT  1149600.0 1786800.0 1159800.0 1800600.0 ;
      RECT  1149600.0 1814400.0 1159800.0 1800600.0 ;
      RECT  1149600.0 1814400.0 1159800.0 1828200.0 ;
      RECT  1149600.0 1842000.0 1159800.0 1828200.0 ;
      RECT  1149600.0 1842000.0 1159800.0 1855800.0 ;
      RECT  1149600.0 1869600.0 1159800.0 1855800.0 ;
      RECT  1149600.0 1869600.0 1159800.0 1883400.0 ;
      RECT  1149600.0 1897200.0 1159800.0 1883400.0 ;
      RECT  1149600.0 1897200.0 1159800.0 1911000.0 ;
      RECT  1149600.0 1924800.0 1159800.0 1911000.0 ;
      RECT  1149600.0 1924800.0 1159800.0 1938600.0 ;
      RECT  1149600.0 1952400.0 1159800.0 1938600.0 ;
      RECT  1149600.0 1952400.0 1159800.0 1966200.0 ;
      RECT  1149600.0 1980000.0 1159800.0 1966200.0 ;
      RECT  1149600.0 1980000.0 1159800.0 1993800.0 ;
      RECT  1149600.0 2007600.0 1159800.0 1993800.0 ;
      RECT  1149600.0 2007600.0 1159800.0 2021400.0 ;
      RECT  1149600.0 2035200.0 1159800.0 2021400.0 ;
      RECT  1149600.0 2035200.0 1159800.0 2049000.0 ;
      RECT  1149600.0 2062800.0 1159800.0 2049000.0 ;
      RECT  1149600.0 2062800.0 1159800.0 2076600.0 ;
      RECT  1149600.0 2090400.0 1159800.0 2076600.0 ;
      RECT  1149600.0 2090400.0 1159800.0 2104200.0 ;
      RECT  1149600.0 2118000.0 1159800.0 2104200.0 ;
      RECT  1149600.0 2118000.0 1159800.0 2131800.0 ;
      RECT  1149600.0 2145600.0 1159800.0 2131800.0 ;
      RECT  1159800.0 379200.0 1170000.0 393000.0 ;
      RECT  1159800.0 406800.0 1170000.0 393000.0 ;
      RECT  1159800.0 406800.0 1170000.0 420600.0 ;
      RECT  1159800.0 434400.0 1170000.0 420600.0 ;
      RECT  1159800.0 434400.0 1170000.0 448200.0 ;
      RECT  1159800.0 462000.0 1170000.0 448200.0 ;
      RECT  1159800.0 462000.0 1170000.0 475800.0 ;
      RECT  1159800.0 489600.0 1170000.0 475800.0 ;
      RECT  1159800.0 489600.0 1170000.0 503400.0 ;
      RECT  1159800.0 517200.0 1170000.0 503400.0 ;
      RECT  1159800.0 517200.0 1170000.0 531000.0 ;
      RECT  1159800.0 544800.0 1170000.0 531000.0 ;
      RECT  1159800.0 544800.0 1170000.0 558600.0 ;
      RECT  1159800.0 572400.0 1170000.0 558600.0 ;
      RECT  1159800.0 572400.0 1170000.0 586200.0 ;
      RECT  1159800.0 600000.0 1170000.0 586200.0 ;
      RECT  1159800.0 600000.0 1170000.0 613800.0 ;
      RECT  1159800.0 627600.0 1170000.0 613800.0 ;
      RECT  1159800.0 627600.0 1170000.0 641400.0 ;
      RECT  1159800.0 655200.0 1170000.0 641400.0 ;
      RECT  1159800.0 655200.0 1170000.0 669000.0 ;
      RECT  1159800.0 682800.0 1170000.0 669000.0 ;
      RECT  1159800.0 682800.0 1170000.0 696600.0 ;
      RECT  1159800.0 710400.0 1170000.0 696600.0 ;
      RECT  1159800.0 710400.0 1170000.0 724200.0 ;
      RECT  1159800.0 738000.0 1170000.0 724200.0 ;
      RECT  1159800.0 738000.0 1170000.0 751800.0 ;
      RECT  1159800.0 765600.0 1170000.0 751800.0 ;
      RECT  1159800.0 765600.0 1170000.0 779400.0 ;
      RECT  1159800.0 793200.0 1170000.0 779400.0 ;
      RECT  1159800.0 793200.0 1170000.0 807000.0 ;
      RECT  1159800.0 820800.0 1170000.0 807000.0 ;
      RECT  1159800.0 820800.0 1170000.0 834600.0 ;
      RECT  1159800.0 848400.0 1170000.0 834600.0 ;
      RECT  1159800.0 848400.0 1170000.0 862200.0 ;
      RECT  1159800.0 876000.0 1170000.0 862200.0 ;
      RECT  1159800.0 876000.0 1170000.0 889800.0 ;
      RECT  1159800.0 903600.0 1170000.0 889800.0 ;
      RECT  1159800.0 903600.0 1170000.0 917400.0 ;
      RECT  1159800.0 931200.0 1170000.0 917400.0 ;
      RECT  1159800.0 931200.0 1170000.0 945000.0 ;
      RECT  1159800.0 958800.0 1170000.0 945000.0 ;
      RECT  1159800.0 958800.0 1170000.0 972600.0 ;
      RECT  1159800.0 986400.0 1170000.0 972600.0 ;
      RECT  1159800.0 986400.0 1170000.0 1000200.0 ;
      RECT  1159800.0 1014000.0 1170000.0 1000200.0 ;
      RECT  1159800.0 1014000.0 1170000.0 1027800.0 ;
      RECT  1159800.0 1041600.0 1170000.0 1027800.0 ;
      RECT  1159800.0 1041600.0 1170000.0 1055400.0 ;
      RECT  1159800.0 1069200.0 1170000.0 1055400.0 ;
      RECT  1159800.0 1069200.0 1170000.0 1083000.0 ;
      RECT  1159800.0 1096800.0 1170000.0 1083000.0 ;
      RECT  1159800.0 1096800.0 1170000.0 1110600.0 ;
      RECT  1159800.0 1124400.0 1170000.0 1110600.0 ;
      RECT  1159800.0 1124400.0 1170000.0 1138200.0 ;
      RECT  1159800.0 1152000.0 1170000.0 1138200.0 ;
      RECT  1159800.0 1152000.0 1170000.0 1165800.0 ;
      RECT  1159800.0 1179600.0 1170000.0 1165800.0 ;
      RECT  1159800.0 1179600.0 1170000.0 1193400.0 ;
      RECT  1159800.0 1207200.0 1170000.0 1193400.0 ;
      RECT  1159800.0 1207200.0 1170000.0 1221000.0 ;
      RECT  1159800.0 1234800.0 1170000.0 1221000.0 ;
      RECT  1159800.0 1234800.0 1170000.0 1248600.0 ;
      RECT  1159800.0 1262400.0 1170000.0 1248600.0 ;
      RECT  1159800.0 1262400.0 1170000.0 1276200.0 ;
      RECT  1159800.0 1290000.0 1170000.0 1276200.0 ;
      RECT  1159800.0 1290000.0 1170000.0 1303800.0 ;
      RECT  1159800.0 1317600.0 1170000.0 1303800.0 ;
      RECT  1159800.0 1317600.0 1170000.0 1331400.0 ;
      RECT  1159800.0 1345200.0 1170000.0 1331400.0 ;
      RECT  1159800.0 1345200.0 1170000.0 1359000.0 ;
      RECT  1159800.0 1372800.0 1170000.0 1359000.0 ;
      RECT  1159800.0 1372800.0 1170000.0 1386600.0 ;
      RECT  1159800.0 1400400.0 1170000.0 1386600.0 ;
      RECT  1159800.0 1400400.0 1170000.0 1414200.0 ;
      RECT  1159800.0 1428000.0 1170000.0 1414200.0 ;
      RECT  1159800.0 1428000.0 1170000.0 1441800.0 ;
      RECT  1159800.0 1455600.0 1170000.0 1441800.0 ;
      RECT  1159800.0 1455600.0 1170000.0 1469400.0 ;
      RECT  1159800.0 1483200.0 1170000.0 1469400.0 ;
      RECT  1159800.0 1483200.0 1170000.0 1497000.0 ;
      RECT  1159800.0 1510800.0 1170000.0 1497000.0 ;
      RECT  1159800.0 1510800.0 1170000.0 1524600.0 ;
      RECT  1159800.0 1538400.0 1170000.0 1524600.0 ;
      RECT  1159800.0 1538400.0 1170000.0 1552200.0 ;
      RECT  1159800.0 1566000.0 1170000.0 1552200.0 ;
      RECT  1159800.0 1566000.0 1170000.0 1579800.0 ;
      RECT  1159800.0 1593600.0 1170000.0 1579800.0 ;
      RECT  1159800.0 1593600.0 1170000.0 1607400.0 ;
      RECT  1159800.0 1621200.0 1170000.0 1607400.0 ;
      RECT  1159800.0 1621200.0 1170000.0 1635000.0 ;
      RECT  1159800.0 1648800.0 1170000.0 1635000.0 ;
      RECT  1159800.0 1648800.0 1170000.0 1662600.0 ;
      RECT  1159800.0 1676400.0 1170000.0 1662600.0 ;
      RECT  1159800.0 1676400.0 1170000.0 1690200.0 ;
      RECT  1159800.0 1704000.0 1170000.0 1690200.0 ;
      RECT  1159800.0 1704000.0 1170000.0 1717800.0 ;
      RECT  1159800.0 1731600.0 1170000.0 1717800.0 ;
      RECT  1159800.0 1731600.0 1170000.0 1745400.0 ;
      RECT  1159800.0 1759200.0 1170000.0 1745400.0 ;
      RECT  1159800.0 1759200.0 1170000.0 1773000.0 ;
      RECT  1159800.0 1786800.0 1170000.0 1773000.0 ;
      RECT  1159800.0 1786800.0 1170000.0 1800600.0 ;
      RECT  1159800.0 1814400.0 1170000.0 1800600.0 ;
      RECT  1159800.0 1814400.0 1170000.0 1828200.0 ;
      RECT  1159800.0 1842000.0 1170000.0 1828200.0 ;
      RECT  1159800.0 1842000.0 1170000.0 1855800.0 ;
      RECT  1159800.0 1869600.0 1170000.0 1855800.0 ;
      RECT  1159800.0 1869600.0 1170000.0 1883400.0 ;
      RECT  1159800.0 1897200.0 1170000.0 1883400.0 ;
      RECT  1159800.0 1897200.0 1170000.0 1911000.0 ;
      RECT  1159800.0 1924800.0 1170000.0 1911000.0 ;
      RECT  1159800.0 1924800.0 1170000.0 1938600.0 ;
      RECT  1159800.0 1952400.0 1170000.0 1938600.0 ;
      RECT  1159800.0 1952400.0 1170000.0 1966200.0 ;
      RECT  1159800.0 1980000.0 1170000.0 1966200.0 ;
      RECT  1159800.0 1980000.0 1170000.0 1993800.0 ;
      RECT  1159800.0 2007600.0 1170000.0 1993800.0 ;
      RECT  1159800.0 2007600.0 1170000.0 2021400.0 ;
      RECT  1159800.0 2035200.0 1170000.0 2021400.0 ;
      RECT  1159800.0 2035200.0 1170000.0 2049000.0 ;
      RECT  1159800.0 2062800.0 1170000.0 2049000.0 ;
      RECT  1159800.0 2062800.0 1170000.0 2076600.0 ;
      RECT  1159800.0 2090400.0 1170000.0 2076600.0 ;
      RECT  1159800.0 2090400.0 1170000.0 2104200.0 ;
      RECT  1159800.0 2118000.0 1170000.0 2104200.0 ;
      RECT  1159800.0 2118000.0 1170000.0 2131800.0 ;
      RECT  1159800.0 2145600.0 1170000.0 2131800.0 ;
      RECT  1170000.0 379200.0 1180200.0 393000.0 ;
      RECT  1170000.0 406800.0 1180200.0 393000.0 ;
      RECT  1170000.0 406800.0 1180200.0 420600.0 ;
      RECT  1170000.0 434400.0 1180200.0 420600.0 ;
      RECT  1170000.0 434400.0 1180200.0 448200.0 ;
      RECT  1170000.0 462000.0 1180200.0 448200.0 ;
      RECT  1170000.0 462000.0 1180200.0 475800.0 ;
      RECT  1170000.0 489600.0 1180200.0 475800.0 ;
      RECT  1170000.0 489600.0 1180200.0 503400.0 ;
      RECT  1170000.0 517200.0 1180200.0 503400.0 ;
      RECT  1170000.0 517200.0 1180200.0 531000.0 ;
      RECT  1170000.0 544800.0 1180200.0 531000.0 ;
      RECT  1170000.0 544800.0 1180200.0 558600.0 ;
      RECT  1170000.0 572400.0 1180200.0 558600.0 ;
      RECT  1170000.0 572400.0 1180200.0 586200.0 ;
      RECT  1170000.0 600000.0 1180200.0 586200.0 ;
      RECT  1170000.0 600000.0 1180200.0 613800.0 ;
      RECT  1170000.0 627600.0 1180200.0 613800.0 ;
      RECT  1170000.0 627600.0 1180200.0 641400.0 ;
      RECT  1170000.0 655200.0 1180200.0 641400.0 ;
      RECT  1170000.0 655200.0 1180200.0 669000.0 ;
      RECT  1170000.0 682800.0 1180200.0 669000.0 ;
      RECT  1170000.0 682800.0 1180200.0 696600.0 ;
      RECT  1170000.0 710400.0 1180200.0 696600.0 ;
      RECT  1170000.0 710400.0 1180200.0 724200.0 ;
      RECT  1170000.0 738000.0 1180200.0 724200.0 ;
      RECT  1170000.0 738000.0 1180200.0 751800.0 ;
      RECT  1170000.0 765600.0 1180200.0 751800.0 ;
      RECT  1170000.0 765600.0 1180200.0 779400.0 ;
      RECT  1170000.0 793200.0 1180200.0 779400.0 ;
      RECT  1170000.0 793200.0 1180200.0 807000.0 ;
      RECT  1170000.0 820800.0 1180200.0 807000.0 ;
      RECT  1170000.0 820800.0 1180200.0 834600.0 ;
      RECT  1170000.0 848400.0 1180200.0 834600.0 ;
      RECT  1170000.0 848400.0 1180200.0 862200.0 ;
      RECT  1170000.0 876000.0 1180200.0 862200.0 ;
      RECT  1170000.0 876000.0 1180200.0 889800.0 ;
      RECT  1170000.0 903600.0 1180200.0 889800.0 ;
      RECT  1170000.0 903600.0 1180200.0 917400.0 ;
      RECT  1170000.0 931200.0 1180200.0 917400.0 ;
      RECT  1170000.0 931200.0 1180200.0 945000.0 ;
      RECT  1170000.0 958800.0 1180200.0 945000.0 ;
      RECT  1170000.0 958800.0 1180200.0 972600.0 ;
      RECT  1170000.0 986400.0 1180200.0 972600.0 ;
      RECT  1170000.0 986400.0 1180200.0 1000200.0 ;
      RECT  1170000.0 1014000.0 1180200.0 1000200.0 ;
      RECT  1170000.0 1014000.0 1180200.0 1027800.0 ;
      RECT  1170000.0 1041600.0 1180200.0 1027800.0 ;
      RECT  1170000.0 1041600.0 1180200.0 1055400.0 ;
      RECT  1170000.0 1069200.0 1180200.0 1055400.0 ;
      RECT  1170000.0 1069200.0 1180200.0 1083000.0 ;
      RECT  1170000.0 1096800.0 1180200.0 1083000.0 ;
      RECT  1170000.0 1096800.0 1180200.0 1110600.0 ;
      RECT  1170000.0 1124400.0 1180200.0 1110600.0 ;
      RECT  1170000.0 1124400.0 1180200.0 1138200.0 ;
      RECT  1170000.0 1152000.0 1180200.0 1138200.0 ;
      RECT  1170000.0 1152000.0 1180200.0 1165800.0 ;
      RECT  1170000.0 1179600.0 1180200.0 1165800.0 ;
      RECT  1170000.0 1179600.0 1180200.0 1193400.0 ;
      RECT  1170000.0 1207200.0 1180200.0 1193400.0 ;
      RECT  1170000.0 1207200.0 1180200.0 1221000.0 ;
      RECT  1170000.0 1234800.0 1180200.0 1221000.0 ;
      RECT  1170000.0 1234800.0 1180200.0 1248600.0 ;
      RECT  1170000.0 1262400.0 1180200.0 1248600.0 ;
      RECT  1170000.0 1262400.0 1180200.0 1276200.0 ;
      RECT  1170000.0 1290000.0 1180200.0 1276200.0 ;
      RECT  1170000.0 1290000.0 1180200.0 1303800.0 ;
      RECT  1170000.0 1317600.0 1180200.0 1303800.0 ;
      RECT  1170000.0 1317600.0 1180200.0 1331400.0 ;
      RECT  1170000.0 1345200.0 1180200.0 1331400.0 ;
      RECT  1170000.0 1345200.0 1180200.0 1359000.0 ;
      RECT  1170000.0 1372800.0 1180200.0 1359000.0 ;
      RECT  1170000.0 1372800.0 1180200.0 1386600.0 ;
      RECT  1170000.0 1400400.0 1180200.0 1386600.0 ;
      RECT  1170000.0 1400400.0 1180200.0 1414200.0 ;
      RECT  1170000.0 1428000.0 1180200.0 1414200.0 ;
      RECT  1170000.0 1428000.0 1180200.0 1441800.0 ;
      RECT  1170000.0 1455600.0 1180200.0 1441800.0 ;
      RECT  1170000.0 1455600.0 1180200.0 1469400.0 ;
      RECT  1170000.0 1483200.0 1180200.0 1469400.0 ;
      RECT  1170000.0 1483200.0 1180200.0 1497000.0 ;
      RECT  1170000.0 1510800.0 1180200.0 1497000.0 ;
      RECT  1170000.0 1510800.0 1180200.0 1524600.0 ;
      RECT  1170000.0 1538400.0 1180200.0 1524600.0 ;
      RECT  1170000.0 1538400.0 1180200.0 1552200.0 ;
      RECT  1170000.0 1566000.0 1180200.0 1552200.0 ;
      RECT  1170000.0 1566000.0 1180200.0 1579800.0 ;
      RECT  1170000.0 1593600.0 1180200.0 1579800.0 ;
      RECT  1170000.0 1593600.0 1180200.0 1607400.0 ;
      RECT  1170000.0 1621200.0 1180200.0 1607400.0 ;
      RECT  1170000.0 1621200.0 1180200.0 1635000.0 ;
      RECT  1170000.0 1648800.0 1180200.0 1635000.0 ;
      RECT  1170000.0 1648800.0 1180200.0 1662600.0 ;
      RECT  1170000.0 1676400.0 1180200.0 1662600.0 ;
      RECT  1170000.0 1676400.0 1180200.0 1690200.0 ;
      RECT  1170000.0 1704000.0 1180200.0 1690200.0 ;
      RECT  1170000.0 1704000.0 1180200.0 1717800.0 ;
      RECT  1170000.0 1731600.0 1180200.0 1717800.0 ;
      RECT  1170000.0 1731600.0 1180200.0 1745400.0 ;
      RECT  1170000.0 1759200.0 1180200.0 1745400.0 ;
      RECT  1170000.0 1759200.0 1180200.0 1773000.0 ;
      RECT  1170000.0 1786800.0 1180200.0 1773000.0 ;
      RECT  1170000.0 1786800.0 1180200.0 1800600.0 ;
      RECT  1170000.0 1814400.0 1180200.0 1800600.0 ;
      RECT  1170000.0 1814400.0 1180200.0 1828200.0 ;
      RECT  1170000.0 1842000.0 1180200.0 1828200.0 ;
      RECT  1170000.0 1842000.0 1180200.0 1855800.0 ;
      RECT  1170000.0 1869600.0 1180200.0 1855800.0 ;
      RECT  1170000.0 1869600.0 1180200.0 1883400.0 ;
      RECT  1170000.0 1897200.0 1180200.0 1883400.0 ;
      RECT  1170000.0 1897200.0 1180200.0 1911000.0 ;
      RECT  1170000.0 1924800.0 1180200.0 1911000.0 ;
      RECT  1170000.0 1924800.0 1180200.0 1938600.0 ;
      RECT  1170000.0 1952400.0 1180200.0 1938600.0 ;
      RECT  1170000.0 1952400.0 1180200.0 1966200.0 ;
      RECT  1170000.0 1980000.0 1180200.0 1966200.0 ;
      RECT  1170000.0 1980000.0 1180200.0 1993800.0 ;
      RECT  1170000.0 2007600.0 1180200.0 1993800.0 ;
      RECT  1170000.0 2007600.0 1180200.0 2021400.0 ;
      RECT  1170000.0 2035200.0 1180200.0 2021400.0 ;
      RECT  1170000.0 2035200.0 1180200.0 2049000.0 ;
      RECT  1170000.0 2062800.0 1180200.0 2049000.0 ;
      RECT  1170000.0 2062800.0 1180200.0 2076600.0 ;
      RECT  1170000.0 2090400.0 1180200.0 2076600.0 ;
      RECT  1170000.0 2090400.0 1180200.0 2104200.0 ;
      RECT  1170000.0 2118000.0 1180200.0 2104200.0 ;
      RECT  1170000.0 2118000.0 1180200.0 2131800.0 ;
      RECT  1170000.0 2145600.0 1180200.0 2131800.0 ;
      RECT  1180200.0 379200.0 1190400.0 393000.0 ;
      RECT  1180200.0 406800.0 1190400.0 393000.0 ;
      RECT  1180200.0 406800.0 1190400.0 420600.0 ;
      RECT  1180200.0 434400.0 1190400.0 420600.0 ;
      RECT  1180200.0 434400.0 1190400.0 448200.0 ;
      RECT  1180200.0 462000.0 1190400.0 448200.0 ;
      RECT  1180200.0 462000.0 1190400.0 475800.0 ;
      RECT  1180200.0 489600.0 1190400.0 475800.0 ;
      RECT  1180200.0 489600.0 1190400.0 503400.0 ;
      RECT  1180200.0 517200.0 1190400.0 503400.0 ;
      RECT  1180200.0 517200.0 1190400.0 531000.0 ;
      RECT  1180200.0 544800.0 1190400.0 531000.0 ;
      RECT  1180200.0 544800.0 1190400.0 558600.0 ;
      RECT  1180200.0 572400.0 1190400.0 558600.0 ;
      RECT  1180200.0 572400.0 1190400.0 586200.0 ;
      RECT  1180200.0 600000.0 1190400.0 586200.0 ;
      RECT  1180200.0 600000.0 1190400.0 613800.0 ;
      RECT  1180200.0 627600.0 1190400.0 613800.0 ;
      RECT  1180200.0 627600.0 1190400.0 641400.0 ;
      RECT  1180200.0 655200.0 1190400.0 641400.0 ;
      RECT  1180200.0 655200.0 1190400.0 669000.0 ;
      RECT  1180200.0 682800.0 1190400.0 669000.0 ;
      RECT  1180200.0 682800.0 1190400.0 696600.0 ;
      RECT  1180200.0 710400.0 1190400.0 696600.0 ;
      RECT  1180200.0 710400.0 1190400.0 724200.0 ;
      RECT  1180200.0 738000.0 1190400.0 724200.0 ;
      RECT  1180200.0 738000.0 1190400.0 751800.0 ;
      RECT  1180200.0 765600.0 1190400.0 751800.0 ;
      RECT  1180200.0 765600.0 1190400.0 779400.0 ;
      RECT  1180200.0 793200.0 1190400.0 779400.0 ;
      RECT  1180200.0 793200.0 1190400.0 807000.0 ;
      RECT  1180200.0 820800.0 1190400.0 807000.0 ;
      RECT  1180200.0 820800.0 1190400.0 834600.0 ;
      RECT  1180200.0 848400.0 1190400.0 834600.0 ;
      RECT  1180200.0 848400.0 1190400.0 862200.0 ;
      RECT  1180200.0 876000.0 1190400.0 862200.0 ;
      RECT  1180200.0 876000.0 1190400.0 889800.0 ;
      RECT  1180200.0 903600.0 1190400.0 889800.0 ;
      RECT  1180200.0 903600.0 1190400.0 917400.0 ;
      RECT  1180200.0 931200.0 1190400.0 917400.0 ;
      RECT  1180200.0 931200.0 1190400.0 945000.0 ;
      RECT  1180200.0 958800.0 1190400.0 945000.0 ;
      RECT  1180200.0 958800.0 1190400.0 972600.0 ;
      RECT  1180200.0 986400.0 1190400.0 972600.0 ;
      RECT  1180200.0 986400.0 1190400.0 1000200.0 ;
      RECT  1180200.0 1014000.0 1190400.0 1000200.0 ;
      RECT  1180200.0 1014000.0 1190400.0 1027800.0 ;
      RECT  1180200.0 1041600.0 1190400.0 1027800.0 ;
      RECT  1180200.0 1041600.0 1190400.0 1055400.0 ;
      RECT  1180200.0 1069200.0 1190400.0 1055400.0 ;
      RECT  1180200.0 1069200.0 1190400.0 1083000.0 ;
      RECT  1180200.0 1096800.0 1190400.0 1083000.0 ;
      RECT  1180200.0 1096800.0 1190400.0 1110600.0 ;
      RECT  1180200.0 1124400.0 1190400.0 1110600.0 ;
      RECT  1180200.0 1124400.0 1190400.0 1138200.0 ;
      RECT  1180200.0 1152000.0 1190400.0 1138200.0 ;
      RECT  1180200.0 1152000.0 1190400.0 1165800.0 ;
      RECT  1180200.0 1179600.0 1190400.0 1165800.0 ;
      RECT  1180200.0 1179600.0 1190400.0 1193400.0 ;
      RECT  1180200.0 1207200.0 1190400.0 1193400.0 ;
      RECT  1180200.0 1207200.0 1190400.0 1221000.0 ;
      RECT  1180200.0 1234800.0 1190400.0 1221000.0 ;
      RECT  1180200.0 1234800.0 1190400.0 1248600.0 ;
      RECT  1180200.0 1262400.0 1190400.0 1248600.0 ;
      RECT  1180200.0 1262400.0 1190400.0 1276200.0 ;
      RECT  1180200.0 1290000.0 1190400.0 1276200.0 ;
      RECT  1180200.0 1290000.0 1190400.0 1303800.0 ;
      RECT  1180200.0 1317600.0 1190400.0 1303800.0 ;
      RECT  1180200.0 1317600.0 1190400.0 1331400.0 ;
      RECT  1180200.0 1345200.0 1190400.0 1331400.0 ;
      RECT  1180200.0 1345200.0 1190400.0 1359000.0 ;
      RECT  1180200.0 1372800.0 1190400.0 1359000.0 ;
      RECT  1180200.0 1372800.0 1190400.0 1386600.0 ;
      RECT  1180200.0 1400400.0 1190400.0 1386600.0 ;
      RECT  1180200.0 1400400.0 1190400.0 1414200.0 ;
      RECT  1180200.0 1428000.0 1190400.0 1414200.0 ;
      RECT  1180200.0 1428000.0 1190400.0 1441800.0 ;
      RECT  1180200.0 1455600.0 1190400.0 1441800.0 ;
      RECT  1180200.0 1455600.0 1190400.0 1469400.0 ;
      RECT  1180200.0 1483200.0 1190400.0 1469400.0 ;
      RECT  1180200.0 1483200.0 1190400.0 1497000.0 ;
      RECT  1180200.0 1510800.0 1190400.0 1497000.0 ;
      RECT  1180200.0 1510800.0 1190400.0 1524600.0 ;
      RECT  1180200.0 1538400.0 1190400.0 1524600.0 ;
      RECT  1180200.0 1538400.0 1190400.0 1552200.0 ;
      RECT  1180200.0 1566000.0 1190400.0 1552200.0 ;
      RECT  1180200.0 1566000.0 1190400.0 1579800.0 ;
      RECT  1180200.0 1593600.0 1190400.0 1579800.0 ;
      RECT  1180200.0 1593600.0 1190400.0 1607400.0 ;
      RECT  1180200.0 1621200.0 1190400.0 1607400.0 ;
      RECT  1180200.0 1621200.0 1190400.0 1635000.0 ;
      RECT  1180200.0 1648800.0 1190400.0 1635000.0 ;
      RECT  1180200.0 1648800.0 1190400.0 1662600.0 ;
      RECT  1180200.0 1676400.0 1190400.0 1662600.0 ;
      RECT  1180200.0 1676400.0 1190400.0 1690200.0 ;
      RECT  1180200.0 1704000.0 1190400.0 1690200.0 ;
      RECT  1180200.0 1704000.0 1190400.0 1717800.0 ;
      RECT  1180200.0 1731600.0 1190400.0 1717800.0 ;
      RECT  1180200.0 1731600.0 1190400.0 1745400.0 ;
      RECT  1180200.0 1759200.0 1190400.0 1745400.0 ;
      RECT  1180200.0 1759200.0 1190400.0 1773000.0 ;
      RECT  1180200.0 1786800.0 1190400.0 1773000.0 ;
      RECT  1180200.0 1786800.0 1190400.0 1800600.0 ;
      RECT  1180200.0 1814400.0 1190400.0 1800600.0 ;
      RECT  1180200.0 1814400.0 1190400.0 1828200.0 ;
      RECT  1180200.0 1842000.0 1190400.0 1828200.0 ;
      RECT  1180200.0 1842000.0 1190400.0 1855800.0 ;
      RECT  1180200.0 1869600.0 1190400.0 1855800.0 ;
      RECT  1180200.0 1869600.0 1190400.0 1883400.0 ;
      RECT  1180200.0 1897200.0 1190400.0 1883400.0 ;
      RECT  1180200.0 1897200.0 1190400.0 1911000.0 ;
      RECT  1180200.0 1924800.0 1190400.0 1911000.0 ;
      RECT  1180200.0 1924800.0 1190400.0 1938600.0 ;
      RECT  1180200.0 1952400.0 1190400.0 1938600.0 ;
      RECT  1180200.0 1952400.0 1190400.0 1966200.0 ;
      RECT  1180200.0 1980000.0 1190400.0 1966200.0 ;
      RECT  1180200.0 1980000.0 1190400.0 1993800.0 ;
      RECT  1180200.0 2007600.0 1190400.0 1993800.0 ;
      RECT  1180200.0 2007600.0 1190400.0 2021400.0 ;
      RECT  1180200.0 2035200.0 1190400.0 2021400.0 ;
      RECT  1180200.0 2035200.0 1190400.0 2049000.0 ;
      RECT  1180200.0 2062800.0 1190400.0 2049000.0 ;
      RECT  1180200.0 2062800.0 1190400.0 2076600.0 ;
      RECT  1180200.0 2090400.0 1190400.0 2076600.0 ;
      RECT  1180200.0 2090400.0 1190400.0 2104200.0 ;
      RECT  1180200.0 2118000.0 1190400.0 2104200.0 ;
      RECT  1180200.0 2118000.0 1190400.0 2131800.0 ;
      RECT  1180200.0 2145600.0 1190400.0 2131800.0 ;
      RECT  1190400.0 379200.0 1200600.0 393000.0 ;
      RECT  1190400.0 406800.0 1200600.0 393000.0 ;
      RECT  1190400.0 406800.0 1200600.0 420600.0 ;
      RECT  1190400.0 434400.0 1200600.0 420600.0 ;
      RECT  1190400.0 434400.0 1200600.0 448200.0 ;
      RECT  1190400.0 462000.0 1200600.0 448200.0 ;
      RECT  1190400.0 462000.0 1200600.0 475800.0 ;
      RECT  1190400.0 489600.0 1200600.0 475800.0 ;
      RECT  1190400.0 489600.0 1200600.0 503400.0 ;
      RECT  1190400.0 517200.0 1200600.0 503400.0 ;
      RECT  1190400.0 517200.0 1200600.0 531000.0 ;
      RECT  1190400.0 544800.0 1200600.0 531000.0 ;
      RECT  1190400.0 544800.0 1200600.0 558600.0 ;
      RECT  1190400.0 572400.0 1200600.0 558600.0 ;
      RECT  1190400.0 572400.0 1200600.0 586200.0 ;
      RECT  1190400.0 600000.0 1200600.0 586200.0 ;
      RECT  1190400.0 600000.0 1200600.0 613800.0 ;
      RECT  1190400.0 627600.0 1200600.0 613800.0 ;
      RECT  1190400.0 627600.0 1200600.0 641400.0 ;
      RECT  1190400.0 655200.0 1200600.0 641400.0 ;
      RECT  1190400.0 655200.0 1200600.0 669000.0 ;
      RECT  1190400.0 682800.0 1200600.0 669000.0 ;
      RECT  1190400.0 682800.0 1200600.0 696600.0 ;
      RECT  1190400.0 710400.0 1200600.0 696600.0 ;
      RECT  1190400.0 710400.0 1200600.0 724200.0 ;
      RECT  1190400.0 738000.0 1200600.0 724200.0 ;
      RECT  1190400.0 738000.0 1200600.0 751800.0 ;
      RECT  1190400.0 765600.0 1200600.0 751800.0 ;
      RECT  1190400.0 765600.0 1200600.0 779400.0 ;
      RECT  1190400.0 793200.0 1200600.0 779400.0 ;
      RECT  1190400.0 793200.0 1200600.0 807000.0 ;
      RECT  1190400.0 820800.0 1200600.0 807000.0 ;
      RECT  1190400.0 820800.0 1200600.0 834600.0 ;
      RECT  1190400.0 848400.0 1200600.0 834600.0 ;
      RECT  1190400.0 848400.0 1200600.0 862200.0 ;
      RECT  1190400.0 876000.0 1200600.0 862200.0 ;
      RECT  1190400.0 876000.0 1200600.0 889800.0 ;
      RECT  1190400.0 903600.0 1200600.0 889800.0 ;
      RECT  1190400.0 903600.0 1200600.0 917400.0 ;
      RECT  1190400.0 931200.0 1200600.0 917400.0 ;
      RECT  1190400.0 931200.0 1200600.0 945000.0 ;
      RECT  1190400.0 958800.0 1200600.0 945000.0 ;
      RECT  1190400.0 958800.0 1200600.0 972600.0 ;
      RECT  1190400.0 986400.0 1200600.0 972600.0 ;
      RECT  1190400.0 986400.0 1200600.0 1000200.0 ;
      RECT  1190400.0 1014000.0 1200600.0 1000200.0 ;
      RECT  1190400.0 1014000.0 1200600.0 1027800.0 ;
      RECT  1190400.0 1041600.0 1200600.0 1027800.0 ;
      RECT  1190400.0 1041600.0 1200600.0 1055400.0 ;
      RECT  1190400.0 1069200.0 1200600.0 1055400.0 ;
      RECT  1190400.0 1069200.0 1200600.0 1083000.0 ;
      RECT  1190400.0 1096800.0 1200600.0 1083000.0 ;
      RECT  1190400.0 1096800.0 1200600.0 1110600.0 ;
      RECT  1190400.0 1124400.0 1200600.0 1110600.0 ;
      RECT  1190400.0 1124400.0 1200600.0 1138200.0 ;
      RECT  1190400.0 1152000.0 1200600.0 1138200.0 ;
      RECT  1190400.0 1152000.0 1200600.0 1165800.0 ;
      RECT  1190400.0 1179600.0 1200600.0 1165800.0 ;
      RECT  1190400.0 1179600.0 1200600.0 1193400.0 ;
      RECT  1190400.0 1207200.0 1200600.0 1193400.0 ;
      RECT  1190400.0 1207200.0 1200600.0 1221000.0 ;
      RECT  1190400.0 1234800.0 1200600.0 1221000.0 ;
      RECT  1190400.0 1234800.0 1200600.0 1248600.0 ;
      RECT  1190400.0 1262400.0 1200600.0 1248600.0 ;
      RECT  1190400.0 1262400.0 1200600.0 1276200.0 ;
      RECT  1190400.0 1290000.0 1200600.0 1276200.0 ;
      RECT  1190400.0 1290000.0 1200600.0 1303800.0 ;
      RECT  1190400.0 1317600.0 1200600.0 1303800.0 ;
      RECT  1190400.0 1317600.0 1200600.0 1331400.0 ;
      RECT  1190400.0 1345200.0 1200600.0 1331400.0 ;
      RECT  1190400.0 1345200.0 1200600.0 1359000.0 ;
      RECT  1190400.0 1372800.0 1200600.0 1359000.0 ;
      RECT  1190400.0 1372800.0 1200600.0 1386600.0 ;
      RECT  1190400.0 1400400.0 1200600.0 1386600.0 ;
      RECT  1190400.0 1400400.0 1200600.0 1414200.0 ;
      RECT  1190400.0 1428000.0 1200600.0 1414200.0 ;
      RECT  1190400.0 1428000.0 1200600.0 1441800.0 ;
      RECT  1190400.0 1455600.0 1200600.0 1441800.0 ;
      RECT  1190400.0 1455600.0 1200600.0 1469400.0 ;
      RECT  1190400.0 1483200.0 1200600.0 1469400.0 ;
      RECT  1190400.0 1483200.0 1200600.0 1497000.0 ;
      RECT  1190400.0 1510800.0 1200600.0 1497000.0 ;
      RECT  1190400.0 1510800.0 1200600.0 1524600.0 ;
      RECT  1190400.0 1538400.0 1200600.0 1524600.0 ;
      RECT  1190400.0 1538400.0 1200600.0 1552200.0 ;
      RECT  1190400.0 1566000.0 1200600.0 1552200.0 ;
      RECT  1190400.0 1566000.0 1200600.0 1579800.0 ;
      RECT  1190400.0 1593600.0 1200600.0 1579800.0 ;
      RECT  1190400.0 1593600.0 1200600.0 1607400.0 ;
      RECT  1190400.0 1621200.0 1200600.0 1607400.0 ;
      RECT  1190400.0 1621200.0 1200600.0 1635000.0 ;
      RECT  1190400.0 1648800.0 1200600.0 1635000.0 ;
      RECT  1190400.0 1648800.0 1200600.0 1662600.0 ;
      RECT  1190400.0 1676400.0 1200600.0 1662600.0 ;
      RECT  1190400.0 1676400.0 1200600.0 1690200.0 ;
      RECT  1190400.0 1704000.0 1200600.0 1690200.0 ;
      RECT  1190400.0 1704000.0 1200600.0 1717800.0 ;
      RECT  1190400.0 1731600.0 1200600.0 1717800.0 ;
      RECT  1190400.0 1731600.0 1200600.0 1745400.0 ;
      RECT  1190400.0 1759200.0 1200600.0 1745400.0 ;
      RECT  1190400.0 1759200.0 1200600.0 1773000.0 ;
      RECT  1190400.0 1786800.0 1200600.0 1773000.0 ;
      RECT  1190400.0 1786800.0 1200600.0 1800600.0 ;
      RECT  1190400.0 1814400.0 1200600.0 1800600.0 ;
      RECT  1190400.0 1814400.0 1200600.0 1828200.0 ;
      RECT  1190400.0 1842000.0 1200600.0 1828200.0 ;
      RECT  1190400.0 1842000.0 1200600.0 1855800.0 ;
      RECT  1190400.0 1869600.0 1200600.0 1855800.0 ;
      RECT  1190400.0 1869600.0 1200600.0 1883400.0 ;
      RECT  1190400.0 1897200.0 1200600.0 1883400.0 ;
      RECT  1190400.0 1897200.0 1200600.0 1911000.0 ;
      RECT  1190400.0 1924800.0 1200600.0 1911000.0 ;
      RECT  1190400.0 1924800.0 1200600.0 1938600.0 ;
      RECT  1190400.0 1952400.0 1200600.0 1938600.0 ;
      RECT  1190400.0 1952400.0 1200600.0 1966200.0 ;
      RECT  1190400.0 1980000.0 1200600.0 1966200.0 ;
      RECT  1190400.0 1980000.0 1200600.0 1993800.0 ;
      RECT  1190400.0 2007600.0 1200600.0 1993800.0 ;
      RECT  1190400.0 2007600.0 1200600.0 2021400.0 ;
      RECT  1190400.0 2035200.0 1200600.0 2021400.0 ;
      RECT  1190400.0 2035200.0 1200600.0 2049000.0 ;
      RECT  1190400.0 2062800.0 1200600.0 2049000.0 ;
      RECT  1190400.0 2062800.0 1200600.0 2076600.0 ;
      RECT  1190400.0 2090400.0 1200600.0 2076600.0 ;
      RECT  1190400.0 2090400.0 1200600.0 2104200.0 ;
      RECT  1190400.0 2118000.0 1200600.0 2104200.0 ;
      RECT  1190400.0 2118000.0 1200600.0 2131800.0 ;
      RECT  1190400.0 2145600.0 1200600.0 2131800.0 ;
      RECT  1200600.0 379200.0 1210800.0 393000.0 ;
      RECT  1200600.0 406800.0 1210800.0 393000.0 ;
      RECT  1200600.0 406800.0 1210800.0 420600.0 ;
      RECT  1200600.0 434400.0 1210800.0 420600.0 ;
      RECT  1200600.0 434400.0 1210800.0 448200.0 ;
      RECT  1200600.0 462000.0 1210800.0 448200.0 ;
      RECT  1200600.0 462000.0 1210800.0 475800.0 ;
      RECT  1200600.0 489600.0 1210800.0 475800.0 ;
      RECT  1200600.0 489600.0 1210800.0 503400.0 ;
      RECT  1200600.0 517200.0 1210800.0 503400.0 ;
      RECT  1200600.0 517200.0 1210800.0 531000.0 ;
      RECT  1200600.0 544800.0 1210800.0 531000.0 ;
      RECT  1200600.0 544800.0 1210800.0 558600.0 ;
      RECT  1200600.0 572400.0 1210800.0 558600.0 ;
      RECT  1200600.0 572400.0 1210800.0 586200.0 ;
      RECT  1200600.0 600000.0 1210800.0 586200.0 ;
      RECT  1200600.0 600000.0 1210800.0 613800.0 ;
      RECT  1200600.0 627600.0 1210800.0 613800.0 ;
      RECT  1200600.0 627600.0 1210800.0 641400.0 ;
      RECT  1200600.0 655200.0 1210800.0 641400.0 ;
      RECT  1200600.0 655200.0 1210800.0 669000.0 ;
      RECT  1200600.0 682800.0 1210800.0 669000.0 ;
      RECT  1200600.0 682800.0 1210800.0 696600.0 ;
      RECT  1200600.0 710400.0 1210800.0 696600.0 ;
      RECT  1200600.0 710400.0 1210800.0 724200.0 ;
      RECT  1200600.0 738000.0 1210800.0 724200.0 ;
      RECT  1200600.0 738000.0 1210800.0 751800.0 ;
      RECT  1200600.0 765600.0 1210800.0 751800.0 ;
      RECT  1200600.0 765600.0 1210800.0 779400.0 ;
      RECT  1200600.0 793200.0 1210800.0 779400.0 ;
      RECT  1200600.0 793200.0 1210800.0 807000.0 ;
      RECT  1200600.0 820800.0 1210800.0 807000.0 ;
      RECT  1200600.0 820800.0 1210800.0 834600.0 ;
      RECT  1200600.0 848400.0 1210800.0 834600.0 ;
      RECT  1200600.0 848400.0 1210800.0 862200.0 ;
      RECT  1200600.0 876000.0 1210800.0 862200.0 ;
      RECT  1200600.0 876000.0 1210800.0 889800.0 ;
      RECT  1200600.0 903600.0 1210800.0 889800.0 ;
      RECT  1200600.0 903600.0 1210800.0 917400.0 ;
      RECT  1200600.0 931200.0 1210800.0 917400.0 ;
      RECT  1200600.0 931200.0 1210800.0 945000.0 ;
      RECT  1200600.0 958800.0 1210800.0 945000.0 ;
      RECT  1200600.0 958800.0 1210800.0 972600.0 ;
      RECT  1200600.0 986400.0 1210800.0 972600.0 ;
      RECT  1200600.0 986400.0 1210800.0 1000200.0 ;
      RECT  1200600.0 1014000.0 1210800.0 1000200.0 ;
      RECT  1200600.0 1014000.0 1210800.0 1027800.0 ;
      RECT  1200600.0 1041600.0 1210800.0 1027800.0 ;
      RECT  1200600.0 1041600.0 1210800.0 1055400.0 ;
      RECT  1200600.0 1069200.0 1210800.0 1055400.0 ;
      RECT  1200600.0 1069200.0 1210800.0 1083000.0 ;
      RECT  1200600.0 1096800.0 1210800.0 1083000.0 ;
      RECT  1200600.0 1096800.0 1210800.0 1110600.0 ;
      RECT  1200600.0 1124400.0 1210800.0 1110600.0 ;
      RECT  1200600.0 1124400.0 1210800.0 1138200.0 ;
      RECT  1200600.0 1152000.0 1210800.0 1138200.0 ;
      RECT  1200600.0 1152000.0 1210800.0 1165800.0 ;
      RECT  1200600.0 1179600.0 1210800.0 1165800.0 ;
      RECT  1200600.0 1179600.0 1210800.0 1193400.0 ;
      RECT  1200600.0 1207200.0 1210800.0 1193400.0 ;
      RECT  1200600.0 1207200.0 1210800.0 1221000.0 ;
      RECT  1200600.0 1234800.0 1210800.0 1221000.0 ;
      RECT  1200600.0 1234800.0 1210800.0 1248600.0 ;
      RECT  1200600.0 1262400.0 1210800.0 1248600.0 ;
      RECT  1200600.0 1262400.0 1210800.0 1276200.0 ;
      RECT  1200600.0 1290000.0 1210800.0 1276200.0 ;
      RECT  1200600.0 1290000.0 1210800.0 1303800.0 ;
      RECT  1200600.0 1317600.0 1210800.0 1303800.0 ;
      RECT  1200600.0 1317600.0 1210800.0 1331400.0 ;
      RECT  1200600.0 1345200.0 1210800.0 1331400.0 ;
      RECT  1200600.0 1345200.0 1210800.0 1359000.0 ;
      RECT  1200600.0 1372800.0 1210800.0 1359000.0 ;
      RECT  1200600.0 1372800.0 1210800.0 1386600.0 ;
      RECT  1200600.0 1400400.0 1210800.0 1386600.0 ;
      RECT  1200600.0 1400400.0 1210800.0 1414200.0 ;
      RECT  1200600.0 1428000.0 1210800.0 1414200.0 ;
      RECT  1200600.0 1428000.0 1210800.0 1441800.0 ;
      RECT  1200600.0 1455600.0 1210800.0 1441800.0 ;
      RECT  1200600.0 1455600.0 1210800.0 1469400.0 ;
      RECT  1200600.0 1483200.0 1210800.0 1469400.0 ;
      RECT  1200600.0 1483200.0 1210800.0 1497000.0 ;
      RECT  1200600.0 1510800.0 1210800.0 1497000.0 ;
      RECT  1200600.0 1510800.0 1210800.0 1524600.0 ;
      RECT  1200600.0 1538400.0 1210800.0 1524600.0 ;
      RECT  1200600.0 1538400.0 1210800.0 1552200.0 ;
      RECT  1200600.0 1566000.0 1210800.0 1552200.0 ;
      RECT  1200600.0 1566000.0 1210800.0 1579800.0 ;
      RECT  1200600.0 1593600.0 1210800.0 1579800.0 ;
      RECT  1200600.0 1593600.0 1210800.0 1607400.0 ;
      RECT  1200600.0 1621200.0 1210800.0 1607400.0 ;
      RECT  1200600.0 1621200.0 1210800.0 1635000.0 ;
      RECT  1200600.0 1648800.0 1210800.0 1635000.0 ;
      RECT  1200600.0 1648800.0 1210800.0 1662600.0 ;
      RECT  1200600.0 1676400.0 1210800.0 1662600.0 ;
      RECT  1200600.0 1676400.0 1210800.0 1690200.0 ;
      RECT  1200600.0 1704000.0 1210800.0 1690200.0 ;
      RECT  1200600.0 1704000.0 1210800.0 1717800.0 ;
      RECT  1200600.0 1731600.0 1210800.0 1717800.0 ;
      RECT  1200600.0 1731600.0 1210800.0 1745400.0 ;
      RECT  1200600.0 1759200.0 1210800.0 1745400.0 ;
      RECT  1200600.0 1759200.0 1210800.0 1773000.0 ;
      RECT  1200600.0 1786800.0 1210800.0 1773000.0 ;
      RECT  1200600.0 1786800.0 1210800.0 1800600.0 ;
      RECT  1200600.0 1814400.0 1210800.0 1800600.0 ;
      RECT  1200600.0 1814400.0 1210800.0 1828200.0 ;
      RECT  1200600.0 1842000.0 1210800.0 1828200.0 ;
      RECT  1200600.0 1842000.0 1210800.0 1855800.0 ;
      RECT  1200600.0 1869600.0 1210800.0 1855800.0 ;
      RECT  1200600.0 1869600.0 1210800.0 1883400.0 ;
      RECT  1200600.0 1897200.0 1210800.0 1883400.0 ;
      RECT  1200600.0 1897200.0 1210800.0 1911000.0 ;
      RECT  1200600.0 1924800.0 1210800.0 1911000.0 ;
      RECT  1200600.0 1924800.0 1210800.0 1938600.0 ;
      RECT  1200600.0 1952400.0 1210800.0 1938600.0 ;
      RECT  1200600.0 1952400.0 1210800.0 1966200.0 ;
      RECT  1200600.0 1980000.0 1210800.0 1966200.0 ;
      RECT  1200600.0 1980000.0 1210800.0 1993800.0 ;
      RECT  1200600.0 2007600.0 1210800.0 1993800.0 ;
      RECT  1200600.0 2007600.0 1210800.0 2021400.0 ;
      RECT  1200600.0 2035200.0 1210800.0 2021400.0 ;
      RECT  1200600.0 2035200.0 1210800.0 2049000.0 ;
      RECT  1200600.0 2062800.0 1210800.0 2049000.0 ;
      RECT  1200600.0 2062800.0 1210800.0 2076600.0 ;
      RECT  1200600.0 2090400.0 1210800.0 2076600.0 ;
      RECT  1200600.0 2090400.0 1210800.0 2104200.0 ;
      RECT  1200600.0 2118000.0 1210800.0 2104200.0 ;
      RECT  1200600.0 2118000.0 1210800.0 2131800.0 ;
      RECT  1200600.0 2145600.0 1210800.0 2131800.0 ;
      RECT  1210800.0 379200.0 1221000.0 393000.0 ;
      RECT  1210800.0 406800.0 1221000.0 393000.0 ;
      RECT  1210800.0 406800.0 1221000.0 420600.0 ;
      RECT  1210800.0 434400.0 1221000.0 420600.0 ;
      RECT  1210800.0 434400.0 1221000.0 448200.0 ;
      RECT  1210800.0 462000.0 1221000.0 448200.0 ;
      RECT  1210800.0 462000.0 1221000.0 475800.0 ;
      RECT  1210800.0 489600.0 1221000.0 475800.0 ;
      RECT  1210800.0 489600.0 1221000.0 503400.0 ;
      RECT  1210800.0 517200.0 1221000.0 503400.0 ;
      RECT  1210800.0 517200.0 1221000.0 531000.0 ;
      RECT  1210800.0 544800.0 1221000.0 531000.0 ;
      RECT  1210800.0 544800.0 1221000.0 558600.0 ;
      RECT  1210800.0 572400.0 1221000.0 558600.0 ;
      RECT  1210800.0 572400.0 1221000.0 586200.0 ;
      RECT  1210800.0 600000.0 1221000.0 586200.0 ;
      RECT  1210800.0 600000.0 1221000.0 613800.0 ;
      RECT  1210800.0 627600.0 1221000.0 613800.0 ;
      RECT  1210800.0 627600.0 1221000.0 641400.0 ;
      RECT  1210800.0 655200.0 1221000.0 641400.0 ;
      RECT  1210800.0 655200.0 1221000.0 669000.0 ;
      RECT  1210800.0 682800.0 1221000.0 669000.0 ;
      RECT  1210800.0 682800.0 1221000.0 696600.0 ;
      RECT  1210800.0 710400.0 1221000.0 696600.0 ;
      RECT  1210800.0 710400.0 1221000.0 724200.0 ;
      RECT  1210800.0 738000.0 1221000.0 724200.0 ;
      RECT  1210800.0 738000.0 1221000.0 751800.0 ;
      RECT  1210800.0 765600.0 1221000.0 751800.0 ;
      RECT  1210800.0 765600.0 1221000.0 779400.0 ;
      RECT  1210800.0 793200.0 1221000.0 779400.0 ;
      RECT  1210800.0 793200.0 1221000.0 807000.0 ;
      RECT  1210800.0 820800.0 1221000.0 807000.0 ;
      RECT  1210800.0 820800.0 1221000.0 834600.0 ;
      RECT  1210800.0 848400.0 1221000.0 834600.0 ;
      RECT  1210800.0 848400.0 1221000.0 862200.0 ;
      RECT  1210800.0 876000.0 1221000.0 862200.0 ;
      RECT  1210800.0 876000.0 1221000.0 889800.0 ;
      RECT  1210800.0 903600.0 1221000.0 889800.0 ;
      RECT  1210800.0 903600.0 1221000.0 917400.0 ;
      RECT  1210800.0 931200.0 1221000.0 917400.0 ;
      RECT  1210800.0 931200.0 1221000.0 945000.0 ;
      RECT  1210800.0 958800.0 1221000.0 945000.0 ;
      RECT  1210800.0 958800.0 1221000.0 972600.0 ;
      RECT  1210800.0 986400.0 1221000.0 972600.0 ;
      RECT  1210800.0 986400.0 1221000.0 1000200.0 ;
      RECT  1210800.0 1014000.0 1221000.0 1000200.0 ;
      RECT  1210800.0 1014000.0 1221000.0 1027800.0 ;
      RECT  1210800.0 1041600.0 1221000.0 1027800.0 ;
      RECT  1210800.0 1041600.0 1221000.0 1055400.0 ;
      RECT  1210800.0 1069200.0 1221000.0 1055400.0 ;
      RECT  1210800.0 1069200.0 1221000.0 1083000.0 ;
      RECT  1210800.0 1096800.0 1221000.0 1083000.0 ;
      RECT  1210800.0 1096800.0 1221000.0 1110600.0 ;
      RECT  1210800.0 1124400.0 1221000.0 1110600.0 ;
      RECT  1210800.0 1124400.0 1221000.0 1138200.0 ;
      RECT  1210800.0 1152000.0 1221000.0 1138200.0 ;
      RECT  1210800.0 1152000.0 1221000.0 1165800.0 ;
      RECT  1210800.0 1179600.0 1221000.0 1165800.0 ;
      RECT  1210800.0 1179600.0 1221000.0 1193400.0 ;
      RECT  1210800.0 1207200.0 1221000.0 1193400.0 ;
      RECT  1210800.0 1207200.0 1221000.0 1221000.0 ;
      RECT  1210800.0 1234800.0 1221000.0 1221000.0 ;
      RECT  1210800.0 1234800.0 1221000.0 1248600.0 ;
      RECT  1210800.0 1262400.0 1221000.0 1248600.0 ;
      RECT  1210800.0 1262400.0 1221000.0 1276200.0 ;
      RECT  1210800.0 1290000.0 1221000.0 1276200.0 ;
      RECT  1210800.0 1290000.0 1221000.0 1303800.0 ;
      RECT  1210800.0 1317600.0 1221000.0 1303800.0 ;
      RECT  1210800.0 1317600.0 1221000.0 1331400.0 ;
      RECT  1210800.0 1345200.0 1221000.0 1331400.0 ;
      RECT  1210800.0 1345200.0 1221000.0 1359000.0 ;
      RECT  1210800.0 1372800.0 1221000.0 1359000.0 ;
      RECT  1210800.0 1372800.0 1221000.0 1386600.0 ;
      RECT  1210800.0 1400400.0 1221000.0 1386600.0 ;
      RECT  1210800.0 1400400.0 1221000.0 1414200.0 ;
      RECT  1210800.0 1428000.0 1221000.0 1414200.0 ;
      RECT  1210800.0 1428000.0 1221000.0 1441800.0 ;
      RECT  1210800.0 1455600.0 1221000.0 1441800.0 ;
      RECT  1210800.0 1455600.0 1221000.0 1469400.0 ;
      RECT  1210800.0 1483200.0 1221000.0 1469400.0 ;
      RECT  1210800.0 1483200.0 1221000.0 1497000.0 ;
      RECT  1210800.0 1510800.0 1221000.0 1497000.0 ;
      RECT  1210800.0 1510800.0 1221000.0 1524600.0 ;
      RECT  1210800.0 1538400.0 1221000.0 1524600.0 ;
      RECT  1210800.0 1538400.0 1221000.0 1552200.0 ;
      RECT  1210800.0 1566000.0 1221000.0 1552200.0 ;
      RECT  1210800.0 1566000.0 1221000.0 1579800.0 ;
      RECT  1210800.0 1593600.0 1221000.0 1579800.0 ;
      RECT  1210800.0 1593600.0 1221000.0 1607400.0 ;
      RECT  1210800.0 1621200.0 1221000.0 1607400.0 ;
      RECT  1210800.0 1621200.0 1221000.0 1635000.0 ;
      RECT  1210800.0 1648800.0 1221000.0 1635000.0 ;
      RECT  1210800.0 1648800.0 1221000.0 1662600.0 ;
      RECT  1210800.0 1676400.0 1221000.0 1662600.0 ;
      RECT  1210800.0 1676400.0 1221000.0 1690200.0 ;
      RECT  1210800.0 1704000.0 1221000.0 1690200.0 ;
      RECT  1210800.0 1704000.0 1221000.0 1717800.0 ;
      RECT  1210800.0 1731600.0 1221000.0 1717800.0 ;
      RECT  1210800.0 1731600.0 1221000.0 1745400.0 ;
      RECT  1210800.0 1759200.0 1221000.0 1745400.0 ;
      RECT  1210800.0 1759200.0 1221000.0 1773000.0 ;
      RECT  1210800.0 1786800.0 1221000.0 1773000.0 ;
      RECT  1210800.0 1786800.0 1221000.0 1800600.0 ;
      RECT  1210800.0 1814400.0 1221000.0 1800600.0 ;
      RECT  1210800.0 1814400.0 1221000.0 1828200.0 ;
      RECT  1210800.0 1842000.0 1221000.0 1828200.0 ;
      RECT  1210800.0 1842000.0 1221000.0 1855800.0 ;
      RECT  1210800.0 1869600.0 1221000.0 1855800.0 ;
      RECT  1210800.0 1869600.0 1221000.0 1883400.0 ;
      RECT  1210800.0 1897200.0 1221000.0 1883400.0 ;
      RECT  1210800.0 1897200.0 1221000.0 1911000.0 ;
      RECT  1210800.0 1924800.0 1221000.0 1911000.0 ;
      RECT  1210800.0 1924800.0 1221000.0 1938600.0 ;
      RECT  1210800.0 1952400.0 1221000.0 1938600.0 ;
      RECT  1210800.0 1952400.0 1221000.0 1966200.0 ;
      RECT  1210800.0 1980000.0 1221000.0 1966200.0 ;
      RECT  1210800.0 1980000.0 1221000.0 1993800.0 ;
      RECT  1210800.0 2007600.0 1221000.0 1993800.0 ;
      RECT  1210800.0 2007600.0 1221000.0 2021400.0 ;
      RECT  1210800.0 2035200.0 1221000.0 2021400.0 ;
      RECT  1210800.0 2035200.0 1221000.0 2049000.0 ;
      RECT  1210800.0 2062800.0 1221000.0 2049000.0 ;
      RECT  1210800.0 2062800.0 1221000.0 2076600.0 ;
      RECT  1210800.0 2090400.0 1221000.0 2076600.0 ;
      RECT  1210800.0 2090400.0 1221000.0 2104200.0 ;
      RECT  1210800.0 2118000.0 1221000.0 2104200.0 ;
      RECT  1210800.0 2118000.0 1221000.0 2131800.0 ;
      RECT  1210800.0 2145600.0 1221000.0 2131800.0 ;
      RECT  1221000.0 379200.0 1231200.0 393000.0 ;
      RECT  1221000.0 406800.0 1231200.0 393000.0 ;
      RECT  1221000.0 406800.0 1231200.0 420600.0 ;
      RECT  1221000.0 434400.0 1231200.0 420600.0 ;
      RECT  1221000.0 434400.0 1231200.0 448200.0 ;
      RECT  1221000.0 462000.0 1231200.0 448200.0 ;
      RECT  1221000.0 462000.0 1231200.0 475800.0 ;
      RECT  1221000.0 489600.0 1231200.0 475800.0 ;
      RECT  1221000.0 489600.0 1231200.0 503400.0 ;
      RECT  1221000.0 517200.0 1231200.0 503400.0 ;
      RECT  1221000.0 517200.0 1231200.0 531000.0 ;
      RECT  1221000.0 544800.0 1231200.0 531000.0 ;
      RECT  1221000.0 544800.0 1231200.0 558600.0 ;
      RECT  1221000.0 572400.0 1231200.0 558600.0 ;
      RECT  1221000.0 572400.0 1231200.0 586200.0 ;
      RECT  1221000.0 600000.0 1231200.0 586200.0 ;
      RECT  1221000.0 600000.0 1231200.0 613800.0 ;
      RECT  1221000.0 627600.0 1231200.0 613800.0 ;
      RECT  1221000.0 627600.0 1231200.0 641400.0 ;
      RECT  1221000.0 655200.0 1231200.0 641400.0 ;
      RECT  1221000.0 655200.0 1231200.0 669000.0 ;
      RECT  1221000.0 682800.0 1231200.0 669000.0 ;
      RECT  1221000.0 682800.0 1231200.0 696600.0 ;
      RECT  1221000.0 710400.0 1231200.0 696600.0 ;
      RECT  1221000.0 710400.0 1231200.0 724200.0 ;
      RECT  1221000.0 738000.0 1231200.0 724200.0 ;
      RECT  1221000.0 738000.0 1231200.0 751800.0 ;
      RECT  1221000.0 765600.0 1231200.0 751800.0 ;
      RECT  1221000.0 765600.0 1231200.0 779400.0 ;
      RECT  1221000.0 793200.0 1231200.0 779400.0 ;
      RECT  1221000.0 793200.0 1231200.0 807000.0 ;
      RECT  1221000.0 820800.0 1231200.0 807000.0 ;
      RECT  1221000.0 820800.0 1231200.0 834600.0 ;
      RECT  1221000.0 848400.0 1231200.0 834600.0 ;
      RECT  1221000.0 848400.0 1231200.0 862200.0 ;
      RECT  1221000.0 876000.0 1231200.0 862200.0 ;
      RECT  1221000.0 876000.0 1231200.0 889800.0 ;
      RECT  1221000.0 903600.0 1231200.0 889800.0 ;
      RECT  1221000.0 903600.0 1231200.0 917400.0 ;
      RECT  1221000.0 931200.0 1231200.0 917400.0 ;
      RECT  1221000.0 931200.0 1231200.0 945000.0 ;
      RECT  1221000.0 958800.0 1231200.0 945000.0 ;
      RECT  1221000.0 958800.0 1231200.0 972600.0 ;
      RECT  1221000.0 986400.0 1231200.0 972600.0 ;
      RECT  1221000.0 986400.0 1231200.0 1000200.0 ;
      RECT  1221000.0 1014000.0 1231200.0 1000200.0 ;
      RECT  1221000.0 1014000.0 1231200.0 1027800.0 ;
      RECT  1221000.0 1041600.0 1231200.0 1027800.0 ;
      RECT  1221000.0 1041600.0 1231200.0 1055400.0 ;
      RECT  1221000.0 1069200.0 1231200.0 1055400.0 ;
      RECT  1221000.0 1069200.0 1231200.0 1083000.0 ;
      RECT  1221000.0 1096800.0 1231200.0 1083000.0 ;
      RECT  1221000.0 1096800.0 1231200.0 1110600.0 ;
      RECT  1221000.0 1124400.0 1231200.0 1110600.0 ;
      RECT  1221000.0 1124400.0 1231200.0 1138200.0 ;
      RECT  1221000.0 1152000.0 1231200.0 1138200.0 ;
      RECT  1221000.0 1152000.0 1231200.0 1165800.0 ;
      RECT  1221000.0 1179600.0 1231200.0 1165800.0 ;
      RECT  1221000.0 1179600.0 1231200.0 1193400.0 ;
      RECT  1221000.0 1207200.0 1231200.0 1193400.0 ;
      RECT  1221000.0 1207200.0 1231200.0 1221000.0 ;
      RECT  1221000.0 1234800.0 1231200.0 1221000.0 ;
      RECT  1221000.0 1234800.0 1231200.0 1248600.0 ;
      RECT  1221000.0 1262400.0 1231200.0 1248600.0 ;
      RECT  1221000.0 1262400.0 1231200.0 1276200.0 ;
      RECT  1221000.0 1290000.0 1231200.0 1276200.0 ;
      RECT  1221000.0 1290000.0 1231200.0 1303800.0 ;
      RECT  1221000.0 1317600.0 1231200.0 1303800.0 ;
      RECT  1221000.0 1317600.0 1231200.0 1331400.0 ;
      RECT  1221000.0 1345200.0 1231200.0 1331400.0 ;
      RECT  1221000.0 1345200.0 1231200.0 1359000.0 ;
      RECT  1221000.0 1372800.0 1231200.0 1359000.0 ;
      RECT  1221000.0 1372800.0 1231200.0 1386600.0 ;
      RECT  1221000.0 1400400.0 1231200.0 1386600.0 ;
      RECT  1221000.0 1400400.0 1231200.0 1414200.0 ;
      RECT  1221000.0 1428000.0 1231200.0 1414200.0 ;
      RECT  1221000.0 1428000.0 1231200.0 1441800.0 ;
      RECT  1221000.0 1455600.0 1231200.0 1441800.0 ;
      RECT  1221000.0 1455600.0 1231200.0 1469400.0 ;
      RECT  1221000.0 1483200.0 1231200.0 1469400.0 ;
      RECT  1221000.0 1483200.0 1231200.0 1497000.0 ;
      RECT  1221000.0 1510800.0 1231200.0 1497000.0 ;
      RECT  1221000.0 1510800.0 1231200.0 1524600.0 ;
      RECT  1221000.0 1538400.0 1231200.0 1524600.0 ;
      RECT  1221000.0 1538400.0 1231200.0 1552200.0 ;
      RECT  1221000.0 1566000.0 1231200.0 1552200.0 ;
      RECT  1221000.0 1566000.0 1231200.0 1579800.0 ;
      RECT  1221000.0 1593600.0 1231200.0 1579800.0 ;
      RECT  1221000.0 1593600.0 1231200.0 1607400.0 ;
      RECT  1221000.0 1621200.0 1231200.0 1607400.0 ;
      RECT  1221000.0 1621200.0 1231200.0 1635000.0 ;
      RECT  1221000.0 1648800.0 1231200.0 1635000.0 ;
      RECT  1221000.0 1648800.0 1231200.0 1662600.0 ;
      RECT  1221000.0 1676400.0 1231200.0 1662600.0 ;
      RECT  1221000.0 1676400.0 1231200.0 1690200.0 ;
      RECT  1221000.0 1704000.0 1231200.0 1690200.0 ;
      RECT  1221000.0 1704000.0 1231200.0 1717800.0 ;
      RECT  1221000.0 1731600.0 1231200.0 1717800.0 ;
      RECT  1221000.0 1731600.0 1231200.0 1745400.0 ;
      RECT  1221000.0 1759200.0 1231200.0 1745400.0 ;
      RECT  1221000.0 1759200.0 1231200.0 1773000.0 ;
      RECT  1221000.0 1786800.0 1231200.0 1773000.0 ;
      RECT  1221000.0 1786800.0 1231200.0 1800600.0 ;
      RECT  1221000.0 1814400.0 1231200.0 1800600.0 ;
      RECT  1221000.0 1814400.0 1231200.0 1828200.0 ;
      RECT  1221000.0 1842000.0 1231200.0 1828200.0 ;
      RECT  1221000.0 1842000.0 1231200.0 1855800.0 ;
      RECT  1221000.0 1869600.0 1231200.0 1855800.0 ;
      RECT  1221000.0 1869600.0 1231200.0 1883400.0 ;
      RECT  1221000.0 1897200.0 1231200.0 1883400.0 ;
      RECT  1221000.0 1897200.0 1231200.0 1911000.0 ;
      RECT  1221000.0 1924800.0 1231200.0 1911000.0 ;
      RECT  1221000.0 1924800.0 1231200.0 1938600.0 ;
      RECT  1221000.0 1952400.0 1231200.0 1938600.0 ;
      RECT  1221000.0 1952400.0 1231200.0 1966200.0 ;
      RECT  1221000.0 1980000.0 1231200.0 1966200.0 ;
      RECT  1221000.0 1980000.0 1231200.0 1993800.0 ;
      RECT  1221000.0 2007600.0 1231200.0 1993800.0 ;
      RECT  1221000.0 2007600.0 1231200.0 2021400.0 ;
      RECT  1221000.0 2035200.0 1231200.0 2021400.0 ;
      RECT  1221000.0 2035200.0 1231200.0 2049000.0 ;
      RECT  1221000.0 2062800.0 1231200.0 2049000.0 ;
      RECT  1221000.0 2062800.0 1231200.0 2076600.0 ;
      RECT  1221000.0 2090400.0 1231200.0 2076600.0 ;
      RECT  1221000.0 2090400.0 1231200.0 2104200.0 ;
      RECT  1221000.0 2118000.0 1231200.0 2104200.0 ;
      RECT  1221000.0 2118000.0 1231200.0 2131800.0 ;
      RECT  1221000.0 2145600.0 1231200.0 2131800.0 ;
      RECT  1231200.0 379200.0 1241400.0 393000.0 ;
      RECT  1231200.0 406800.0 1241400.0 393000.0 ;
      RECT  1231200.0 406800.0 1241400.0 420600.0 ;
      RECT  1231200.0 434400.0 1241400.0 420600.0 ;
      RECT  1231200.0 434400.0 1241400.0 448200.0 ;
      RECT  1231200.0 462000.0 1241400.0 448200.0 ;
      RECT  1231200.0 462000.0 1241400.0 475800.0 ;
      RECT  1231200.0 489600.0 1241400.0 475800.0 ;
      RECT  1231200.0 489600.0 1241400.0 503400.0 ;
      RECT  1231200.0 517200.0 1241400.0 503400.0 ;
      RECT  1231200.0 517200.0 1241400.0 531000.0 ;
      RECT  1231200.0 544800.0 1241400.0 531000.0 ;
      RECT  1231200.0 544800.0 1241400.0 558600.0 ;
      RECT  1231200.0 572400.0 1241400.0 558600.0 ;
      RECT  1231200.0 572400.0 1241400.0 586200.0 ;
      RECT  1231200.0 600000.0 1241400.0 586200.0 ;
      RECT  1231200.0 600000.0 1241400.0 613800.0 ;
      RECT  1231200.0 627600.0 1241400.0 613800.0 ;
      RECT  1231200.0 627600.0 1241400.0 641400.0 ;
      RECT  1231200.0 655200.0 1241400.0 641400.0 ;
      RECT  1231200.0 655200.0 1241400.0 669000.0 ;
      RECT  1231200.0 682800.0 1241400.0 669000.0 ;
      RECT  1231200.0 682800.0 1241400.0 696600.0 ;
      RECT  1231200.0 710400.0 1241400.0 696600.0 ;
      RECT  1231200.0 710400.0 1241400.0 724200.0 ;
      RECT  1231200.0 738000.0 1241400.0 724200.0 ;
      RECT  1231200.0 738000.0 1241400.0 751800.0 ;
      RECT  1231200.0 765600.0 1241400.0 751800.0 ;
      RECT  1231200.0 765600.0 1241400.0 779400.0 ;
      RECT  1231200.0 793200.0 1241400.0 779400.0 ;
      RECT  1231200.0 793200.0 1241400.0 807000.0 ;
      RECT  1231200.0 820800.0 1241400.0 807000.0 ;
      RECT  1231200.0 820800.0 1241400.0 834600.0 ;
      RECT  1231200.0 848400.0 1241400.0 834600.0 ;
      RECT  1231200.0 848400.0 1241400.0 862200.0 ;
      RECT  1231200.0 876000.0 1241400.0 862200.0 ;
      RECT  1231200.0 876000.0 1241400.0 889800.0 ;
      RECT  1231200.0 903600.0 1241400.0 889800.0 ;
      RECT  1231200.0 903600.0 1241400.0 917400.0 ;
      RECT  1231200.0 931200.0 1241400.0 917400.0 ;
      RECT  1231200.0 931200.0 1241400.0 945000.0 ;
      RECT  1231200.0 958800.0 1241400.0 945000.0 ;
      RECT  1231200.0 958800.0 1241400.0 972600.0 ;
      RECT  1231200.0 986400.0 1241400.0 972600.0 ;
      RECT  1231200.0 986400.0 1241400.0 1000200.0 ;
      RECT  1231200.0 1014000.0 1241400.0 1000200.0 ;
      RECT  1231200.0 1014000.0 1241400.0 1027800.0 ;
      RECT  1231200.0 1041600.0 1241400.0 1027800.0 ;
      RECT  1231200.0 1041600.0 1241400.0 1055400.0 ;
      RECT  1231200.0 1069200.0 1241400.0 1055400.0 ;
      RECT  1231200.0 1069200.0 1241400.0 1083000.0 ;
      RECT  1231200.0 1096800.0 1241400.0 1083000.0 ;
      RECT  1231200.0 1096800.0 1241400.0 1110600.0 ;
      RECT  1231200.0 1124400.0 1241400.0 1110600.0 ;
      RECT  1231200.0 1124400.0 1241400.0 1138200.0 ;
      RECT  1231200.0 1152000.0 1241400.0 1138200.0 ;
      RECT  1231200.0 1152000.0 1241400.0 1165800.0 ;
      RECT  1231200.0 1179600.0 1241400.0 1165800.0 ;
      RECT  1231200.0 1179600.0 1241400.0 1193400.0 ;
      RECT  1231200.0 1207200.0 1241400.0 1193400.0 ;
      RECT  1231200.0 1207200.0 1241400.0 1221000.0 ;
      RECT  1231200.0 1234800.0 1241400.0 1221000.0 ;
      RECT  1231200.0 1234800.0 1241400.0 1248600.0 ;
      RECT  1231200.0 1262400.0 1241400.0 1248600.0 ;
      RECT  1231200.0 1262400.0 1241400.0 1276200.0 ;
      RECT  1231200.0 1290000.0 1241400.0 1276200.0 ;
      RECT  1231200.0 1290000.0 1241400.0 1303800.0 ;
      RECT  1231200.0 1317600.0 1241400.0 1303800.0 ;
      RECT  1231200.0 1317600.0 1241400.0 1331400.0 ;
      RECT  1231200.0 1345200.0 1241400.0 1331400.0 ;
      RECT  1231200.0 1345200.0 1241400.0 1359000.0 ;
      RECT  1231200.0 1372800.0 1241400.0 1359000.0 ;
      RECT  1231200.0 1372800.0 1241400.0 1386600.0 ;
      RECT  1231200.0 1400400.0 1241400.0 1386600.0 ;
      RECT  1231200.0 1400400.0 1241400.0 1414200.0 ;
      RECT  1231200.0 1428000.0 1241400.0 1414200.0 ;
      RECT  1231200.0 1428000.0 1241400.0 1441800.0 ;
      RECT  1231200.0 1455600.0 1241400.0 1441800.0 ;
      RECT  1231200.0 1455600.0 1241400.0 1469400.0 ;
      RECT  1231200.0 1483200.0 1241400.0 1469400.0 ;
      RECT  1231200.0 1483200.0 1241400.0 1497000.0 ;
      RECT  1231200.0 1510800.0 1241400.0 1497000.0 ;
      RECT  1231200.0 1510800.0 1241400.0 1524600.0 ;
      RECT  1231200.0 1538400.0 1241400.0 1524600.0 ;
      RECT  1231200.0 1538400.0 1241400.0 1552200.0 ;
      RECT  1231200.0 1566000.0 1241400.0 1552200.0 ;
      RECT  1231200.0 1566000.0 1241400.0 1579800.0 ;
      RECT  1231200.0 1593600.0 1241400.0 1579800.0 ;
      RECT  1231200.0 1593600.0 1241400.0 1607400.0 ;
      RECT  1231200.0 1621200.0 1241400.0 1607400.0 ;
      RECT  1231200.0 1621200.0 1241400.0 1635000.0 ;
      RECT  1231200.0 1648800.0 1241400.0 1635000.0 ;
      RECT  1231200.0 1648800.0 1241400.0 1662600.0 ;
      RECT  1231200.0 1676400.0 1241400.0 1662600.0 ;
      RECT  1231200.0 1676400.0 1241400.0 1690200.0 ;
      RECT  1231200.0 1704000.0 1241400.0 1690200.0 ;
      RECT  1231200.0 1704000.0 1241400.0 1717800.0 ;
      RECT  1231200.0 1731600.0 1241400.0 1717800.0 ;
      RECT  1231200.0 1731600.0 1241400.0 1745400.0 ;
      RECT  1231200.0 1759200.0 1241400.0 1745400.0 ;
      RECT  1231200.0 1759200.0 1241400.0 1773000.0 ;
      RECT  1231200.0 1786800.0 1241400.0 1773000.0 ;
      RECT  1231200.0 1786800.0 1241400.0 1800600.0 ;
      RECT  1231200.0 1814400.0 1241400.0 1800600.0 ;
      RECT  1231200.0 1814400.0 1241400.0 1828200.0 ;
      RECT  1231200.0 1842000.0 1241400.0 1828200.0 ;
      RECT  1231200.0 1842000.0 1241400.0 1855800.0 ;
      RECT  1231200.0 1869600.0 1241400.0 1855800.0 ;
      RECT  1231200.0 1869600.0 1241400.0 1883400.0 ;
      RECT  1231200.0 1897200.0 1241400.0 1883400.0 ;
      RECT  1231200.0 1897200.0 1241400.0 1911000.0 ;
      RECT  1231200.0 1924800.0 1241400.0 1911000.0 ;
      RECT  1231200.0 1924800.0 1241400.0 1938600.0 ;
      RECT  1231200.0 1952400.0 1241400.0 1938600.0 ;
      RECT  1231200.0 1952400.0 1241400.0 1966200.0 ;
      RECT  1231200.0 1980000.0 1241400.0 1966200.0 ;
      RECT  1231200.0 1980000.0 1241400.0 1993800.0 ;
      RECT  1231200.0 2007600.0 1241400.0 1993800.0 ;
      RECT  1231200.0 2007600.0 1241400.0 2021400.0 ;
      RECT  1231200.0 2035200.0 1241400.0 2021400.0 ;
      RECT  1231200.0 2035200.0 1241400.0 2049000.0 ;
      RECT  1231200.0 2062800.0 1241400.0 2049000.0 ;
      RECT  1231200.0 2062800.0 1241400.0 2076600.0 ;
      RECT  1231200.0 2090400.0 1241400.0 2076600.0 ;
      RECT  1231200.0 2090400.0 1241400.0 2104200.0 ;
      RECT  1231200.0 2118000.0 1241400.0 2104200.0 ;
      RECT  1231200.0 2118000.0 1241400.0 2131800.0 ;
      RECT  1231200.0 2145600.0 1241400.0 2131800.0 ;
      RECT  1241400.0 379200.0 1251600.0 393000.0 ;
      RECT  1241400.0 406800.0 1251600.0 393000.0 ;
      RECT  1241400.0 406800.0 1251600.0 420600.0 ;
      RECT  1241400.0 434400.0 1251600.0 420600.0 ;
      RECT  1241400.0 434400.0 1251600.0 448200.0 ;
      RECT  1241400.0 462000.0 1251600.0 448200.0 ;
      RECT  1241400.0 462000.0 1251600.0 475800.0 ;
      RECT  1241400.0 489600.0 1251600.0 475800.0 ;
      RECT  1241400.0 489600.0 1251600.0 503400.0 ;
      RECT  1241400.0 517200.0 1251600.0 503400.0 ;
      RECT  1241400.0 517200.0 1251600.0 531000.0 ;
      RECT  1241400.0 544800.0 1251600.0 531000.0 ;
      RECT  1241400.0 544800.0 1251600.0 558600.0 ;
      RECT  1241400.0 572400.0 1251600.0 558600.0 ;
      RECT  1241400.0 572400.0 1251600.0 586200.0 ;
      RECT  1241400.0 600000.0 1251600.0 586200.0 ;
      RECT  1241400.0 600000.0 1251600.0 613800.0 ;
      RECT  1241400.0 627600.0 1251600.0 613800.0 ;
      RECT  1241400.0 627600.0 1251600.0 641400.0 ;
      RECT  1241400.0 655200.0 1251600.0 641400.0 ;
      RECT  1241400.0 655200.0 1251600.0 669000.0 ;
      RECT  1241400.0 682800.0 1251600.0 669000.0 ;
      RECT  1241400.0 682800.0 1251600.0 696600.0 ;
      RECT  1241400.0 710400.0 1251600.0 696600.0 ;
      RECT  1241400.0 710400.0 1251600.0 724200.0 ;
      RECT  1241400.0 738000.0 1251600.0 724200.0 ;
      RECT  1241400.0 738000.0 1251600.0 751800.0 ;
      RECT  1241400.0 765600.0 1251600.0 751800.0 ;
      RECT  1241400.0 765600.0 1251600.0 779400.0 ;
      RECT  1241400.0 793200.0 1251600.0 779400.0 ;
      RECT  1241400.0 793200.0 1251600.0 807000.0 ;
      RECT  1241400.0 820800.0 1251600.0 807000.0 ;
      RECT  1241400.0 820800.0 1251600.0 834600.0 ;
      RECT  1241400.0 848400.0 1251600.0 834600.0 ;
      RECT  1241400.0 848400.0 1251600.0 862200.0 ;
      RECT  1241400.0 876000.0 1251600.0 862200.0 ;
      RECT  1241400.0 876000.0 1251600.0 889800.0 ;
      RECT  1241400.0 903600.0 1251600.0 889800.0 ;
      RECT  1241400.0 903600.0 1251600.0 917400.0 ;
      RECT  1241400.0 931200.0 1251600.0 917400.0 ;
      RECT  1241400.0 931200.0 1251600.0 945000.0 ;
      RECT  1241400.0 958800.0 1251600.0 945000.0 ;
      RECT  1241400.0 958800.0 1251600.0 972600.0 ;
      RECT  1241400.0 986400.0 1251600.0 972600.0 ;
      RECT  1241400.0 986400.0 1251600.0 1000200.0 ;
      RECT  1241400.0 1014000.0 1251600.0 1000200.0 ;
      RECT  1241400.0 1014000.0 1251600.0 1027800.0 ;
      RECT  1241400.0 1041600.0 1251600.0 1027800.0 ;
      RECT  1241400.0 1041600.0 1251600.0 1055400.0 ;
      RECT  1241400.0 1069200.0 1251600.0 1055400.0 ;
      RECT  1241400.0 1069200.0 1251600.0 1083000.0 ;
      RECT  1241400.0 1096800.0 1251600.0 1083000.0 ;
      RECT  1241400.0 1096800.0 1251600.0 1110600.0 ;
      RECT  1241400.0 1124400.0 1251600.0 1110600.0 ;
      RECT  1241400.0 1124400.0 1251600.0 1138200.0 ;
      RECT  1241400.0 1152000.0 1251600.0 1138200.0 ;
      RECT  1241400.0 1152000.0 1251600.0 1165800.0 ;
      RECT  1241400.0 1179600.0 1251600.0 1165800.0 ;
      RECT  1241400.0 1179600.0 1251600.0 1193400.0 ;
      RECT  1241400.0 1207200.0 1251600.0 1193400.0 ;
      RECT  1241400.0 1207200.0 1251600.0 1221000.0 ;
      RECT  1241400.0 1234800.0 1251600.0 1221000.0 ;
      RECT  1241400.0 1234800.0 1251600.0 1248600.0 ;
      RECT  1241400.0 1262400.0 1251600.0 1248600.0 ;
      RECT  1241400.0 1262400.0 1251600.0 1276200.0 ;
      RECT  1241400.0 1290000.0 1251600.0 1276200.0 ;
      RECT  1241400.0 1290000.0 1251600.0 1303800.0 ;
      RECT  1241400.0 1317600.0 1251600.0 1303800.0 ;
      RECT  1241400.0 1317600.0 1251600.0 1331400.0 ;
      RECT  1241400.0 1345200.0 1251600.0 1331400.0 ;
      RECT  1241400.0 1345200.0 1251600.0 1359000.0 ;
      RECT  1241400.0 1372800.0 1251600.0 1359000.0 ;
      RECT  1241400.0 1372800.0 1251600.0 1386600.0 ;
      RECT  1241400.0 1400400.0 1251600.0 1386600.0 ;
      RECT  1241400.0 1400400.0 1251600.0 1414200.0 ;
      RECT  1241400.0 1428000.0 1251600.0 1414200.0 ;
      RECT  1241400.0 1428000.0 1251600.0 1441800.0 ;
      RECT  1241400.0 1455600.0 1251600.0 1441800.0 ;
      RECT  1241400.0 1455600.0 1251600.0 1469400.0 ;
      RECT  1241400.0 1483200.0 1251600.0 1469400.0 ;
      RECT  1241400.0 1483200.0 1251600.0 1497000.0 ;
      RECT  1241400.0 1510800.0 1251600.0 1497000.0 ;
      RECT  1241400.0 1510800.0 1251600.0 1524600.0 ;
      RECT  1241400.0 1538400.0 1251600.0 1524600.0 ;
      RECT  1241400.0 1538400.0 1251600.0 1552200.0 ;
      RECT  1241400.0 1566000.0 1251600.0 1552200.0 ;
      RECT  1241400.0 1566000.0 1251600.0 1579800.0 ;
      RECT  1241400.0 1593600.0 1251600.0 1579800.0 ;
      RECT  1241400.0 1593600.0 1251600.0 1607400.0 ;
      RECT  1241400.0 1621200.0 1251600.0 1607400.0 ;
      RECT  1241400.0 1621200.0 1251600.0 1635000.0 ;
      RECT  1241400.0 1648800.0 1251600.0 1635000.0 ;
      RECT  1241400.0 1648800.0 1251600.0 1662600.0 ;
      RECT  1241400.0 1676400.0 1251600.0 1662600.0 ;
      RECT  1241400.0 1676400.0 1251600.0 1690200.0 ;
      RECT  1241400.0 1704000.0 1251600.0 1690200.0 ;
      RECT  1241400.0 1704000.0 1251600.0 1717800.0 ;
      RECT  1241400.0 1731600.0 1251600.0 1717800.0 ;
      RECT  1241400.0 1731600.0 1251600.0 1745400.0 ;
      RECT  1241400.0 1759200.0 1251600.0 1745400.0 ;
      RECT  1241400.0 1759200.0 1251600.0 1773000.0 ;
      RECT  1241400.0 1786800.0 1251600.0 1773000.0 ;
      RECT  1241400.0 1786800.0 1251600.0 1800600.0 ;
      RECT  1241400.0 1814400.0 1251600.0 1800600.0 ;
      RECT  1241400.0 1814400.0 1251600.0 1828200.0 ;
      RECT  1241400.0 1842000.0 1251600.0 1828200.0 ;
      RECT  1241400.0 1842000.0 1251600.0 1855800.0 ;
      RECT  1241400.0 1869600.0 1251600.0 1855800.0 ;
      RECT  1241400.0 1869600.0 1251600.0 1883400.0 ;
      RECT  1241400.0 1897200.0 1251600.0 1883400.0 ;
      RECT  1241400.0 1897200.0 1251600.0 1911000.0 ;
      RECT  1241400.0 1924800.0 1251600.0 1911000.0 ;
      RECT  1241400.0 1924800.0 1251600.0 1938600.0 ;
      RECT  1241400.0 1952400.0 1251600.0 1938600.0 ;
      RECT  1241400.0 1952400.0 1251600.0 1966200.0 ;
      RECT  1241400.0 1980000.0 1251600.0 1966200.0 ;
      RECT  1241400.0 1980000.0 1251600.0 1993800.0 ;
      RECT  1241400.0 2007600.0 1251600.0 1993800.0 ;
      RECT  1241400.0 2007600.0 1251600.0 2021400.0 ;
      RECT  1241400.0 2035200.0 1251600.0 2021400.0 ;
      RECT  1241400.0 2035200.0 1251600.0 2049000.0 ;
      RECT  1241400.0 2062800.0 1251600.0 2049000.0 ;
      RECT  1241400.0 2062800.0 1251600.0 2076600.0 ;
      RECT  1241400.0 2090400.0 1251600.0 2076600.0 ;
      RECT  1241400.0 2090400.0 1251600.0 2104200.0 ;
      RECT  1241400.0 2118000.0 1251600.0 2104200.0 ;
      RECT  1241400.0 2118000.0 1251600.0 2131800.0 ;
      RECT  1241400.0 2145600.0 1251600.0 2131800.0 ;
      RECT  1251600.0 379200.0 1261800.0 393000.0 ;
      RECT  1251600.0 406800.0 1261800.0 393000.0 ;
      RECT  1251600.0 406800.0 1261800.0 420600.0 ;
      RECT  1251600.0 434400.0 1261800.0 420600.0 ;
      RECT  1251600.0 434400.0 1261800.0 448200.0 ;
      RECT  1251600.0 462000.0 1261800.0 448200.0 ;
      RECT  1251600.0 462000.0 1261800.0 475800.0 ;
      RECT  1251600.0 489600.0 1261800.0 475800.0 ;
      RECT  1251600.0 489600.0 1261800.0 503400.0 ;
      RECT  1251600.0 517200.0 1261800.0 503400.0 ;
      RECT  1251600.0 517200.0 1261800.0 531000.0 ;
      RECT  1251600.0 544800.0 1261800.0 531000.0 ;
      RECT  1251600.0 544800.0 1261800.0 558600.0 ;
      RECT  1251600.0 572400.0 1261800.0 558600.0 ;
      RECT  1251600.0 572400.0 1261800.0 586200.0 ;
      RECT  1251600.0 600000.0 1261800.0 586200.0 ;
      RECT  1251600.0 600000.0 1261800.0 613800.0 ;
      RECT  1251600.0 627600.0 1261800.0 613800.0 ;
      RECT  1251600.0 627600.0 1261800.0 641400.0 ;
      RECT  1251600.0 655200.0 1261800.0 641400.0 ;
      RECT  1251600.0 655200.0 1261800.0 669000.0 ;
      RECT  1251600.0 682800.0 1261800.0 669000.0 ;
      RECT  1251600.0 682800.0 1261800.0 696600.0 ;
      RECT  1251600.0 710400.0 1261800.0 696600.0 ;
      RECT  1251600.0 710400.0 1261800.0 724200.0 ;
      RECT  1251600.0 738000.0 1261800.0 724200.0 ;
      RECT  1251600.0 738000.0 1261800.0 751800.0 ;
      RECT  1251600.0 765600.0 1261800.0 751800.0 ;
      RECT  1251600.0 765600.0 1261800.0 779400.0 ;
      RECT  1251600.0 793200.0 1261800.0 779400.0 ;
      RECT  1251600.0 793200.0 1261800.0 807000.0 ;
      RECT  1251600.0 820800.0 1261800.0 807000.0 ;
      RECT  1251600.0 820800.0 1261800.0 834600.0 ;
      RECT  1251600.0 848400.0 1261800.0 834600.0 ;
      RECT  1251600.0 848400.0 1261800.0 862200.0 ;
      RECT  1251600.0 876000.0 1261800.0 862200.0 ;
      RECT  1251600.0 876000.0 1261800.0 889800.0 ;
      RECT  1251600.0 903600.0 1261800.0 889800.0 ;
      RECT  1251600.0 903600.0 1261800.0 917400.0 ;
      RECT  1251600.0 931200.0 1261800.0 917400.0 ;
      RECT  1251600.0 931200.0 1261800.0 945000.0 ;
      RECT  1251600.0 958800.0 1261800.0 945000.0 ;
      RECT  1251600.0 958800.0 1261800.0 972600.0 ;
      RECT  1251600.0 986400.0 1261800.0 972600.0 ;
      RECT  1251600.0 986400.0 1261800.0 1000200.0 ;
      RECT  1251600.0 1014000.0 1261800.0 1000200.0 ;
      RECT  1251600.0 1014000.0 1261800.0 1027800.0 ;
      RECT  1251600.0 1041600.0 1261800.0 1027800.0 ;
      RECT  1251600.0 1041600.0 1261800.0 1055400.0 ;
      RECT  1251600.0 1069200.0 1261800.0 1055400.0 ;
      RECT  1251600.0 1069200.0 1261800.0 1083000.0 ;
      RECT  1251600.0 1096800.0 1261800.0 1083000.0 ;
      RECT  1251600.0 1096800.0 1261800.0 1110600.0 ;
      RECT  1251600.0 1124400.0 1261800.0 1110600.0 ;
      RECT  1251600.0 1124400.0 1261800.0 1138200.0 ;
      RECT  1251600.0 1152000.0 1261800.0 1138200.0 ;
      RECT  1251600.0 1152000.0 1261800.0 1165800.0 ;
      RECT  1251600.0 1179600.0 1261800.0 1165800.0 ;
      RECT  1251600.0 1179600.0 1261800.0 1193400.0 ;
      RECT  1251600.0 1207200.0 1261800.0 1193400.0 ;
      RECT  1251600.0 1207200.0 1261800.0 1221000.0 ;
      RECT  1251600.0 1234800.0 1261800.0 1221000.0 ;
      RECT  1251600.0 1234800.0 1261800.0 1248600.0 ;
      RECT  1251600.0 1262400.0 1261800.0 1248600.0 ;
      RECT  1251600.0 1262400.0 1261800.0 1276200.0 ;
      RECT  1251600.0 1290000.0 1261800.0 1276200.0 ;
      RECT  1251600.0 1290000.0 1261800.0 1303800.0 ;
      RECT  1251600.0 1317600.0 1261800.0 1303800.0 ;
      RECT  1251600.0 1317600.0 1261800.0 1331400.0 ;
      RECT  1251600.0 1345200.0 1261800.0 1331400.0 ;
      RECT  1251600.0 1345200.0 1261800.0 1359000.0 ;
      RECT  1251600.0 1372800.0 1261800.0 1359000.0 ;
      RECT  1251600.0 1372800.0 1261800.0 1386600.0 ;
      RECT  1251600.0 1400400.0 1261800.0 1386600.0 ;
      RECT  1251600.0 1400400.0 1261800.0 1414200.0 ;
      RECT  1251600.0 1428000.0 1261800.0 1414200.0 ;
      RECT  1251600.0 1428000.0 1261800.0 1441800.0 ;
      RECT  1251600.0 1455600.0 1261800.0 1441800.0 ;
      RECT  1251600.0 1455600.0 1261800.0 1469400.0 ;
      RECT  1251600.0 1483200.0 1261800.0 1469400.0 ;
      RECT  1251600.0 1483200.0 1261800.0 1497000.0 ;
      RECT  1251600.0 1510800.0 1261800.0 1497000.0 ;
      RECT  1251600.0 1510800.0 1261800.0 1524600.0 ;
      RECT  1251600.0 1538400.0 1261800.0 1524600.0 ;
      RECT  1251600.0 1538400.0 1261800.0 1552200.0 ;
      RECT  1251600.0 1566000.0 1261800.0 1552200.0 ;
      RECT  1251600.0 1566000.0 1261800.0 1579800.0 ;
      RECT  1251600.0 1593600.0 1261800.0 1579800.0 ;
      RECT  1251600.0 1593600.0 1261800.0 1607400.0 ;
      RECT  1251600.0 1621200.0 1261800.0 1607400.0 ;
      RECT  1251600.0 1621200.0 1261800.0 1635000.0 ;
      RECT  1251600.0 1648800.0 1261800.0 1635000.0 ;
      RECT  1251600.0 1648800.0 1261800.0 1662600.0 ;
      RECT  1251600.0 1676400.0 1261800.0 1662600.0 ;
      RECT  1251600.0 1676400.0 1261800.0 1690200.0 ;
      RECT  1251600.0 1704000.0 1261800.0 1690200.0 ;
      RECT  1251600.0 1704000.0 1261800.0 1717800.0 ;
      RECT  1251600.0 1731600.0 1261800.0 1717800.0 ;
      RECT  1251600.0 1731600.0 1261800.0 1745400.0 ;
      RECT  1251600.0 1759200.0 1261800.0 1745400.0 ;
      RECT  1251600.0 1759200.0 1261800.0 1773000.0 ;
      RECT  1251600.0 1786800.0 1261800.0 1773000.0 ;
      RECT  1251600.0 1786800.0 1261800.0 1800600.0 ;
      RECT  1251600.0 1814400.0 1261800.0 1800600.0 ;
      RECT  1251600.0 1814400.0 1261800.0 1828200.0 ;
      RECT  1251600.0 1842000.0 1261800.0 1828200.0 ;
      RECT  1251600.0 1842000.0 1261800.0 1855800.0 ;
      RECT  1251600.0 1869600.0 1261800.0 1855800.0 ;
      RECT  1251600.0 1869600.0 1261800.0 1883400.0 ;
      RECT  1251600.0 1897200.0 1261800.0 1883400.0 ;
      RECT  1251600.0 1897200.0 1261800.0 1911000.0 ;
      RECT  1251600.0 1924800.0 1261800.0 1911000.0 ;
      RECT  1251600.0 1924800.0 1261800.0 1938600.0 ;
      RECT  1251600.0 1952400.0 1261800.0 1938600.0 ;
      RECT  1251600.0 1952400.0 1261800.0 1966200.0 ;
      RECT  1251600.0 1980000.0 1261800.0 1966200.0 ;
      RECT  1251600.0 1980000.0 1261800.0 1993800.0 ;
      RECT  1251600.0 2007600.0 1261800.0 1993800.0 ;
      RECT  1251600.0 2007600.0 1261800.0 2021400.0 ;
      RECT  1251600.0 2035200.0 1261800.0 2021400.0 ;
      RECT  1251600.0 2035200.0 1261800.0 2049000.0 ;
      RECT  1251600.0 2062800.0 1261800.0 2049000.0 ;
      RECT  1251600.0 2062800.0 1261800.0 2076600.0 ;
      RECT  1251600.0 2090400.0 1261800.0 2076600.0 ;
      RECT  1251600.0 2090400.0 1261800.0 2104200.0 ;
      RECT  1251600.0 2118000.0 1261800.0 2104200.0 ;
      RECT  1251600.0 2118000.0 1261800.0 2131800.0 ;
      RECT  1251600.0 2145600.0 1261800.0 2131800.0 ;
      RECT  1261800.0 379200.0 1272000.0 393000.0 ;
      RECT  1261800.0 406800.0 1272000.0 393000.0 ;
      RECT  1261800.0 406800.0 1272000.0 420600.0 ;
      RECT  1261800.0 434400.0 1272000.0 420600.0 ;
      RECT  1261800.0 434400.0 1272000.0 448200.0 ;
      RECT  1261800.0 462000.0 1272000.0 448200.0 ;
      RECT  1261800.0 462000.0 1272000.0 475800.0 ;
      RECT  1261800.0 489600.0 1272000.0 475800.0 ;
      RECT  1261800.0 489600.0 1272000.0 503400.0 ;
      RECT  1261800.0 517200.0 1272000.0 503400.0 ;
      RECT  1261800.0 517200.0 1272000.0 531000.0 ;
      RECT  1261800.0 544800.0 1272000.0 531000.0 ;
      RECT  1261800.0 544800.0 1272000.0 558600.0 ;
      RECT  1261800.0 572400.0 1272000.0 558600.0 ;
      RECT  1261800.0 572400.0 1272000.0 586200.0 ;
      RECT  1261800.0 600000.0 1272000.0 586200.0 ;
      RECT  1261800.0 600000.0 1272000.0 613800.0 ;
      RECT  1261800.0 627600.0 1272000.0 613800.0 ;
      RECT  1261800.0 627600.0 1272000.0 641400.0 ;
      RECT  1261800.0 655200.0 1272000.0 641400.0 ;
      RECT  1261800.0 655200.0 1272000.0 669000.0 ;
      RECT  1261800.0 682800.0 1272000.0 669000.0 ;
      RECT  1261800.0 682800.0 1272000.0 696600.0 ;
      RECT  1261800.0 710400.0 1272000.0 696600.0 ;
      RECT  1261800.0 710400.0 1272000.0 724200.0 ;
      RECT  1261800.0 738000.0 1272000.0 724200.0 ;
      RECT  1261800.0 738000.0 1272000.0 751800.0 ;
      RECT  1261800.0 765600.0 1272000.0 751800.0 ;
      RECT  1261800.0 765600.0 1272000.0 779400.0 ;
      RECT  1261800.0 793200.0 1272000.0 779400.0 ;
      RECT  1261800.0 793200.0 1272000.0 807000.0 ;
      RECT  1261800.0 820800.0 1272000.0 807000.0 ;
      RECT  1261800.0 820800.0 1272000.0 834600.0 ;
      RECT  1261800.0 848400.0 1272000.0 834600.0 ;
      RECT  1261800.0 848400.0 1272000.0 862200.0 ;
      RECT  1261800.0 876000.0 1272000.0 862200.0 ;
      RECT  1261800.0 876000.0 1272000.0 889800.0 ;
      RECT  1261800.0 903600.0 1272000.0 889800.0 ;
      RECT  1261800.0 903600.0 1272000.0 917400.0 ;
      RECT  1261800.0 931200.0 1272000.0 917400.0 ;
      RECT  1261800.0 931200.0 1272000.0 945000.0 ;
      RECT  1261800.0 958800.0 1272000.0 945000.0 ;
      RECT  1261800.0 958800.0 1272000.0 972600.0 ;
      RECT  1261800.0 986400.0 1272000.0 972600.0 ;
      RECT  1261800.0 986400.0 1272000.0 1000200.0 ;
      RECT  1261800.0 1014000.0 1272000.0 1000200.0 ;
      RECT  1261800.0 1014000.0 1272000.0 1027800.0 ;
      RECT  1261800.0 1041600.0 1272000.0 1027800.0 ;
      RECT  1261800.0 1041600.0 1272000.0 1055400.0 ;
      RECT  1261800.0 1069200.0 1272000.0 1055400.0 ;
      RECT  1261800.0 1069200.0 1272000.0 1083000.0 ;
      RECT  1261800.0 1096800.0 1272000.0 1083000.0 ;
      RECT  1261800.0 1096800.0 1272000.0 1110600.0 ;
      RECT  1261800.0 1124400.0 1272000.0 1110600.0 ;
      RECT  1261800.0 1124400.0 1272000.0 1138200.0 ;
      RECT  1261800.0 1152000.0 1272000.0 1138200.0 ;
      RECT  1261800.0 1152000.0 1272000.0 1165800.0 ;
      RECT  1261800.0 1179600.0 1272000.0 1165800.0 ;
      RECT  1261800.0 1179600.0 1272000.0 1193400.0 ;
      RECT  1261800.0 1207200.0 1272000.0 1193400.0 ;
      RECT  1261800.0 1207200.0 1272000.0 1221000.0 ;
      RECT  1261800.0 1234800.0 1272000.0 1221000.0 ;
      RECT  1261800.0 1234800.0 1272000.0 1248600.0 ;
      RECT  1261800.0 1262400.0 1272000.0 1248600.0 ;
      RECT  1261800.0 1262400.0 1272000.0 1276200.0 ;
      RECT  1261800.0 1290000.0 1272000.0 1276200.0 ;
      RECT  1261800.0 1290000.0 1272000.0 1303800.0 ;
      RECT  1261800.0 1317600.0 1272000.0 1303800.0 ;
      RECT  1261800.0 1317600.0 1272000.0 1331400.0 ;
      RECT  1261800.0 1345200.0 1272000.0 1331400.0 ;
      RECT  1261800.0 1345200.0 1272000.0 1359000.0 ;
      RECT  1261800.0 1372800.0 1272000.0 1359000.0 ;
      RECT  1261800.0 1372800.0 1272000.0 1386600.0 ;
      RECT  1261800.0 1400400.0 1272000.0 1386600.0 ;
      RECT  1261800.0 1400400.0 1272000.0 1414200.0 ;
      RECT  1261800.0 1428000.0 1272000.0 1414200.0 ;
      RECT  1261800.0 1428000.0 1272000.0 1441800.0 ;
      RECT  1261800.0 1455600.0 1272000.0 1441800.0 ;
      RECT  1261800.0 1455600.0 1272000.0 1469400.0 ;
      RECT  1261800.0 1483200.0 1272000.0 1469400.0 ;
      RECT  1261800.0 1483200.0 1272000.0 1497000.0 ;
      RECT  1261800.0 1510800.0 1272000.0 1497000.0 ;
      RECT  1261800.0 1510800.0 1272000.0 1524600.0 ;
      RECT  1261800.0 1538400.0 1272000.0 1524600.0 ;
      RECT  1261800.0 1538400.0 1272000.0 1552200.0 ;
      RECT  1261800.0 1566000.0 1272000.0 1552200.0 ;
      RECT  1261800.0 1566000.0 1272000.0 1579800.0 ;
      RECT  1261800.0 1593600.0 1272000.0 1579800.0 ;
      RECT  1261800.0 1593600.0 1272000.0 1607400.0 ;
      RECT  1261800.0 1621200.0 1272000.0 1607400.0 ;
      RECT  1261800.0 1621200.0 1272000.0 1635000.0 ;
      RECT  1261800.0 1648800.0 1272000.0 1635000.0 ;
      RECT  1261800.0 1648800.0 1272000.0 1662600.0 ;
      RECT  1261800.0 1676400.0 1272000.0 1662600.0 ;
      RECT  1261800.0 1676400.0 1272000.0 1690200.0 ;
      RECT  1261800.0 1704000.0 1272000.0 1690200.0 ;
      RECT  1261800.0 1704000.0 1272000.0 1717800.0 ;
      RECT  1261800.0 1731600.0 1272000.0 1717800.0 ;
      RECT  1261800.0 1731600.0 1272000.0 1745400.0 ;
      RECT  1261800.0 1759200.0 1272000.0 1745400.0 ;
      RECT  1261800.0 1759200.0 1272000.0 1773000.0 ;
      RECT  1261800.0 1786800.0 1272000.0 1773000.0 ;
      RECT  1261800.0 1786800.0 1272000.0 1800600.0 ;
      RECT  1261800.0 1814400.0 1272000.0 1800600.0 ;
      RECT  1261800.0 1814400.0 1272000.0 1828200.0 ;
      RECT  1261800.0 1842000.0 1272000.0 1828200.0 ;
      RECT  1261800.0 1842000.0 1272000.0 1855800.0 ;
      RECT  1261800.0 1869600.0 1272000.0 1855800.0 ;
      RECT  1261800.0 1869600.0 1272000.0 1883400.0 ;
      RECT  1261800.0 1897200.0 1272000.0 1883400.0 ;
      RECT  1261800.0 1897200.0 1272000.0 1911000.0 ;
      RECT  1261800.0 1924800.0 1272000.0 1911000.0 ;
      RECT  1261800.0 1924800.0 1272000.0 1938600.0 ;
      RECT  1261800.0 1952400.0 1272000.0 1938600.0 ;
      RECT  1261800.0 1952400.0 1272000.0 1966200.0 ;
      RECT  1261800.0 1980000.0 1272000.0 1966200.0 ;
      RECT  1261800.0 1980000.0 1272000.0 1993800.0 ;
      RECT  1261800.0 2007600.0 1272000.0 1993800.0 ;
      RECT  1261800.0 2007600.0 1272000.0 2021400.0 ;
      RECT  1261800.0 2035200.0 1272000.0 2021400.0 ;
      RECT  1261800.0 2035200.0 1272000.0 2049000.0 ;
      RECT  1261800.0 2062800.0 1272000.0 2049000.0 ;
      RECT  1261800.0 2062800.0 1272000.0 2076600.0 ;
      RECT  1261800.0 2090400.0 1272000.0 2076600.0 ;
      RECT  1261800.0 2090400.0 1272000.0 2104200.0 ;
      RECT  1261800.0 2118000.0 1272000.0 2104200.0 ;
      RECT  1261800.0 2118000.0 1272000.0 2131800.0 ;
      RECT  1261800.0 2145600.0 1272000.0 2131800.0 ;
      RECT  1272000.0 379200.0 1282200.0 393000.0 ;
      RECT  1272000.0 406800.0 1282200.0 393000.0 ;
      RECT  1272000.0 406800.0 1282200.0 420600.0 ;
      RECT  1272000.0 434400.0 1282200.0 420600.0 ;
      RECT  1272000.0 434400.0 1282200.0 448200.0 ;
      RECT  1272000.0 462000.0 1282200.0 448200.0 ;
      RECT  1272000.0 462000.0 1282200.0 475800.0 ;
      RECT  1272000.0 489600.0 1282200.0 475800.0 ;
      RECT  1272000.0 489600.0 1282200.0 503400.0 ;
      RECT  1272000.0 517200.0 1282200.0 503400.0 ;
      RECT  1272000.0 517200.0 1282200.0 531000.0 ;
      RECT  1272000.0 544800.0 1282200.0 531000.0 ;
      RECT  1272000.0 544800.0 1282200.0 558600.0 ;
      RECT  1272000.0 572400.0 1282200.0 558600.0 ;
      RECT  1272000.0 572400.0 1282200.0 586200.0 ;
      RECT  1272000.0 600000.0 1282200.0 586200.0 ;
      RECT  1272000.0 600000.0 1282200.0 613800.0 ;
      RECT  1272000.0 627600.0 1282200.0 613800.0 ;
      RECT  1272000.0 627600.0 1282200.0 641400.0 ;
      RECT  1272000.0 655200.0 1282200.0 641400.0 ;
      RECT  1272000.0 655200.0 1282200.0 669000.0 ;
      RECT  1272000.0 682800.0 1282200.0 669000.0 ;
      RECT  1272000.0 682800.0 1282200.0 696600.0 ;
      RECT  1272000.0 710400.0 1282200.0 696600.0 ;
      RECT  1272000.0 710400.0 1282200.0 724200.0 ;
      RECT  1272000.0 738000.0 1282200.0 724200.0 ;
      RECT  1272000.0 738000.0 1282200.0 751800.0 ;
      RECT  1272000.0 765600.0 1282200.0 751800.0 ;
      RECT  1272000.0 765600.0 1282200.0 779400.0 ;
      RECT  1272000.0 793200.0 1282200.0 779400.0 ;
      RECT  1272000.0 793200.0 1282200.0 807000.0 ;
      RECT  1272000.0 820800.0 1282200.0 807000.0 ;
      RECT  1272000.0 820800.0 1282200.0 834600.0 ;
      RECT  1272000.0 848400.0 1282200.0 834600.0 ;
      RECT  1272000.0 848400.0 1282200.0 862200.0 ;
      RECT  1272000.0 876000.0 1282200.0 862200.0 ;
      RECT  1272000.0 876000.0 1282200.0 889800.0 ;
      RECT  1272000.0 903600.0 1282200.0 889800.0 ;
      RECT  1272000.0 903600.0 1282200.0 917400.0 ;
      RECT  1272000.0 931200.0 1282200.0 917400.0 ;
      RECT  1272000.0 931200.0 1282200.0 945000.0 ;
      RECT  1272000.0 958800.0 1282200.0 945000.0 ;
      RECT  1272000.0 958800.0 1282200.0 972600.0 ;
      RECT  1272000.0 986400.0 1282200.0 972600.0 ;
      RECT  1272000.0 986400.0 1282200.0 1000200.0 ;
      RECT  1272000.0 1014000.0 1282200.0 1000200.0 ;
      RECT  1272000.0 1014000.0 1282200.0 1027800.0 ;
      RECT  1272000.0 1041600.0 1282200.0 1027800.0 ;
      RECT  1272000.0 1041600.0 1282200.0 1055400.0 ;
      RECT  1272000.0 1069200.0 1282200.0 1055400.0 ;
      RECT  1272000.0 1069200.0 1282200.0 1083000.0 ;
      RECT  1272000.0 1096800.0 1282200.0 1083000.0 ;
      RECT  1272000.0 1096800.0 1282200.0 1110600.0 ;
      RECT  1272000.0 1124400.0 1282200.0 1110600.0 ;
      RECT  1272000.0 1124400.0 1282200.0 1138200.0 ;
      RECT  1272000.0 1152000.0 1282200.0 1138200.0 ;
      RECT  1272000.0 1152000.0 1282200.0 1165800.0 ;
      RECT  1272000.0 1179600.0 1282200.0 1165800.0 ;
      RECT  1272000.0 1179600.0 1282200.0 1193400.0 ;
      RECT  1272000.0 1207200.0 1282200.0 1193400.0 ;
      RECT  1272000.0 1207200.0 1282200.0 1221000.0 ;
      RECT  1272000.0 1234800.0 1282200.0 1221000.0 ;
      RECT  1272000.0 1234800.0 1282200.0 1248600.0 ;
      RECT  1272000.0 1262400.0 1282200.0 1248600.0 ;
      RECT  1272000.0 1262400.0 1282200.0 1276200.0 ;
      RECT  1272000.0 1290000.0 1282200.0 1276200.0 ;
      RECT  1272000.0 1290000.0 1282200.0 1303800.0 ;
      RECT  1272000.0 1317600.0 1282200.0 1303800.0 ;
      RECT  1272000.0 1317600.0 1282200.0 1331400.0 ;
      RECT  1272000.0 1345200.0 1282200.0 1331400.0 ;
      RECT  1272000.0 1345200.0 1282200.0 1359000.0 ;
      RECT  1272000.0 1372800.0 1282200.0 1359000.0 ;
      RECT  1272000.0 1372800.0 1282200.0 1386600.0 ;
      RECT  1272000.0 1400400.0 1282200.0 1386600.0 ;
      RECT  1272000.0 1400400.0 1282200.0 1414200.0 ;
      RECT  1272000.0 1428000.0 1282200.0 1414200.0 ;
      RECT  1272000.0 1428000.0 1282200.0 1441800.0 ;
      RECT  1272000.0 1455600.0 1282200.0 1441800.0 ;
      RECT  1272000.0 1455600.0 1282200.0 1469400.0 ;
      RECT  1272000.0 1483200.0 1282200.0 1469400.0 ;
      RECT  1272000.0 1483200.0 1282200.0 1497000.0 ;
      RECT  1272000.0 1510800.0 1282200.0 1497000.0 ;
      RECT  1272000.0 1510800.0 1282200.0 1524600.0 ;
      RECT  1272000.0 1538400.0 1282200.0 1524600.0 ;
      RECT  1272000.0 1538400.0 1282200.0 1552200.0 ;
      RECT  1272000.0 1566000.0 1282200.0 1552200.0 ;
      RECT  1272000.0 1566000.0 1282200.0 1579800.0 ;
      RECT  1272000.0 1593600.0 1282200.0 1579800.0 ;
      RECT  1272000.0 1593600.0 1282200.0 1607400.0 ;
      RECT  1272000.0 1621200.0 1282200.0 1607400.0 ;
      RECT  1272000.0 1621200.0 1282200.0 1635000.0 ;
      RECT  1272000.0 1648800.0 1282200.0 1635000.0 ;
      RECT  1272000.0 1648800.0 1282200.0 1662600.0 ;
      RECT  1272000.0 1676400.0 1282200.0 1662600.0 ;
      RECT  1272000.0 1676400.0 1282200.0 1690200.0 ;
      RECT  1272000.0 1704000.0 1282200.0 1690200.0 ;
      RECT  1272000.0 1704000.0 1282200.0 1717800.0 ;
      RECT  1272000.0 1731600.0 1282200.0 1717800.0 ;
      RECT  1272000.0 1731600.0 1282200.0 1745400.0 ;
      RECT  1272000.0 1759200.0 1282200.0 1745400.0 ;
      RECT  1272000.0 1759200.0 1282200.0 1773000.0 ;
      RECT  1272000.0 1786800.0 1282200.0 1773000.0 ;
      RECT  1272000.0 1786800.0 1282200.0 1800600.0 ;
      RECT  1272000.0 1814400.0 1282200.0 1800600.0 ;
      RECT  1272000.0 1814400.0 1282200.0 1828200.0 ;
      RECT  1272000.0 1842000.0 1282200.0 1828200.0 ;
      RECT  1272000.0 1842000.0 1282200.0 1855800.0 ;
      RECT  1272000.0 1869600.0 1282200.0 1855800.0 ;
      RECT  1272000.0 1869600.0 1282200.0 1883400.0 ;
      RECT  1272000.0 1897200.0 1282200.0 1883400.0 ;
      RECT  1272000.0 1897200.0 1282200.0 1911000.0 ;
      RECT  1272000.0 1924800.0 1282200.0 1911000.0 ;
      RECT  1272000.0 1924800.0 1282200.0 1938600.0 ;
      RECT  1272000.0 1952400.0 1282200.0 1938600.0 ;
      RECT  1272000.0 1952400.0 1282200.0 1966200.0 ;
      RECT  1272000.0 1980000.0 1282200.0 1966200.0 ;
      RECT  1272000.0 1980000.0 1282200.0 1993800.0 ;
      RECT  1272000.0 2007600.0 1282200.0 1993800.0 ;
      RECT  1272000.0 2007600.0 1282200.0 2021400.0 ;
      RECT  1272000.0 2035200.0 1282200.0 2021400.0 ;
      RECT  1272000.0 2035200.0 1282200.0 2049000.0 ;
      RECT  1272000.0 2062800.0 1282200.0 2049000.0 ;
      RECT  1272000.0 2062800.0 1282200.0 2076600.0 ;
      RECT  1272000.0 2090400.0 1282200.0 2076600.0 ;
      RECT  1272000.0 2090400.0 1282200.0 2104200.0 ;
      RECT  1272000.0 2118000.0 1282200.0 2104200.0 ;
      RECT  1272000.0 2118000.0 1282200.0 2131800.0 ;
      RECT  1272000.0 2145600.0 1282200.0 2131800.0 ;
      RECT  1282200.0 379200.0 1292400.0 393000.0 ;
      RECT  1282200.0 406800.0 1292400.0 393000.0 ;
      RECT  1282200.0 406800.0 1292400.0 420600.0 ;
      RECT  1282200.0 434400.0 1292400.0 420600.0 ;
      RECT  1282200.0 434400.0 1292400.0 448200.0 ;
      RECT  1282200.0 462000.0 1292400.0 448200.0 ;
      RECT  1282200.0 462000.0 1292400.0 475800.0 ;
      RECT  1282200.0 489600.0 1292400.0 475800.0 ;
      RECT  1282200.0 489600.0 1292400.0 503400.0 ;
      RECT  1282200.0 517200.0 1292400.0 503400.0 ;
      RECT  1282200.0 517200.0 1292400.0 531000.0 ;
      RECT  1282200.0 544800.0 1292400.0 531000.0 ;
      RECT  1282200.0 544800.0 1292400.0 558600.0 ;
      RECT  1282200.0 572400.0 1292400.0 558600.0 ;
      RECT  1282200.0 572400.0 1292400.0 586200.0 ;
      RECT  1282200.0 600000.0 1292400.0 586200.0 ;
      RECT  1282200.0 600000.0 1292400.0 613800.0 ;
      RECT  1282200.0 627600.0 1292400.0 613800.0 ;
      RECT  1282200.0 627600.0 1292400.0 641400.0 ;
      RECT  1282200.0 655200.0 1292400.0 641400.0 ;
      RECT  1282200.0 655200.0 1292400.0 669000.0 ;
      RECT  1282200.0 682800.0 1292400.0 669000.0 ;
      RECT  1282200.0 682800.0 1292400.0 696600.0 ;
      RECT  1282200.0 710400.0 1292400.0 696600.0 ;
      RECT  1282200.0 710400.0 1292400.0 724200.0 ;
      RECT  1282200.0 738000.0 1292400.0 724200.0 ;
      RECT  1282200.0 738000.0 1292400.0 751800.0 ;
      RECT  1282200.0 765600.0 1292400.0 751800.0 ;
      RECT  1282200.0 765600.0 1292400.0 779400.0 ;
      RECT  1282200.0 793200.0 1292400.0 779400.0 ;
      RECT  1282200.0 793200.0 1292400.0 807000.0 ;
      RECT  1282200.0 820800.0 1292400.0 807000.0 ;
      RECT  1282200.0 820800.0 1292400.0 834600.0 ;
      RECT  1282200.0 848400.0 1292400.0 834600.0 ;
      RECT  1282200.0 848400.0 1292400.0 862200.0 ;
      RECT  1282200.0 876000.0 1292400.0 862200.0 ;
      RECT  1282200.0 876000.0 1292400.0 889800.0 ;
      RECT  1282200.0 903600.0 1292400.0 889800.0 ;
      RECT  1282200.0 903600.0 1292400.0 917400.0 ;
      RECT  1282200.0 931200.0 1292400.0 917400.0 ;
      RECT  1282200.0 931200.0 1292400.0 945000.0 ;
      RECT  1282200.0 958800.0 1292400.0 945000.0 ;
      RECT  1282200.0 958800.0 1292400.0 972600.0 ;
      RECT  1282200.0 986400.0 1292400.0 972600.0 ;
      RECT  1282200.0 986400.0 1292400.0 1000200.0 ;
      RECT  1282200.0 1014000.0 1292400.0 1000200.0 ;
      RECT  1282200.0 1014000.0 1292400.0 1027800.0 ;
      RECT  1282200.0 1041600.0 1292400.0 1027800.0 ;
      RECT  1282200.0 1041600.0 1292400.0 1055400.0 ;
      RECT  1282200.0 1069200.0 1292400.0 1055400.0 ;
      RECT  1282200.0 1069200.0 1292400.0 1083000.0 ;
      RECT  1282200.0 1096800.0 1292400.0 1083000.0 ;
      RECT  1282200.0 1096800.0 1292400.0 1110600.0 ;
      RECT  1282200.0 1124400.0 1292400.0 1110600.0 ;
      RECT  1282200.0 1124400.0 1292400.0 1138200.0 ;
      RECT  1282200.0 1152000.0 1292400.0 1138200.0 ;
      RECT  1282200.0 1152000.0 1292400.0 1165800.0 ;
      RECT  1282200.0 1179600.0 1292400.0 1165800.0 ;
      RECT  1282200.0 1179600.0 1292400.0 1193400.0 ;
      RECT  1282200.0 1207200.0 1292400.0 1193400.0 ;
      RECT  1282200.0 1207200.0 1292400.0 1221000.0 ;
      RECT  1282200.0 1234800.0 1292400.0 1221000.0 ;
      RECT  1282200.0 1234800.0 1292400.0 1248600.0 ;
      RECT  1282200.0 1262400.0 1292400.0 1248600.0 ;
      RECT  1282200.0 1262400.0 1292400.0 1276200.0 ;
      RECT  1282200.0 1290000.0 1292400.0 1276200.0 ;
      RECT  1282200.0 1290000.0 1292400.0 1303800.0 ;
      RECT  1282200.0 1317600.0 1292400.0 1303800.0 ;
      RECT  1282200.0 1317600.0 1292400.0 1331400.0 ;
      RECT  1282200.0 1345200.0 1292400.0 1331400.0 ;
      RECT  1282200.0 1345200.0 1292400.0 1359000.0 ;
      RECT  1282200.0 1372800.0 1292400.0 1359000.0 ;
      RECT  1282200.0 1372800.0 1292400.0 1386600.0 ;
      RECT  1282200.0 1400400.0 1292400.0 1386600.0 ;
      RECT  1282200.0 1400400.0 1292400.0 1414200.0 ;
      RECT  1282200.0 1428000.0 1292400.0 1414200.0 ;
      RECT  1282200.0 1428000.0 1292400.0 1441800.0 ;
      RECT  1282200.0 1455600.0 1292400.0 1441800.0 ;
      RECT  1282200.0 1455600.0 1292400.0 1469400.0 ;
      RECT  1282200.0 1483200.0 1292400.0 1469400.0 ;
      RECT  1282200.0 1483200.0 1292400.0 1497000.0 ;
      RECT  1282200.0 1510800.0 1292400.0 1497000.0 ;
      RECT  1282200.0 1510800.0 1292400.0 1524600.0 ;
      RECT  1282200.0 1538400.0 1292400.0 1524600.0 ;
      RECT  1282200.0 1538400.0 1292400.0 1552200.0 ;
      RECT  1282200.0 1566000.0 1292400.0 1552200.0 ;
      RECT  1282200.0 1566000.0 1292400.0 1579800.0 ;
      RECT  1282200.0 1593600.0 1292400.0 1579800.0 ;
      RECT  1282200.0 1593600.0 1292400.0 1607400.0 ;
      RECT  1282200.0 1621200.0 1292400.0 1607400.0 ;
      RECT  1282200.0 1621200.0 1292400.0 1635000.0 ;
      RECT  1282200.0 1648800.0 1292400.0 1635000.0 ;
      RECT  1282200.0 1648800.0 1292400.0 1662600.0 ;
      RECT  1282200.0 1676400.0 1292400.0 1662600.0 ;
      RECT  1282200.0 1676400.0 1292400.0 1690200.0 ;
      RECT  1282200.0 1704000.0 1292400.0 1690200.0 ;
      RECT  1282200.0 1704000.0 1292400.0 1717800.0 ;
      RECT  1282200.0 1731600.0 1292400.0 1717800.0 ;
      RECT  1282200.0 1731600.0 1292400.0 1745400.0 ;
      RECT  1282200.0 1759200.0 1292400.0 1745400.0 ;
      RECT  1282200.0 1759200.0 1292400.0 1773000.0 ;
      RECT  1282200.0 1786800.0 1292400.0 1773000.0 ;
      RECT  1282200.0 1786800.0 1292400.0 1800600.0 ;
      RECT  1282200.0 1814400.0 1292400.0 1800600.0 ;
      RECT  1282200.0 1814400.0 1292400.0 1828200.0 ;
      RECT  1282200.0 1842000.0 1292400.0 1828200.0 ;
      RECT  1282200.0 1842000.0 1292400.0 1855800.0 ;
      RECT  1282200.0 1869600.0 1292400.0 1855800.0 ;
      RECT  1282200.0 1869600.0 1292400.0 1883400.0 ;
      RECT  1282200.0 1897200.0 1292400.0 1883400.0 ;
      RECT  1282200.0 1897200.0 1292400.0 1911000.0 ;
      RECT  1282200.0 1924800.0 1292400.0 1911000.0 ;
      RECT  1282200.0 1924800.0 1292400.0 1938600.0 ;
      RECT  1282200.0 1952400.0 1292400.0 1938600.0 ;
      RECT  1282200.0 1952400.0 1292400.0 1966200.0 ;
      RECT  1282200.0 1980000.0 1292400.0 1966200.0 ;
      RECT  1282200.0 1980000.0 1292400.0 1993800.0 ;
      RECT  1282200.0 2007600.0 1292400.0 1993800.0 ;
      RECT  1282200.0 2007600.0 1292400.0 2021400.0 ;
      RECT  1282200.0 2035200.0 1292400.0 2021400.0 ;
      RECT  1282200.0 2035200.0 1292400.0 2049000.0 ;
      RECT  1282200.0 2062800.0 1292400.0 2049000.0 ;
      RECT  1282200.0 2062800.0 1292400.0 2076600.0 ;
      RECT  1282200.0 2090400.0 1292400.0 2076600.0 ;
      RECT  1282200.0 2090400.0 1292400.0 2104200.0 ;
      RECT  1282200.0 2118000.0 1292400.0 2104200.0 ;
      RECT  1282200.0 2118000.0 1292400.0 2131800.0 ;
      RECT  1282200.0 2145600.0 1292400.0 2131800.0 ;
      RECT  1292400.0 379200.0 1302600.0 393000.0 ;
      RECT  1292400.0 406800.0 1302600.0 393000.0 ;
      RECT  1292400.0 406800.0 1302600.0 420600.0 ;
      RECT  1292400.0 434400.0 1302600.0 420600.0 ;
      RECT  1292400.0 434400.0 1302600.0 448200.0 ;
      RECT  1292400.0 462000.0 1302600.0 448200.0 ;
      RECT  1292400.0 462000.0 1302600.0 475800.0 ;
      RECT  1292400.0 489600.0 1302600.0 475800.0 ;
      RECT  1292400.0 489600.0 1302600.0 503400.0 ;
      RECT  1292400.0 517200.0 1302600.0 503400.0 ;
      RECT  1292400.0 517200.0 1302600.0 531000.0 ;
      RECT  1292400.0 544800.0 1302600.0 531000.0 ;
      RECT  1292400.0 544800.0 1302600.0 558600.0 ;
      RECT  1292400.0 572400.0 1302600.0 558600.0 ;
      RECT  1292400.0 572400.0 1302600.0 586200.0 ;
      RECT  1292400.0 600000.0 1302600.0 586200.0 ;
      RECT  1292400.0 600000.0 1302600.0 613800.0 ;
      RECT  1292400.0 627600.0 1302600.0 613800.0 ;
      RECT  1292400.0 627600.0 1302600.0 641400.0 ;
      RECT  1292400.0 655200.0 1302600.0 641400.0 ;
      RECT  1292400.0 655200.0 1302600.0 669000.0 ;
      RECT  1292400.0 682800.0 1302600.0 669000.0 ;
      RECT  1292400.0 682800.0 1302600.0 696600.0 ;
      RECT  1292400.0 710400.0 1302600.0 696600.0 ;
      RECT  1292400.0 710400.0 1302600.0 724200.0 ;
      RECT  1292400.0 738000.0 1302600.0 724200.0 ;
      RECT  1292400.0 738000.0 1302600.0 751800.0 ;
      RECT  1292400.0 765600.0 1302600.0 751800.0 ;
      RECT  1292400.0 765600.0 1302600.0 779400.0 ;
      RECT  1292400.0 793200.0 1302600.0 779400.0 ;
      RECT  1292400.0 793200.0 1302600.0 807000.0 ;
      RECT  1292400.0 820800.0 1302600.0 807000.0 ;
      RECT  1292400.0 820800.0 1302600.0 834600.0 ;
      RECT  1292400.0 848400.0 1302600.0 834600.0 ;
      RECT  1292400.0 848400.0 1302600.0 862200.0 ;
      RECT  1292400.0 876000.0 1302600.0 862200.0 ;
      RECT  1292400.0 876000.0 1302600.0 889800.0 ;
      RECT  1292400.0 903600.0 1302600.0 889800.0 ;
      RECT  1292400.0 903600.0 1302600.0 917400.0 ;
      RECT  1292400.0 931200.0 1302600.0 917400.0 ;
      RECT  1292400.0 931200.0 1302600.0 945000.0 ;
      RECT  1292400.0 958800.0 1302600.0 945000.0 ;
      RECT  1292400.0 958800.0 1302600.0 972600.0 ;
      RECT  1292400.0 986400.0 1302600.0 972600.0 ;
      RECT  1292400.0 986400.0 1302600.0 1000200.0 ;
      RECT  1292400.0 1014000.0 1302600.0 1000200.0 ;
      RECT  1292400.0 1014000.0 1302600.0 1027800.0 ;
      RECT  1292400.0 1041600.0 1302600.0 1027800.0 ;
      RECT  1292400.0 1041600.0 1302600.0 1055400.0 ;
      RECT  1292400.0 1069200.0 1302600.0 1055400.0 ;
      RECT  1292400.0 1069200.0 1302600.0 1083000.0 ;
      RECT  1292400.0 1096800.0 1302600.0 1083000.0 ;
      RECT  1292400.0 1096800.0 1302600.0 1110600.0 ;
      RECT  1292400.0 1124400.0 1302600.0 1110600.0 ;
      RECT  1292400.0 1124400.0 1302600.0 1138200.0 ;
      RECT  1292400.0 1152000.0 1302600.0 1138200.0 ;
      RECT  1292400.0 1152000.0 1302600.0 1165800.0 ;
      RECT  1292400.0 1179600.0 1302600.0 1165800.0 ;
      RECT  1292400.0 1179600.0 1302600.0 1193400.0 ;
      RECT  1292400.0 1207200.0 1302600.0 1193400.0 ;
      RECT  1292400.0 1207200.0 1302600.0 1221000.0 ;
      RECT  1292400.0 1234800.0 1302600.0 1221000.0 ;
      RECT  1292400.0 1234800.0 1302600.0 1248600.0 ;
      RECT  1292400.0 1262400.0 1302600.0 1248600.0 ;
      RECT  1292400.0 1262400.0 1302600.0 1276200.0 ;
      RECT  1292400.0 1290000.0 1302600.0 1276200.0 ;
      RECT  1292400.0 1290000.0 1302600.0 1303800.0 ;
      RECT  1292400.0 1317600.0 1302600.0 1303800.0 ;
      RECT  1292400.0 1317600.0 1302600.0 1331400.0 ;
      RECT  1292400.0 1345200.0 1302600.0 1331400.0 ;
      RECT  1292400.0 1345200.0 1302600.0 1359000.0 ;
      RECT  1292400.0 1372800.0 1302600.0 1359000.0 ;
      RECT  1292400.0 1372800.0 1302600.0 1386600.0 ;
      RECT  1292400.0 1400400.0 1302600.0 1386600.0 ;
      RECT  1292400.0 1400400.0 1302600.0 1414200.0 ;
      RECT  1292400.0 1428000.0 1302600.0 1414200.0 ;
      RECT  1292400.0 1428000.0 1302600.0 1441800.0 ;
      RECT  1292400.0 1455600.0 1302600.0 1441800.0 ;
      RECT  1292400.0 1455600.0 1302600.0 1469400.0 ;
      RECT  1292400.0 1483200.0 1302600.0 1469400.0 ;
      RECT  1292400.0 1483200.0 1302600.0 1497000.0 ;
      RECT  1292400.0 1510800.0 1302600.0 1497000.0 ;
      RECT  1292400.0 1510800.0 1302600.0 1524600.0 ;
      RECT  1292400.0 1538400.0 1302600.0 1524600.0 ;
      RECT  1292400.0 1538400.0 1302600.0 1552200.0 ;
      RECT  1292400.0 1566000.0 1302600.0 1552200.0 ;
      RECT  1292400.0 1566000.0 1302600.0 1579800.0 ;
      RECT  1292400.0 1593600.0 1302600.0 1579800.0 ;
      RECT  1292400.0 1593600.0 1302600.0 1607400.0 ;
      RECT  1292400.0 1621200.0 1302600.0 1607400.0 ;
      RECT  1292400.0 1621200.0 1302600.0 1635000.0 ;
      RECT  1292400.0 1648800.0 1302600.0 1635000.0 ;
      RECT  1292400.0 1648800.0 1302600.0 1662600.0 ;
      RECT  1292400.0 1676400.0 1302600.0 1662600.0 ;
      RECT  1292400.0 1676400.0 1302600.0 1690200.0 ;
      RECT  1292400.0 1704000.0 1302600.0 1690200.0 ;
      RECT  1292400.0 1704000.0 1302600.0 1717800.0 ;
      RECT  1292400.0 1731600.0 1302600.0 1717800.0 ;
      RECT  1292400.0 1731600.0 1302600.0 1745400.0 ;
      RECT  1292400.0 1759200.0 1302600.0 1745400.0 ;
      RECT  1292400.0 1759200.0 1302600.0 1773000.0 ;
      RECT  1292400.0 1786800.0 1302600.0 1773000.0 ;
      RECT  1292400.0 1786800.0 1302600.0 1800600.0 ;
      RECT  1292400.0 1814400.0 1302600.0 1800600.0 ;
      RECT  1292400.0 1814400.0 1302600.0 1828200.0 ;
      RECT  1292400.0 1842000.0 1302600.0 1828200.0 ;
      RECT  1292400.0 1842000.0 1302600.0 1855800.0 ;
      RECT  1292400.0 1869600.0 1302600.0 1855800.0 ;
      RECT  1292400.0 1869600.0 1302600.0 1883400.0 ;
      RECT  1292400.0 1897200.0 1302600.0 1883400.0 ;
      RECT  1292400.0 1897200.0 1302600.0 1911000.0 ;
      RECT  1292400.0 1924800.0 1302600.0 1911000.0 ;
      RECT  1292400.0 1924800.0 1302600.0 1938600.0 ;
      RECT  1292400.0 1952400.0 1302600.0 1938600.0 ;
      RECT  1292400.0 1952400.0 1302600.0 1966200.0 ;
      RECT  1292400.0 1980000.0 1302600.0 1966200.0 ;
      RECT  1292400.0 1980000.0 1302600.0 1993800.0 ;
      RECT  1292400.0 2007600.0 1302600.0 1993800.0 ;
      RECT  1292400.0 2007600.0 1302600.0 2021400.0 ;
      RECT  1292400.0 2035200.0 1302600.0 2021400.0 ;
      RECT  1292400.0 2035200.0 1302600.0 2049000.0 ;
      RECT  1292400.0 2062800.0 1302600.0 2049000.0 ;
      RECT  1292400.0 2062800.0 1302600.0 2076600.0 ;
      RECT  1292400.0 2090400.0 1302600.0 2076600.0 ;
      RECT  1292400.0 2090400.0 1302600.0 2104200.0 ;
      RECT  1292400.0 2118000.0 1302600.0 2104200.0 ;
      RECT  1292400.0 2118000.0 1302600.0 2131800.0 ;
      RECT  1292400.0 2145600.0 1302600.0 2131800.0 ;
      RECT  1302600.0 379200.0 1312800.0 393000.0 ;
      RECT  1302600.0 406800.0 1312800.0 393000.0 ;
      RECT  1302600.0 406800.0 1312800.0 420600.0 ;
      RECT  1302600.0 434400.0 1312800.0 420600.0 ;
      RECT  1302600.0 434400.0 1312800.0 448200.0 ;
      RECT  1302600.0 462000.0 1312800.0 448200.0 ;
      RECT  1302600.0 462000.0 1312800.0 475800.0 ;
      RECT  1302600.0 489600.0 1312800.0 475800.0 ;
      RECT  1302600.0 489600.0 1312800.0 503400.0 ;
      RECT  1302600.0 517200.0 1312800.0 503400.0 ;
      RECT  1302600.0 517200.0 1312800.0 531000.0 ;
      RECT  1302600.0 544800.0 1312800.0 531000.0 ;
      RECT  1302600.0 544800.0 1312800.0 558600.0 ;
      RECT  1302600.0 572400.0 1312800.0 558600.0 ;
      RECT  1302600.0 572400.0 1312800.0 586200.0 ;
      RECT  1302600.0 600000.0 1312800.0 586200.0 ;
      RECT  1302600.0 600000.0 1312800.0 613800.0 ;
      RECT  1302600.0 627600.0 1312800.0 613800.0 ;
      RECT  1302600.0 627600.0 1312800.0 641400.0 ;
      RECT  1302600.0 655200.0 1312800.0 641400.0 ;
      RECT  1302600.0 655200.0 1312800.0 669000.0 ;
      RECT  1302600.0 682800.0 1312800.0 669000.0 ;
      RECT  1302600.0 682800.0 1312800.0 696600.0 ;
      RECT  1302600.0 710400.0 1312800.0 696600.0 ;
      RECT  1302600.0 710400.0 1312800.0 724200.0 ;
      RECT  1302600.0 738000.0 1312800.0 724200.0 ;
      RECT  1302600.0 738000.0 1312800.0 751800.0 ;
      RECT  1302600.0 765600.0 1312800.0 751800.0 ;
      RECT  1302600.0 765600.0 1312800.0 779400.0 ;
      RECT  1302600.0 793200.0 1312800.0 779400.0 ;
      RECT  1302600.0 793200.0 1312800.0 807000.0 ;
      RECT  1302600.0 820800.0 1312800.0 807000.0 ;
      RECT  1302600.0 820800.0 1312800.0 834600.0 ;
      RECT  1302600.0 848400.0 1312800.0 834600.0 ;
      RECT  1302600.0 848400.0 1312800.0 862200.0 ;
      RECT  1302600.0 876000.0 1312800.0 862200.0 ;
      RECT  1302600.0 876000.0 1312800.0 889800.0 ;
      RECT  1302600.0 903600.0 1312800.0 889800.0 ;
      RECT  1302600.0 903600.0 1312800.0 917400.0 ;
      RECT  1302600.0 931200.0 1312800.0 917400.0 ;
      RECT  1302600.0 931200.0 1312800.0 945000.0 ;
      RECT  1302600.0 958800.0 1312800.0 945000.0 ;
      RECT  1302600.0 958800.0 1312800.0 972600.0 ;
      RECT  1302600.0 986400.0 1312800.0 972600.0 ;
      RECT  1302600.0 986400.0 1312800.0 1000200.0 ;
      RECT  1302600.0 1014000.0 1312800.0 1000200.0 ;
      RECT  1302600.0 1014000.0 1312800.0 1027800.0 ;
      RECT  1302600.0 1041600.0 1312800.0 1027800.0 ;
      RECT  1302600.0 1041600.0 1312800.0 1055400.0 ;
      RECT  1302600.0 1069200.0 1312800.0 1055400.0 ;
      RECT  1302600.0 1069200.0 1312800.0 1083000.0 ;
      RECT  1302600.0 1096800.0 1312800.0 1083000.0 ;
      RECT  1302600.0 1096800.0 1312800.0 1110600.0 ;
      RECT  1302600.0 1124400.0 1312800.0 1110600.0 ;
      RECT  1302600.0 1124400.0 1312800.0 1138200.0 ;
      RECT  1302600.0 1152000.0 1312800.0 1138200.0 ;
      RECT  1302600.0 1152000.0 1312800.0 1165800.0 ;
      RECT  1302600.0 1179600.0 1312800.0 1165800.0 ;
      RECT  1302600.0 1179600.0 1312800.0 1193400.0 ;
      RECT  1302600.0 1207200.0 1312800.0 1193400.0 ;
      RECT  1302600.0 1207200.0 1312800.0 1221000.0 ;
      RECT  1302600.0 1234800.0 1312800.0 1221000.0 ;
      RECT  1302600.0 1234800.0 1312800.0 1248600.0 ;
      RECT  1302600.0 1262400.0 1312800.0 1248600.0 ;
      RECT  1302600.0 1262400.0 1312800.0 1276200.0 ;
      RECT  1302600.0 1290000.0 1312800.0 1276200.0 ;
      RECT  1302600.0 1290000.0 1312800.0 1303800.0 ;
      RECT  1302600.0 1317600.0 1312800.0 1303800.0 ;
      RECT  1302600.0 1317600.0 1312800.0 1331400.0 ;
      RECT  1302600.0 1345200.0 1312800.0 1331400.0 ;
      RECT  1302600.0 1345200.0 1312800.0 1359000.0 ;
      RECT  1302600.0 1372800.0 1312800.0 1359000.0 ;
      RECT  1302600.0 1372800.0 1312800.0 1386600.0 ;
      RECT  1302600.0 1400400.0 1312800.0 1386600.0 ;
      RECT  1302600.0 1400400.0 1312800.0 1414200.0 ;
      RECT  1302600.0 1428000.0 1312800.0 1414200.0 ;
      RECT  1302600.0 1428000.0 1312800.0 1441800.0 ;
      RECT  1302600.0 1455600.0 1312800.0 1441800.0 ;
      RECT  1302600.0 1455600.0 1312800.0 1469400.0 ;
      RECT  1302600.0 1483200.0 1312800.0 1469400.0 ;
      RECT  1302600.0 1483200.0 1312800.0 1497000.0 ;
      RECT  1302600.0 1510800.0 1312800.0 1497000.0 ;
      RECT  1302600.0 1510800.0 1312800.0 1524600.0 ;
      RECT  1302600.0 1538400.0 1312800.0 1524600.0 ;
      RECT  1302600.0 1538400.0 1312800.0 1552200.0 ;
      RECT  1302600.0 1566000.0 1312800.0 1552200.0 ;
      RECT  1302600.0 1566000.0 1312800.0 1579800.0 ;
      RECT  1302600.0 1593600.0 1312800.0 1579800.0 ;
      RECT  1302600.0 1593600.0 1312800.0 1607400.0 ;
      RECT  1302600.0 1621200.0 1312800.0 1607400.0 ;
      RECT  1302600.0 1621200.0 1312800.0 1635000.0 ;
      RECT  1302600.0 1648800.0 1312800.0 1635000.0 ;
      RECT  1302600.0 1648800.0 1312800.0 1662600.0 ;
      RECT  1302600.0 1676400.0 1312800.0 1662600.0 ;
      RECT  1302600.0 1676400.0 1312800.0 1690200.0 ;
      RECT  1302600.0 1704000.0 1312800.0 1690200.0 ;
      RECT  1302600.0 1704000.0 1312800.0 1717800.0 ;
      RECT  1302600.0 1731600.0 1312800.0 1717800.0 ;
      RECT  1302600.0 1731600.0 1312800.0 1745400.0 ;
      RECT  1302600.0 1759200.0 1312800.0 1745400.0 ;
      RECT  1302600.0 1759200.0 1312800.0 1773000.0 ;
      RECT  1302600.0 1786800.0 1312800.0 1773000.0 ;
      RECT  1302600.0 1786800.0 1312800.0 1800600.0 ;
      RECT  1302600.0 1814400.0 1312800.0 1800600.0 ;
      RECT  1302600.0 1814400.0 1312800.0 1828200.0 ;
      RECT  1302600.0 1842000.0 1312800.0 1828200.0 ;
      RECT  1302600.0 1842000.0 1312800.0 1855800.0 ;
      RECT  1302600.0 1869600.0 1312800.0 1855800.0 ;
      RECT  1302600.0 1869600.0 1312800.0 1883400.0 ;
      RECT  1302600.0 1897200.0 1312800.0 1883400.0 ;
      RECT  1302600.0 1897200.0 1312800.0 1911000.0 ;
      RECT  1302600.0 1924800.0 1312800.0 1911000.0 ;
      RECT  1302600.0 1924800.0 1312800.0 1938600.0 ;
      RECT  1302600.0 1952400.0 1312800.0 1938600.0 ;
      RECT  1302600.0 1952400.0 1312800.0 1966200.0 ;
      RECT  1302600.0 1980000.0 1312800.0 1966200.0 ;
      RECT  1302600.0 1980000.0 1312800.0 1993800.0 ;
      RECT  1302600.0 2007600.0 1312800.0 1993800.0 ;
      RECT  1302600.0 2007600.0 1312800.0 2021400.0 ;
      RECT  1302600.0 2035200.0 1312800.0 2021400.0 ;
      RECT  1302600.0 2035200.0 1312800.0 2049000.0 ;
      RECT  1302600.0 2062800.0 1312800.0 2049000.0 ;
      RECT  1302600.0 2062800.0 1312800.0 2076600.0 ;
      RECT  1302600.0 2090400.0 1312800.0 2076600.0 ;
      RECT  1302600.0 2090400.0 1312800.0 2104200.0 ;
      RECT  1302600.0 2118000.0 1312800.0 2104200.0 ;
      RECT  1302600.0 2118000.0 1312800.0 2131800.0 ;
      RECT  1302600.0 2145600.0 1312800.0 2131800.0 ;
      RECT  1312800.0 379200.0 1323000.0 393000.0 ;
      RECT  1312800.0 406800.0 1323000.0 393000.0 ;
      RECT  1312800.0 406800.0 1323000.0 420600.0 ;
      RECT  1312800.0 434400.0 1323000.0 420600.0 ;
      RECT  1312800.0 434400.0 1323000.0 448200.0 ;
      RECT  1312800.0 462000.0 1323000.0 448200.0 ;
      RECT  1312800.0 462000.0 1323000.0 475800.0 ;
      RECT  1312800.0 489600.0 1323000.0 475800.0 ;
      RECT  1312800.0 489600.0 1323000.0 503400.0 ;
      RECT  1312800.0 517200.0 1323000.0 503400.0 ;
      RECT  1312800.0 517200.0 1323000.0 531000.0 ;
      RECT  1312800.0 544800.0 1323000.0 531000.0 ;
      RECT  1312800.0 544800.0 1323000.0 558600.0 ;
      RECT  1312800.0 572400.0 1323000.0 558600.0 ;
      RECT  1312800.0 572400.0 1323000.0 586200.0 ;
      RECT  1312800.0 600000.0 1323000.0 586200.0 ;
      RECT  1312800.0 600000.0 1323000.0 613800.0 ;
      RECT  1312800.0 627600.0 1323000.0 613800.0 ;
      RECT  1312800.0 627600.0 1323000.0 641400.0 ;
      RECT  1312800.0 655200.0 1323000.0 641400.0 ;
      RECT  1312800.0 655200.0 1323000.0 669000.0 ;
      RECT  1312800.0 682800.0 1323000.0 669000.0 ;
      RECT  1312800.0 682800.0 1323000.0 696600.0 ;
      RECT  1312800.0 710400.0 1323000.0 696600.0 ;
      RECT  1312800.0 710400.0 1323000.0 724200.0 ;
      RECT  1312800.0 738000.0 1323000.0 724200.0 ;
      RECT  1312800.0 738000.0 1323000.0 751800.0 ;
      RECT  1312800.0 765600.0 1323000.0 751800.0 ;
      RECT  1312800.0 765600.0 1323000.0 779400.0 ;
      RECT  1312800.0 793200.0 1323000.0 779400.0 ;
      RECT  1312800.0 793200.0 1323000.0 807000.0 ;
      RECT  1312800.0 820800.0 1323000.0 807000.0 ;
      RECT  1312800.0 820800.0 1323000.0 834600.0 ;
      RECT  1312800.0 848400.0 1323000.0 834600.0 ;
      RECT  1312800.0 848400.0 1323000.0 862200.0 ;
      RECT  1312800.0 876000.0 1323000.0 862200.0 ;
      RECT  1312800.0 876000.0 1323000.0 889800.0 ;
      RECT  1312800.0 903600.0 1323000.0 889800.0 ;
      RECT  1312800.0 903600.0 1323000.0 917400.0 ;
      RECT  1312800.0 931200.0 1323000.0 917400.0 ;
      RECT  1312800.0 931200.0 1323000.0 945000.0 ;
      RECT  1312800.0 958800.0 1323000.0 945000.0 ;
      RECT  1312800.0 958800.0 1323000.0 972600.0 ;
      RECT  1312800.0 986400.0 1323000.0 972600.0 ;
      RECT  1312800.0 986400.0 1323000.0 1000200.0 ;
      RECT  1312800.0 1014000.0 1323000.0 1000200.0 ;
      RECT  1312800.0 1014000.0 1323000.0 1027800.0 ;
      RECT  1312800.0 1041600.0 1323000.0 1027800.0 ;
      RECT  1312800.0 1041600.0 1323000.0 1055400.0 ;
      RECT  1312800.0 1069200.0 1323000.0 1055400.0 ;
      RECT  1312800.0 1069200.0 1323000.0 1083000.0 ;
      RECT  1312800.0 1096800.0 1323000.0 1083000.0 ;
      RECT  1312800.0 1096800.0 1323000.0 1110600.0 ;
      RECT  1312800.0 1124400.0 1323000.0 1110600.0 ;
      RECT  1312800.0 1124400.0 1323000.0 1138200.0 ;
      RECT  1312800.0 1152000.0 1323000.0 1138200.0 ;
      RECT  1312800.0 1152000.0 1323000.0 1165800.0 ;
      RECT  1312800.0 1179600.0 1323000.0 1165800.0 ;
      RECT  1312800.0 1179600.0 1323000.0 1193400.0 ;
      RECT  1312800.0 1207200.0 1323000.0 1193400.0 ;
      RECT  1312800.0 1207200.0 1323000.0 1221000.0 ;
      RECT  1312800.0 1234800.0 1323000.0 1221000.0 ;
      RECT  1312800.0 1234800.0 1323000.0 1248600.0 ;
      RECT  1312800.0 1262400.0 1323000.0 1248600.0 ;
      RECT  1312800.0 1262400.0 1323000.0 1276200.0 ;
      RECT  1312800.0 1290000.0 1323000.0 1276200.0 ;
      RECT  1312800.0 1290000.0 1323000.0 1303800.0 ;
      RECT  1312800.0 1317600.0 1323000.0 1303800.0 ;
      RECT  1312800.0 1317600.0 1323000.0 1331400.0 ;
      RECT  1312800.0 1345200.0 1323000.0 1331400.0 ;
      RECT  1312800.0 1345200.0 1323000.0 1359000.0 ;
      RECT  1312800.0 1372800.0 1323000.0 1359000.0 ;
      RECT  1312800.0 1372800.0 1323000.0 1386600.0 ;
      RECT  1312800.0 1400400.0 1323000.0 1386600.0 ;
      RECT  1312800.0 1400400.0 1323000.0 1414200.0 ;
      RECT  1312800.0 1428000.0 1323000.0 1414200.0 ;
      RECT  1312800.0 1428000.0 1323000.0 1441800.0 ;
      RECT  1312800.0 1455600.0 1323000.0 1441800.0 ;
      RECT  1312800.0 1455600.0 1323000.0 1469400.0 ;
      RECT  1312800.0 1483200.0 1323000.0 1469400.0 ;
      RECT  1312800.0 1483200.0 1323000.0 1497000.0 ;
      RECT  1312800.0 1510800.0 1323000.0 1497000.0 ;
      RECT  1312800.0 1510800.0 1323000.0 1524600.0 ;
      RECT  1312800.0 1538400.0 1323000.0 1524600.0 ;
      RECT  1312800.0 1538400.0 1323000.0 1552200.0 ;
      RECT  1312800.0 1566000.0 1323000.0 1552200.0 ;
      RECT  1312800.0 1566000.0 1323000.0 1579800.0 ;
      RECT  1312800.0 1593600.0 1323000.0 1579800.0 ;
      RECT  1312800.0 1593600.0 1323000.0 1607400.0 ;
      RECT  1312800.0 1621200.0 1323000.0 1607400.0 ;
      RECT  1312800.0 1621200.0 1323000.0 1635000.0 ;
      RECT  1312800.0 1648800.0 1323000.0 1635000.0 ;
      RECT  1312800.0 1648800.0 1323000.0 1662600.0 ;
      RECT  1312800.0 1676400.0 1323000.0 1662600.0 ;
      RECT  1312800.0 1676400.0 1323000.0 1690200.0 ;
      RECT  1312800.0 1704000.0 1323000.0 1690200.0 ;
      RECT  1312800.0 1704000.0 1323000.0 1717800.0 ;
      RECT  1312800.0 1731600.0 1323000.0 1717800.0 ;
      RECT  1312800.0 1731600.0 1323000.0 1745400.0 ;
      RECT  1312800.0 1759200.0 1323000.0 1745400.0 ;
      RECT  1312800.0 1759200.0 1323000.0 1773000.0 ;
      RECT  1312800.0 1786800.0 1323000.0 1773000.0 ;
      RECT  1312800.0 1786800.0 1323000.0 1800600.0 ;
      RECT  1312800.0 1814400.0 1323000.0 1800600.0 ;
      RECT  1312800.0 1814400.0 1323000.0 1828200.0 ;
      RECT  1312800.0 1842000.0 1323000.0 1828200.0 ;
      RECT  1312800.0 1842000.0 1323000.0 1855800.0 ;
      RECT  1312800.0 1869600.0 1323000.0 1855800.0 ;
      RECT  1312800.0 1869600.0 1323000.0 1883400.0 ;
      RECT  1312800.0 1897200.0 1323000.0 1883400.0 ;
      RECT  1312800.0 1897200.0 1323000.0 1911000.0 ;
      RECT  1312800.0 1924800.0 1323000.0 1911000.0 ;
      RECT  1312800.0 1924800.0 1323000.0 1938600.0 ;
      RECT  1312800.0 1952400.0 1323000.0 1938600.0 ;
      RECT  1312800.0 1952400.0 1323000.0 1966200.0 ;
      RECT  1312800.0 1980000.0 1323000.0 1966200.0 ;
      RECT  1312800.0 1980000.0 1323000.0 1993800.0 ;
      RECT  1312800.0 2007600.0 1323000.0 1993800.0 ;
      RECT  1312800.0 2007600.0 1323000.0 2021400.0 ;
      RECT  1312800.0 2035200.0 1323000.0 2021400.0 ;
      RECT  1312800.0 2035200.0 1323000.0 2049000.0 ;
      RECT  1312800.0 2062800.0 1323000.0 2049000.0 ;
      RECT  1312800.0 2062800.0 1323000.0 2076600.0 ;
      RECT  1312800.0 2090400.0 1323000.0 2076600.0 ;
      RECT  1312800.0 2090400.0 1323000.0 2104200.0 ;
      RECT  1312800.0 2118000.0 1323000.0 2104200.0 ;
      RECT  1312800.0 2118000.0 1323000.0 2131800.0 ;
      RECT  1312800.0 2145600.0 1323000.0 2131800.0 ;
      RECT  1323000.0 379200.0 1333200.0 393000.0 ;
      RECT  1323000.0 406800.0 1333200.0 393000.0 ;
      RECT  1323000.0 406800.0 1333200.0 420600.0 ;
      RECT  1323000.0 434400.0 1333200.0 420600.0 ;
      RECT  1323000.0 434400.0 1333200.0 448200.0 ;
      RECT  1323000.0 462000.0 1333200.0 448200.0 ;
      RECT  1323000.0 462000.0 1333200.0 475800.0 ;
      RECT  1323000.0 489600.0 1333200.0 475800.0 ;
      RECT  1323000.0 489600.0 1333200.0 503400.0 ;
      RECT  1323000.0 517200.0 1333200.0 503400.0 ;
      RECT  1323000.0 517200.0 1333200.0 531000.0 ;
      RECT  1323000.0 544800.0 1333200.0 531000.0 ;
      RECT  1323000.0 544800.0 1333200.0 558600.0 ;
      RECT  1323000.0 572400.0 1333200.0 558600.0 ;
      RECT  1323000.0 572400.0 1333200.0 586200.0 ;
      RECT  1323000.0 600000.0 1333200.0 586200.0 ;
      RECT  1323000.0 600000.0 1333200.0 613800.0 ;
      RECT  1323000.0 627600.0 1333200.0 613800.0 ;
      RECT  1323000.0 627600.0 1333200.0 641400.0 ;
      RECT  1323000.0 655200.0 1333200.0 641400.0 ;
      RECT  1323000.0 655200.0 1333200.0 669000.0 ;
      RECT  1323000.0 682800.0 1333200.0 669000.0 ;
      RECT  1323000.0 682800.0 1333200.0 696600.0 ;
      RECT  1323000.0 710400.0 1333200.0 696600.0 ;
      RECT  1323000.0 710400.0 1333200.0 724200.0 ;
      RECT  1323000.0 738000.0 1333200.0 724200.0 ;
      RECT  1323000.0 738000.0 1333200.0 751800.0 ;
      RECT  1323000.0 765600.0 1333200.0 751800.0 ;
      RECT  1323000.0 765600.0 1333200.0 779400.0 ;
      RECT  1323000.0 793200.0 1333200.0 779400.0 ;
      RECT  1323000.0 793200.0 1333200.0 807000.0 ;
      RECT  1323000.0 820800.0 1333200.0 807000.0 ;
      RECT  1323000.0 820800.0 1333200.0 834600.0 ;
      RECT  1323000.0 848400.0 1333200.0 834600.0 ;
      RECT  1323000.0 848400.0 1333200.0 862200.0 ;
      RECT  1323000.0 876000.0 1333200.0 862200.0 ;
      RECT  1323000.0 876000.0 1333200.0 889800.0 ;
      RECT  1323000.0 903600.0 1333200.0 889800.0 ;
      RECT  1323000.0 903600.0 1333200.0 917400.0 ;
      RECT  1323000.0 931200.0 1333200.0 917400.0 ;
      RECT  1323000.0 931200.0 1333200.0 945000.0 ;
      RECT  1323000.0 958800.0 1333200.0 945000.0 ;
      RECT  1323000.0 958800.0 1333200.0 972600.0 ;
      RECT  1323000.0 986400.0 1333200.0 972600.0 ;
      RECT  1323000.0 986400.0 1333200.0 1000200.0 ;
      RECT  1323000.0 1014000.0 1333200.0 1000200.0 ;
      RECT  1323000.0 1014000.0 1333200.0 1027800.0 ;
      RECT  1323000.0 1041600.0 1333200.0 1027800.0 ;
      RECT  1323000.0 1041600.0 1333200.0 1055400.0 ;
      RECT  1323000.0 1069200.0 1333200.0 1055400.0 ;
      RECT  1323000.0 1069200.0 1333200.0 1083000.0 ;
      RECT  1323000.0 1096800.0 1333200.0 1083000.0 ;
      RECT  1323000.0 1096800.0 1333200.0 1110600.0 ;
      RECT  1323000.0 1124400.0 1333200.0 1110600.0 ;
      RECT  1323000.0 1124400.0 1333200.0 1138200.0 ;
      RECT  1323000.0 1152000.0 1333200.0 1138200.0 ;
      RECT  1323000.0 1152000.0 1333200.0 1165800.0 ;
      RECT  1323000.0 1179600.0 1333200.0 1165800.0 ;
      RECT  1323000.0 1179600.0 1333200.0 1193400.0 ;
      RECT  1323000.0 1207200.0 1333200.0 1193400.0 ;
      RECT  1323000.0 1207200.0 1333200.0 1221000.0 ;
      RECT  1323000.0 1234800.0 1333200.0 1221000.0 ;
      RECT  1323000.0 1234800.0 1333200.0 1248600.0 ;
      RECT  1323000.0 1262400.0 1333200.0 1248600.0 ;
      RECT  1323000.0 1262400.0 1333200.0 1276200.0 ;
      RECT  1323000.0 1290000.0 1333200.0 1276200.0 ;
      RECT  1323000.0 1290000.0 1333200.0 1303800.0 ;
      RECT  1323000.0 1317600.0 1333200.0 1303800.0 ;
      RECT  1323000.0 1317600.0 1333200.0 1331400.0 ;
      RECT  1323000.0 1345200.0 1333200.0 1331400.0 ;
      RECT  1323000.0 1345200.0 1333200.0 1359000.0 ;
      RECT  1323000.0 1372800.0 1333200.0 1359000.0 ;
      RECT  1323000.0 1372800.0 1333200.0 1386600.0 ;
      RECT  1323000.0 1400400.0 1333200.0 1386600.0 ;
      RECT  1323000.0 1400400.0 1333200.0 1414200.0 ;
      RECT  1323000.0 1428000.0 1333200.0 1414200.0 ;
      RECT  1323000.0 1428000.0 1333200.0 1441800.0 ;
      RECT  1323000.0 1455600.0 1333200.0 1441800.0 ;
      RECT  1323000.0 1455600.0 1333200.0 1469400.0 ;
      RECT  1323000.0 1483200.0 1333200.0 1469400.0 ;
      RECT  1323000.0 1483200.0 1333200.0 1497000.0 ;
      RECT  1323000.0 1510800.0 1333200.0 1497000.0 ;
      RECT  1323000.0 1510800.0 1333200.0 1524600.0 ;
      RECT  1323000.0 1538400.0 1333200.0 1524600.0 ;
      RECT  1323000.0 1538400.0 1333200.0 1552200.0 ;
      RECT  1323000.0 1566000.0 1333200.0 1552200.0 ;
      RECT  1323000.0 1566000.0 1333200.0 1579800.0 ;
      RECT  1323000.0 1593600.0 1333200.0 1579800.0 ;
      RECT  1323000.0 1593600.0 1333200.0 1607400.0 ;
      RECT  1323000.0 1621200.0 1333200.0 1607400.0 ;
      RECT  1323000.0 1621200.0 1333200.0 1635000.0 ;
      RECT  1323000.0 1648800.0 1333200.0 1635000.0 ;
      RECT  1323000.0 1648800.0 1333200.0 1662600.0 ;
      RECT  1323000.0 1676400.0 1333200.0 1662600.0 ;
      RECT  1323000.0 1676400.0 1333200.0 1690200.0 ;
      RECT  1323000.0 1704000.0 1333200.0 1690200.0 ;
      RECT  1323000.0 1704000.0 1333200.0 1717800.0 ;
      RECT  1323000.0 1731600.0 1333200.0 1717800.0 ;
      RECT  1323000.0 1731600.0 1333200.0 1745400.0 ;
      RECT  1323000.0 1759200.0 1333200.0 1745400.0 ;
      RECT  1323000.0 1759200.0 1333200.0 1773000.0 ;
      RECT  1323000.0 1786800.0 1333200.0 1773000.0 ;
      RECT  1323000.0 1786800.0 1333200.0 1800600.0 ;
      RECT  1323000.0 1814400.0 1333200.0 1800600.0 ;
      RECT  1323000.0 1814400.0 1333200.0 1828200.0 ;
      RECT  1323000.0 1842000.0 1333200.0 1828200.0 ;
      RECT  1323000.0 1842000.0 1333200.0 1855800.0 ;
      RECT  1323000.0 1869600.0 1333200.0 1855800.0 ;
      RECT  1323000.0 1869600.0 1333200.0 1883400.0 ;
      RECT  1323000.0 1897200.0 1333200.0 1883400.0 ;
      RECT  1323000.0 1897200.0 1333200.0 1911000.0 ;
      RECT  1323000.0 1924800.0 1333200.0 1911000.0 ;
      RECT  1323000.0 1924800.0 1333200.0 1938600.0 ;
      RECT  1323000.0 1952400.0 1333200.0 1938600.0 ;
      RECT  1323000.0 1952400.0 1333200.0 1966200.0 ;
      RECT  1323000.0 1980000.0 1333200.0 1966200.0 ;
      RECT  1323000.0 1980000.0 1333200.0 1993800.0 ;
      RECT  1323000.0 2007600.0 1333200.0 1993800.0 ;
      RECT  1323000.0 2007600.0 1333200.0 2021400.0 ;
      RECT  1323000.0 2035200.0 1333200.0 2021400.0 ;
      RECT  1323000.0 2035200.0 1333200.0 2049000.0 ;
      RECT  1323000.0 2062800.0 1333200.0 2049000.0 ;
      RECT  1323000.0 2062800.0 1333200.0 2076600.0 ;
      RECT  1323000.0 2090400.0 1333200.0 2076600.0 ;
      RECT  1323000.0 2090400.0 1333200.0 2104200.0 ;
      RECT  1323000.0 2118000.0 1333200.0 2104200.0 ;
      RECT  1323000.0 2118000.0 1333200.0 2131800.0 ;
      RECT  1323000.0 2145600.0 1333200.0 2131800.0 ;
      RECT  1333200.0 379200.0 1343400.0 393000.0 ;
      RECT  1333200.0 406800.0 1343400.0 393000.0 ;
      RECT  1333200.0 406800.0 1343400.0 420600.0 ;
      RECT  1333200.0 434400.0 1343400.0 420600.0 ;
      RECT  1333200.0 434400.0 1343400.0 448200.0 ;
      RECT  1333200.0 462000.0 1343400.0 448200.0 ;
      RECT  1333200.0 462000.0 1343400.0 475800.0 ;
      RECT  1333200.0 489600.0 1343400.0 475800.0 ;
      RECT  1333200.0 489600.0 1343400.0 503400.0 ;
      RECT  1333200.0 517200.0 1343400.0 503400.0 ;
      RECT  1333200.0 517200.0 1343400.0 531000.0 ;
      RECT  1333200.0 544800.0 1343400.0 531000.0 ;
      RECT  1333200.0 544800.0 1343400.0 558600.0 ;
      RECT  1333200.0 572400.0 1343400.0 558600.0 ;
      RECT  1333200.0 572400.0 1343400.0 586200.0 ;
      RECT  1333200.0 600000.0 1343400.0 586200.0 ;
      RECT  1333200.0 600000.0 1343400.0 613800.0 ;
      RECT  1333200.0 627600.0 1343400.0 613800.0 ;
      RECT  1333200.0 627600.0 1343400.0 641400.0 ;
      RECT  1333200.0 655200.0 1343400.0 641400.0 ;
      RECT  1333200.0 655200.0 1343400.0 669000.0 ;
      RECT  1333200.0 682800.0 1343400.0 669000.0 ;
      RECT  1333200.0 682800.0 1343400.0 696600.0 ;
      RECT  1333200.0 710400.0 1343400.0 696600.0 ;
      RECT  1333200.0 710400.0 1343400.0 724200.0 ;
      RECT  1333200.0 738000.0 1343400.0 724200.0 ;
      RECT  1333200.0 738000.0 1343400.0 751800.0 ;
      RECT  1333200.0 765600.0 1343400.0 751800.0 ;
      RECT  1333200.0 765600.0 1343400.0 779400.0 ;
      RECT  1333200.0 793200.0 1343400.0 779400.0 ;
      RECT  1333200.0 793200.0 1343400.0 807000.0 ;
      RECT  1333200.0 820800.0 1343400.0 807000.0 ;
      RECT  1333200.0 820800.0 1343400.0 834600.0 ;
      RECT  1333200.0 848400.0 1343400.0 834600.0 ;
      RECT  1333200.0 848400.0 1343400.0 862200.0 ;
      RECT  1333200.0 876000.0 1343400.0 862200.0 ;
      RECT  1333200.0 876000.0 1343400.0 889800.0 ;
      RECT  1333200.0 903600.0 1343400.0 889800.0 ;
      RECT  1333200.0 903600.0 1343400.0 917400.0 ;
      RECT  1333200.0 931200.0 1343400.0 917400.0 ;
      RECT  1333200.0 931200.0 1343400.0 945000.0 ;
      RECT  1333200.0 958800.0 1343400.0 945000.0 ;
      RECT  1333200.0 958800.0 1343400.0 972600.0 ;
      RECT  1333200.0 986400.0 1343400.0 972600.0 ;
      RECT  1333200.0 986400.0 1343400.0 1000200.0 ;
      RECT  1333200.0 1014000.0 1343400.0 1000200.0 ;
      RECT  1333200.0 1014000.0 1343400.0 1027800.0 ;
      RECT  1333200.0 1041600.0 1343400.0 1027800.0 ;
      RECT  1333200.0 1041600.0 1343400.0 1055400.0 ;
      RECT  1333200.0 1069200.0 1343400.0 1055400.0 ;
      RECT  1333200.0 1069200.0 1343400.0 1083000.0 ;
      RECT  1333200.0 1096800.0 1343400.0 1083000.0 ;
      RECT  1333200.0 1096800.0 1343400.0 1110600.0 ;
      RECT  1333200.0 1124400.0 1343400.0 1110600.0 ;
      RECT  1333200.0 1124400.0 1343400.0 1138200.0 ;
      RECT  1333200.0 1152000.0 1343400.0 1138200.0 ;
      RECT  1333200.0 1152000.0 1343400.0 1165800.0 ;
      RECT  1333200.0 1179600.0 1343400.0 1165800.0 ;
      RECT  1333200.0 1179600.0 1343400.0 1193400.0 ;
      RECT  1333200.0 1207200.0 1343400.0 1193400.0 ;
      RECT  1333200.0 1207200.0 1343400.0 1221000.0 ;
      RECT  1333200.0 1234800.0 1343400.0 1221000.0 ;
      RECT  1333200.0 1234800.0 1343400.0 1248600.0 ;
      RECT  1333200.0 1262400.0 1343400.0 1248600.0 ;
      RECT  1333200.0 1262400.0 1343400.0 1276200.0 ;
      RECT  1333200.0 1290000.0 1343400.0 1276200.0 ;
      RECT  1333200.0 1290000.0 1343400.0 1303800.0 ;
      RECT  1333200.0 1317600.0 1343400.0 1303800.0 ;
      RECT  1333200.0 1317600.0 1343400.0 1331400.0 ;
      RECT  1333200.0 1345200.0 1343400.0 1331400.0 ;
      RECT  1333200.0 1345200.0 1343400.0 1359000.0 ;
      RECT  1333200.0 1372800.0 1343400.0 1359000.0 ;
      RECT  1333200.0 1372800.0 1343400.0 1386600.0 ;
      RECT  1333200.0 1400400.0 1343400.0 1386600.0 ;
      RECT  1333200.0 1400400.0 1343400.0 1414200.0 ;
      RECT  1333200.0 1428000.0 1343400.0 1414200.0 ;
      RECT  1333200.0 1428000.0 1343400.0 1441800.0 ;
      RECT  1333200.0 1455600.0 1343400.0 1441800.0 ;
      RECT  1333200.0 1455600.0 1343400.0 1469400.0 ;
      RECT  1333200.0 1483200.0 1343400.0 1469400.0 ;
      RECT  1333200.0 1483200.0 1343400.0 1497000.0 ;
      RECT  1333200.0 1510800.0 1343400.0 1497000.0 ;
      RECT  1333200.0 1510800.0 1343400.0 1524600.0 ;
      RECT  1333200.0 1538400.0 1343400.0 1524600.0 ;
      RECT  1333200.0 1538400.0 1343400.0 1552200.0 ;
      RECT  1333200.0 1566000.0 1343400.0 1552200.0 ;
      RECT  1333200.0 1566000.0 1343400.0 1579800.0 ;
      RECT  1333200.0 1593600.0 1343400.0 1579800.0 ;
      RECT  1333200.0 1593600.0 1343400.0 1607400.0 ;
      RECT  1333200.0 1621200.0 1343400.0 1607400.0 ;
      RECT  1333200.0 1621200.0 1343400.0 1635000.0 ;
      RECT  1333200.0 1648800.0 1343400.0 1635000.0 ;
      RECT  1333200.0 1648800.0 1343400.0 1662600.0 ;
      RECT  1333200.0 1676400.0 1343400.0 1662600.0 ;
      RECT  1333200.0 1676400.0 1343400.0 1690200.0 ;
      RECT  1333200.0 1704000.0 1343400.0 1690200.0 ;
      RECT  1333200.0 1704000.0 1343400.0 1717800.0 ;
      RECT  1333200.0 1731600.0 1343400.0 1717800.0 ;
      RECT  1333200.0 1731600.0 1343400.0 1745400.0 ;
      RECT  1333200.0 1759200.0 1343400.0 1745400.0 ;
      RECT  1333200.0 1759200.0 1343400.0 1773000.0 ;
      RECT  1333200.0 1786800.0 1343400.0 1773000.0 ;
      RECT  1333200.0 1786800.0 1343400.0 1800600.0 ;
      RECT  1333200.0 1814400.0 1343400.0 1800600.0 ;
      RECT  1333200.0 1814400.0 1343400.0 1828200.0 ;
      RECT  1333200.0 1842000.0 1343400.0 1828200.0 ;
      RECT  1333200.0 1842000.0 1343400.0 1855800.0 ;
      RECT  1333200.0 1869600.0 1343400.0 1855800.0 ;
      RECT  1333200.0 1869600.0 1343400.0 1883400.0 ;
      RECT  1333200.0 1897200.0 1343400.0 1883400.0 ;
      RECT  1333200.0 1897200.0 1343400.0 1911000.0 ;
      RECT  1333200.0 1924800.0 1343400.0 1911000.0 ;
      RECT  1333200.0 1924800.0 1343400.0 1938600.0 ;
      RECT  1333200.0 1952400.0 1343400.0 1938600.0 ;
      RECT  1333200.0 1952400.0 1343400.0 1966200.0 ;
      RECT  1333200.0 1980000.0 1343400.0 1966200.0 ;
      RECT  1333200.0 1980000.0 1343400.0 1993800.0 ;
      RECT  1333200.0 2007600.0 1343400.0 1993800.0 ;
      RECT  1333200.0 2007600.0 1343400.0 2021400.0 ;
      RECT  1333200.0 2035200.0 1343400.0 2021400.0 ;
      RECT  1333200.0 2035200.0 1343400.0 2049000.0 ;
      RECT  1333200.0 2062800.0 1343400.0 2049000.0 ;
      RECT  1333200.0 2062800.0 1343400.0 2076600.0 ;
      RECT  1333200.0 2090400.0 1343400.0 2076600.0 ;
      RECT  1333200.0 2090400.0 1343400.0 2104200.0 ;
      RECT  1333200.0 2118000.0 1343400.0 2104200.0 ;
      RECT  1333200.0 2118000.0 1343400.0 2131800.0 ;
      RECT  1333200.0 2145600.0 1343400.0 2131800.0 ;
      RECT  1343400.0 379200.0 1353600.0 393000.0 ;
      RECT  1343400.0 406800.0 1353600.0 393000.0 ;
      RECT  1343400.0 406800.0 1353600.0 420600.0 ;
      RECT  1343400.0 434400.0 1353600.0 420600.0 ;
      RECT  1343400.0 434400.0 1353600.0 448200.0 ;
      RECT  1343400.0 462000.0 1353600.0 448200.0 ;
      RECT  1343400.0 462000.0 1353600.0 475800.0 ;
      RECT  1343400.0 489600.0 1353600.0 475800.0 ;
      RECT  1343400.0 489600.0 1353600.0 503400.0 ;
      RECT  1343400.0 517200.0 1353600.0 503400.0 ;
      RECT  1343400.0 517200.0 1353600.0 531000.0 ;
      RECT  1343400.0 544800.0 1353600.0 531000.0 ;
      RECT  1343400.0 544800.0 1353600.0 558600.0 ;
      RECT  1343400.0 572400.0 1353600.0 558600.0 ;
      RECT  1343400.0 572400.0 1353600.0 586200.0 ;
      RECT  1343400.0 600000.0 1353600.0 586200.0 ;
      RECT  1343400.0 600000.0 1353600.0 613800.0 ;
      RECT  1343400.0 627600.0 1353600.0 613800.0 ;
      RECT  1343400.0 627600.0 1353600.0 641400.0 ;
      RECT  1343400.0 655200.0 1353600.0 641400.0 ;
      RECT  1343400.0 655200.0 1353600.0 669000.0 ;
      RECT  1343400.0 682800.0 1353600.0 669000.0 ;
      RECT  1343400.0 682800.0 1353600.0 696600.0 ;
      RECT  1343400.0 710400.0 1353600.0 696600.0 ;
      RECT  1343400.0 710400.0 1353600.0 724200.0 ;
      RECT  1343400.0 738000.0 1353600.0 724200.0 ;
      RECT  1343400.0 738000.0 1353600.0 751800.0 ;
      RECT  1343400.0 765600.0 1353600.0 751800.0 ;
      RECT  1343400.0 765600.0 1353600.0 779400.0 ;
      RECT  1343400.0 793200.0 1353600.0 779400.0 ;
      RECT  1343400.0 793200.0 1353600.0 807000.0 ;
      RECT  1343400.0 820800.0 1353600.0 807000.0 ;
      RECT  1343400.0 820800.0 1353600.0 834600.0 ;
      RECT  1343400.0 848400.0 1353600.0 834600.0 ;
      RECT  1343400.0 848400.0 1353600.0 862200.0 ;
      RECT  1343400.0 876000.0 1353600.0 862200.0 ;
      RECT  1343400.0 876000.0 1353600.0 889800.0 ;
      RECT  1343400.0 903600.0 1353600.0 889800.0 ;
      RECT  1343400.0 903600.0 1353600.0 917400.0 ;
      RECT  1343400.0 931200.0 1353600.0 917400.0 ;
      RECT  1343400.0 931200.0 1353600.0 945000.0 ;
      RECT  1343400.0 958800.0 1353600.0 945000.0 ;
      RECT  1343400.0 958800.0 1353600.0 972600.0 ;
      RECT  1343400.0 986400.0 1353600.0 972600.0 ;
      RECT  1343400.0 986400.0 1353600.0 1000200.0 ;
      RECT  1343400.0 1014000.0 1353600.0 1000200.0 ;
      RECT  1343400.0 1014000.0 1353600.0 1027800.0 ;
      RECT  1343400.0 1041600.0 1353600.0 1027800.0 ;
      RECT  1343400.0 1041600.0 1353600.0 1055400.0 ;
      RECT  1343400.0 1069200.0 1353600.0 1055400.0 ;
      RECT  1343400.0 1069200.0 1353600.0 1083000.0 ;
      RECT  1343400.0 1096800.0 1353600.0 1083000.0 ;
      RECT  1343400.0 1096800.0 1353600.0 1110600.0 ;
      RECT  1343400.0 1124400.0 1353600.0 1110600.0 ;
      RECT  1343400.0 1124400.0 1353600.0 1138200.0 ;
      RECT  1343400.0 1152000.0 1353600.0 1138200.0 ;
      RECT  1343400.0 1152000.0 1353600.0 1165800.0 ;
      RECT  1343400.0 1179600.0 1353600.0 1165800.0 ;
      RECT  1343400.0 1179600.0 1353600.0 1193400.0 ;
      RECT  1343400.0 1207200.0 1353600.0 1193400.0 ;
      RECT  1343400.0 1207200.0 1353600.0 1221000.0 ;
      RECT  1343400.0 1234800.0 1353600.0 1221000.0 ;
      RECT  1343400.0 1234800.0 1353600.0 1248600.0 ;
      RECT  1343400.0 1262400.0 1353600.0 1248600.0 ;
      RECT  1343400.0 1262400.0 1353600.0 1276200.0 ;
      RECT  1343400.0 1290000.0 1353600.0 1276200.0 ;
      RECT  1343400.0 1290000.0 1353600.0 1303800.0 ;
      RECT  1343400.0 1317600.0 1353600.0 1303800.0 ;
      RECT  1343400.0 1317600.0 1353600.0 1331400.0 ;
      RECT  1343400.0 1345200.0 1353600.0 1331400.0 ;
      RECT  1343400.0 1345200.0 1353600.0 1359000.0 ;
      RECT  1343400.0 1372800.0 1353600.0 1359000.0 ;
      RECT  1343400.0 1372800.0 1353600.0 1386600.0 ;
      RECT  1343400.0 1400400.0 1353600.0 1386600.0 ;
      RECT  1343400.0 1400400.0 1353600.0 1414200.0 ;
      RECT  1343400.0 1428000.0 1353600.0 1414200.0 ;
      RECT  1343400.0 1428000.0 1353600.0 1441800.0 ;
      RECT  1343400.0 1455600.0 1353600.0 1441800.0 ;
      RECT  1343400.0 1455600.0 1353600.0 1469400.0 ;
      RECT  1343400.0 1483200.0 1353600.0 1469400.0 ;
      RECT  1343400.0 1483200.0 1353600.0 1497000.0 ;
      RECT  1343400.0 1510800.0 1353600.0 1497000.0 ;
      RECT  1343400.0 1510800.0 1353600.0 1524600.0 ;
      RECT  1343400.0 1538400.0 1353600.0 1524600.0 ;
      RECT  1343400.0 1538400.0 1353600.0 1552200.0 ;
      RECT  1343400.0 1566000.0 1353600.0 1552200.0 ;
      RECT  1343400.0 1566000.0 1353600.0 1579800.0 ;
      RECT  1343400.0 1593600.0 1353600.0 1579800.0 ;
      RECT  1343400.0 1593600.0 1353600.0 1607400.0 ;
      RECT  1343400.0 1621200.0 1353600.0 1607400.0 ;
      RECT  1343400.0 1621200.0 1353600.0 1635000.0 ;
      RECT  1343400.0 1648800.0 1353600.0 1635000.0 ;
      RECT  1343400.0 1648800.0 1353600.0 1662600.0 ;
      RECT  1343400.0 1676400.0 1353600.0 1662600.0 ;
      RECT  1343400.0 1676400.0 1353600.0 1690200.0 ;
      RECT  1343400.0 1704000.0 1353600.0 1690200.0 ;
      RECT  1343400.0 1704000.0 1353600.0 1717800.0 ;
      RECT  1343400.0 1731600.0 1353600.0 1717800.0 ;
      RECT  1343400.0 1731600.0 1353600.0 1745400.0 ;
      RECT  1343400.0 1759200.0 1353600.0 1745400.0 ;
      RECT  1343400.0 1759200.0 1353600.0 1773000.0 ;
      RECT  1343400.0 1786800.0 1353600.0 1773000.0 ;
      RECT  1343400.0 1786800.0 1353600.0 1800600.0 ;
      RECT  1343400.0 1814400.0 1353600.0 1800600.0 ;
      RECT  1343400.0 1814400.0 1353600.0 1828200.0 ;
      RECT  1343400.0 1842000.0 1353600.0 1828200.0 ;
      RECT  1343400.0 1842000.0 1353600.0 1855800.0 ;
      RECT  1343400.0 1869600.0 1353600.0 1855800.0 ;
      RECT  1343400.0 1869600.0 1353600.0 1883400.0 ;
      RECT  1343400.0 1897200.0 1353600.0 1883400.0 ;
      RECT  1343400.0 1897200.0 1353600.0 1911000.0 ;
      RECT  1343400.0 1924800.0 1353600.0 1911000.0 ;
      RECT  1343400.0 1924800.0 1353600.0 1938600.0 ;
      RECT  1343400.0 1952400.0 1353600.0 1938600.0 ;
      RECT  1343400.0 1952400.0 1353600.0 1966200.0 ;
      RECT  1343400.0 1980000.0 1353600.0 1966200.0 ;
      RECT  1343400.0 1980000.0 1353600.0 1993800.0 ;
      RECT  1343400.0 2007600.0 1353600.0 1993800.0 ;
      RECT  1343400.0 2007600.0 1353600.0 2021400.0 ;
      RECT  1343400.0 2035200.0 1353600.0 2021400.0 ;
      RECT  1343400.0 2035200.0 1353600.0 2049000.0 ;
      RECT  1343400.0 2062800.0 1353600.0 2049000.0 ;
      RECT  1343400.0 2062800.0 1353600.0 2076600.0 ;
      RECT  1343400.0 2090400.0 1353600.0 2076600.0 ;
      RECT  1343400.0 2090400.0 1353600.0 2104200.0 ;
      RECT  1343400.0 2118000.0 1353600.0 2104200.0 ;
      RECT  1343400.0 2118000.0 1353600.0 2131800.0 ;
      RECT  1343400.0 2145600.0 1353600.0 2131800.0 ;
      RECT  1353600.0 379200.0 1363800.0 393000.0 ;
      RECT  1353600.0 406800.0 1363800.0 393000.0 ;
      RECT  1353600.0 406800.0 1363800.0 420600.0 ;
      RECT  1353600.0 434400.0 1363800.0 420600.0 ;
      RECT  1353600.0 434400.0 1363800.0 448200.0 ;
      RECT  1353600.0 462000.0 1363800.0 448200.0 ;
      RECT  1353600.0 462000.0 1363800.0 475800.0 ;
      RECT  1353600.0 489600.0 1363800.0 475800.0 ;
      RECT  1353600.0 489600.0 1363800.0 503400.0 ;
      RECT  1353600.0 517200.0 1363800.0 503400.0 ;
      RECT  1353600.0 517200.0 1363800.0 531000.0 ;
      RECT  1353600.0 544800.0 1363800.0 531000.0 ;
      RECT  1353600.0 544800.0 1363800.0 558600.0 ;
      RECT  1353600.0 572400.0 1363800.0 558600.0 ;
      RECT  1353600.0 572400.0 1363800.0 586200.0 ;
      RECT  1353600.0 600000.0 1363800.0 586200.0 ;
      RECT  1353600.0 600000.0 1363800.0 613800.0 ;
      RECT  1353600.0 627600.0 1363800.0 613800.0 ;
      RECT  1353600.0 627600.0 1363800.0 641400.0 ;
      RECT  1353600.0 655200.0 1363800.0 641400.0 ;
      RECT  1353600.0 655200.0 1363800.0 669000.0 ;
      RECT  1353600.0 682800.0 1363800.0 669000.0 ;
      RECT  1353600.0 682800.0 1363800.0 696600.0 ;
      RECT  1353600.0 710400.0 1363800.0 696600.0 ;
      RECT  1353600.0 710400.0 1363800.0 724200.0 ;
      RECT  1353600.0 738000.0 1363800.0 724200.0 ;
      RECT  1353600.0 738000.0 1363800.0 751800.0 ;
      RECT  1353600.0 765600.0 1363800.0 751800.0 ;
      RECT  1353600.0 765600.0 1363800.0 779400.0 ;
      RECT  1353600.0 793200.0 1363800.0 779400.0 ;
      RECT  1353600.0 793200.0 1363800.0 807000.0 ;
      RECT  1353600.0 820800.0 1363800.0 807000.0 ;
      RECT  1353600.0 820800.0 1363800.0 834600.0 ;
      RECT  1353600.0 848400.0 1363800.0 834600.0 ;
      RECT  1353600.0 848400.0 1363800.0 862200.0 ;
      RECT  1353600.0 876000.0 1363800.0 862200.0 ;
      RECT  1353600.0 876000.0 1363800.0 889800.0 ;
      RECT  1353600.0 903600.0 1363800.0 889800.0 ;
      RECT  1353600.0 903600.0 1363800.0 917400.0 ;
      RECT  1353600.0 931200.0 1363800.0 917400.0 ;
      RECT  1353600.0 931200.0 1363800.0 945000.0 ;
      RECT  1353600.0 958800.0 1363800.0 945000.0 ;
      RECT  1353600.0 958800.0 1363800.0 972600.0 ;
      RECT  1353600.0 986400.0 1363800.0 972600.0 ;
      RECT  1353600.0 986400.0 1363800.0 1000200.0 ;
      RECT  1353600.0 1014000.0 1363800.0 1000200.0 ;
      RECT  1353600.0 1014000.0 1363800.0 1027800.0 ;
      RECT  1353600.0 1041600.0 1363800.0 1027800.0 ;
      RECT  1353600.0 1041600.0 1363800.0 1055400.0 ;
      RECT  1353600.0 1069200.0 1363800.0 1055400.0 ;
      RECT  1353600.0 1069200.0 1363800.0 1083000.0 ;
      RECT  1353600.0 1096800.0 1363800.0 1083000.0 ;
      RECT  1353600.0 1096800.0 1363800.0 1110600.0 ;
      RECT  1353600.0 1124400.0 1363800.0 1110600.0 ;
      RECT  1353600.0 1124400.0 1363800.0 1138200.0 ;
      RECT  1353600.0 1152000.0 1363800.0 1138200.0 ;
      RECT  1353600.0 1152000.0 1363800.0 1165800.0 ;
      RECT  1353600.0 1179600.0 1363800.0 1165800.0 ;
      RECT  1353600.0 1179600.0 1363800.0 1193400.0 ;
      RECT  1353600.0 1207200.0 1363800.0 1193400.0 ;
      RECT  1353600.0 1207200.0 1363800.0 1221000.0 ;
      RECT  1353600.0 1234800.0 1363800.0 1221000.0 ;
      RECT  1353600.0 1234800.0 1363800.0 1248600.0 ;
      RECT  1353600.0 1262400.0 1363800.0 1248600.0 ;
      RECT  1353600.0 1262400.0 1363800.0 1276200.0 ;
      RECT  1353600.0 1290000.0 1363800.0 1276200.0 ;
      RECT  1353600.0 1290000.0 1363800.0 1303800.0 ;
      RECT  1353600.0 1317600.0 1363800.0 1303800.0 ;
      RECT  1353600.0 1317600.0 1363800.0 1331400.0 ;
      RECT  1353600.0 1345200.0 1363800.0 1331400.0 ;
      RECT  1353600.0 1345200.0 1363800.0 1359000.0 ;
      RECT  1353600.0 1372800.0 1363800.0 1359000.0 ;
      RECT  1353600.0 1372800.0 1363800.0 1386600.0 ;
      RECT  1353600.0 1400400.0 1363800.0 1386600.0 ;
      RECT  1353600.0 1400400.0 1363800.0 1414200.0 ;
      RECT  1353600.0 1428000.0 1363800.0 1414200.0 ;
      RECT  1353600.0 1428000.0 1363800.0 1441800.0 ;
      RECT  1353600.0 1455600.0 1363800.0 1441800.0 ;
      RECT  1353600.0 1455600.0 1363800.0 1469400.0 ;
      RECT  1353600.0 1483200.0 1363800.0 1469400.0 ;
      RECT  1353600.0 1483200.0 1363800.0 1497000.0 ;
      RECT  1353600.0 1510800.0 1363800.0 1497000.0 ;
      RECT  1353600.0 1510800.0 1363800.0 1524600.0 ;
      RECT  1353600.0 1538400.0 1363800.0 1524600.0 ;
      RECT  1353600.0 1538400.0 1363800.0 1552200.0 ;
      RECT  1353600.0 1566000.0 1363800.0 1552200.0 ;
      RECT  1353600.0 1566000.0 1363800.0 1579800.0 ;
      RECT  1353600.0 1593600.0 1363800.0 1579800.0 ;
      RECT  1353600.0 1593600.0 1363800.0 1607400.0 ;
      RECT  1353600.0 1621200.0 1363800.0 1607400.0 ;
      RECT  1353600.0 1621200.0 1363800.0 1635000.0 ;
      RECT  1353600.0 1648800.0 1363800.0 1635000.0 ;
      RECT  1353600.0 1648800.0 1363800.0 1662600.0 ;
      RECT  1353600.0 1676400.0 1363800.0 1662600.0 ;
      RECT  1353600.0 1676400.0 1363800.0 1690200.0 ;
      RECT  1353600.0 1704000.0 1363800.0 1690200.0 ;
      RECT  1353600.0 1704000.0 1363800.0 1717800.0 ;
      RECT  1353600.0 1731600.0 1363800.0 1717800.0 ;
      RECT  1353600.0 1731600.0 1363800.0 1745400.0 ;
      RECT  1353600.0 1759200.0 1363800.0 1745400.0 ;
      RECT  1353600.0 1759200.0 1363800.0 1773000.0 ;
      RECT  1353600.0 1786800.0 1363800.0 1773000.0 ;
      RECT  1353600.0 1786800.0 1363800.0 1800600.0 ;
      RECT  1353600.0 1814400.0 1363800.0 1800600.0 ;
      RECT  1353600.0 1814400.0 1363800.0 1828200.0 ;
      RECT  1353600.0 1842000.0 1363800.0 1828200.0 ;
      RECT  1353600.0 1842000.0 1363800.0 1855800.0 ;
      RECT  1353600.0 1869600.0 1363800.0 1855800.0 ;
      RECT  1353600.0 1869600.0 1363800.0 1883400.0 ;
      RECT  1353600.0 1897200.0 1363800.0 1883400.0 ;
      RECT  1353600.0 1897200.0 1363800.0 1911000.0 ;
      RECT  1353600.0 1924800.0 1363800.0 1911000.0 ;
      RECT  1353600.0 1924800.0 1363800.0 1938600.0 ;
      RECT  1353600.0 1952400.0 1363800.0 1938600.0 ;
      RECT  1353600.0 1952400.0 1363800.0 1966200.0 ;
      RECT  1353600.0 1980000.0 1363800.0 1966200.0 ;
      RECT  1353600.0 1980000.0 1363800.0 1993800.0 ;
      RECT  1353600.0 2007600.0 1363800.0 1993800.0 ;
      RECT  1353600.0 2007600.0 1363800.0 2021400.0 ;
      RECT  1353600.0 2035200.0 1363800.0 2021400.0 ;
      RECT  1353600.0 2035200.0 1363800.0 2049000.0 ;
      RECT  1353600.0 2062800.0 1363800.0 2049000.0 ;
      RECT  1353600.0 2062800.0 1363800.0 2076600.0 ;
      RECT  1353600.0 2090400.0 1363800.0 2076600.0 ;
      RECT  1353600.0 2090400.0 1363800.0 2104200.0 ;
      RECT  1353600.0 2118000.0 1363800.0 2104200.0 ;
      RECT  1353600.0 2118000.0 1363800.0 2131800.0 ;
      RECT  1353600.0 2145600.0 1363800.0 2131800.0 ;
      RECT  1363800.0 379200.0 1374000.0 393000.0 ;
      RECT  1363800.0 406800.0 1374000.0 393000.0 ;
      RECT  1363800.0 406800.0 1374000.0 420600.0 ;
      RECT  1363800.0 434400.0 1374000.0 420600.0 ;
      RECT  1363800.0 434400.0 1374000.0 448200.0 ;
      RECT  1363800.0 462000.0 1374000.0 448200.0 ;
      RECT  1363800.0 462000.0 1374000.0 475800.0 ;
      RECT  1363800.0 489600.0 1374000.0 475800.0 ;
      RECT  1363800.0 489600.0 1374000.0 503400.0 ;
      RECT  1363800.0 517200.0 1374000.0 503400.0 ;
      RECT  1363800.0 517200.0 1374000.0 531000.0 ;
      RECT  1363800.0 544800.0 1374000.0 531000.0 ;
      RECT  1363800.0 544800.0 1374000.0 558600.0 ;
      RECT  1363800.0 572400.0 1374000.0 558600.0 ;
      RECT  1363800.0 572400.0 1374000.0 586200.0 ;
      RECT  1363800.0 600000.0 1374000.0 586200.0 ;
      RECT  1363800.0 600000.0 1374000.0 613800.0 ;
      RECT  1363800.0 627600.0 1374000.0 613800.0 ;
      RECT  1363800.0 627600.0 1374000.0 641400.0 ;
      RECT  1363800.0 655200.0 1374000.0 641400.0 ;
      RECT  1363800.0 655200.0 1374000.0 669000.0 ;
      RECT  1363800.0 682800.0 1374000.0 669000.0 ;
      RECT  1363800.0 682800.0 1374000.0 696600.0 ;
      RECT  1363800.0 710400.0 1374000.0 696600.0 ;
      RECT  1363800.0 710400.0 1374000.0 724200.0 ;
      RECT  1363800.0 738000.0 1374000.0 724200.0 ;
      RECT  1363800.0 738000.0 1374000.0 751800.0 ;
      RECT  1363800.0 765600.0 1374000.0 751800.0 ;
      RECT  1363800.0 765600.0 1374000.0 779400.0 ;
      RECT  1363800.0 793200.0 1374000.0 779400.0 ;
      RECT  1363800.0 793200.0 1374000.0 807000.0 ;
      RECT  1363800.0 820800.0 1374000.0 807000.0 ;
      RECT  1363800.0 820800.0 1374000.0 834600.0 ;
      RECT  1363800.0 848400.0 1374000.0 834600.0 ;
      RECT  1363800.0 848400.0 1374000.0 862200.0 ;
      RECT  1363800.0 876000.0 1374000.0 862200.0 ;
      RECT  1363800.0 876000.0 1374000.0 889800.0 ;
      RECT  1363800.0 903600.0 1374000.0 889800.0 ;
      RECT  1363800.0 903600.0 1374000.0 917400.0 ;
      RECT  1363800.0 931200.0 1374000.0 917400.0 ;
      RECT  1363800.0 931200.0 1374000.0 945000.0 ;
      RECT  1363800.0 958800.0 1374000.0 945000.0 ;
      RECT  1363800.0 958800.0 1374000.0 972600.0 ;
      RECT  1363800.0 986400.0 1374000.0 972600.0 ;
      RECT  1363800.0 986400.0 1374000.0 1000200.0 ;
      RECT  1363800.0 1014000.0 1374000.0 1000200.0 ;
      RECT  1363800.0 1014000.0 1374000.0 1027800.0 ;
      RECT  1363800.0 1041600.0 1374000.0 1027800.0 ;
      RECT  1363800.0 1041600.0 1374000.0 1055400.0 ;
      RECT  1363800.0 1069200.0 1374000.0 1055400.0 ;
      RECT  1363800.0 1069200.0 1374000.0 1083000.0 ;
      RECT  1363800.0 1096800.0 1374000.0 1083000.0 ;
      RECT  1363800.0 1096800.0 1374000.0 1110600.0 ;
      RECT  1363800.0 1124400.0 1374000.0 1110600.0 ;
      RECT  1363800.0 1124400.0 1374000.0 1138200.0 ;
      RECT  1363800.0 1152000.0 1374000.0 1138200.0 ;
      RECT  1363800.0 1152000.0 1374000.0 1165800.0 ;
      RECT  1363800.0 1179600.0 1374000.0 1165800.0 ;
      RECT  1363800.0 1179600.0 1374000.0 1193400.0 ;
      RECT  1363800.0 1207200.0 1374000.0 1193400.0 ;
      RECT  1363800.0 1207200.0 1374000.0 1221000.0 ;
      RECT  1363800.0 1234800.0 1374000.0 1221000.0 ;
      RECT  1363800.0 1234800.0 1374000.0 1248600.0 ;
      RECT  1363800.0 1262400.0 1374000.0 1248600.0 ;
      RECT  1363800.0 1262400.0 1374000.0 1276200.0 ;
      RECT  1363800.0 1290000.0 1374000.0 1276200.0 ;
      RECT  1363800.0 1290000.0 1374000.0 1303800.0 ;
      RECT  1363800.0 1317600.0 1374000.0 1303800.0 ;
      RECT  1363800.0 1317600.0 1374000.0 1331400.0 ;
      RECT  1363800.0 1345200.0 1374000.0 1331400.0 ;
      RECT  1363800.0 1345200.0 1374000.0 1359000.0 ;
      RECT  1363800.0 1372800.0 1374000.0 1359000.0 ;
      RECT  1363800.0 1372800.0 1374000.0 1386600.0 ;
      RECT  1363800.0 1400400.0 1374000.0 1386600.0 ;
      RECT  1363800.0 1400400.0 1374000.0 1414200.0 ;
      RECT  1363800.0 1428000.0 1374000.0 1414200.0 ;
      RECT  1363800.0 1428000.0 1374000.0 1441800.0 ;
      RECT  1363800.0 1455600.0 1374000.0 1441800.0 ;
      RECT  1363800.0 1455600.0 1374000.0 1469400.0 ;
      RECT  1363800.0 1483200.0 1374000.0 1469400.0 ;
      RECT  1363800.0 1483200.0 1374000.0 1497000.0 ;
      RECT  1363800.0 1510800.0 1374000.0 1497000.0 ;
      RECT  1363800.0 1510800.0 1374000.0 1524600.0 ;
      RECT  1363800.0 1538400.0 1374000.0 1524600.0 ;
      RECT  1363800.0 1538400.0 1374000.0 1552200.0 ;
      RECT  1363800.0 1566000.0 1374000.0 1552200.0 ;
      RECT  1363800.0 1566000.0 1374000.0 1579800.0 ;
      RECT  1363800.0 1593600.0 1374000.0 1579800.0 ;
      RECT  1363800.0 1593600.0 1374000.0 1607400.0 ;
      RECT  1363800.0 1621200.0 1374000.0 1607400.0 ;
      RECT  1363800.0 1621200.0 1374000.0 1635000.0 ;
      RECT  1363800.0 1648800.0 1374000.0 1635000.0 ;
      RECT  1363800.0 1648800.0 1374000.0 1662600.0 ;
      RECT  1363800.0 1676400.0 1374000.0 1662600.0 ;
      RECT  1363800.0 1676400.0 1374000.0 1690200.0 ;
      RECT  1363800.0 1704000.0 1374000.0 1690200.0 ;
      RECT  1363800.0 1704000.0 1374000.0 1717800.0 ;
      RECT  1363800.0 1731600.0 1374000.0 1717800.0 ;
      RECT  1363800.0 1731600.0 1374000.0 1745400.0 ;
      RECT  1363800.0 1759200.0 1374000.0 1745400.0 ;
      RECT  1363800.0 1759200.0 1374000.0 1773000.0 ;
      RECT  1363800.0 1786800.0 1374000.0 1773000.0 ;
      RECT  1363800.0 1786800.0 1374000.0 1800600.0 ;
      RECT  1363800.0 1814400.0 1374000.0 1800600.0 ;
      RECT  1363800.0 1814400.0 1374000.0 1828200.0 ;
      RECT  1363800.0 1842000.0 1374000.0 1828200.0 ;
      RECT  1363800.0 1842000.0 1374000.0 1855800.0 ;
      RECT  1363800.0 1869600.0 1374000.0 1855800.0 ;
      RECT  1363800.0 1869600.0 1374000.0 1883400.0 ;
      RECT  1363800.0 1897200.0 1374000.0 1883400.0 ;
      RECT  1363800.0 1897200.0 1374000.0 1911000.0 ;
      RECT  1363800.0 1924800.0 1374000.0 1911000.0 ;
      RECT  1363800.0 1924800.0 1374000.0 1938600.0 ;
      RECT  1363800.0 1952400.0 1374000.0 1938600.0 ;
      RECT  1363800.0 1952400.0 1374000.0 1966200.0 ;
      RECT  1363800.0 1980000.0 1374000.0 1966200.0 ;
      RECT  1363800.0 1980000.0 1374000.0 1993800.0 ;
      RECT  1363800.0 2007600.0 1374000.0 1993800.0 ;
      RECT  1363800.0 2007600.0 1374000.0 2021400.0 ;
      RECT  1363800.0 2035200.0 1374000.0 2021400.0 ;
      RECT  1363800.0 2035200.0 1374000.0 2049000.0 ;
      RECT  1363800.0 2062800.0 1374000.0 2049000.0 ;
      RECT  1363800.0 2062800.0 1374000.0 2076600.0 ;
      RECT  1363800.0 2090400.0 1374000.0 2076600.0 ;
      RECT  1363800.0 2090400.0 1374000.0 2104200.0 ;
      RECT  1363800.0 2118000.0 1374000.0 2104200.0 ;
      RECT  1363800.0 2118000.0 1374000.0 2131800.0 ;
      RECT  1363800.0 2145600.0 1374000.0 2131800.0 ;
      RECT  1374000.0 379200.0 1384200.0 393000.0 ;
      RECT  1374000.0 406800.0 1384200.0 393000.0 ;
      RECT  1374000.0 406800.0 1384200.0 420600.0 ;
      RECT  1374000.0 434400.0 1384200.0 420600.0 ;
      RECT  1374000.0 434400.0 1384200.0 448200.0 ;
      RECT  1374000.0 462000.0 1384200.0 448200.0 ;
      RECT  1374000.0 462000.0 1384200.0 475800.0 ;
      RECT  1374000.0 489600.0 1384200.0 475800.0 ;
      RECT  1374000.0 489600.0 1384200.0 503400.0 ;
      RECT  1374000.0 517200.0 1384200.0 503400.0 ;
      RECT  1374000.0 517200.0 1384200.0 531000.0 ;
      RECT  1374000.0 544800.0 1384200.0 531000.0 ;
      RECT  1374000.0 544800.0 1384200.0 558600.0 ;
      RECT  1374000.0 572400.0 1384200.0 558600.0 ;
      RECT  1374000.0 572400.0 1384200.0 586200.0 ;
      RECT  1374000.0 600000.0 1384200.0 586200.0 ;
      RECT  1374000.0 600000.0 1384200.0 613800.0 ;
      RECT  1374000.0 627600.0 1384200.0 613800.0 ;
      RECT  1374000.0 627600.0 1384200.0 641400.0 ;
      RECT  1374000.0 655200.0 1384200.0 641400.0 ;
      RECT  1374000.0 655200.0 1384200.0 669000.0 ;
      RECT  1374000.0 682800.0 1384200.0 669000.0 ;
      RECT  1374000.0 682800.0 1384200.0 696600.0 ;
      RECT  1374000.0 710400.0 1384200.0 696600.0 ;
      RECT  1374000.0 710400.0 1384200.0 724200.0 ;
      RECT  1374000.0 738000.0 1384200.0 724200.0 ;
      RECT  1374000.0 738000.0 1384200.0 751800.0 ;
      RECT  1374000.0 765600.0 1384200.0 751800.0 ;
      RECT  1374000.0 765600.0 1384200.0 779400.0 ;
      RECT  1374000.0 793200.0 1384200.0 779400.0 ;
      RECT  1374000.0 793200.0 1384200.0 807000.0 ;
      RECT  1374000.0 820800.0 1384200.0 807000.0 ;
      RECT  1374000.0 820800.0 1384200.0 834600.0 ;
      RECT  1374000.0 848400.0 1384200.0 834600.0 ;
      RECT  1374000.0 848400.0 1384200.0 862200.0 ;
      RECT  1374000.0 876000.0 1384200.0 862200.0 ;
      RECT  1374000.0 876000.0 1384200.0 889800.0 ;
      RECT  1374000.0 903600.0 1384200.0 889800.0 ;
      RECT  1374000.0 903600.0 1384200.0 917400.0 ;
      RECT  1374000.0 931200.0 1384200.0 917400.0 ;
      RECT  1374000.0 931200.0 1384200.0 945000.0 ;
      RECT  1374000.0 958800.0 1384200.0 945000.0 ;
      RECT  1374000.0 958800.0 1384200.0 972600.0 ;
      RECT  1374000.0 986400.0 1384200.0 972600.0 ;
      RECT  1374000.0 986400.0 1384200.0 1000200.0 ;
      RECT  1374000.0 1014000.0 1384200.0 1000200.0 ;
      RECT  1374000.0 1014000.0 1384200.0 1027800.0 ;
      RECT  1374000.0 1041600.0 1384200.0 1027800.0 ;
      RECT  1374000.0 1041600.0 1384200.0 1055400.0 ;
      RECT  1374000.0 1069200.0 1384200.0 1055400.0 ;
      RECT  1374000.0 1069200.0 1384200.0 1083000.0 ;
      RECT  1374000.0 1096800.0 1384200.0 1083000.0 ;
      RECT  1374000.0 1096800.0 1384200.0 1110600.0 ;
      RECT  1374000.0 1124400.0 1384200.0 1110600.0 ;
      RECT  1374000.0 1124400.0 1384200.0 1138200.0 ;
      RECT  1374000.0 1152000.0 1384200.0 1138200.0 ;
      RECT  1374000.0 1152000.0 1384200.0 1165800.0 ;
      RECT  1374000.0 1179600.0 1384200.0 1165800.0 ;
      RECT  1374000.0 1179600.0 1384200.0 1193400.0 ;
      RECT  1374000.0 1207200.0 1384200.0 1193400.0 ;
      RECT  1374000.0 1207200.0 1384200.0 1221000.0 ;
      RECT  1374000.0 1234800.0 1384200.0 1221000.0 ;
      RECT  1374000.0 1234800.0 1384200.0 1248600.0 ;
      RECT  1374000.0 1262400.0 1384200.0 1248600.0 ;
      RECT  1374000.0 1262400.0 1384200.0 1276200.0 ;
      RECT  1374000.0 1290000.0 1384200.0 1276200.0 ;
      RECT  1374000.0 1290000.0 1384200.0 1303800.0 ;
      RECT  1374000.0 1317600.0 1384200.0 1303800.0 ;
      RECT  1374000.0 1317600.0 1384200.0 1331400.0 ;
      RECT  1374000.0 1345200.0 1384200.0 1331400.0 ;
      RECT  1374000.0 1345200.0 1384200.0 1359000.0 ;
      RECT  1374000.0 1372800.0 1384200.0 1359000.0 ;
      RECT  1374000.0 1372800.0 1384200.0 1386600.0 ;
      RECT  1374000.0 1400400.0 1384200.0 1386600.0 ;
      RECT  1374000.0 1400400.0 1384200.0 1414200.0 ;
      RECT  1374000.0 1428000.0 1384200.0 1414200.0 ;
      RECT  1374000.0 1428000.0 1384200.0 1441800.0 ;
      RECT  1374000.0 1455600.0 1384200.0 1441800.0 ;
      RECT  1374000.0 1455600.0 1384200.0 1469400.0 ;
      RECT  1374000.0 1483200.0 1384200.0 1469400.0 ;
      RECT  1374000.0 1483200.0 1384200.0 1497000.0 ;
      RECT  1374000.0 1510800.0 1384200.0 1497000.0 ;
      RECT  1374000.0 1510800.0 1384200.0 1524600.0 ;
      RECT  1374000.0 1538400.0 1384200.0 1524600.0 ;
      RECT  1374000.0 1538400.0 1384200.0 1552200.0 ;
      RECT  1374000.0 1566000.0 1384200.0 1552200.0 ;
      RECT  1374000.0 1566000.0 1384200.0 1579800.0 ;
      RECT  1374000.0 1593600.0 1384200.0 1579800.0 ;
      RECT  1374000.0 1593600.0 1384200.0 1607400.0 ;
      RECT  1374000.0 1621200.0 1384200.0 1607400.0 ;
      RECT  1374000.0 1621200.0 1384200.0 1635000.0 ;
      RECT  1374000.0 1648800.0 1384200.0 1635000.0 ;
      RECT  1374000.0 1648800.0 1384200.0 1662600.0 ;
      RECT  1374000.0 1676400.0 1384200.0 1662600.0 ;
      RECT  1374000.0 1676400.0 1384200.0 1690200.0 ;
      RECT  1374000.0 1704000.0 1384200.0 1690200.0 ;
      RECT  1374000.0 1704000.0 1384200.0 1717800.0 ;
      RECT  1374000.0 1731600.0 1384200.0 1717800.0 ;
      RECT  1374000.0 1731600.0 1384200.0 1745400.0 ;
      RECT  1374000.0 1759200.0 1384200.0 1745400.0 ;
      RECT  1374000.0 1759200.0 1384200.0 1773000.0 ;
      RECT  1374000.0 1786800.0 1384200.0 1773000.0 ;
      RECT  1374000.0 1786800.0 1384200.0 1800600.0 ;
      RECT  1374000.0 1814400.0 1384200.0 1800600.0 ;
      RECT  1374000.0 1814400.0 1384200.0 1828200.0 ;
      RECT  1374000.0 1842000.0 1384200.0 1828200.0 ;
      RECT  1374000.0 1842000.0 1384200.0 1855800.0 ;
      RECT  1374000.0 1869600.0 1384200.0 1855800.0 ;
      RECT  1374000.0 1869600.0 1384200.0 1883400.0 ;
      RECT  1374000.0 1897200.0 1384200.0 1883400.0 ;
      RECT  1374000.0 1897200.0 1384200.0 1911000.0 ;
      RECT  1374000.0 1924800.0 1384200.0 1911000.0 ;
      RECT  1374000.0 1924800.0 1384200.0 1938600.0 ;
      RECT  1374000.0 1952400.0 1384200.0 1938600.0 ;
      RECT  1374000.0 1952400.0 1384200.0 1966200.0 ;
      RECT  1374000.0 1980000.0 1384200.0 1966200.0 ;
      RECT  1374000.0 1980000.0 1384200.0 1993800.0 ;
      RECT  1374000.0 2007600.0 1384200.0 1993800.0 ;
      RECT  1374000.0 2007600.0 1384200.0 2021400.0 ;
      RECT  1374000.0 2035200.0 1384200.0 2021400.0 ;
      RECT  1374000.0 2035200.0 1384200.0 2049000.0 ;
      RECT  1374000.0 2062800.0 1384200.0 2049000.0 ;
      RECT  1374000.0 2062800.0 1384200.0 2076600.0 ;
      RECT  1374000.0 2090400.0 1384200.0 2076600.0 ;
      RECT  1374000.0 2090400.0 1384200.0 2104200.0 ;
      RECT  1374000.0 2118000.0 1384200.0 2104200.0 ;
      RECT  1374000.0 2118000.0 1384200.0 2131800.0 ;
      RECT  1374000.0 2145600.0 1384200.0 2131800.0 ;
      RECT  1384200.0 379200.0 1394400.0 393000.0 ;
      RECT  1384200.0 406800.0 1394400.0 393000.0 ;
      RECT  1384200.0 406800.0 1394400.0 420600.0 ;
      RECT  1384200.0 434400.0 1394400.0 420600.0 ;
      RECT  1384200.0 434400.0 1394400.0 448200.0 ;
      RECT  1384200.0 462000.0 1394400.0 448200.0 ;
      RECT  1384200.0 462000.0 1394400.0 475800.0 ;
      RECT  1384200.0 489600.0 1394400.0 475800.0 ;
      RECT  1384200.0 489600.0 1394400.0 503400.0 ;
      RECT  1384200.0 517200.0 1394400.0 503400.0 ;
      RECT  1384200.0 517200.0 1394400.0 531000.0 ;
      RECT  1384200.0 544800.0 1394400.0 531000.0 ;
      RECT  1384200.0 544800.0 1394400.0 558600.0 ;
      RECT  1384200.0 572400.0 1394400.0 558600.0 ;
      RECT  1384200.0 572400.0 1394400.0 586200.0 ;
      RECT  1384200.0 600000.0 1394400.0 586200.0 ;
      RECT  1384200.0 600000.0 1394400.0 613800.0 ;
      RECT  1384200.0 627600.0 1394400.0 613800.0 ;
      RECT  1384200.0 627600.0 1394400.0 641400.0 ;
      RECT  1384200.0 655200.0 1394400.0 641400.0 ;
      RECT  1384200.0 655200.0 1394400.0 669000.0 ;
      RECT  1384200.0 682800.0 1394400.0 669000.0 ;
      RECT  1384200.0 682800.0 1394400.0 696600.0 ;
      RECT  1384200.0 710400.0 1394400.0 696600.0 ;
      RECT  1384200.0 710400.0 1394400.0 724200.0 ;
      RECT  1384200.0 738000.0 1394400.0 724200.0 ;
      RECT  1384200.0 738000.0 1394400.0 751800.0 ;
      RECT  1384200.0 765600.0 1394400.0 751800.0 ;
      RECT  1384200.0 765600.0 1394400.0 779400.0 ;
      RECT  1384200.0 793200.0 1394400.0 779400.0 ;
      RECT  1384200.0 793200.0 1394400.0 807000.0 ;
      RECT  1384200.0 820800.0 1394400.0 807000.0 ;
      RECT  1384200.0 820800.0 1394400.0 834600.0 ;
      RECT  1384200.0 848400.0 1394400.0 834600.0 ;
      RECT  1384200.0 848400.0 1394400.0 862200.0 ;
      RECT  1384200.0 876000.0 1394400.0 862200.0 ;
      RECT  1384200.0 876000.0 1394400.0 889800.0 ;
      RECT  1384200.0 903600.0 1394400.0 889800.0 ;
      RECT  1384200.0 903600.0 1394400.0 917400.0 ;
      RECT  1384200.0 931200.0 1394400.0 917400.0 ;
      RECT  1384200.0 931200.0 1394400.0 945000.0 ;
      RECT  1384200.0 958800.0 1394400.0 945000.0 ;
      RECT  1384200.0 958800.0 1394400.0 972600.0 ;
      RECT  1384200.0 986400.0 1394400.0 972600.0 ;
      RECT  1384200.0 986400.0 1394400.0 1000200.0 ;
      RECT  1384200.0 1014000.0 1394400.0 1000200.0 ;
      RECT  1384200.0 1014000.0 1394400.0 1027800.0 ;
      RECT  1384200.0 1041600.0 1394400.0 1027800.0 ;
      RECT  1384200.0 1041600.0 1394400.0 1055400.0 ;
      RECT  1384200.0 1069200.0 1394400.0 1055400.0 ;
      RECT  1384200.0 1069200.0 1394400.0 1083000.0 ;
      RECT  1384200.0 1096800.0 1394400.0 1083000.0 ;
      RECT  1384200.0 1096800.0 1394400.0 1110600.0 ;
      RECT  1384200.0 1124400.0 1394400.0 1110600.0 ;
      RECT  1384200.0 1124400.0 1394400.0 1138200.0 ;
      RECT  1384200.0 1152000.0 1394400.0 1138200.0 ;
      RECT  1384200.0 1152000.0 1394400.0 1165800.0 ;
      RECT  1384200.0 1179600.0 1394400.0 1165800.0 ;
      RECT  1384200.0 1179600.0 1394400.0 1193400.0 ;
      RECT  1384200.0 1207200.0 1394400.0 1193400.0 ;
      RECT  1384200.0 1207200.0 1394400.0 1221000.0 ;
      RECT  1384200.0 1234800.0 1394400.0 1221000.0 ;
      RECT  1384200.0 1234800.0 1394400.0 1248600.0 ;
      RECT  1384200.0 1262400.0 1394400.0 1248600.0 ;
      RECT  1384200.0 1262400.0 1394400.0 1276200.0 ;
      RECT  1384200.0 1290000.0 1394400.0 1276200.0 ;
      RECT  1384200.0 1290000.0 1394400.0 1303800.0 ;
      RECT  1384200.0 1317600.0 1394400.0 1303800.0 ;
      RECT  1384200.0 1317600.0 1394400.0 1331400.0 ;
      RECT  1384200.0 1345200.0 1394400.0 1331400.0 ;
      RECT  1384200.0 1345200.0 1394400.0 1359000.0 ;
      RECT  1384200.0 1372800.0 1394400.0 1359000.0 ;
      RECT  1384200.0 1372800.0 1394400.0 1386600.0 ;
      RECT  1384200.0 1400400.0 1394400.0 1386600.0 ;
      RECT  1384200.0 1400400.0 1394400.0 1414200.0 ;
      RECT  1384200.0 1428000.0 1394400.0 1414200.0 ;
      RECT  1384200.0 1428000.0 1394400.0 1441800.0 ;
      RECT  1384200.0 1455600.0 1394400.0 1441800.0 ;
      RECT  1384200.0 1455600.0 1394400.0 1469400.0 ;
      RECT  1384200.0 1483200.0 1394400.0 1469400.0 ;
      RECT  1384200.0 1483200.0 1394400.0 1497000.0 ;
      RECT  1384200.0 1510800.0 1394400.0 1497000.0 ;
      RECT  1384200.0 1510800.0 1394400.0 1524600.0 ;
      RECT  1384200.0 1538400.0 1394400.0 1524600.0 ;
      RECT  1384200.0 1538400.0 1394400.0 1552200.0 ;
      RECT  1384200.0 1566000.0 1394400.0 1552200.0 ;
      RECT  1384200.0 1566000.0 1394400.0 1579800.0 ;
      RECT  1384200.0 1593600.0 1394400.0 1579800.0 ;
      RECT  1384200.0 1593600.0 1394400.0 1607400.0 ;
      RECT  1384200.0 1621200.0 1394400.0 1607400.0 ;
      RECT  1384200.0 1621200.0 1394400.0 1635000.0 ;
      RECT  1384200.0 1648800.0 1394400.0 1635000.0 ;
      RECT  1384200.0 1648800.0 1394400.0 1662600.0 ;
      RECT  1384200.0 1676400.0 1394400.0 1662600.0 ;
      RECT  1384200.0 1676400.0 1394400.0 1690200.0 ;
      RECT  1384200.0 1704000.0 1394400.0 1690200.0 ;
      RECT  1384200.0 1704000.0 1394400.0 1717800.0 ;
      RECT  1384200.0 1731600.0 1394400.0 1717800.0 ;
      RECT  1384200.0 1731600.0 1394400.0 1745400.0 ;
      RECT  1384200.0 1759200.0 1394400.0 1745400.0 ;
      RECT  1384200.0 1759200.0 1394400.0 1773000.0 ;
      RECT  1384200.0 1786800.0 1394400.0 1773000.0 ;
      RECT  1384200.0 1786800.0 1394400.0 1800600.0 ;
      RECT  1384200.0 1814400.0 1394400.0 1800600.0 ;
      RECT  1384200.0 1814400.0 1394400.0 1828200.0 ;
      RECT  1384200.0 1842000.0 1394400.0 1828200.0 ;
      RECT  1384200.0 1842000.0 1394400.0 1855800.0 ;
      RECT  1384200.0 1869600.0 1394400.0 1855800.0 ;
      RECT  1384200.0 1869600.0 1394400.0 1883400.0 ;
      RECT  1384200.0 1897200.0 1394400.0 1883400.0 ;
      RECT  1384200.0 1897200.0 1394400.0 1911000.0 ;
      RECT  1384200.0 1924800.0 1394400.0 1911000.0 ;
      RECT  1384200.0 1924800.0 1394400.0 1938600.0 ;
      RECT  1384200.0 1952400.0 1394400.0 1938600.0 ;
      RECT  1384200.0 1952400.0 1394400.0 1966200.0 ;
      RECT  1384200.0 1980000.0 1394400.0 1966200.0 ;
      RECT  1384200.0 1980000.0 1394400.0 1993800.0 ;
      RECT  1384200.0 2007600.0 1394400.0 1993800.0 ;
      RECT  1384200.0 2007600.0 1394400.0 2021400.0 ;
      RECT  1384200.0 2035200.0 1394400.0 2021400.0 ;
      RECT  1384200.0 2035200.0 1394400.0 2049000.0 ;
      RECT  1384200.0 2062800.0 1394400.0 2049000.0 ;
      RECT  1384200.0 2062800.0 1394400.0 2076600.0 ;
      RECT  1384200.0 2090400.0 1394400.0 2076600.0 ;
      RECT  1384200.0 2090400.0 1394400.0 2104200.0 ;
      RECT  1384200.0 2118000.0 1394400.0 2104200.0 ;
      RECT  1384200.0 2118000.0 1394400.0 2131800.0 ;
      RECT  1384200.0 2145600.0 1394400.0 2131800.0 ;
      RECT  1394400.0 379200.0 1404600.0 393000.0 ;
      RECT  1394400.0 406800.0 1404600.0 393000.0 ;
      RECT  1394400.0 406800.0 1404600.0 420600.0 ;
      RECT  1394400.0 434400.0 1404600.0 420600.0 ;
      RECT  1394400.0 434400.0 1404600.0 448200.0 ;
      RECT  1394400.0 462000.0 1404600.0 448200.0 ;
      RECT  1394400.0 462000.0 1404600.0 475800.0 ;
      RECT  1394400.0 489600.0 1404600.0 475800.0 ;
      RECT  1394400.0 489600.0 1404600.0 503400.0 ;
      RECT  1394400.0 517200.0 1404600.0 503400.0 ;
      RECT  1394400.0 517200.0 1404600.0 531000.0 ;
      RECT  1394400.0 544800.0 1404600.0 531000.0 ;
      RECT  1394400.0 544800.0 1404600.0 558600.0 ;
      RECT  1394400.0 572400.0 1404600.0 558600.0 ;
      RECT  1394400.0 572400.0 1404600.0 586200.0 ;
      RECT  1394400.0 600000.0 1404600.0 586200.0 ;
      RECT  1394400.0 600000.0 1404600.0 613800.0 ;
      RECT  1394400.0 627600.0 1404600.0 613800.0 ;
      RECT  1394400.0 627600.0 1404600.0 641400.0 ;
      RECT  1394400.0 655200.0 1404600.0 641400.0 ;
      RECT  1394400.0 655200.0 1404600.0 669000.0 ;
      RECT  1394400.0 682800.0 1404600.0 669000.0 ;
      RECT  1394400.0 682800.0 1404600.0 696600.0 ;
      RECT  1394400.0 710400.0 1404600.0 696600.0 ;
      RECT  1394400.0 710400.0 1404600.0 724200.0 ;
      RECT  1394400.0 738000.0 1404600.0 724200.0 ;
      RECT  1394400.0 738000.0 1404600.0 751800.0 ;
      RECT  1394400.0 765600.0 1404600.0 751800.0 ;
      RECT  1394400.0 765600.0 1404600.0 779400.0 ;
      RECT  1394400.0 793200.0 1404600.0 779400.0 ;
      RECT  1394400.0 793200.0 1404600.0 807000.0 ;
      RECT  1394400.0 820800.0 1404600.0 807000.0 ;
      RECT  1394400.0 820800.0 1404600.0 834600.0 ;
      RECT  1394400.0 848400.0 1404600.0 834600.0 ;
      RECT  1394400.0 848400.0 1404600.0 862200.0 ;
      RECT  1394400.0 876000.0 1404600.0 862200.0 ;
      RECT  1394400.0 876000.0 1404600.0 889800.0 ;
      RECT  1394400.0 903600.0 1404600.0 889800.0 ;
      RECT  1394400.0 903600.0 1404600.0 917400.0 ;
      RECT  1394400.0 931200.0 1404600.0 917400.0 ;
      RECT  1394400.0 931200.0 1404600.0 945000.0 ;
      RECT  1394400.0 958800.0 1404600.0 945000.0 ;
      RECT  1394400.0 958800.0 1404600.0 972600.0 ;
      RECT  1394400.0 986400.0 1404600.0 972600.0 ;
      RECT  1394400.0 986400.0 1404600.0 1000200.0 ;
      RECT  1394400.0 1014000.0 1404600.0 1000200.0 ;
      RECT  1394400.0 1014000.0 1404600.0 1027800.0 ;
      RECT  1394400.0 1041600.0 1404600.0 1027800.0 ;
      RECT  1394400.0 1041600.0 1404600.0 1055400.0 ;
      RECT  1394400.0 1069200.0 1404600.0 1055400.0 ;
      RECT  1394400.0 1069200.0 1404600.0 1083000.0 ;
      RECT  1394400.0 1096800.0 1404600.0 1083000.0 ;
      RECT  1394400.0 1096800.0 1404600.0 1110600.0 ;
      RECT  1394400.0 1124400.0 1404600.0 1110600.0 ;
      RECT  1394400.0 1124400.0 1404600.0 1138200.0 ;
      RECT  1394400.0 1152000.0 1404600.0 1138200.0 ;
      RECT  1394400.0 1152000.0 1404600.0 1165800.0 ;
      RECT  1394400.0 1179600.0 1404600.0 1165800.0 ;
      RECT  1394400.0 1179600.0 1404600.0 1193400.0 ;
      RECT  1394400.0 1207200.0 1404600.0 1193400.0 ;
      RECT  1394400.0 1207200.0 1404600.0 1221000.0 ;
      RECT  1394400.0 1234800.0 1404600.0 1221000.0 ;
      RECT  1394400.0 1234800.0 1404600.0 1248600.0 ;
      RECT  1394400.0 1262400.0 1404600.0 1248600.0 ;
      RECT  1394400.0 1262400.0 1404600.0 1276200.0 ;
      RECT  1394400.0 1290000.0 1404600.0 1276200.0 ;
      RECT  1394400.0 1290000.0 1404600.0 1303800.0 ;
      RECT  1394400.0 1317600.0 1404600.0 1303800.0 ;
      RECT  1394400.0 1317600.0 1404600.0 1331400.0 ;
      RECT  1394400.0 1345200.0 1404600.0 1331400.0 ;
      RECT  1394400.0 1345200.0 1404600.0 1359000.0 ;
      RECT  1394400.0 1372800.0 1404600.0 1359000.0 ;
      RECT  1394400.0 1372800.0 1404600.0 1386600.0 ;
      RECT  1394400.0 1400400.0 1404600.0 1386600.0 ;
      RECT  1394400.0 1400400.0 1404600.0 1414200.0 ;
      RECT  1394400.0 1428000.0 1404600.0 1414200.0 ;
      RECT  1394400.0 1428000.0 1404600.0 1441800.0 ;
      RECT  1394400.0 1455600.0 1404600.0 1441800.0 ;
      RECT  1394400.0 1455600.0 1404600.0 1469400.0 ;
      RECT  1394400.0 1483200.0 1404600.0 1469400.0 ;
      RECT  1394400.0 1483200.0 1404600.0 1497000.0 ;
      RECT  1394400.0 1510800.0 1404600.0 1497000.0 ;
      RECT  1394400.0 1510800.0 1404600.0 1524600.0 ;
      RECT  1394400.0 1538400.0 1404600.0 1524600.0 ;
      RECT  1394400.0 1538400.0 1404600.0 1552200.0 ;
      RECT  1394400.0 1566000.0 1404600.0 1552200.0 ;
      RECT  1394400.0 1566000.0 1404600.0 1579800.0 ;
      RECT  1394400.0 1593600.0 1404600.0 1579800.0 ;
      RECT  1394400.0 1593600.0 1404600.0 1607400.0 ;
      RECT  1394400.0 1621200.0 1404600.0 1607400.0 ;
      RECT  1394400.0 1621200.0 1404600.0 1635000.0 ;
      RECT  1394400.0 1648800.0 1404600.0 1635000.0 ;
      RECT  1394400.0 1648800.0 1404600.0 1662600.0 ;
      RECT  1394400.0 1676400.0 1404600.0 1662600.0 ;
      RECT  1394400.0 1676400.0 1404600.0 1690200.0 ;
      RECT  1394400.0 1704000.0 1404600.0 1690200.0 ;
      RECT  1394400.0 1704000.0 1404600.0 1717800.0 ;
      RECT  1394400.0 1731600.0 1404600.0 1717800.0 ;
      RECT  1394400.0 1731600.0 1404600.0 1745400.0 ;
      RECT  1394400.0 1759200.0 1404600.0 1745400.0 ;
      RECT  1394400.0 1759200.0 1404600.0 1773000.0 ;
      RECT  1394400.0 1786800.0 1404600.0 1773000.0 ;
      RECT  1394400.0 1786800.0 1404600.0 1800600.0 ;
      RECT  1394400.0 1814400.0 1404600.0 1800600.0 ;
      RECT  1394400.0 1814400.0 1404600.0 1828200.0 ;
      RECT  1394400.0 1842000.0 1404600.0 1828200.0 ;
      RECT  1394400.0 1842000.0 1404600.0 1855800.0 ;
      RECT  1394400.0 1869600.0 1404600.0 1855800.0 ;
      RECT  1394400.0 1869600.0 1404600.0 1883400.0 ;
      RECT  1394400.0 1897200.0 1404600.0 1883400.0 ;
      RECT  1394400.0 1897200.0 1404600.0 1911000.0 ;
      RECT  1394400.0 1924800.0 1404600.0 1911000.0 ;
      RECT  1394400.0 1924800.0 1404600.0 1938600.0 ;
      RECT  1394400.0 1952400.0 1404600.0 1938600.0 ;
      RECT  1394400.0 1952400.0 1404600.0 1966200.0 ;
      RECT  1394400.0 1980000.0 1404600.0 1966200.0 ;
      RECT  1394400.0 1980000.0 1404600.0 1993800.0 ;
      RECT  1394400.0 2007600.0 1404600.0 1993800.0 ;
      RECT  1394400.0 2007600.0 1404600.0 2021400.0 ;
      RECT  1394400.0 2035200.0 1404600.0 2021400.0 ;
      RECT  1394400.0 2035200.0 1404600.0 2049000.0 ;
      RECT  1394400.0 2062800.0 1404600.0 2049000.0 ;
      RECT  1394400.0 2062800.0 1404600.0 2076600.0 ;
      RECT  1394400.0 2090400.0 1404600.0 2076600.0 ;
      RECT  1394400.0 2090400.0 1404600.0 2104200.0 ;
      RECT  1394400.0 2118000.0 1404600.0 2104200.0 ;
      RECT  1394400.0 2118000.0 1404600.0 2131800.0 ;
      RECT  1394400.0 2145600.0 1404600.0 2131800.0 ;
      RECT  1404600.0 379200.0 1414800.0 393000.0 ;
      RECT  1404600.0 406800.0 1414800.0 393000.0 ;
      RECT  1404600.0 406800.0 1414800.0 420600.0 ;
      RECT  1404600.0 434400.0 1414800.0 420600.0 ;
      RECT  1404600.0 434400.0 1414800.0 448200.0 ;
      RECT  1404600.0 462000.0 1414800.0 448200.0 ;
      RECT  1404600.0 462000.0 1414800.0 475800.0 ;
      RECT  1404600.0 489600.0 1414800.0 475800.0 ;
      RECT  1404600.0 489600.0 1414800.0 503400.0 ;
      RECT  1404600.0 517200.0 1414800.0 503400.0 ;
      RECT  1404600.0 517200.0 1414800.0 531000.0 ;
      RECT  1404600.0 544800.0 1414800.0 531000.0 ;
      RECT  1404600.0 544800.0 1414800.0 558600.0 ;
      RECT  1404600.0 572400.0 1414800.0 558600.0 ;
      RECT  1404600.0 572400.0 1414800.0 586200.0 ;
      RECT  1404600.0 600000.0 1414800.0 586200.0 ;
      RECT  1404600.0 600000.0 1414800.0 613800.0 ;
      RECT  1404600.0 627600.0 1414800.0 613800.0 ;
      RECT  1404600.0 627600.0 1414800.0 641400.0 ;
      RECT  1404600.0 655200.0 1414800.0 641400.0 ;
      RECT  1404600.0 655200.0 1414800.0 669000.0 ;
      RECT  1404600.0 682800.0 1414800.0 669000.0 ;
      RECT  1404600.0 682800.0 1414800.0 696600.0 ;
      RECT  1404600.0 710400.0 1414800.0 696600.0 ;
      RECT  1404600.0 710400.0 1414800.0 724200.0 ;
      RECT  1404600.0 738000.0 1414800.0 724200.0 ;
      RECT  1404600.0 738000.0 1414800.0 751800.0 ;
      RECT  1404600.0 765600.0 1414800.0 751800.0 ;
      RECT  1404600.0 765600.0 1414800.0 779400.0 ;
      RECT  1404600.0 793200.0 1414800.0 779400.0 ;
      RECT  1404600.0 793200.0 1414800.0 807000.0 ;
      RECT  1404600.0 820800.0 1414800.0 807000.0 ;
      RECT  1404600.0 820800.0 1414800.0 834600.0 ;
      RECT  1404600.0 848400.0 1414800.0 834600.0 ;
      RECT  1404600.0 848400.0 1414800.0 862200.0 ;
      RECT  1404600.0 876000.0 1414800.0 862200.0 ;
      RECT  1404600.0 876000.0 1414800.0 889800.0 ;
      RECT  1404600.0 903600.0 1414800.0 889800.0 ;
      RECT  1404600.0 903600.0 1414800.0 917400.0 ;
      RECT  1404600.0 931200.0 1414800.0 917400.0 ;
      RECT  1404600.0 931200.0 1414800.0 945000.0 ;
      RECT  1404600.0 958800.0 1414800.0 945000.0 ;
      RECT  1404600.0 958800.0 1414800.0 972600.0 ;
      RECT  1404600.0 986400.0 1414800.0 972600.0 ;
      RECT  1404600.0 986400.0 1414800.0 1000200.0 ;
      RECT  1404600.0 1014000.0 1414800.0 1000200.0 ;
      RECT  1404600.0 1014000.0 1414800.0 1027800.0 ;
      RECT  1404600.0 1041600.0 1414800.0 1027800.0 ;
      RECT  1404600.0 1041600.0 1414800.0 1055400.0 ;
      RECT  1404600.0 1069200.0 1414800.0 1055400.0 ;
      RECT  1404600.0 1069200.0 1414800.0 1083000.0 ;
      RECT  1404600.0 1096800.0 1414800.0 1083000.0 ;
      RECT  1404600.0 1096800.0 1414800.0 1110600.0 ;
      RECT  1404600.0 1124400.0 1414800.0 1110600.0 ;
      RECT  1404600.0 1124400.0 1414800.0 1138200.0 ;
      RECT  1404600.0 1152000.0 1414800.0 1138200.0 ;
      RECT  1404600.0 1152000.0 1414800.0 1165800.0 ;
      RECT  1404600.0 1179600.0 1414800.0 1165800.0 ;
      RECT  1404600.0 1179600.0 1414800.0 1193400.0 ;
      RECT  1404600.0 1207200.0 1414800.0 1193400.0 ;
      RECT  1404600.0 1207200.0 1414800.0 1221000.0 ;
      RECT  1404600.0 1234800.0 1414800.0 1221000.0 ;
      RECT  1404600.0 1234800.0 1414800.0 1248600.0 ;
      RECT  1404600.0 1262400.0 1414800.0 1248600.0 ;
      RECT  1404600.0 1262400.0 1414800.0 1276200.0 ;
      RECT  1404600.0 1290000.0 1414800.0 1276200.0 ;
      RECT  1404600.0 1290000.0 1414800.0 1303800.0 ;
      RECT  1404600.0 1317600.0 1414800.0 1303800.0 ;
      RECT  1404600.0 1317600.0 1414800.0 1331400.0 ;
      RECT  1404600.0 1345200.0 1414800.0 1331400.0 ;
      RECT  1404600.0 1345200.0 1414800.0 1359000.0 ;
      RECT  1404600.0 1372800.0 1414800.0 1359000.0 ;
      RECT  1404600.0 1372800.0 1414800.0 1386600.0 ;
      RECT  1404600.0 1400400.0 1414800.0 1386600.0 ;
      RECT  1404600.0 1400400.0 1414800.0 1414200.0 ;
      RECT  1404600.0 1428000.0 1414800.0 1414200.0 ;
      RECT  1404600.0 1428000.0 1414800.0 1441800.0 ;
      RECT  1404600.0 1455600.0 1414800.0 1441800.0 ;
      RECT  1404600.0 1455600.0 1414800.0 1469400.0 ;
      RECT  1404600.0 1483200.0 1414800.0 1469400.0 ;
      RECT  1404600.0 1483200.0 1414800.0 1497000.0 ;
      RECT  1404600.0 1510800.0 1414800.0 1497000.0 ;
      RECT  1404600.0 1510800.0 1414800.0 1524600.0 ;
      RECT  1404600.0 1538400.0 1414800.0 1524600.0 ;
      RECT  1404600.0 1538400.0 1414800.0 1552200.0 ;
      RECT  1404600.0 1566000.0 1414800.0 1552200.0 ;
      RECT  1404600.0 1566000.0 1414800.0 1579800.0 ;
      RECT  1404600.0 1593600.0 1414800.0 1579800.0 ;
      RECT  1404600.0 1593600.0 1414800.0 1607400.0 ;
      RECT  1404600.0 1621200.0 1414800.0 1607400.0 ;
      RECT  1404600.0 1621200.0 1414800.0 1635000.0 ;
      RECT  1404600.0 1648800.0 1414800.0 1635000.0 ;
      RECT  1404600.0 1648800.0 1414800.0 1662600.0 ;
      RECT  1404600.0 1676400.0 1414800.0 1662600.0 ;
      RECT  1404600.0 1676400.0 1414800.0 1690200.0 ;
      RECT  1404600.0 1704000.0 1414800.0 1690200.0 ;
      RECT  1404600.0 1704000.0 1414800.0 1717800.0 ;
      RECT  1404600.0 1731600.0 1414800.0 1717800.0 ;
      RECT  1404600.0 1731600.0 1414800.0 1745400.0 ;
      RECT  1404600.0 1759200.0 1414800.0 1745400.0 ;
      RECT  1404600.0 1759200.0 1414800.0 1773000.0 ;
      RECT  1404600.0 1786800.0 1414800.0 1773000.0 ;
      RECT  1404600.0 1786800.0 1414800.0 1800600.0 ;
      RECT  1404600.0 1814400.0 1414800.0 1800600.0 ;
      RECT  1404600.0 1814400.0 1414800.0 1828200.0 ;
      RECT  1404600.0 1842000.0 1414800.0 1828200.0 ;
      RECT  1404600.0 1842000.0 1414800.0 1855800.0 ;
      RECT  1404600.0 1869600.0 1414800.0 1855800.0 ;
      RECT  1404600.0 1869600.0 1414800.0 1883400.0 ;
      RECT  1404600.0 1897200.0 1414800.0 1883400.0 ;
      RECT  1404600.0 1897200.0 1414800.0 1911000.0 ;
      RECT  1404600.0 1924800.0 1414800.0 1911000.0 ;
      RECT  1404600.0 1924800.0 1414800.0 1938600.0 ;
      RECT  1404600.0 1952400.0 1414800.0 1938600.0 ;
      RECT  1404600.0 1952400.0 1414800.0 1966200.0 ;
      RECT  1404600.0 1980000.0 1414800.0 1966200.0 ;
      RECT  1404600.0 1980000.0 1414800.0 1993800.0 ;
      RECT  1404600.0 2007600.0 1414800.0 1993800.0 ;
      RECT  1404600.0 2007600.0 1414800.0 2021400.0 ;
      RECT  1404600.0 2035200.0 1414800.0 2021400.0 ;
      RECT  1404600.0 2035200.0 1414800.0 2049000.0 ;
      RECT  1404600.0 2062800.0 1414800.0 2049000.0 ;
      RECT  1404600.0 2062800.0 1414800.0 2076600.0 ;
      RECT  1404600.0 2090400.0 1414800.0 2076600.0 ;
      RECT  1404600.0 2090400.0 1414800.0 2104200.0 ;
      RECT  1404600.0 2118000.0 1414800.0 2104200.0 ;
      RECT  1404600.0 2118000.0 1414800.0 2131800.0 ;
      RECT  1404600.0 2145600.0 1414800.0 2131800.0 ;
      RECT  1414800.0 379200.0 1425000.0 393000.0 ;
      RECT  1414800.0 406800.0 1425000.0 393000.0 ;
      RECT  1414800.0 406800.0 1425000.0 420600.0 ;
      RECT  1414800.0 434400.0 1425000.0 420600.0 ;
      RECT  1414800.0 434400.0 1425000.0 448200.0 ;
      RECT  1414800.0 462000.0 1425000.0 448200.0 ;
      RECT  1414800.0 462000.0 1425000.0 475800.0 ;
      RECT  1414800.0 489600.0 1425000.0 475800.0 ;
      RECT  1414800.0 489600.0 1425000.0 503400.0 ;
      RECT  1414800.0 517200.0 1425000.0 503400.0 ;
      RECT  1414800.0 517200.0 1425000.0 531000.0 ;
      RECT  1414800.0 544800.0 1425000.0 531000.0 ;
      RECT  1414800.0 544800.0 1425000.0 558600.0 ;
      RECT  1414800.0 572400.0 1425000.0 558600.0 ;
      RECT  1414800.0 572400.0 1425000.0 586200.0 ;
      RECT  1414800.0 600000.0 1425000.0 586200.0 ;
      RECT  1414800.0 600000.0 1425000.0 613800.0 ;
      RECT  1414800.0 627600.0 1425000.0 613800.0 ;
      RECT  1414800.0 627600.0 1425000.0 641400.0 ;
      RECT  1414800.0 655200.0 1425000.0 641400.0 ;
      RECT  1414800.0 655200.0 1425000.0 669000.0 ;
      RECT  1414800.0 682800.0 1425000.0 669000.0 ;
      RECT  1414800.0 682800.0 1425000.0 696600.0 ;
      RECT  1414800.0 710400.0 1425000.0 696600.0 ;
      RECT  1414800.0 710400.0 1425000.0 724200.0 ;
      RECT  1414800.0 738000.0 1425000.0 724200.0 ;
      RECT  1414800.0 738000.0 1425000.0 751800.0 ;
      RECT  1414800.0 765600.0 1425000.0 751800.0 ;
      RECT  1414800.0 765600.0 1425000.0 779400.0 ;
      RECT  1414800.0 793200.0 1425000.0 779400.0 ;
      RECT  1414800.0 793200.0 1425000.0 807000.0 ;
      RECT  1414800.0 820800.0 1425000.0 807000.0 ;
      RECT  1414800.0 820800.0 1425000.0 834600.0 ;
      RECT  1414800.0 848400.0 1425000.0 834600.0 ;
      RECT  1414800.0 848400.0 1425000.0 862200.0 ;
      RECT  1414800.0 876000.0 1425000.0 862200.0 ;
      RECT  1414800.0 876000.0 1425000.0 889800.0 ;
      RECT  1414800.0 903600.0 1425000.0 889800.0 ;
      RECT  1414800.0 903600.0 1425000.0 917400.0 ;
      RECT  1414800.0 931200.0 1425000.0 917400.0 ;
      RECT  1414800.0 931200.0 1425000.0 945000.0 ;
      RECT  1414800.0 958800.0 1425000.0 945000.0 ;
      RECT  1414800.0 958800.0 1425000.0 972600.0 ;
      RECT  1414800.0 986400.0 1425000.0 972600.0 ;
      RECT  1414800.0 986400.0 1425000.0 1000200.0 ;
      RECT  1414800.0 1014000.0 1425000.0 1000200.0 ;
      RECT  1414800.0 1014000.0 1425000.0 1027800.0 ;
      RECT  1414800.0 1041600.0 1425000.0 1027800.0 ;
      RECT  1414800.0 1041600.0 1425000.0 1055400.0 ;
      RECT  1414800.0 1069200.0 1425000.0 1055400.0 ;
      RECT  1414800.0 1069200.0 1425000.0 1083000.0 ;
      RECT  1414800.0 1096800.0 1425000.0 1083000.0 ;
      RECT  1414800.0 1096800.0 1425000.0 1110600.0 ;
      RECT  1414800.0 1124400.0 1425000.0 1110600.0 ;
      RECT  1414800.0 1124400.0 1425000.0 1138200.0 ;
      RECT  1414800.0 1152000.0 1425000.0 1138200.0 ;
      RECT  1414800.0 1152000.0 1425000.0 1165800.0 ;
      RECT  1414800.0 1179600.0 1425000.0 1165800.0 ;
      RECT  1414800.0 1179600.0 1425000.0 1193400.0 ;
      RECT  1414800.0 1207200.0 1425000.0 1193400.0 ;
      RECT  1414800.0 1207200.0 1425000.0 1221000.0 ;
      RECT  1414800.0 1234800.0 1425000.0 1221000.0 ;
      RECT  1414800.0 1234800.0 1425000.0 1248600.0 ;
      RECT  1414800.0 1262400.0 1425000.0 1248600.0 ;
      RECT  1414800.0 1262400.0 1425000.0 1276200.0 ;
      RECT  1414800.0 1290000.0 1425000.0 1276200.0 ;
      RECT  1414800.0 1290000.0 1425000.0 1303800.0 ;
      RECT  1414800.0 1317600.0 1425000.0 1303800.0 ;
      RECT  1414800.0 1317600.0 1425000.0 1331400.0 ;
      RECT  1414800.0 1345200.0 1425000.0 1331400.0 ;
      RECT  1414800.0 1345200.0 1425000.0 1359000.0 ;
      RECT  1414800.0 1372800.0 1425000.0 1359000.0 ;
      RECT  1414800.0 1372800.0 1425000.0 1386600.0 ;
      RECT  1414800.0 1400400.0 1425000.0 1386600.0 ;
      RECT  1414800.0 1400400.0 1425000.0 1414200.0 ;
      RECT  1414800.0 1428000.0 1425000.0 1414200.0 ;
      RECT  1414800.0 1428000.0 1425000.0 1441800.0 ;
      RECT  1414800.0 1455600.0 1425000.0 1441800.0 ;
      RECT  1414800.0 1455600.0 1425000.0 1469400.0 ;
      RECT  1414800.0 1483200.0 1425000.0 1469400.0 ;
      RECT  1414800.0 1483200.0 1425000.0 1497000.0 ;
      RECT  1414800.0 1510800.0 1425000.0 1497000.0 ;
      RECT  1414800.0 1510800.0 1425000.0 1524600.0 ;
      RECT  1414800.0 1538400.0 1425000.0 1524600.0 ;
      RECT  1414800.0 1538400.0 1425000.0 1552200.0 ;
      RECT  1414800.0 1566000.0 1425000.0 1552200.0 ;
      RECT  1414800.0 1566000.0 1425000.0 1579800.0 ;
      RECT  1414800.0 1593600.0 1425000.0 1579800.0 ;
      RECT  1414800.0 1593600.0 1425000.0 1607400.0 ;
      RECT  1414800.0 1621200.0 1425000.0 1607400.0 ;
      RECT  1414800.0 1621200.0 1425000.0 1635000.0 ;
      RECT  1414800.0 1648800.0 1425000.0 1635000.0 ;
      RECT  1414800.0 1648800.0 1425000.0 1662600.0 ;
      RECT  1414800.0 1676400.0 1425000.0 1662600.0 ;
      RECT  1414800.0 1676400.0 1425000.0 1690200.0 ;
      RECT  1414800.0 1704000.0 1425000.0 1690200.0 ;
      RECT  1414800.0 1704000.0 1425000.0 1717800.0 ;
      RECT  1414800.0 1731600.0 1425000.0 1717800.0 ;
      RECT  1414800.0 1731600.0 1425000.0 1745400.0 ;
      RECT  1414800.0 1759200.0 1425000.0 1745400.0 ;
      RECT  1414800.0 1759200.0 1425000.0 1773000.0 ;
      RECT  1414800.0 1786800.0 1425000.0 1773000.0 ;
      RECT  1414800.0 1786800.0 1425000.0 1800600.0 ;
      RECT  1414800.0 1814400.0 1425000.0 1800600.0 ;
      RECT  1414800.0 1814400.0 1425000.0 1828200.0 ;
      RECT  1414800.0 1842000.0 1425000.0 1828200.0 ;
      RECT  1414800.0 1842000.0 1425000.0 1855800.0 ;
      RECT  1414800.0 1869600.0 1425000.0 1855800.0 ;
      RECT  1414800.0 1869600.0 1425000.0 1883400.0 ;
      RECT  1414800.0 1897200.0 1425000.0 1883400.0 ;
      RECT  1414800.0 1897200.0 1425000.0 1911000.0 ;
      RECT  1414800.0 1924800.0 1425000.0 1911000.0 ;
      RECT  1414800.0 1924800.0 1425000.0 1938600.0 ;
      RECT  1414800.0 1952400.0 1425000.0 1938600.0 ;
      RECT  1414800.0 1952400.0 1425000.0 1966200.0 ;
      RECT  1414800.0 1980000.0 1425000.0 1966200.0 ;
      RECT  1414800.0 1980000.0 1425000.0 1993800.0 ;
      RECT  1414800.0 2007600.0 1425000.0 1993800.0 ;
      RECT  1414800.0 2007600.0 1425000.0 2021400.0 ;
      RECT  1414800.0 2035200.0 1425000.0 2021400.0 ;
      RECT  1414800.0 2035200.0 1425000.0 2049000.0 ;
      RECT  1414800.0 2062800.0 1425000.0 2049000.0 ;
      RECT  1414800.0 2062800.0 1425000.0 2076600.0 ;
      RECT  1414800.0 2090400.0 1425000.0 2076600.0 ;
      RECT  1414800.0 2090400.0 1425000.0 2104200.0 ;
      RECT  1414800.0 2118000.0 1425000.0 2104200.0 ;
      RECT  1414800.0 2118000.0 1425000.0 2131800.0 ;
      RECT  1414800.0 2145600.0 1425000.0 2131800.0 ;
      RECT  1425000.0 379200.0 1435200.0 393000.0 ;
      RECT  1425000.0 406800.0 1435200.0 393000.0 ;
      RECT  1425000.0 406800.0 1435200.0 420600.0 ;
      RECT  1425000.0 434400.0 1435200.0 420600.0 ;
      RECT  1425000.0 434400.0 1435200.0 448200.0 ;
      RECT  1425000.0 462000.0 1435200.0 448200.0 ;
      RECT  1425000.0 462000.0 1435200.0 475800.0 ;
      RECT  1425000.0 489600.0 1435200.0 475800.0 ;
      RECT  1425000.0 489600.0 1435200.0 503400.0 ;
      RECT  1425000.0 517200.0 1435200.0 503400.0 ;
      RECT  1425000.0 517200.0 1435200.0 531000.0 ;
      RECT  1425000.0 544800.0 1435200.0 531000.0 ;
      RECT  1425000.0 544800.0 1435200.0 558600.0 ;
      RECT  1425000.0 572400.0 1435200.0 558600.0 ;
      RECT  1425000.0 572400.0 1435200.0 586200.0 ;
      RECT  1425000.0 600000.0 1435200.0 586200.0 ;
      RECT  1425000.0 600000.0 1435200.0 613800.0 ;
      RECT  1425000.0 627600.0 1435200.0 613800.0 ;
      RECT  1425000.0 627600.0 1435200.0 641400.0 ;
      RECT  1425000.0 655200.0 1435200.0 641400.0 ;
      RECT  1425000.0 655200.0 1435200.0 669000.0 ;
      RECT  1425000.0 682800.0 1435200.0 669000.0 ;
      RECT  1425000.0 682800.0 1435200.0 696600.0 ;
      RECT  1425000.0 710400.0 1435200.0 696600.0 ;
      RECT  1425000.0 710400.0 1435200.0 724200.0 ;
      RECT  1425000.0 738000.0 1435200.0 724200.0 ;
      RECT  1425000.0 738000.0 1435200.0 751800.0 ;
      RECT  1425000.0 765600.0 1435200.0 751800.0 ;
      RECT  1425000.0 765600.0 1435200.0 779400.0 ;
      RECT  1425000.0 793200.0 1435200.0 779400.0 ;
      RECT  1425000.0 793200.0 1435200.0 807000.0 ;
      RECT  1425000.0 820800.0 1435200.0 807000.0 ;
      RECT  1425000.0 820800.0 1435200.0 834600.0 ;
      RECT  1425000.0 848400.0 1435200.0 834600.0 ;
      RECT  1425000.0 848400.0 1435200.0 862200.0 ;
      RECT  1425000.0 876000.0 1435200.0 862200.0 ;
      RECT  1425000.0 876000.0 1435200.0 889800.0 ;
      RECT  1425000.0 903600.0 1435200.0 889800.0 ;
      RECT  1425000.0 903600.0 1435200.0 917400.0 ;
      RECT  1425000.0 931200.0 1435200.0 917400.0 ;
      RECT  1425000.0 931200.0 1435200.0 945000.0 ;
      RECT  1425000.0 958800.0 1435200.0 945000.0 ;
      RECT  1425000.0 958800.0 1435200.0 972600.0 ;
      RECT  1425000.0 986400.0 1435200.0 972600.0 ;
      RECT  1425000.0 986400.0 1435200.0 1000200.0 ;
      RECT  1425000.0 1014000.0 1435200.0 1000200.0 ;
      RECT  1425000.0 1014000.0 1435200.0 1027800.0 ;
      RECT  1425000.0 1041600.0 1435200.0 1027800.0 ;
      RECT  1425000.0 1041600.0 1435200.0 1055400.0 ;
      RECT  1425000.0 1069200.0 1435200.0 1055400.0 ;
      RECT  1425000.0 1069200.0 1435200.0 1083000.0 ;
      RECT  1425000.0 1096800.0 1435200.0 1083000.0 ;
      RECT  1425000.0 1096800.0 1435200.0 1110600.0 ;
      RECT  1425000.0 1124400.0 1435200.0 1110600.0 ;
      RECT  1425000.0 1124400.0 1435200.0 1138200.0 ;
      RECT  1425000.0 1152000.0 1435200.0 1138200.0 ;
      RECT  1425000.0 1152000.0 1435200.0 1165800.0 ;
      RECT  1425000.0 1179600.0 1435200.0 1165800.0 ;
      RECT  1425000.0 1179600.0 1435200.0 1193400.0 ;
      RECT  1425000.0 1207200.0 1435200.0 1193400.0 ;
      RECT  1425000.0 1207200.0 1435200.0 1221000.0 ;
      RECT  1425000.0 1234800.0 1435200.0 1221000.0 ;
      RECT  1425000.0 1234800.0 1435200.0 1248600.0 ;
      RECT  1425000.0 1262400.0 1435200.0 1248600.0 ;
      RECT  1425000.0 1262400.0 1435200.0 1276200.0 ;
      RECT  1425000.0 1290000.0 1435200.0 1276200.0 ;
      RECT  1425000.0 1290000.0 1435200.0 1303800.0 ;
      RECT  1425000.0 1317600.0 1435200.0 1303800.0 ;
      RECT  1425000.0 1317600.0 1435200.0 1331400.0 ;
      RECT  1425000.0 1345200.0 1435200.0 1331400.0 ;
      RECT  1425000.0 1345200.0 1435200.0 1359000.0 ;
      RECT  1425000.0 1372800.0 1435200.0 1359000.0 ;
      RECT  1425000.0 1372800.0 1435200.0 1386600.0 ;
      RECT  1425000.0 1400400.0 1435200.0 1386600.0 ;
      RECT  1425000.0 1400400.0 1435200.0 1414200.0 ;
      RECT  1425000.0 1428000.0 1435200.0 1414200.0 ;
      RECT  1425000.0 1428000.0 1435200.0 1441800.0 ;
      RECT  1425000.0 1455600.0 1435200.0 1441800.0 ;
      RECT  1425000.0 1455600.0 1435200.0 1469400.0 ;
      RECT  1425000.0 1483200.0 1435200.0 1469400.0 ;
      RECT  1425000.0 1483200.0 1435200.0 1497000.0 ;
      RECT  1425000.0 1510800.0 1435200.0 1497000.0 ;
      RECT  1425000.0 1510800.0 1435200.0 1524600.0 ;
      RECT  1425000.0 1538400.0 1435200.0 1524600.0 ;
      RECT  1425000.0 1538400.0 1435200.0 1552200.0 ;
      RECT  1425000.0 1566000.0 1435200.0 1552200.0 ;
      RECT  1425000.0 1566000.0 1435200.0 1579800.0 ;
      RECT  1425000.0 1593600.0 1435200.0 1579800.0 ;
      RECT  1425000.0 1593600.0 1435200.0 1607400.0 ;
      RECT  1425000.0 1621200.0 1435200.0 1607400.0 ;
      RECT  1425000.0 1621200.0 1435200.0 1635000.0 ;
      RECT  1425000.0 1648800.0 1435200.0 1635000.0 ;
      RECT  1425000.0 1648800.0 1435200.0 1662600.0 ;
      RECT  1425000.0 1676400.0 1435200.0 1662600.0 ;
      RECT  1425000.0 1676400.0 1435200.0 1690200.0 ;
      RECT  1425000.0 1704000.0 1435200.0 1690200.0 ;
      RECT  1425000.0 1704000.0 1435200.0 1717800.0 ;
      RECT  1425000.0 1731600.0 1435200.0 1717800.0 ;
      RECT  1425000.0 1731600.0 1435200.0 1745400.0 ;
      RECT  1425000.0 1759200.0 1435200.0 1745400.0 ;
      RECT  1425000.0 1759200.0 1435200.0 1773000.0 ;
      RECT  1425000.0 1786800.0 1435200.0 1773000.0 ;
      RECT  1425000.0 1786800.0 1435200.0 1800600.0 ;
      RECT  1425000.0 1814400.0 1435200.0 1800600.0 ;
      RECT  1425000.0 1814400.0 1435200.0 1828200.0 ;
      RECT  1425000.0 1842000.0 1435200.0 1828200.0 ;
      RECT  1425000.0 1842000.0 1435200.0 1855800.0 ;
      RECT  1425000.0 1869600.0 1435200.0 1855800.0 ;
      RECT  1425000.0 1869600.0 1435200.0 1883400.0 ;
      RECT  1425000.0 1897200.0 1435200.0 1883400.0 ;
      RECT  1425000.0 1897200.0 1435200.0 1911000.0 ;
      RECT  1425000.0 1924800.0 1435200.0 1911000.0 ;
      RECT  1425000.0 1924800.0 1435200.0 1938600.0 ;
      RECT  1425000.0 1952400.0 1435200.0 1938600.0 ;
      RECT  1425000.0 1952400.0 1435200.0 1966200.0 ;
      RECT  1425000.0 1980000.0 1435200.0 1966200.0 ;
      RECT  1425000.0 1980000.0 1435200.0 1993800.0 ;
      RECT  1425000.0 2007600.0 1435200.0 1993800.0 ;
      RECT  1425000.0 2007600.0 1435200.0 2021400.0 ;
      RECT  1425000.0 2035200.0 1435200.0 2021400.0 ;
      RECT  1425000.0 2035200.0 1435200.0 2049000.0 ;
      RECT  1425000.0 2062800.0 1435200.0 2049000.0 ;
      RECT  1425000.0 2062800.0 1435200.0 2076600.0 ;
      RECT  1425000.0 2090400.0 1435200.0 2076600.0 ;
      RECT  1425000.0 2090400.0 1435200.0 2104200.0 ;
      RECT  1425000.0 2118000.0 1435200.0 2104200.0 ;
      RECT  1425000.0 2118000.0 1435200.0 2131800.0 ;
      RECT  1425000.0 2145600.0 1435200.0 2131800.0 ;
      RECT  1435200.0 379200.0 1445400.0 393000.0 ;
      RECT  1435200.0 406800.0 1445400.0 393000.0 ;
      RECT  1435200.0 406800.0 1445400.0 420600.0 ;
      RECT  1435200.0 434400.0 1445400.0 420600.0 ;
      RECT  1435200.0 434400.0 1445400.0 448200.0 ;
      RECT  1435200.0 462000.0 1445400.0 448200.0 ;
      RECT  1435200.0 462000.0 1445400.0 475800.0 ;
      RECT  1435200.0 489600.0 1445400.0 475800.0 ;
      RECT  1435200.0 489600.0 1445400.0 503400.0 ;
      RECT  1435200.0 517200.0 1445400.0 503400.0 ;
      RECT  1435200.0 517200.0 1445400.0 531000.0 ;
      RECT  1435200.0 544800.0 1445400.0 531000.0 ;
      RECT  1435200.0 544800.0 1445400.0 558600.0 ;
      RECT  1435200.0 572400.0 1445400.0 558600.0 ;
      RECT  1435200.0 572400.0 1445400.0 586200.0 ;
      RECT  1435200.0 600000.0 1445400.0 586200.0 ;
      RECT  1435200.0 600000.0 1445400.0 613800.0 ;
      RECT  1435200.0 627600.0 1445400.0 613800.0 ;
      RECT  1435200.0 627600.0 1445400.0 641400.0 ;
      RECT  1435200.0 655200.0 1445400.0 641400.0 ;
      RECT  1435200.0 655200.0 1445400.0 669000.0 ;
      RECT  1435200.0 682800.0 1445400.0 669000.0 ;
      RECT  1435200.0 682800.0 1445400.0 696600.0 ;
      RECT  1435200.0 710400.0 1445400.0 696600.0 ;
      RECT  1435200.0 710400.0 1445400.0 724200.0 ;
      RECT  1435200.0 738000.0 1445400.0 724200.0 ;
      RECT  1435200.0 738000.0 1445400.0 751800.0 ;
      RECT  1435200.0 765600.0 1445400.0 751800.0 ;
      RECT  1435200.0 765600.0 1445400.0 779400.0 ;
      RECT  1435200.0 793200.0 1445400.0 779400.0 ;
      RECT  1435200.0 793200.0 1445400.0 807000.0 ;
      RECT  1435200.0 820800.0 1445400.0 807000.0 ;
      RECT  1435200.0 820800.0 1445400.0 834600.0 ;
      RECT  1435200.0 848400.0 1445400.0 834600.0 ;
      RECT  1435200.0 848400.0 1445400.0 862200.0 ;
      RECT  1435200.0 876000.0 1445400.0 862200.0 ;
      RECT  1435200.0 876000.0 1445400.0 889800.0 ;
      RECT  1435200.0 903600.0 1445400.0 889800.0 ;
      RECT  1435200.0 903600.0 1445400.0 917400.0 ;
      RECT  1435200.0 931200.0 1445400.0 917400.0 ;
      RECT  1435200.0 931200.0 1445400.0 945000.0 ;
      RECT  1435200.0 958800.0 1445400.0 945000.0 ;
      RECT  1435200.0 958800.0 1445400.0 972600.0 ;
      RECT  1435200.0 986400.0 1445400.0 972600.0 ;
      RECT  1435200.0 986400.0 1445400.0 1000200.0 ;
      RECT  1435200.0 1014000.0 1445400.0 1000200.0 ;
      RECT  1435200.0 1014000.0 1445400.0 1027800.0 ;
      RECT  1435200.0 1041600.0 1445400.0 1027800.0 ;
      RECT  1435200.0 1041600.0 1445400.0 1055400.0 ;
      RECT  1435200.0 1069200.0 1445400.0 1055400.0 ;
      RECT  1435200.0 1069200.0 1445400.0 1083000.0 ;
      RECT  1435200.0 1096800.0 1445400.0 1083000.0 ;
      RECT  1435200.0 1096800.0 1445400.0 1110600.0 ;
      RECT  1435200.0 1124400.0 1445400.0 1110600.0 ;
      RECT  1435200.0 1124400.0 1445400.0 1138200.0 ;
      RECT  1435200.0 1152000.0 1445400.0 1138200.0 ;
      RECT  1435200.0 1152000.0 1445400.0 1165800.0 ;
      RECT  1435200.0 1179600.0 1445400.0 1165800.0 ;
      RECT  1435200.0 1179600.0 1445400.0 1193400.0 ;
      RECT  1435200.0 1207200.0 1445400.0 1193400.0 ;
      RECT  1435200.0 1207200.0 1445400.0 1221000.0 ;
      RECT  1435200.0 1234800.0 1445400.0 1221000.0 ;
      RECT  1435200.0 1234800.0 1445400.0 1248600.0 ;
      RECT  1435200.0 1262400.0 1445400.0 1248600.0 ;
      RECT  1435200.0 1262400.0 1445400.0 1276200.0 ;
      RECT  1435200.0 1290000.0 1445400.0 1276200.0 ;
      RECT  1435200.0 1290000.0 1445400.0 1303800.0 ;
      RECT  1435200.0 1317600.0 1445400.0 1303800.0 ;
      RECT  1435200.0 1317600.0 1445400.0 1331400.0 ;
      RECT  1435200.0 1345200.0 1445400.0 1331400.0 ;
      RECT  1435200.0 1345200.0 1445400.0 1359000.0 ;
      RECT  1435200.0 1372800.0 1445400.0 1359000.0 ;
      RECT  1435200.0 1372800.0 1445400.0 1386600.0 ;
      RECT  1435200.0 1400400.0 1445400.0 1386600.0 ;
      RECT  1435200.0 1400400.0 1445400.0 1414200.0 ;
      RECT  1435200.0 1428000.0 1445400.0 1414200.0 ;
      RECT  1435200.0 1428000.0 1445400.0 1441800.0 ;
      RECT  1435200.0 1455600.0 1445400.0 1441800.0 ;
      RECT  1435200.0 1455600.0 1445400.0 1469400.0 ;
      RECT  1435200.0 1483200.0 1445400.0 1469400.0 ;
      RECT  1435200.0 1483200.0 1445400.0 1497000.0 ;
      RECT  1435200.0 1510800.0 1445400.0 1497000.0 ;
      RECT  1435200.0 1510800.0 1445400.0 1524600.0 ;
      RECT  1435200.0 1538400.0 1445400.0 1524600.0 ;
      RECT  1435200.0 1538400.0 1445400.0 1552200.0 ;
      RECT  1435200.0 1566000.0 1445400.0 1552200.0 ;
      RECT  1435200.0 1566000.0 1445400.0 1579800.0 ;
      RECT  1435200.0 1593600.0 1445400.0 1579800.0 ;
      RECT  1435200.0 1593600.0 1445400.0 1607400.0 ;
      RECT  1435200.0 1621200.0 1445400.0 1607400.0 ;
      RECT  1435200.0 1621200.0 1445400.0 1635000.0 ;
      RECT  1435200.0 1648800.0 1445400.0 1635000.0 ;
      RECT  1435200.0 1648800.0 1445400.0 1662600.0 ;
      RECT  1435200.0 1676400.0 1445400.0 1662600.0 ;
      RECT  1435200.0 1676400.0 1445400.0 1690200.0 ;
      RECT  1435200.0 1704000.0 1445400.0 1690200.0 ;
      RECT  1435200.0 1704000.0 1445400.0 1717800.0 ;
      RECT  1435200.0 1731600.0 1445400.0 1717800.0 ;
      RECT  1435200.0 1731600.0 1445400.0 1745400.0 ;
      RECT  1435200.0 1759200.0 1445400.0 1745400.0 ;
      RECT  1435200.0 1759200.0 1445400.0 1773000.0 ;
      RECT  1435200.0 1786800.0 1445400.0 1773000.0 ;
      RECT  1435200.0 1786800.0 1445400.0 1800600.0 ;
      RECT  1435200.0 1814400.0 1445400.0 1800600.0 ;
      RECT  1435200.0 1814400.0 1445400.0 1828200.0 ;
      RECT  1435200.0 1842000.0 1445400.0 1828200.0 ;
      RECT  1435200.0 1842000.0 1445400.0 1855800.0 ;
      RECT  1435200.0 1869600.0 1445400.0 1855800.0 ;
      RECT  1435200.0 1869600.0 1445400.0 1883400.0 ;
      RECT  1435200.0 1897200.0 1445400.0 1883400.0 ;
      RECT  1435200.0 1897200.0 1445400.0 1911000.0 ;
      RECT  1435200.0 1924800.0 1445400.0 1911000.0 ;
      RECT  1435200.0 1924800.0 1445400.0 1938600.0 ;
      RECT  1435200.0 1952400.0 1445400.0 1938600.0 ;
      RECT  1435200.0 1952400.0 1445400.0 1966200.0 ;
      RECT  1435200.0 1980000.0 1445400.0 1966200.0 ;
      RECT  1435200.0 1980000.0 1445400.0 1993800.0 ;
      RECT  1435200.0 2007600.0 1445400.0 1993800.0 ;
      RECT  1435200.0 2007600.0 1445400.0 2021400.0 ;
      RECT  1435200.0 2035200.0 1445400.0 2021400.0 ;
      RECT  1435200.0 2035200.0 1445400.0 2049000.0 ;
      RECT  1435200.0 2062800.0 1445400.0 2049000.0 ;
      RECT  1435200.0 2062800.0 1445400.0 2076600.0 ;
      RECT  1435200.0 2090400.0 1445400.0 2076600.0 ;
      RECT  1435200.0 2090400.0 1445400.0 2104200.0 ;
      RECT  1435200.0 2118000.0 1445400.0 2104200.0 ;
      RECT  1435200.0 2118000.0 1445400.0 2131800.0 ;
      RECT  1435200.0 2145600.0 1445400.0 2131800.0 ;
      RECT  1445400.0 379200.0 1455600.0 393000.0 ;
      RECT  1445400.0 406800.0 1455600.0 393000.0 ;
      RECT  1445400.0 406800.0 1455600.0 420600.0 ;
      RECT  1445400.0 434400.0 1455600.0 420600.0 ;
      RECT  1445400.0 434400.0 1455600.0 448200.0 ;
      RECT  1445400.0 462000.0 1455600.0 448200.0 ;
      RECT  1445400.0 462000.0 1455600.0 475800.0 ;
      RECT  1445400.0 489600.0 1455600.0 475800.0 ;
      RECT  1445400.0 489600.0 1455600.0 503400.0 ;
      RECT  1445400.0 517200.0 1455600.0 503400.0 ;
      RECT  1445400.0 517200.0 1455600.0 531000.0 ;
      RECT  1445400.0 544800.0 1455600.0 531000.0 ;
      RECT  1445400.0 544800.0 1455600.0 558600.0 ;
      RECT  1445400.0 572400.0 1455600.0 558600.0 ;
      RECT  1445400.0 572400.0 1455600.0 586200.0 ;
      RECT  1445400.0 600000.0 1455600.0 586200.0 ;
      RECT  1445400.0 600000.0 1455600.0 613800.0 ;
      RECT  1445400.0 627600.0 1455600.0 613800.0 ;
      RECT  1445400.0 627600.0 1455600.0 641400.0 ;
      RECT  1445400.0 655200.0 1455600.0 641400.0 ;
      RECT  1445400.0 655200.0 1455600.0 669000.0 ;
      RECT  1445400.0 682800.0 1455600.0 669000.0 ;
      RECT  1445400.0 682800.0 1455600.0 696600.0 ;
      RECT  1445400.0 710400.0 1455600.0 696600.0 ;
      RECT  1445400.0 710400.0 1455600.0 724200.0 ;
      RECT  1445400.0 738000.0 1455600.0 724200.0 ;
      RECT  1445400.0 738000.0 1455600.0 751800.0 ;
      RECT  1445400.0 765600.0 1455600.0 751800.0 ;
      RECT  1445400.0 765600.0 1455600.0 779400.0 ;
      RECT  1445400.0 793200.0 1455600.0 779400.0 ;
      RECT  1445400.0 793200.0 1455600.0 807000.0 ;
      RECT  1445400.0 820800.0 1455600.0 807000.0 ;
      RECT  1445400.0 820800.0 1455600.0 834600.0 ;
      RECT  1445400.0 848400.0 1455600.0 834600.0 ;
      RECT  1445400.0 848400.0 1455600.0 862200.0 ;
      RECT  1445400.0 876000.0 1455600.0 862200.0 ;
      RECT  1445400.0 876000.0 1455600.0 889800.0 ;
      RECT  1445400.0 903600.0 1455600.0 889800.0 ;
      RECT  1445400.0 903600.0 1455600.0 917400.0 ;
      RECT  1445400.0 931200.0 1455600.0 917400.0 ;
      RECT  1445400.0 931200.0 1455600.0 945000.0 ;
      RECT  1445400.0 958800.0 1455600.0 945000.0 ;
      RECT  1445400.0 958800.0 1455600.0 972600.0 ;
      RECT  1445400.0 986400.0 1455600.0 972600.0 ;
      RECT  1445400.0 986400.0 1455600.0 1000200.0 ;
      RECT  1445400.0 1014000.0 1455600.0 1000200.0 ;
      RECT  1445400.0 1014000.0 1455600.0 1027800.0 ;
      RECT  1445400.0 1041600.0 1455600.0 1027800.0 ;
      RECT  1445400.0 1041600.0 1455600.0 1055400.0 ;
      RECT  1445400.0 1069200.0 1455600.0 1055400.0 ;
      RECT  1445400.0 1069200.0 1455600.0 1083000.0 ;
      RECT  1445400.0 1096800.0 1455600.0 1083000.0 ;
      RECT  1445400.0 1096800.0 1455600.0 1110600.0 ;
      RECT  1445400.0 1124400.0 1455600.0 1110600.0 ;
      RECT  1445400.0 1124400.0 1455600.0 1138200.0 ;
      RECT  1445400.0 1152000.0 1455600.0 1138200.0 ;
      RECT  1445400.0 1152000.0 1455600.0 1165800.0 ;
      RECT  1445400.0 1179600.0 1455600.0 1165800.0 ;
      RECT  1445400.0 1179600.0 1455600.0 1193400.0 ;
      RECT  1445400.0 1207200.0 1455600.0 1193400.0 ;
      RECT  1445400.0 1207200.0 1455600.0 1221000.0 ;
      RECT  1445400.0 1234800.0 1455600.0 1221000.0 ;
      RECT  1445400.0 1234800.0 1455600.0 1248600.0 ;
      RECT  1445400.0 1262400.0 1455600.0 1248600.0 ;
      RECT  1445400.0 1262400.0 1455600.0 1276200.0 ;
      RECT  1445400.0 1290000.0 1455600.0 1276200.0 ;
      RECT  1445400.0 1290000.0 1455600.0 1303800.0 ;
      RECT  1445400.0 1317600.0 1455600.0 1303800.0 ;
      RECT  1445400.0 1317600.0 1455600.0 1331400.0 ;
      RECT  1445400.0 1345200.0 1455600.0 1331400.0 ;
      RECT  1445400.0 1345200.0 1455600.0 1359000.0 ;
      RECT  1445400.0 1372800.0 1455600.0 1359000.0 ;
      RECT  1445400.0 1372800.0 1455600.0 1386600.0 ;
      RECT  1445400.0 1400400.0 1455600.0 1386600.0 ;
      RECT  1445400.0 1400400.0 1455600.0 1414200.0 ;
      RECT  1445400.0 1428000.0 1455600.0 1414200.0 ;
      RECT  1445400.0 1428000.0 1455600.0 1441800.0 ;
      RECT  1445400.0 1455600.0 1455600.0 1441800.0 ;
      RECT  1445400.0 1455600.0 1455600.0 1469400.0 ;
      RECT  1445400.0 1483200.0 1455600.0 1469400.0 ;
      RECT  1445400.0 1483200.0 1455600.0 1497000.0 ;
      RECT  1445400.0 1510800.0 1455600.0 1497000.0 ;
      RECT  1445400.0 1510800.0 1455600.0 1524600.0 ;
      RECT  1445400.0 1538400.0 1455600.0 1524600.0 ;
      RECT  1445400.0 1538400.0 1455600.0 1552200.0 ;
      RECT  1445400.0 1566000.0 1455600.0 1552200.0 ;
      RECT  1445400.0 1566000.0 1455600.0 1579800.0 ;
      RECT  1445400.0 1593600.0 1455600.0 1579800.0 ;
      RECT  1445400.0 1593600.0 1455600.0 1607400.0 ;
      RECT  1445400.0 1621200.0 1455600.0 1607400.0 ;
      RECT  1445400.0 1621200.0 1455600.0 1635000.0 ;
      RECT  1445400.0 1648800.0 1455600.0 1635000.0 ;
      RECT  1445400.0 1648800.0 1455600.0 1662600.0 ;
      RECT  1445400.0 1676400.0 1455600.0 1662600.0 ;
      RECT  1445400.0 1676400.0 1455600.0 1690200.0 ;
      RECT  1445400.0 1704000.0 1455600.0 1690200.0 ;
      RECT  1445400.0 1704000.0 1455600.0 1717800.0 ;
      RECT  1445400.0 1731600.0 1455600.0 1717800.0 ;
      RECT  1445400.0 1731600.0 1455600.0 1745400.0 ;
      RECT  1445400.0 1759200.0 1455600.0 1745400.0 ;
      RECT  1445400.0 1759200.0 1455600.0 1773000.0 ;
      RECT  1445400.0 1786800.0 1455600.0 1773000.0 ;
      RECT  1445400.0 1786800.0 1455600.0 1800600.0 ;
      RECT  1445400.0 1814400.0 1455600.0 1800600.0 ;
      RECT  1445400.0 1814400.0 1455600.0 1828200.0 ;
      RECT  1445400.0 1842000.0 1455600.0 1828200.0 ;
      RECT  1445400.0 1842000.0 1455600.0 1855800.0 ;
      RECT  1445400.0 1869600.0 1455600.0 1855800.0 ;
      RECT  1445400.0 1869600.0 1455600.0 1883400.0 ;
      RECT  1445400.0 1897200.0 1455600.0 1883400.0 ;
      RECT  1445400.0 1897200.0 1455600.0 1911000.0 ;
      RECT  1445400.0 1924800.0 1455600.0 1911000.0 ;
      RECT  1445400.0 1924800.0 1455600.0 1938600.0 ;
      RECT  1445400.0 1952400.0 1455600.0 1938600.0 ;
      RECT  1445400.0 1952400.0 1455600.0 1966200.0 ;
      RECT  1445400.0 1980000.0 1455600.0 1966200.0 ;
      RECT  1445400.0 1980000.0 1455600.0 1993800.0 ;
      RECT  1445400.0 2007600.0 1455600.0 1993800.0 ;
      RECT  1445400.0 2007600.0 1455600.0 2021400.0 ;
      RECT  1445400.0 2035200.0 1455600.0 2021400.0 ;
      RECT  1445400.0 2035200.0 1455600.0 2049000.0 ;
      RECT  1445400.0 2062800.0 1455600.0 2049000.0 ;
      RECT  1445400.0 2062800.0 1455600.0 2076600.0 ;
      RECT  1445400.0 2090400.0 1455600.0 2076600.0 ;
      RECT  1445400.0 2090400.0 1455600.0 2104200.0 ;
      RECT  1445400.0 2118000.0 1455600.0 2104200.0 ;
      RECT  1445400.0 2118000.0 1455600.0 2131800.0 ;
      RECT  1445400.0 2145600.0 1455600.0 2131800.0 ;
      RECT  1455600.0 379200.0 1465800.0 393000.0 ;
      RECT  1455600.0 406800.0 1465800.0 393000.0 ;
      RECT  1455600.0 406800.0 1465800.0 420600.0 ;
      RECT  1455600.0 434400.0 1465800.0 420600.0 ;
      RECT  1455600.0 434400.0 1465800.0 448200.0 ;
      RECT  1455600.0 462000.0 1465800.0 448200.0 ;
      RECT  1455600.0 462000.0 1465800.0 475800.0 ;
      RECT  1455600.0 489600.0 1465800.0 475800.0 ;
      RECT  1455600.0 489600.0 1465800.0 503400.0 ;
      RECT  1455600.0 517200.0 1465800.0 503400.0 ;
      RECT  1455600.0 517200.0 1465800.0 531000.0 ;
      RECT  1455600.0 544800.0 1465800.0 531000.0 ;
      RECT  1455600.0 544800.0 1465800.0 558600.0 ;
      RECT  1455600.0 572400.0 1465800.0 558600.0 ;
      RECT  1455600.0 572400.0 1465800.0 586200.0 ;
      RECT  1455600.0 600000.0 1465800.0 586200.0 ;
      RECT  1455600.0 600000.0 1465800.0 613800.0 ;
      RECT  1455600.0 627600.0 1465800.0 613800.0 ;
      RECT  1455600.0 627600.0 1465800.0 641400.0 ;
      RECT  1455600.0 655200.0 1465800.0 641400.0 ;
      RECT  1455600.0 655200.0 1465800.0 669000.0 ;
      RECT  1455600.0 682800.0 1465800.0 669000.0 ;
      RECT  1455600.0 682800.0 1465800.0 696600.0 ;
      RECT  1455600.0 710400.0 1465800.0 696600.0 ;
      RECT  1455600.0 710400.0 1465800.0 724200.0 ;
      RECT  1455600.0 738000.0 1465800.0 724200.0 ;
      RECT  1455600.0 738000.0 1465800.0 751800.0 ;
      RECT  1455600.0 765600.0 1465800.0 751800.0 ;
      RECT  1455600.0 765600.0 1465800.0 779400.0 ;
      RECT  1455600.0 793200.0 1465800.0 779400.0 ;
      RECT  1455600.0 793200.0 1465800.0 807000.0 ;
      RECT  1455600.0 820800.0 1465800.0 807000.0 ;
      RECT  1455600.0 820800.0 1465800.0 834600.0 ;
      RECT  1455600.0 848400.0 1465800.0 834600.0 ;
      RECT  1455600.0 848400.0 1465800.0 862200.0 ;
      RECT  1455600.0 876000.0 1465800.0 862200.0 ;
      RECT  1455600.0 876000.0 1465800.0 889800.0 ;
      RECT  1455600.0 903600.0 1465800.0 889800.0 ;
      RECT  1455600.0 903600.0 1465800.0 917400.0 ;
      RECT  1455600.0 931200.0 1465800.0 917400.0 ;
      RECT  1455600.0 931200.0 1465800.0 945000.0 ;
      RECT  1455600.0 958800.0 1465800.0 945000.0 ;
      RECT  1455600.0 958800.0 1465800.0 972600.0 ;
      RECT  1455600.0 986400.0 1465800.0 972600.0 ;
      RECT  1455600.0 986400.0 1465800.0 1000200.0 ;
      RECT  1455600.0 1014000.0 1465800.0 1000200.0 ;
      RECT  1455600.0 1014000.0 1465800.0 1027800.0 ;
      RECT  1455600.0 1041600.0 1465800.0 1027800.0 ;
      RECT  1455600.0 1041600.0 1465800.0 1055400.0 ;
      RECT  1455600.0 1069200.0 1465800.0 1055400.0 ;
      RECT  1455600.0 1069200.0 1465800.0 1083000.0 ;
      RECT  1455600.0 1096800.0 1465800.0 1083000.0 ;
      RECT  1455600.0 1096800.0 1465800.0 1110600.0 ;
      RECT  1455600.0 1124400.0 1465800.0 1110600.0 ;
      RECT  1455600.0 1124400.0 1465800.0 1138200.0 ;
      RECT  1455600.0 1152000.0 1465800.0 1138200.0 ;
      RECT  1455600.0 1152000.0 1465800.0 1165800.0 ;
      RECT  1455600.0 1179600.0 1465800.0 1165800.0 ;
      RECT  1455600.0 1179600.0 1465800.0 1193400.0 ;
      RECT  1455600.0 1207200.0 1465800.0 1193400.0 ;
      RECT  1455600.0 1207200.0 1465800.0 1221000.0 ;
      RECT  1455600.0 1234800.0 1465800.0 1221000.0 ;
      RECT  1455600.0 1234800.0 1465800.0 1248600.0 ;
      RECT  1455600.0 1262400.0 1465800.0 1248600.0 ;
      RECT  1455600.0 1262400.0 1465800.0 1276200.0 ;
      RECT  1455600.0 1290000.0 1465800.0 1276200.0 ;
      RECT  1455600.0 1290000.0 1465800.0 1303800.0 ;
      RECT  1455600.0 1317600.0 1465800.0 1303800.0 ;
      RECT  1455600.0 1317600.0 1465800.0 1331400.0 ;
      RECT  1455600.0 1345200.0 1465800.0 1331400.0 ;
      RECT  1455600.0 1345200.0 1465800.0 1359000.0 ;
      RECT  1455600.0 1372800.0 1465800.0 1359000.0 ;
      RECT  1455600.0 1372800.0 1465800.0 1386600.0 ;
      RECT  1455600.0 1400400.0 1465800.0 1386600.0 ;
      RECT  1455600.0 1400400.0 1465800.0 1414200.0 ;
      RECT  1455600.0 1428000.0 1465800.0 1414200.0 ;
      RECT  1455600.0 1428000.0 1465800.0 1441800.0 ;
      RECT  1455600.0 1455600.0 1465800.0 1441800.0 ;
      RECT  1455600.0 1455600.0 1465800.0 1469400.0 ;
      RECT  1455600.0 1483200.0 1465800.0 1469400.0 ;
      RECT  1455600.0 1483200.0 1465800.0 1497000.0 ;
      RECT  1455600.0 1510800.0 1465800.0 1497000.0 ;
      RECT  1455600.0 1510800.0 1465800.0 1524600.0 ;
      RECT  1455600.0 1538400.0 1465800.0 1524600.0 ;
      RECT  1455600.0 1538400.0 1465800.0 1552200.0 ;
      RECT  1455600.0 1566000.0 1465800.0 1552200.0 ;
      RECT  1455600.0 1566000.0 1465800.0 1579800.0 ;
      RECT  1455600.0 1593600.0 1465800.0 1579800.0 ;
      RECT  1455600.0 1593600.0 1465800.0 1607400.0 ;
      RECT  1455600.0 1621200.0 1465800.0 1607400.0 ;
      RECT  1455600.0 1621200.0 1465800.0 1635000.0 ;
      RECT  1455600.0 1648800.0 1465800.0 1635000.0 ;
      RECT  1455600.0 1648800.0 1465800.0 1662600.0 ;
      RECT  1455600.0 1676400.0 1465800.0 1662600.0 ;
      RECT  1455600.0 1676400.0 1465800.0 1690200.0 ;
      RECT  1455600.0 1704000.0 1465800.0 1690200.0 ;
      RECT  1455600.0 1704000.0 1465800.0 1717800.0 ;
      RECT  1455600.0 1731600.0 1465800.0 1717800.0 ;
      RECT  1455600.0 1731600.0 1465800.0 1745400.0 ;
      RECT  1455600.0 1759200.0 1465800.0 1745400.0 ;
      RECT  1455600.0 1759200.0 1465800.0 1773000.0 ;
      RECT  1455600.0 1786800.0 1465800.0 1773000.0 ;
      RECT  1455600.0 1786800.0 1465800.0 1800600.0 ;
      RECT  1455600.0 1814400.0 1465800.0 1800600.0 ;
      RECT  1455600.0 1814400.0 1465800.0 1828200.0 ;
      RECT  1455600.0 1842000.0 1465800.0 1828200.0 ;
      RECT  1455600.0 1842000.0 1465800.0 1855800.0 ;
      RECT  1455600.0 1869600.0 1465800.0 1855800.0 ;
      RECT  1455600.0 1869600.0 1465800.0 1883400.0 ;
      RECT  1455600.0 1897200.0 1465800.0 1883400.0 ;
      RECT  1455600.0 1897200.0 1465800.0 1911000.0 ;
      RECT  1455600.0 1924800.0 1465800.0 1911000.0 ;
      RECT  1455600.0 1924800.0 1465800.0 1938600.0 ;
      RECT  1455600.0 1952400.0 1465800.0 1938600.0 ;
      RECT  1455600.0 1952400.0 1465800.0 1966200.0 ;
      RECT  1455600.0 1980000.0 1465800.0 1966200.0 ;
      RECT  1455600.0 1980000.0 1465800.0 1993800.0 ;
      RECT  1455600.0 2007600.0 1465800.0 1993800.0 ;
      RECT  1455600.0 2007600.0 1465800.0 2021400.0 ;
      RECT  1455600.0 2035200.0 1465800.0 2021400.0 ;
      RECT  1455600.0 2035200.0 1465800.0 2049000.0 ;
      RECT  1455600.0 2062800.0 1465800.0 2049000.0 ;
      RECT  1455600.0 2062800.0 1465800.0 2076600.0 ;
      RECT  1455600.0 2090400.0 1465800.0 2076600.0 ;
      RECT  1455600.0 2090400.0 1465800.0 2104200.0 ;
      RECT  1455600.0 2118000.0 1465800.0 2104200.0 ;
      RECT  1455600.0 2118000.0 1465800.0 2131800.0 ;
      RECT  1455600.0 2145600.0 1465800.0 2131800.0 ;
      RECT  1465800.0 379200.0 1476000.0 393000.0 ;
      RECT  1465800.0 406800.0 1476000.0 393000.0 ;
      RECT  1465800.0 406800.0 1476000.0 420600.0 ;
      RECT  1465800.0 434400.0 1476000.0 420600.0 ;
      RECT  1465800.0 434400.0 1476000.0 448200.0 ;
      RECT  1465800.0 462000.0 1476000.0 448200.0 ;
      RECT  1465800.0 462000.0 1476000.0 475800.0 ;
      RECT  1465800.0 489600.0 1476000.0 475800.0 ;
      RECT  1465800.0 489600.0 1476000.0 503400.0 ;
      RECT  1465800.0 517200.0 1476000.0 503400.0 ;
      RECT  1465800.0 517200.0 1476000.0 531000.0 ;
      RECT  1465800.0 544800.0 1476000.0 531000.0 ;
      RECT  1465800.0 544800.0 1476000.0 558600.0 ;
      RECT  1465800.0 572400.0 1476000.0 558600.0 ;
      RECT  1465800.0 572400.0 1476000.0 586200.0 ;
      RECT  1465800.0 600000.0 1476000.0 586200.0 ;
      RECT  1465800.0 600000.0 1476000.0 613800.0 ;
      RECT  1465800.0 627600.0 1476000.0 613800.0 ;
      RECT  1465800.0 627600.0 1476000.0 641400.0 ;
      RECT  1465800.0 655200.0 1476000.0 641400.0 ;
      RECT  1465800.0 655200.0 1476000.0 669000.0 ;
      RECT  1465800.0 682800.0 1476000.0 669000.0 ;
      RECT  1465800.0 682800.0 1476000.0 696600.0 ;
      RECT  1465800.0 710400.0 1476000.0 696600.0 ;
      RECT  1465800.0 710400.0 1476000.0 724200.0 ;
      RECT  1465800.0 738000.0 1476000.0 724200.0 ;
      RECT  1465800.0 738000.0 1476000.0 751800.0 ;
      RECT  1465800.0 765600.0 1476000.0 751800.0 ;
      RECT  1465800.0 765600.0 1476000.0 779400.0 ;
      RECT  1465800.0 793200.0 1476000.0 779400.0 ;
      RECT  1465800.0 793200.0 1476000.0 807000.0 ;
      RECT  1465800.0 820800.0 1476000.0 807000.0 ;
      RECT  1465800.0 820800.0 1476000.0 834600.0 ;
      RECT  1465800.0 848400.0 1476000.0 834600.0 ;
      RECT  1465800.0 848400.0 1476000.0 862200.0 ;
      RECT  1465800.0 876000.0 1476000.0 862200.0 ;
      RECT  1465800.0 876000.0 1476000.0 889800.0 ;
      RECT  1465800.0 903600.0 1476000.0 889800.0 ;
      RECT  1465800.0 903600.0 1476000.0 917400.0 ;
      RECT  1465800.0 931200.0 1476000.0 917400.0 ;
      RECT  1465800.0 931200.0 1476000.0 945000.0 ;
      RECT  1465800.0 958800.0 1476000.0 945000.0 ;
      RECT  1465800.0 958800.0 1476000.0 972600.0 ;
      RECT  1465800.0 986400.0 1476000.0 972600.0 ;
      RECT  1465800.0 986400.0 1476000.0 1000200.0 ;
      RECT  1465800.0 1014000.0 1476000.0 1000200.0 ;
      RECT  1465800.0 1014000.0 1476000.0 1027800.0 ;
      RECT  1465800.0 1041600.0 1476000.0 1027800.0 ;
      RECT  1465800.0 1041600.0 1476000.0 1055400.0 ;
      RECT  1465800.0 1069200.0 1476000.0 1055400.0 ;
      RECT  1465800.0 1069200.0 1476000.0 1083000.0 ;
      RECT  1465800.0 1096800.0 1476000.0 1083000.0 ;
      RECT  1465800.0 1096800.0 1476000.0 1110600.0 ;
      RECT  1465800.0 1124400.0 1476000.0 1110600.0 ;
      RECT  1465800.0 1124400.0 1476000.0 1138200.0 ;
      RECT  1465800.0 1152000.0 1476000.0 1138200.0 ;
      RECT  1465800.0 1152000.0 1476000.0 1165800.0 ;
      RECT  1465800.0 1179600.0 1476000.0 1165800.0 ;
      RECT  1465800.0 1179600.0 1476000.0 1193400.0 ;
      RECT  1465800.0 1207200.0 1476000.0 1193400.0 ;
      RECT  1465800.0 1207200.0 1476000.0 1221000.0 ;
      RECT  1465800.0 1234800.0 1476000.0 1221000.0 ;
      RECT  1465800.0 1234800.0 1476000.0 1248600.0 ;
      RECT  1465800.0 1262400.0 1476000.0 1248600.0 ;
      RECT  1465800.0 1262400.0 1476000.0 1276200.0 ;
      RECT  1465800.0 1290000.0 1476000.0 1276200.0 ;
      RECT  1465800.0 1290000.0 1476000.0 1303800.0 ;
      RECT  1465800.0 1317600.0 1476000.0 1303800.0 ;
      RECT  1465800.0 1317600.0 1476000.0 1331400.0 ;
      RECT  1465800.0 1345200.0 1476000.0 1331400.0 ;
      RECT  1465800.0 1345200.0 1476000.0 1359000.0 ;
      RECT  1465800.0 1372800.0 1476000.0 1359000.0 ;
      RECT  1465800.0 1372800.0 1476000.0 1386600.0 ;
      RECT  1465800.0 1400400.0 1476000.0 1386600.0 ;
      RECT  1465800.0 1400400.0 1476000.0 1414200.0 ;
      RECT  1465800.0 1428000.0 1476000.0 1414200.0 ;
      RECT  1465800.0 1428000.0 1476000.0 1441800.0 ;
      RECT  1465800.0 1455600.0 1476000.0 1441800.0 ;
      RECT  1465800.0 1455600.0 1476000.0 1469400.0 ;
      RECT  1465800.0 1483200.0 1476000.0 1469400.0 ;
      RECT  1465800.0 1483200.0 1476000.0 1497000.0 ;
      RECT  1465800.0 1510800.0 1476000.0 1497000.0 ;
      RECT  1465800.0 1510800.0 1476000.0 1524600.0 ;
      RECT  1465800.0 1538400.0 1476000.0 1524600.0 ;
      RECT  1465800.0 1538400.0 1476000.0 1552200.0 ;
      RECT  1465800.0 1566000.0 1476000.0 1552200.0 ;
      RECT  1465800.0 1566000.0 1476000.0 1579800.0 ;
      RECT  1465800.0 1593600.0 1476000.0 1579800.0 ;
      RECT  1465800.0 1593600.0 1476000.0 1607400.0 ;
      RECT  1465800.0 1621200.0 1476000.0 1607400.0 ;
      RECT  1465800.0 1621200.0 1476000.0 1635000.0 ;
      RECT  1465800.0 1648800.0 1476000.0 1635000.0 ;
      RECT  1465800.0 1648800.0 1476000.0 1662600.0 ;
      RECT  1465800.0 1676400.0 1476000.0 1662600.0 ;
      RECT  1465800.0 1676400.0 1476000.0 1690200.0 ;
      RECT  1465800.0 1704000.0 1476000.0 1690200.0 ;
      RECT  1465800.0 1704000.0 1476000.0 1717800.0 ;
      RECT  1465800.0 1731600.0 1476000.0 1717800.0 ;
      RECT  1465800.0 1731600.0 1476000.0 1745400.0 ;
      RECT  1465800.0 1759200.0 1476000.0 1745400.0 ;
      RECT  1465800.0 1759200.0 1476000.0 1773000.0 ;
      RECT  1465800.0 1786800.0 1476000.0 1773000.0 ;
      RECT  1465800.0 1786800.0 1476000.0 1800600.0 ;
      RECT  1465800.0 1814400.0 1476000.0 1800600.0 ;
      RECT  1465800.0 1814400.0 1476000.0 1828200.0 ;
      RECT  1465800.0 1842000.0 1476000.0 1828200.0 ;
      RECT  1465800.0 1842000.0 1476000.0 1855800.0 ;
      RECT  1465800.0 1869600.0 1476000.0 1855800.0 ;
      RECT  1465800.0 1869600.0 1476000.0 1883400.0 ;
      RECT  1465800.0 1897200.0 1476000.0 1883400.0 ;
      RECT  1465800.0 1897200.0 1476000.0 1911000.0 ;
      RECT  1465800.0 1924800.0 1476000.0 1911000.0 ;
      RECT  1465800.0 1924800.0 1476000.0 1938600.0 ;
      RECT  1465800.0 1952400.0 1476000.0 1938600.0 ;
      RECT  1465800.0 1952400.0 1476000.0 1966200.0 ;
      RECT  1465800.0 1980000.0 1476000.0 1966200.0 ;
      RECT  1465800.0 1980000.0 1476000.0 1993800.0 ;
      RECT  1465800.0 2007600.0 1476000.0 1993800.0 ;
      RECT  1465800.0 2007600.0 1476000.0 2021400.0 ;
      RECT  1465800.0 2035200.0 1476000.0 2021400.0 ;
      RECT  1465800.0 2035200.0 1476000.0 2049000.0 ;
      RECT  1465800.0 2062800.0 1476000.0 2049000.0 ;
      RECT  1465800.0 2062800.0 1476000.0 2076600.0 ;
      RECT  1465800.0 2090400.0 1476000.0 2076600.0 ;
      RECT  1465800.0 2090400.0 1476000.0 2104200.0 ;
      RECT  1465800.0 2118000.0 1476000.0 2104200.0 ;
      RECT  1465800.0 2118000.0 1476000.0 2131800.0 ;
      RECT  1465800.0 2145600.0 1476000.0 2131800.0 ;
      RECT  1476000.0 379200.0 1486200.0 393000.0 ;
      RECT  1476000.0 406800.0 1486200.0 393000.0 ;
      RECT  1476000.0 406800.0 1486200.0 420600.0 ;
      RECT  1476000.0 434400.0 1486200.0 420600.0 ;
      RECT  1476000.0 434400.0 1486200.0 448200.0 ;
      RECT  1476000.0 462000.0 1486200.0 448200.0 ;
      RECT  1476000.0 462000.0 1486200.0 475800.0 ;
      RECT  1476000.0 489600.0 1486200.0 475800.0 ;
      RECT  1476000.0 489600.0 1486200.0 503400.0 ;
      RECT  1476000.0 517200.0 1486200.0 503400.0 ;
      RECT  1476000.0 517200.0 1486200.0 531000.0 ;
      RECT  1476000.0 544800.0 1486200.0 531000.0 ;
      RECT  1476000.0 544800.0 1486200.0 558600.0 ;
      RECT  1476000.0 572400.0 1486200.0 558600.0 ;
      RECT  1476000.0 572400.0 1486200.0 586200.0 ;
      RECT  1476000.0 600000.0 1486200.0 586200.0 ;
      RECT  1476000.0 600000.0 1486200.0 613800.0 ;
      RECT  1476000.0 627600.0 1486200.0 613800.0 ;
      RECT  1476000.0 627600.0 1486200.0 641400.0 ;
      RECT  1476000.0 655200.0 1486200.0 641400.0 ;
      RECT  1476000.0 655200.0 1486200.0 669000.0 ;
      RECT  1476000.0 682800.0 1486200.0 669000.0 ;
      RECT  1476000.0 682800.0 1486200.0 696600.0 ;
      RECT  1476000.0 710400.0 1486200.0 696600.0 ;
      RECT  1476000.0 710400.0 1486200.0 724200.0 ;
      RECT  1476000.0 738000.0 1486200.0 724200.0 ;
      RECT  1476000.0 738000.0 1486200.0 751800.0 ;
      RECT  1476000.0 765600.0 1486200.0 751800.0 ;
      RECT  1476000.0 765600.0 1486200.0 779400.0 ;
      RECT  1476000.0 793200.0 1486200.0 779400.0 ;
      RECT  1476000.0 793200.0 1486200.0 807000.0 ;
      RECT  1476000.0 820800.0 1486200.0 807000.0 ;
      RECT  1476000.0 820800.0 1486200.0 834600.0 ;
      RECT  1476000.0 848400.0 1486200.0 834600.0 ;
      RECT  1476000.0 848400.0 1486200.0 862200.0 ;
      RECT  1476000.0 876000.0 1486200.0 862200.0 ;
      RECT  1476000.0 876000.0 1486200.0 889800.0 ;
      RECT  1476000.0 903600.0 1486200.0 889800.0 ;
      RECT  1476000.0 903600.0 1486200.0 917400.0 ;
      RECT  1476000.0 931200.0 1486200.0 917400.0 ;
      RECT  1476000.0 931200.0 1486200.0 945000.0 ;
      RECT  1476000.0 958800.0 1486200.0 945000.0 ;
      RECT  1476000.0 958800.0 1486200.0 972600.0 ;
      RECT  1476000.0 986400.0 1486200.0 972600.0 ;
      RECT  1476000.0 986400.0 1486200.0 1000200.0 ;
      RECT  1476000.0 1014000.0 1486200.0 1000200.0 ;
      RECT  1476000.0 1014000.0 1486200.0 1027800.0 ;
      RECT  1476000.0 1041600.0 1486200.0 1027800.0 ;
      RECT  1476000.0 1041600.0 1486200.0 1055400.0 ;
      RECT  1476000.0 1069200.0 1486200.0 1055400.0 ;
      RECT  1476000.0 1069200.0 1486200.0 1083000.0 ;
      RECT  1476000.0 1096800.0 1486200.0 1083000.0 ;
      RECT  1476000.0 1096800.0 1486200.0 1110600.0 ;
      RECT  1476000.0 1124400.0 1486200.0 1110600.0 ;
      RECT  1476000.0 1124400.0 1486200.0 1138200.0 ;
      RECT  1476000.0 1152000.0 1486200.0 1138200.0 ;
      RECT  1476000.0 1152000.0 1486200.0 1165800.0 ;
      RECT  1476000.0 1179600.0 1486200.0 1165800.0 ;
      RECT  1476000.0 1179600.0 1486200.0 1193400.0 ;
      RECT  1476000.0 1207200.0 1486200.0 1193400.0 ;
      RECT  1476000.0 1207200.0 1486200.0 1221000.0 ;
      RECT  1476000.0 1234800.0 1486200.0 1221000.0 ;
      RECT  1476000.0 1234800.0 1486200.0 1248600.0 ;
      RECT  1476000.0 1262400.0 1486200.0 1248600.0 ;
      RECT  1476000.0 1262400.0 1486200.0 1276200.0 ;
      RECT  1476000.0 1290000.0 1486200.0 1276200.0 ;
      RECT  1476000.0 1290000.0 1486200.0 1303800.0 ;
      RECT  1476000.0 1317600.0 1486200.0 1303800.0 ;
      RECT  1476000.0 1317600.0 1486200.0 1331400.0 ;
      RECT  1476000.0 1345200.0 1486200.0 1331400.0 ;
      RECT  1476000.0 1345200.0 1486200.0 1359000.0 ;
      RECT  1476000.0 1372800.0 1486200.0 1359000.0 ;
      RECT  1476000.0 1372800.0 1486200.0 1386600.0 ;
      RECT  1476000.0 1400400.0 1486200.0 1386600.0 ;
      RECT  1476000.0 1400400.0 1486200.0 1414200.0 ;
      RECT  1476000.0 1428000.0 1486200.0 1414200.0 ;
      RECT  1476000.0 1428000.0 1486200.0 1441800.0 ;
      RECT  1476000.0 1455600.0 1486200.0 1441800.0 ;
      RECT  1476000.0 1455600.0 1486200.0 1469400.0 ;
      RECT  1476000.0 1483200.0 1486200.0 1469400.0 ;
      RECT  1476000.0 1483200.0 1486200.0 1497000.0 ;
      RECT  1476000.0 1510800.0 1486200.0 1497000.0 ;
      RECT  1476000.0 1510800.0 1486200.0 1524600.0 ;
      RECT  1476000.0 1538400.0 1486200.0 1524600.0 ;
      RECT  1476000.0 1538400.0 1486200.0 1552200.0 ;
      RECT  1476000.0 1566000.0 1486200.0 1552200.0 ;
      RECT  1476000.0 1566000.0 1486200.0 1579800.0 ;
      RECT  1476000.0 1593600.0 1486200.0 1579800.0 ;
      RECT  1476000.0 1593600.0 1486200.0 1607400.0 ;
      RECT  1476000.0 1621200.0 1486200.0 1607400.0 ;
      RECT  1476000.0 1621200.0 1486200.0 1635000.0 ;
      RECT  1476000.0 1648800.0 1486200.0 1635000.0 ;
      RECT  1476000.0 1648800.0 1486200.0 1662600.0 ;
      RECT  1476000.0 1676400.0 1486200.0 1662600.0 ;
      RECT  1476000.0 1676400.0 1486200.0 1690200.0 ;
      RECT  1476000.0 1704000.0 1486200.0 1690200.0 ;
      RECT  1476000.0 1704000.0 1486200.0 1717800.0 ;
      RECT  1476000.0 1731600.0 1486200.0 1717800.0 ;
      RECT  1476000.0 1731600.0 1486200.0 1745400.0 ;
      RECT  1476000.0 1759200.0 1486200.0 1745400.0 ;
      RECT  1476000.0 1759200.0 1486200.0 1773000.0 ;
      RECT  1476000.0 1786800.0 1486200.0 1773000.0 ;
      RECT  1476000.0 1786800.0 1486200.0 1800600.0 ;
      RECT  1476000.0 1814400.0 1486200.0 1800600.0 ;
      RECT  1476000.0 1814400.0 1486200.0 1828200.0 ;
      RECT  1476000.0 1842000.0 1486200.0 1828200.0 ;
      RECT  1476000.0 1842000.0 1486200.0 1855800.0 ;
      RECT  1476000.0 1869600.0 1486200.0 1855800.0 ;
      RECT  1476000.0 1869600.0 1486200.0 1883400.0 ;
      RECT  1476000.0 1897200.0 1486200.0 1883400.0 ;
      RECT  1476000.0 1897200.0 1486200.0 1911000.0 ;
      RECT  1476000.0 1924800.0 1486200.0 1911000.0 ;
      RECT  1476000.0 1924800.0 1486200.0 1938600.0 ;
      RECT  1476000.0 1952400.0 1486200.0 1938600.0 ;
      RECT  1476000.0 1952400.0 1486200.0 1966200.0 ;
      RECT  1476000.0 1980000.0 1486200.0 1966200.0 ;
      RECT  1476000.0 1980000.0 1486200.0 1993800.0 ;
      RECT  1476000.0 2007600.0 1486200.0 1993800.0 ;
      RECT  1476000.0 2007600.0 1486200.0 2021400.0 ;
      RECT  1476000.0 2035200.0 1486200.0 2021400.0 ;
      RECT  1476000.0 2035200.0 1486200.0 2049000.0 ;
      RECT  1476000.0 2062800.0 1486200.0 2049000.0 ;
      RECT  1476000.0 2062800.0 1486200.0 2076600.0 ;
      RECT  1476000.0 2090400.0 1486200.0 2076600.0 ;
      RECT  1476000.0 2090400.0 1486200.0 2104200.0 ;
      RECT  1476000.0 2118000.0 1486200.0 2104200.0 ;
      RECT  1476000.0 2118000.0 1486200.0 2131800.0 ;
      RECT  1476000.0 2145600.0 1486200.0 2131800.0 ;
      RECT  1486200.0 379200.0 1496400.0 393000.0 ;
      RECT  1486200.0 406800.0 1496400.0 393000.0 ;
      RECT  1486200.0 406800.0 1496400.0 420600.0 ;
      RECT  1486200.0 434400.0 1496400.0 420600.0 ;
      RECT  1486200.0 434400.0 1496400.0 448200.0 ;
      RECT  1486200.0 462000.0 1496400.0 448200.0 ;
      RECT  1486200.0 462000.0 1496400.0 475800.0 ;
      RECT  1486200.0 489600.0 1496400.0 475800.0 ;
      RECT  1486200.0 489600.0 1496400.0 503400.0 ;
      RECT  1486200.0 517200.0 1496400.0 503400.0 ;
      RECT  1486200.0 517200.0 1496400.0 531000.0 ;
      RECT  1486200.0 544800.0 1496400.0 531000.0 ;
      RECT  1486200.0 544800.0 1496400.0 558600.0 ;
      RECT  1486200.0 572400.0 1496400.0 558600.0 ;
      RECT  1486200.0 572400.0 1496400.0 586200.0 ;
      RECT  1486200.0 600000.0 1496400.0 586200.0 ;
      RECT  1486200.0 600000.0 1496400.0 613800.0 ;
      RECT  1486200.0 627600.0 1496400.0 613800.0 ;
      RECT  1486200.0 627600.0 1496400.0 641400.0 ;
      RECT  1486200.0 655200.0 1496400.0 641400.0 ;
      RECT  1486200.0 655200.0 1496400.0 669000.0 ;
      RECT  1486200.0 682800.0 1496400.0 669000.0 ;
      RECT  1486200.0 682800.0 1496400.0 696600.0 ;
      RECT  1486200.0 710400.0 1496400.0 696600.0 ;
      RECT  1486200.0 710400.0 1496400.0 724200.0 ;
      RECT  1486200.0 738000.0 1496400.0 724200.0 ;
      RECT  1486200.0 738000.0 1496400.0 751800.0 ;
      RECT  1486200.0 765600.0 1496400.0 751800.0 ;
      RECT  1486200.0 765600.0 1496400.0 779400.0 ;
      RECT  1486200.0 793200.0 1496400.0 779400.0 ;
      RECT  1486200.0 793200.0 1496400.0 807000.0 ;
      RECT  1486200.0 820800.0 1496400.0 807000.0 ;
      RECT  1486200.0 820800.0 1496400.0 834600.0 ;
      RECT  1486200.0 848400.0 1496400.0 834600.0 ;
      RECT  1486200.0 848400.0 1496400.0 862200.0 ;
      RECT  1486200.0 876000.0 1496400.0 862200.0 ;
      RECT  1486200.0 876000.0 1496400.0 889800.0 ;
      RECT  1486200.0 903600.0 1496400.0 889800.0 ;
      RECT  1486200.0 903600.0 1496400.0 917400.0 ;
      RECT  1486200.0 931200.0 1496400.0 917400.0 ;
      RECT  1486200.0 931200.0 1496400.0 945000.0 ;
      RECT  1486200.0 958800.0 1496400.0 945000.0 ;
      RECT  1486200.0 958800.0 1496400.0 972600.0 ;
      RECT  1486200.0 986400.0 1496400.0 972600.0 ;
      RECT  1486200.0 986400.0 1496400.0 1000200.0 ;
      RECT  1486200.0 1014000.0 1496400.0 1000200.0 ;
      RECT  1486200.0 1014000.0 1496400.0 1027800.0 ;
      RECT  1486200.0 1041600.0 1496400.0 1027800.0 ;
      RECT  1486200.0 1041600.0 1496400.0 1055400.0 ;
      RECT  1486200.0 1069200.0 1496400.0 1055400.0 ;
      RECT  1486200.0 1069200.0 1496400.0 1083000.0 ;
      RECT  1486200.0 1096800.0 1496400.0 1083000.0 ;
      RECT  1486200.0 1096800.0 1496400.0 1110600.0 ;
      RECT  1486200.0 1124400.0 1496400.0 1110600.0 ;
      RECT  1486200.0 1124400.0 1496400.0 1138200.0 ;
      RECT  1486200.0 1152000.0 1496400.0 1138200.0 ;
      RECT  1486200.0 1152000.0 1496400.0 1165800.0 ;
      RECT  1486200.0 1179600.0 1496400.0 1165800.0 ;
      RECT  1486200.0 1179600.0 1496400.0 1193400.0 ;
      RECT  1486200.0 1207200.0 1496400.0 1193400.0 ;
      RECT  1486200.0 1207200.0 1496400.0 1221000.0 ;
      RECT  1486200.0 1234800.0 1496400.0 1221000.0 ;
      RECT  1486200.0 1234800.0 1496400.0 1248600.0 ;
      RECT  1486200.0 1262400.0 1496400.0 1248600.0 ;
      RECT  1486200.0 1262400.0 1496400.0 1276200.0 ;
      RECT  1486200.0 1290000.0 1496400.0 1276200.0 ;
      RECT  1486200.0 1290000.0 1496400.0 1303800.0 ;
      RECT  1486200.0 1317600.0 1496400.0 1303800.0 ;
      RECT  1486200.0 1317600.0 1496400.0 1331400.0 ;
      RECT  1486200.0 1345200.0 1496400.0 1331400.0 ;
      RECT  1486200.0 1345200.0 1496400.0 1359000.0 ;
      RECT  1486200.0 1372800.0 1496400.0 1359000.0 ;
      RECT  1486200.0 1372800.0 1496400.0 1386600.0 ;
      RECT  1486200.0 1400400.0 1496400.0 1386600.0 ;
      RECT  1486200.0 1400400.0 1496400.0 1414200.0 ;
      RECT  1486200.0 1428000.0 1496400.0 1414200.0 ;
      RECT  1486200.0 1428000.0 1496400.0 1441800.0 ;
      RECT  1486200.0 1455600.0 1496400.0 1441800.0 ;
      RECT  1486200.0 1455600.0 1496400.0 1469400.0 ;
      RECT  1486200.0 1483200.0 1496400.0 1469400.0 ;
      RECT  1486200.0 1483200.0 1496400.0 1497000.0 ;
      RECT  1486200.0 1510800.0 1496400.0 1497000.0 ;
      RECT  1486200.0 1510800.0 1496400.0 1524600.0 ;
      RECT  1486200.0 1538400.0 1496400.0 1524600.0 ;
      RECT  1486200.0 1538400.0 1496400.0 1552200.0 ;
      RECT  1486200.0 1566000.0 1496400.0 1552200.0 ;
      RECT  1486200.0 1566000.0 1496400.0 1579800.0 ;
      RECT  1486200.0 1593600.0 1496400.0 1579800.0 ;
      RECT  1486200.0 1593600.0 1496400.0 1607400.0 ;
      RECT  1486200.0 1621200.0 1496400.0 1607400.0 ;
      RECT  1486200.0 1621200.0 1496400.0 1635000.0 ;
      RECT  1486200.0 1648800.0 1496400.0 1635000.0 ;
      RECT  1486200.0 1648800.0 1496400.0 1662600.0 ;
      RECT  1486200.0 1676400.0 1496400.0 1662600.0 ;
      RECT  1486200.0 1676400.0 1496400.0 1690200.0 ;
      RECT  1486200.0 1704000.0 1496400.0 1690200.0 ;
      RECT  1486200.0 1704000.0 1496400.0 1717800.0 ;
      RECT  1486200.0 1731600.0 1496400.0 1717800.0 ;
      RECT  1486200.0 1731600.0 1496400.0 1745400.0 ;
      RECT  1486200.0 1759200.0 1496400.0 1745400.0 ;
      RECT  1486200.0 1759200.0 1496400.0 1773000.0 ;
      RECT  1486200.0 1786800.0 1496400.0 1773000.0 ;
      RECT  1486200.0 1786800.0 1496400.0 1800600.0 ;
      RECT  1486200.0 1814400.0 1496400.0 1800600.0 ;
      RECT  1486200.0 1814400.0 1496400.0 1828200.0 ;
      RECT  1486200.0 1842000.0 1496400.0 1828200.0 ;
      RECT  1486200.0 1842000.0 1496400.0 1855800.0 ;
      RECT  1486200.0 1869600.0 1496400.0 1855800.0 ;
      RECT  1486200.0 1869600.0 1496400.0 1883400.0 ;
      RECT  1486200.0 1897200.0 1496400.0 1883400.0 ;
      RECT  1486200.0 1897200.0 1496400.0 1911000.0 ;
      RECT  1486200.0 1924800.0 1496400.0 1911000.0 ;
      RECT  1486200.0 1924800.0 1496400.0 1938600.0 ;
      RECT  1486200.0 1952400.0 1496400.0 1938600.0 ;
      RECT  1486200.0 1952400.0 1496400.0 1966200.0 ;
      RECT  1486200.0 1980000.0 1496400.0 1966200.0 ;
      RECT  1486200.0 1980000.0 1496400.0 1993800.0 ;
      RECT  1486200.0 2007600.0 1496400.0 1993800.0 ;
      RECT  1486200.0 2007600.0 1496400.0 2021400.0 ;
      RECT  1486200.0 2035200.0 1496400.0 2021400.0 ;
      RECT  1486200.0 2035200.0 1496400.0 2049000.0 ;
      RECT  1486200.0 2062800.0 1496400.0 2049000.0 ;
      RECT  1486200.0 2062800.0 1496400.0 2076600.0 ;
      RECT  1486200.0 2090400.0 1496400.0 2076600.0 ;
      RECT  1486200.0 2090400.0 1496400.0 2104200.0 ;
      RECT  1486200.0 2118000.0 1496400.0 2104200.0 ;
      RECT  1486200.0 2118000.0 1496400.0 2131800.0 ;
      RECT  1486200.0 2145600.0 1496400.0 2131800.0 ;
      RECT  1496400.0 379200.0 1506600.0 393000.0 ;
      RECT  1496400.0 406800.0 1506600.0 393000.0 ;
      RECT  1496400.0 406800.0 1506600.0 420600.0 ;
      RECT  1496400.0 434400.0 1506600.0 420600.0 ;
      RECT  1496400.0 434400.0 1506600.0 448200.0 ;
      RECT  1496400.0 462000.0 1506600.0 448200.0 ;
      RECT  1496400.0 462000.0 1506600.0 475800.0 ;
      RECT  1496400.0 489600.0 1506600.0 475800.0 ;
      RECT  1496400.0 489600.0 1506600.0 503400.0 ;
      RECT  1496400.0 517200.0 1506600.0 503400.0 ;
      RECT  1496400.0 517200.0 1506600.0 531000.0 ;
      RECT  1496400.0 544800.0 1506600.0 531000.0 ;
      RECT  1496400.0 544800.0 1506600.0 558600.0 ;
      RECT  1496400.0 572400.0 1506600.0 558600.0 ;
      RECT  1496400.0 572400.0 1506600.0 586200.0 ;
      RECT  1496400.0 600000.0 1506600.0 586200.0 ;
      RECT  1496400.0 600000.0 1506600.0 613800.0 ;
      RECT  1496400.0 627600.0 1506600.0 613800.0 ;
      RECT  1496400.0 627600.0 1506600.0 641400.0 ;
      RECT  1496400.0 655200.0 1506600.0 641400.0 ;
      RECT  1496400.0 655200.0 1506600.0 669000.0 ;
      RECT  1496400.0 682800.0 1506600.0 669000.0 ;
      RECT  1496400.0 682800.0 1506600.0 696600.0 ;
      RECT  1496400.0 710400.0 1506600.0 696600.0 ;
      RECT  1496400.0 710400.0 1506600.0 724200.0 ;
      RECT  1496400.0 738000.0 1506600.0 724200.0 ;
      RECT  1496400.0 738000.0 1506600.0 751800.0 ;
      RECT  1496400.0 765600.0 1506600.0 751800.0 ;
      RECT  1496400.0 765600.0 1506600.0 779400.0 ;
      RECT  1496400.0 793200.0 1506600.0 779400.0 ;
      RECT  1496400.0 793200.0 1506600.0 807000.0 ;
      RECT  1496400.0 820800.0 1506600.0 807000.0 ;
      RECT  1496400.0 820800.0 1506600.0 834600.0 ;
      RECT  1496400.0 848400.0 1506600.0 834600.0 ;
      RECT  1496400.0 848400.0 1506600.0 862200.0 ;
      RECT  1496400.0 876000.0 1506600.0 862200.0 ;
      RECT  1496400.0 876000.0 1506600.0 889800.0 ;
      RECT  1496400.0 903600.0 1506600.0 889800.0 ;
      RECT  1496400.0 903600.0 1506600.0 917400.0 ;
      RECT  1496400.0 931200.0 1506600.0 917400.0 ;
      RECT  1496400.0 931200.0 1506600.0 945000.0 ;
      RECT  1496400.0 958800.0 1506600.0 945000.0 ;
      RECT  1496400.0 958800.0 1506600.0 972600.0 ;
      RECT  1496400.0 986400.0 1506600.0 972600.0 ;
      RECT  1496400.0 986400.0 1506600.0 1000200.0 ;
      RECT  1496400.0 1014000.0 1506600.0 1000200.0 ;
      RECT  1496400.0 1014000.0 1506600.0 1027800.0 ;
      RECT  1496400.0 1041600.0 1506600.0 1027800.0 ;
      RECT  1496400.0 1041600.0 1506600.0 1055400.0 ;
      RECT  1496400.0 1069200.0 1506600.0 1055400.0 ;
      RECT  1496400.0 1069200.0 1506600.0 1083000.0 ;
      RECT  1496400.0 1096800.0 1506600.0 1083000.0 ;
      RECT  1496400.0 1096800.0 1506600.0 1110600.0 ;
      RECT  1496400.0 1124400.0 1506600.0 1110600.0 ;
      RECT  1496400.0 1124400.0 1506600.0 1138200.0 ;
      RECT  1496400.0 1152000.0 1506600.0 1138200.0 ;
      RECT  1496400.0 1152000.0 1506600.0 1165800.0 ;
      RECT  1496400.0 1179600.0 1506600.0 1165800.0 ;
      RECT  1496400.0 1179600.0 1506600.0 1193400.0 ;
      RECT  1496400.0 1207200.0 1506600.0 1193400.0 ;
      RECT  1496400.0 1207200.0 1506600.0 1221000.0 ;
      RECT  1496400.0 1234800.0 1506600.0 1221000.0 ;
      RECT  1496400.0 1234800.0 1506600.0 1248600.0 ;
      RECT  1496400.0 1262400.0 1506600.0 1248600.0 ;
      RECT  1496400.0 1262400.0 1506600.0 1276200.0 ;
      RECT  1496400.0 1290000.0 1506600.0 1276200.0 ;
      RECT  1496400.0 1290000.0 1506600.0 1303800.0 ;
      RECT  1496400.0 1317600.0 1506600.0 1303800.0 ;
      RECT  1496400.0 1317600.0 1506600.0 1331400.0 ;
      RECT  1496400.0 1345200.0 1506600.0 1331400.0 ;
      RECT  1496400.0 1345200.0 1506600.0 1359000.0 ;
      RECT  1496400.0 1372800.0 1506600.0 1359000.0 ;
      RECT  1496400.0 1372800.0 1506600.0 1386600.0 ;
      RECT  1496400.0 1400400.0 1506600.0 1386600.0 ;
      RECT  1496400.0 1400400.0 1506600.0 1414200.0 ;
      RECT  1496400.0 1428000.0 1506600.0 1414200.0 ;
      RECT  1496400.0 1428000.0 1506600.0 1441800.0 ;
      RECT  1496400.0 1455600.0 1506600.0 1441800.0 ;
      RECT  1496400.0 1455600.0 1506600.0 1469400.0 ;
      RECT  1496400.0 1483200.0 1506600.0 1469400.0 ;
      RECT  1496400.0 1483200.0 1506600.0 1497000.0 ;
      RECT  1496400.0 1510800.0 1506600.0 1497000.0 ;
      RECT  1496400.0 1510800.0 1506600.0 1524600.0 ;
      RECT  1496400.0 1538400.0 1506600.0 1524600.0 ;
      RECT  1496400.0 1538400.0 1506600.0 1552200.0 ;
      RECT  1496400.0 1566000.0 1506600.0 1552200.0 ;
      RECT  1496400.0 1566000.0 1506600.0 1579800.0 ;
      RECT  1496400.0 1593600.0 1506600.0 1579800.0 ;
      RECT  1496400.0 1593600.0 1506600.0 1607400.0 ;
      RECT  1496400.0 1621200.0 1506600.0 1607400.0 ;
      RECT  1496400.0 1621200.0 1506600.0 1635000.0 ;
      RECT  1496400.0 1648800.0 1506600.0 1635000.0 ;
      RECT  1496400.0 1648800.0 1506600.0 1662600.0 ;
      RECT  1496400.0 1676400.0 1506600.0 1662600.0 ;
      RECT  1496400.0 1676400.0 1506600.0 1690200.0 ;
      RECT  1496400.0 1704000.0 1506600.0 1690200.0 ;
      RECT  1496400.0 1704000.0 1506600.0 1717800.0 ;
      RECT  1496400.0 1731600.0 1506600.0 1717800.0 ;
      RECT  1496400.0 1731600.0 1506600.0 1745400.0 ;
      RECT  1496400.0 1759200.0 1506600.0 1745400.0 ;
      RECT  1496400.0 1759200.0 1506600.0 1773000.0 ;
      RECT  1496400.0 1786800.0 1506600.0 1773000.0 ;
      RECT  1496400.0 1786800.0 1506600.0 1800600.0 ;
      RECT  1496400.0 1814400.0 1506600.0 1800600.0 ;
      RECT  1496400.0 1814400.0 1506600.0 1828200.0 ;
      RECT  1496400.0 1842000.0 1506600.0 1828200.0 ;
      RECT  1496400.0 1842000.0 1506600.0 1855800.0 ;
      RECT  1496400.0 1869600.0 1506600.0 1855800.0 ;
      RECT  1496400.0 1869600.0 1506600.0 1883400.0 ;
      RECT  1496400.0 1897200.0 1506600.0 1883400.0 ;
      RECT  1496400.0 1897200.0 1506600.0 1911000.0 ;
      RECT  1496400.0 1924800.0 1506600.0 1911000.0 ;
      RECT  1496400.0 1924800.0 1506600.0 1938600.0 ;
      RECT  1496400.0 1952400.0 1506600.0 1938600.0 ;
      RECT  1496400.0 1952400.0 1506600.0 1966200.0 ;
      RECT  1496400.0 1980000.0 1506600.0 1966200.0 ;
      RECT  1496400.0 1980000.0 1506600.0 1993800.0 ;
      RECT  1496400.0 2007600.0 1506600.0 1993800.0 ;
      RECT  1496400.0 2007600.0 1506600.0 2021400.0 ;
      RECT  1496400.0 2035200.0 1506600.0 2021400.0 ;
      RECT  1496400.0 2035200.0 1506600.0 2049000.0 ;
      RECT  1496400.0 2062800.0 1506600.0 2049000.0 ;
      RECT  1496400.0 2062800.0 1506600.0 2076600.0 ;
      RECT  1496400.0 2090400.0 1506600.0 2076600.0 ;
      RECT  1496400.0 2090400.0 1506600.0 2104200.0 ;
      RECT  1496400.0 2118000.0 1506600.0 2104200.0 ;
      RECT  1496400.0 2118000.0 1506600.0 2131800.0 ;
      RECT  1496400.0 2145600.0 1506600.0 2131800.0 ;
      RECT  1506600.0 379200.0 1516800.0 393000.0 ;
      RECT  1506600.0 406800.0 1516800.0 393000.0 ;
      RECT  1506600.0 406800.0 1516800.0 420600.0 ;
      RECT  1506600.0 434400.0 1516800.0 420600.0 ;
      RECT  1506600.0 434400.0 1516800.0 448200.0 ;
      RECT  1506600.0 462000.0 1516800.0 448200.0 ;
      RECT  1506600.0 462000.0 1516800.0 475800.0 ;
      RECT  1506600.0 489600.0 1516800.0 475800.0 ;
      RECT  1506600.0 489600.0 1516800.0 503400.0 ;
      RECT  1506600.0 517200.0 1516800.0 503400.0 ;
      RECT  1506600.0 517200.0 1516800.0 531000.0 ;
      RECT  1506600.0 544800.0 1516800.0 531000.0 ;
      RECT  1506600.0 544800.0 1516800.0 558600.0 ;
      RECT  1506600.0 572400.0 1516800.0 558600.0 ;
      RECT  1506600.0 572400.0 1516800.0 586200.0 ;
      RECT  1506600.0 600000.0 1516800.0 586200.0 ;
      RECT  1506600.0 600000.0 1516800.0 613800.0 ;
      RECT  1506600.0 627600.0 1516800.0 613800.0 ;
      RECT  1506600.0 627600.0 1516800.0 641400.0 ;
      RECT  1506600.0 655200.0 1516800.0 641400.0 ;
      RECT  1506600.0 655200.0 1516800.0 669000.0 ;
      RECT  1506600.0 682800.0 1516800.0 669000.0 ;
      RECT  1506600.0 682800.0 1516800.0 696600.0 ;
      RECT  1506600.0 710400.0 1516800.0 696600.0 ;
      RECT  1506600.0 710400.0 1516800.0 724200.0 ;
      RECT  1506600.0 738000.0 1516800.0 724200.0 ;
      RECT  1506600.0 738000.0 1516800.0 751800.0 ;
      RECT  1506600.0 765600.0 1516800.0 751800.0 ;
      RECT  1506600.0 765600.0 1516800.0 779400.0 ;
      RECT  1506600.0 793200.0 1516800.0 779400.0 ;
      RECT  1506600.0 793200.0 1516800.0 807000.0 ;
      RECT  1506600.0 820800.0 1516800.0 807000.0 ;
      RECT  1506600.0 820800.0 1516800.0 834600.0 ;
      RECT  1506600.0 848400.0 1516800.0 834600.0 ;
      RECT  1506600.0 848400.0 1516800.0 862200.0 ;
      RECT  1506600.0 876000.0 1516800.0 862200.0 ;
      RECT  1506600.0 876000.0 1516800.0 889800.0 ;
      RECT  1506600.0 903600.0 1516800.0 889800.0 ;
      RECT  1506600.0 903600.0 1516800.0 917400.0 ;
      RECT  1506600.0 931200.0 1516800.0 917400.0 ;
      RECT  1506600.0 931200.0 1516800.0 945000.0 ;
      RECT  1506600.0 958800.0 1516800.0 945000.0 ;
      RECT  1506600.0 958800.0 1516800.0 972600.0 ;
      RECT  1506600.0 986400.0 1516800.0 972600.0 ;
      RECT  1506600.0 986400.0 1516800.0 1000200.0 ;
      RECT  1506600.0 1014000.0 1516800.0 1000200.0 ;
      RECT  1506600.0 1014000.0 1516800.0 1027800.0 ;
      RECT  1506600.0 1041600.0 1516800.0 1027800.0 ;
      RECT  1506600.0 1041600.0 1516800.0 1055400.0 ;
      RECT  1506600.0 1069200.0 1516800.0 1055400.0 ;
      RECT  1506600.0 1069200.0 1516800.0 1083000.0 ;
      RECT  1506600.0 1096800.0 1516800.0 1083000.0 ;
      RECT  1506600.0 1096800.0 1516800.0 1110600.0 ;
      RECT  1506600.0 1124400.0 1516800.0 1110600.0 ;
      RECT  1506600.0 1124400.0 1516800.0 1138200.0 ;
      RECT  1506600.0 1152000.0 1516800.0 1138200.0 ;
      RECT  1506600.0 1152000.0 1516800.0 1165800.0 ;
      RECT  1506600.0 1179600.0 1516800.0 1165800.0 ;
      RECT  1506600.0 1179600.0 1516800.0 1193400.0 ;
      RECT  1506600.0 1207200.0 1516800.0 1193400.0 ;
      RECT  1506600.0 1207200.0 1516800.0 1221000.0 ;
      RECT  1506600.0 1234800.0 1516800.0 1221000.0 ;
      RECT  1506600.0 1234800.0 1516800.0 1248600.0 ;
      RECT  1506600.0 1262400.0 1516800.0 1248600.0 ;
      RECT  1506600.0 1262400.0 1516800.0 1276200.0 ;
      RECT  1506600.0 1290000.0 1516800.0 1276200.0 ;
      RECT  1506600.0 1290000.0 1516800.0 1303800.0 ;
      RECT  1506600.0 1317600.0 1516800.0 1303800.0 ;
      RECT  1506600.0 1317600.0 1516800.0 1331400.0 ;
      RECT  1506600.0 1345200.0 1516800.0 1331400.0 ;
      RECT  1506600.0 1345200.0 1516800.0 1359000.0 ;
      RECT  1506600.0 1372800.0 1516800.0 1359000.0 ;
      RECT  1506600.0 1372800.0 1516800.0 1386600.0 ;
      RECT  1506600.0 1400400.0 1516800.0 1386600.0 ;
      RECT  1506600.0 1400400.0 1516800.0 1414200.0 ;
      RECT  1506600.0 1428000.0 1516800.0 1414200.0 ;
      RECT  1506600.0 1428000.0 1516800.0 1441800.0 ;
      RECT  1506600.0 1455600.0 1516800.0 1441800.0 ;
      RECT  1506600.0 1455600.0 1516800.0 1469400.0 ;
      RECT  1506600.0 1483200.0 1516800.0 1469400.0 ;
      RECT  1506600.0 1483200.0 1516800.0 1497000.0 ;
      RECT  1506600.0 1510800.0 1516800.0 1497000.0 ;
      RECT  1506600.0 1510800.0 1516800.0 1524600.0 ;
      RECT  1506600.0 1538400.0 1516800.0 1524600.0 ;
      RECT  1506600.0 1538400.0 1516800.0 1552200.0 ;
      RECT  1506600.0 1566000.0 1516800.0 1552200.0 ;
      RECT  1506600.0 1566000.0 1516800.0 1579800.0 ;
      RECT  1506600.0 1593600.0 1516800.0 1579800.0 ;
      RECT  1506600.0 1593600.0 1516800.0 1607400.0 ;
      RECT  1506600.0 1621200.0 1516800.0 1607400.0 ;
      RECT  1506600.0 1621200.0 1516800.0 1635000.0 ;
      RECT  1506600.0 1648800.0 1516800.0 1635000.0 ;
      RECT  1506600.0 1648800.0 1516800.0 1662600.0 ;
      RECT  1506600.0 1676400.0 1516800.0 1662600.0 ;
      RECT  1506600.0 1676400.0 1516800.0 1690200.0 ;
      RECT  1506600.0 1704000.0 1516800.0 1690200.0 ;
      RECT  1506600.0 1704000.0 1516800.0 1717800.0 ;
      RECT  1506600.0 1731600.0 1516800.0 1717800.0 ;
      RECT  1506600.0 1731600.0 1516800.0 1745400.0 ;
      RECT  1506600.0 1759200.0 1516800.0 1745400.0 ;
      RECT  1506600.0 1759200.0 1516800.0 1773000.0 ;
      RECT  1506600.0 1786800.0 1516800.0 1773000.0 ;
      RECT  1506600.0 1786800.0 1516800.0 1800600.0 ;
      RECT  1506600.0 1814400.0 1516800.0 1800600.0 ;
      RECT  1506600.0 1814400.0 1516800.0 1828200.0 ;
      RECT  1506600.0 1842000.0 1516800.0 1828200.0 ;
      RECT  1506600.0 1842000.0 1516800.0 1855800.0 ;
      RECT  1506600.0 1869600.0 1516800.0 1855800.0 ;
      RECT  1506600.0 1869600.0 1516800.0 1883400.0 ;
      RECT  1506600.0 1897200.0 1516800.0 1883400.0 ;
      RECT  1506600.0 1897200.0 1516800.0 1911000.0 ;
      RECT  1506600.0 1924800.0 1516800.0 1911000.0 ;
      RECT  1506600.0 1924800.0 1516800.0 1938600.0 ;
      RECT  1506600.0 1952400.0 1516800.0 1938600.0 ;
      RECT  1506600.0 1952400.0 1516800.0 1966200.0 ;
      RECT  1506600.0 1980000.0 1516800.0 1966200.0 ;
      RECT  1506600.0 1980000.0 1516800.0 1993800.0 ;
      RECT  1506600.0 2007600.0 1516800.0 1993800.0 ;
      RECT  1506600.0 2007600.0 1516800.0 2021400.0 ;
      RECT  1506600.0 2035200.0 1516800.0 2021400.0 ;
      RECT  1506600.0 2035200.0 1516800.0 2049000.0 ;
      RECT  1506600.0 2062800.0 1516800.0 2049000.0 ;
      RECT  1506600.0 2062800.0 1516800.0 2076600.0 ;
      RECT  1506600.0 2090400.0 1516800.0 2076600.0 ;
      RECT  1506600.0 2090400.0 1516800.0 2104200.0 ;
      RECT  1506600.0 2118000.0 1516800.0 2104200.0 ;
      RECT  1506600.0 2118000.0 1516800.0 2131800.0 ;
      RECT  1506600.0 2145600.0 1516800.0 2131800.0 ;
      RECT  1516800.0 379200.0 1527000.0 393000.0 ;
      RECT  1516800.0 406800.0 1527000.0 393000.0 ;
      RECT  1516800.0 406800.0 1527000.0 420600.0 ;
      RECT  1516800.0 434400.0 1527000.0 420600.0 ;
      RECT  1516800.0 434400.0 1527000.0 448200.0 ;
      RECT  1516800.0 462000.0 1527000.0 448200.0 ;
      RECT  1516800.0 462000.0 1527000.0 475800.0 ;
      RECT  1516800.0 489600.0 1527000.0 475800.0 ;
      RECT  1516800.0 489600.0 1527000.0 503400.0 ;
      RECT  1516800.0 517200.0 1527000.0 503400.0 ;
      RECT  1516800.0 517200.0 1527000.0 531000.0 ;
      RECT  1516800.0 544800.0 1527000.0 531000.0 ;
      RECT  1516800.0 544800.0 1527000.0 558600.0 ;
      RECT  1516800.0 572400.0 1527000.0 558600.0 ;
      RECT  1516800.0 572400.0 1527000.0 586200.0 ;
      RECT  1516800.0 600000.0 1527000.0 586200.0 ;
      RECT  1516800.0 600000.0 1527000.0 613800.0 ;
      RECT  1516800.0 627600.0 1527000.0 613800.0 ;
      RECT  1516800.0 627600.0 1527000.0 641400.0 ;
      RECT  1516800.0 655200.0 1527000.0 641400.0 ;
      RECT  1516800.0 655200.0 1527000.0 669000.0 ;
      RECT  1516800.0 682800.0 1527000.0 669000.0 ;
      RECT  1516800.0 682800.0 1527000.0 696600.0 ;
      RECT  1516800.0 710400.0 1527000.0 696600.0 ;
      RECT  1516800.0 710400.0 1527000.0 724200.0 ;
      RECT  1516800.0 738000.0 1527000.0 724200.0 ;
      RECT  1516800.0 738000.0 1527000.0 751800.0 ;
      RECT  1516800.0 765600.0 1527000.0 751800.0 ;
      RECT  1516800.0 765600.0 1527000.0 779400.0 ;
      RECT  1516800.0 793200.0 1527000.0 779400.0 ;
      RECT  1516800.0 793200.0 1527000.0 807000.0 ;
      RECT  1516800.0 820800.0 1527000.0 807000.0 ;
      RECT  1516800.0 820800.0 1527000.0 834600.0 ;
      RECT  1516800.0 848400.0 1527000.0 834600.0 ;
      RECT  1516800.0 848400.0 1527000.0 862200.0 ;
      RECT  1516800.0 876000.0 1527000.0 862200.0 ;
      RECT  1516800.0 876000.0 1527000.0 889800.0 ;
      RECT  1516800.0 903600.0 1527000.0 889800.0 ;
      RECT  1516800.0 903600.0 1527000.0 917400.0 ;
      RECT  1516800.0 931200.0 1527000.0 917400.0 ;
      RECT  1516800.0 931200.0 1527000.0 945000.0 ;
      RECT  1516800.0 958800.0 1527000.0 945000.0 ;
      RECT  1516800.0 958800.0 1527000.0 972600.0 ;
      RECT  1516800.0 986400.0 1527000.0 972600.0 ;
      RECT  1516800.0 986400.0 1527000.0 1000200.0 ;
      RECT  1516800.0 1014000.0 1527000.0 1000200.0 ;
      RECT  1516800.0 1014000.0 1527000.0 1027800.0 ;
      RECT  1516800.0 1041600.0 1527000.0 1027800.0 ;
      RECT  1516800.0 1041600.0 1527000.0 1055400.0 ;
      RECT  1516800.0 1069200.0 1527000.0 1055400.0 ;
      RECT  1516800.0 1069200.0 1527000.0 1083000.0 ;
      RECT  1516800.0 1096800.0 1527000.0 1083000.0 ;
      RECT  1516800.0 1096800.0 1527000.0 1110600.0 ;
      RECT  1516800.0 1124400.0 1527000.0 1110600.0 ;
      RECT  1516800.0 1124400.0 1527000.0 1138200.0 ;
      RECT  1516800.0 1152000.0 1527000.0 1138200.0 ;
      RECT  1516800.0 1152000.0 1527000.0 1165800.0 ;
      RECT  1516800.0 1179600.0 1527000.0 1165800.0 ;
      RECT  1516800.0 1179600.0 1527000.0 1193400.0 ;
      RECT  1516800.0 1207200.0 1527000.0 1193400.0 ;
      RECT  1516800.0 1207200.0 1527000.0 1221000.0 ;
      RECT  1516800.0 1234800.0 1527000.0 1221000.0 ;
      RECT  1516800.0 1234800.0 1527000.0 1248600.0 ;
      RECT  1516800.0 1262400.0 1527000.0 1248600.0 ;
      RECT  1516800.0 1262400.0 1527000.0 1276200.0 ;
      RECT  1516800.0 1290000.0 1527000.0 1276200.0 ;
      RECT  1516800.0 1290000.0 1527000.0 1303800.0 ;
      RECT  1516800.0 1317600.0 1527000.0 1303800.0 ;
      RECT  1516800.0 1317600.0 1527000.0 1331400.0 ;
      RECT  1516800.0 1345200.0 1527000.0 1331400.0 ;
      RECT  1516800.0 1345200.0 1527000.0 1359000.0 ;
      RECT  1516800.0 1372800.0 1527000.0 1359000.0 ;
      RECT  1516800.0 1372800.0 1527000.0 1386600.0 ;
      RECT  1516800.0 1400400.0 1527000.0 1386600.0 ;
      RECT  1516800.0 1400400.0 1527000.0 1414200.0 ;
      RECT  1516800.0 1428000.0 1527000.0 1414200.0 ;
      RECT  1516800.0 1428000.0 1527000.0 1441800.0 ;
      RECT  1516800.0 1455600.0 1527000.0 1441800.0 ;
      RECT  1516800.0 1455600.0 1527000.0 1469400.0 ;
      RECT  1516800.0 1483200.0 1527000.0 1469400.0 ;
      RECT  1516800.0 1483200.0 1527000.0 1497000.0 ;
      RECT  1516800.0 1510800.0 1527000.0 1497000.0 ;
      RECT  1516800.0 1510800.0 1527000.0 1524600.0 ;
      RECT  1516800.0 1538400.0 1527000.0 1524600.0 ;
      RECT  1516800.0 1538400.0 1527000.0 1552200.0 ;
      RECT  1516800.0 1566000.0 1527000.0 1552200.0 ;
      RECT  1516800.0 1566000.0 1527000.0 1579800.0 ;
      RECT  1516800.0 1593600.0 1527000.0 1579800.0 ;
      RECT  1516800.0 1593600.0 1527000.0 1607400.0 ;
      RECT  1516800.0 1621200.0 1527000.0 1607400.0 ;
      RECT  1516800.0 1621200.0 1527000.0 1635000.0 ;
      RECT  1516800.0 1648800.0 1527000.0 1635000.0 ;
      RECT  1516800.0 1648800.0 1527000.0 1662600.0 ;
      RECT  1516800.0 1676400.0 1527000.0 1662600.0 ;
      RECT  1516800.0 1676400.0 1527000.0 1690200.0 ;
      RECT  1516800.0 1704000.0 1527000.0 1690200.0 ;
      RECT  1516800.0 1704000.0 1527000.0 1717800.0 ;
      RECT  1516800.0 1731600.0 1527000.0 1717800.0 ;
      RECT  1516800.0 1731600.0 1527000.0 1745400.0 ;
      RECT  1516800.0 1759200.0 1527000.0 1745400.0 ;
      RECT  1516800.0 1759200.0 1527000.0 1773000.0 ;
      RECT  1516800.0 1786800.0 1527000.0 1773000.0 ;
      RECT  1516800.0 1786800.0 1527000.0 1800600.0 ;
      RECT  1516800.0 1814400.0 1527000.0 1800600.0 ;
      RECT  1516800.0 1814400.0 1527000.0 1828200.0 ;
      RECT  1516800.0 1842000.0 1527000.0 1828200.0 ;
      RECT  1516800.0 1842000.0 1527000.0 1855800.0 ;
      RECT  1516800.0 1869600.0 1527000.0 1855800.0 ;
      RECT  1516800.0 1869600.0 1527000.0 1883400.0 ;
      RECT  1516800.0 1897200.0 1527000.0 1883400.0 ;
      RECT  1516800.0 1897200.0 1527000.0 1911000.0 ;
      RECT  1516800.0 1924800.0 1527000.0 1911000.0 ;
      RECT  1516800.0 1924800.0 1527000.0 1938600.0 ;
      RECT  1516800.0 1952400.0 1527000.0 1938600.0 ;
      RECT  1516800.0 1952400.0 1527000.0 1966200.0 ;
      RECT  1516800.0 1980000.0 1527000.0 1966200.0 ;
      RECT  1516800.0 1980000.0 1527000.0 1993800.0 ;
      RECT  1516800.0 2007600.0 1527000.0 1993800.0 ;
      RECT  1516800.0 2007600.0 1527000.0 2021400.0 ;
      RECT  1516800.0 2035200.0 1527000.0 2021400.0 ;
      RECT  1516800.0 2035200.0 1527000.0 2049000.0 ;
      RECT  1516800.0 2062800.0 1527000.0 2049000.0 ;
      RECT  1516800.0 2062800.0 1527000.0 2076600.0 ;
      RECT  1516800.0 2090400.0 1527000.0 2076600.0 ;
      RECT  1516800.0 2090400.0 1527000.0 2104200.0 ;
      RECT  1516800.0 2118000.0 1527000.0 2104200.0 ;
      RECT  1516800.0 2118000.0 1527000.0 2131800.0 ;
      RECT  1516800.0 2145600.0 1527000.0 2131800.0 ;
      RECT  224400.0 379800.0 225600.0 2149200.0 ;
      RECT  227400.0 378600.0 228600.0 2148000.0 ;
      RECT  234600.0 379800.0 235800.0 2149200.0 ;
      RECT  237600.0 378600.0 238800.0 2148000.0 ;
      RECT  244800.0 379800.0 246000.0 2149200.0 ;
      RECT  247800.0 378600.0 249000.0 2148000.0 ;
      RECT  255000.0 379800.0 256200.0 2149200.0 ;
      RECT  258000.0 378600.0 259200.0 2148000.0 ;
      RECT  265200.0 379800.0 266400.0 2149200.0 ;
      RECT  268200.0 378600.0 269400.0 2148000.0 ;
      RECT  275400.0 379800.0 276600.0 2149200.0 ;
      RECT  278400.0 378600.0 279600.0 2148000.0 ;
      RECT  285600.0 379800.0 286800.0 2149200.0 ;
      RECT  288600.0 378600.0 289800.0 2148000.0 ;
      RECT  295800.0 379800.0 297000.0 2149200.0 ;
      RECT  298800.0 378600.0 300000.0 2148000.0 ;
      RECT  306000.0 379800.0 307200.0 2149200.0 ;
      RECT  309000.0 378600.0 310200.0 2148000.0 ;
      RECT  316200.0 379800.0 317400.0 2149200.0 ;
      RECT  319200.0 378600.0 320400.0 2148000.0 ;
      RECT  326400.0 379800.0 327600.0 2149200.0 ;
      RECT  329400.0 378600.0 330600.0 2148000.0 ;
      RECT  336600.0 379800.0 337800.0 2149200.0 ;
      RECT  339600.0 378600.0 340800.0 2148000.0 ;
      RECT  346800.0 379800.0 348000.0 2149200.0 ;
      RECT  349800.0 378600.0 351000.0 2148000.0 ;
      RECT  357000.0 379800.0 358200.0 2149200.0 ;
      RECT  360000.0 378600.0 361200.0 2148000.0 ;
      RECT  367200.0 379800.0 368400.0 2149200.0 ;
      RECT  370200.0 378600.0 371400.0 2148000.0 ;
      RECT  377400.0 379800.0 378600.0 2149200.0 ;
      RECT  380400.0 378600.0 381600.0 2148000.0 ;
      RECT  387600.0 379800.0 388800.0 2149200.0 ;
      RECT  390600.0 378600.0 391800.0 2148000.0 ;
      RECT  397800.0 379800.0 399000.0 2149200.0 ;
      RECT  400800.0 378600.0 402000.0 2148000.0 ;
      RECT  408000.0 379800.0 409200.0 2149200.0 ;
      RECT  411000.0 378600.0 412200.0 2148000.0 ;
      RECT  418200.0 379800.0 419400.0 2149200.0 ;
      RECT  421200.0 378600.0 422400.0 2148000.0 ;
      RECT  428400.0 379800.0 429600.0 2149200.0 ;
      RECT  431400.0 378600.0 432600.0 2148000.0 ;
      RECT  438600.0 379800.0 439800.0 2149200.0 ;
      RECT  441600.0 378600.0 442800.0 2148000.0 ;
      RECT  448800.0 379800.0 450000.0 2149200.0 ;
      RECT  451800.0 378600.0 453000.0 2148000.0 ;
      RECT  459000.0 379800.0 460200.0 2149200.0 ;
      RECT  462000.0 378600.0 463200.0 2148000.0 ;
      RECT  469200.0 379800.0 470400.0 2149200.0 ;
      RECT  472200.0 378600.0 473400.0 2148000.0 ;
      RECT  479400.0 379800.0 480600.0 2149200.0 ;
      RECT  482400.0 378600.0 483600.0 2148000.0 ;
      RECT  489600.0 379800.0 490800.0 2149200.0 ;
      RECT  492600.0 378600.0 493800.0 2148000.0 ;
      RECT  499800.0 379800.0 501000.0 2149200.0 ;
      RECT  502800.0 378600.0 504000.0 2148000.0 ;
      RECT  510000.0 379800.0 511200.0 2149200.0 ;
      RECT  513000.0 378600.0 514200.0 2148000.0 ;
      RECT  520200.0 379800.0 521400.0 2149200.0 ;
      RECT  523200.0 378600.0 524400.0 2148000.0 ;
      RECT  530400.0 379800.0 531600.0 2149200.0 ;
      RECT  533400.0 378600.0 534600.0 2148000.0 ;
      RECT  540600.0 379800.0 541800.0 2149200.0 ;
      RECT  543600.0 378600.0 544800.0 2148000.0 ;
      RECT  550800.0 379800.0 552000.0 2149200.0 ;
      RECT  553800.0 378600.0 555000.0 2148000.0 ;
      RECT  561000.0 379800.0 562200.0 2149200.0 ;
      RECT  564000.0 378600.0 565200.0 2148000.0 ;
      RECT  571200.0 379800.0 572400.0 2149200.0 ;
      RECT  574200.0 378600.0 575400.0 2148000.0 ;
      RECT  581400.0 379800.0 582600.0 2149200.0 ;
      RECT  584400.0 378600.0 585600.0 2148000.0 ;
      RECT  591600.0 379800.0 592800.0 2149200.0 ;
      RECT  594600.0 378600.0 595800.0 2148000.0 ;
      RECT  601800.0 379800.0 603000.0 2149200.0 ;
      RECT  604800.0 378600.0 606000.0 2148000.0 ;
      RECT  612000.0 379800.0 613200.0 2149200.0 ;
      RECT  615000.0 378600.0 616200.0 2148000.0 ;
      RECT  622200.0 379800.0 623400.0 2149200.0 ;
      RECT  625200.0 378600.0 626400.0 2148000.0 ;
      RECT  632400.0 379800.0 633600.0 2149200.0 ;
      RECT  635400.0 378600.0 636600.0 2148000.0 ;
      RECT  642600.0 379800.0 643800.0 2149200.0 ;
      RECT  645600.0 378600.0 646800.0 2148000.0 ;
      RECT  652800.0 379800.0 654000.0 2149200.0 ;
      RECT  655800.0 378600.0 657000.0 2148000.0 ;
      RECT  663000.0 379800.0 664200.0 2149200.0 ;
      RECT  666000.0 378600.0 667200.0 2148000.0 ;
      RECT  673200.0 379800.0 674400.0 2149200.0 ;
      RECT  676200.0 378600.0 677400.0 2148000.0 ;
      RECT  683400.0 379800.0 684600.0 2149200.0 ;
      RECT  686400.0 378600.0 687600.0 2148000.0 ;
      RECT  693600.0 379800.0 694800.0 2149200.0 ;
      RECT  696600.0 378600.0 697800.0 2148000.0 ;
      RECT  703800.0 379800.0 705000.0 2149200.0 ;
      RECT  706800.0 378600.0 708000.0 2148000.0 ;
      RECT  714000.0 379800.0 715200.0 2149200.0 ;
      RECT  717000.0 378600.0 718200.0 2148000.0 ;
      RECT  724200.0 379800.0 725400.0 2149200.0 ;
      RECT  727200.0 378600.0 728400.0 2148000.0 ;
      RECT  734400.0 379800.0 735600.0 2149200.0 ;
      RECT  737400.0 378600.0 738600.0 2148000.0 ;
      RECT  744600.0 379800.0 745800.0 2149200.0 ;
      RECT  747600.0 378600.0 748800.0 2148000.0 ;
      RECT  754800.0 379800.0 756000.0 2149200.0 ;
      RECT  757800.0 378600.0 759000.0 2148000.0 ;
      RECT  765000.0 379800.0 766200.0 2149200.0 ;
      RECT  768000.0 378600.0 769200.0 2148000.0 ;
      RECT  775200.0 379800.0 776400.0 2149200.0 ;
      RECT  778200.0 378600.0 779400.0 2148000.0 ;
      RECT  785400.0 379800.0 786600.0 2149200.0 ;
      RECT  788400.0 378600.0 789600.0 2148000.0 ;
      RECT  795600.0 379800.0 796800.0 2149200.0 ;
      RECT  798600.0 378600.0 799800.0 2148000.0 ;
      RECT  805800.0 379800.0 807000.0 2149200.0 ;
      RECT  808800.0 378600.0 810000.0 2148000.0 ;
      RECT  816000.0 379800.0 817200.0 2149200.0 ;
      RECT  819000.0 378600.0 820200.0 2148000.0 ;
      RECT  826200.0 379800.0 827400.0 2149200.0 ;
      RECT  829200.0 378600.0 830400.0 2148000.0 ;
      RECT  836400.0 379800.0 837600.0 2149200.0 ;
      RECT  839400.0 378600.0 840600.0 2148000.0 ;
      RECT  846600.0 379800.0 847800.0 2149200.0 ;
      RECT  849600.0 378600.0 850800.0 2148000.0 ;
      RECT  856800.0 379800.0 858000.0 2149200.0 ;
      RECT  859800.0 378600.0 861000.0 2148000.0 ;
      RECT  867000.0 379800.0 868200.0 2149200.0 ;
      RECT  870000.0 378600.0 871200.0 2148000.0 ;
      RECT  877200.0 379800.0 878400.0 2149200.0 ;
      RECT  880200.0 378600.0 881400.0 2148000.0 ;
      RECT  887400.0 379800.0 888600.0 2149200.0 ;
      RECT  890400.0 378600.0 891600.0 2148000.0 ;
      RECT  897600.0 379800.0 898800.0 2149200.0 ;
      RECT  900600.0 378600.0 901800.0 2148000.0 ;
      RECT  907800.0 379800.0 909000.0 2149200.0 ;
      RECT  910800.0 378600.0 912000.0 2148000.0 ;
      RECT  918000.0 379800.0 919200.0 2149200.0 ;
      RECT  921000.0 378600.0 922200.0 2148000.0 ;
      RECT  928200.0 379800.0 929400.0 2149200.0 ;
      RECT  931200.0 378600.0 932400.0 2148000.0 ;
      RECT  938400.0 379800.0 939600.0 2149200.0 ;
      RECT  941400.0 378600.0 942600.0 2148000.0 ;
      RECT  948600.0 379800.0 949800.0 2149200.0 ;
      RECT  951600.0 378600.0 952800.0 2148000.0 ;
      RECT  958800.0 379800.0 960000.0 2149200.0 ;
      RECT  961800.0 378600.0 963000.0 2148000.0 ;
      RECT  969000.0 379800.0 970200.0 2149200.0 ;
      RECT  972000.0 378600.0 973200.0 2148000.0 ;
      RECT  979200.0 379800.0 980400.0 2149200.0 ;
      RECT  982200.0 378600.0 983400.0 2148000.0 ;
      RECT  989400.0 379800.0 990600.0 2149200.0 ;
      RECT  992400.0 378600.0 993600.0 2148000.0 ;
      RECT  999600.0 379800.0 1000800.0 2149200.0 ;
      RECT  1002600.0 378600.0 1003800.0 2148000.0 ;
      RECT  1009800.0 379800.0 1011000.0 2149200.0 ;
      RECT  1012800.0 378600.0 1014000.0 2148000.0 ;
      RECT  1020000.0 379800.0 1021200.0 2149200.0 ;
      RECT  1023000.0 378600.0 1024200.0 2148000.0 ;
      RECT  1030200.0 379800.0 1031400.0 2149200.0 ;
      RECT  1033200.0 378600.0 1034400.0 2148000.0 ;
      RECT  1040400.0 379800.0 1041600.0 2149200.0 ;
      RECT  1043400.0 378600.0 1044600.0 2148000.0 ;
      RECT  1050600.0 379800.0 1051800.0 2149200.0 ;
      RECT  1053600.0 378600.0 1054800.0 2148000.0 ;
      RECT  1060800.0 379800.0 1062000.0 2149200.0 ;
      RECT  1063800.0 378600.0 1065000.0 2148000.0 ;
      RECT  1071000.0 379800.0 1072200.0 2149200.0 ;
      RECT  1074000.0 378600.0 1075200.0 2148000.0 ;
      RECT  1081200.0 379800.0 1082400.0 2149200.0 ;
      RECT  1084200.0 378600.0 1085400.0 2148000.0 ;
      RECT  1091400.0 379800.0 1092600.0 2149200.0 ;
      RECT  1094400.0 378600.0 1095600.0 2148000.0 ;
      RECT  1101600.0 379800.0 1102800.0 2149200.0 ;
      RECT  1104600.0 378600.0 1105800.0 2148000.0 ;
      RECT  1111800.0 379800.0 1113000.0 2149200.0 ;
      RECT  1114800.0 378600.0 1116000.0 2148000.0 ;
      RECT  1122000.0 379800.0 1123200.0 2149200.0 ;
      RECT  1125000.0 378600.0 1126200.0 2148000.0 ;
      RECT  1132200.0 379800.0 1133400.0 2149200.0 ;
      RECT  1135200.0 378600.0 1136400.0 2148000.0 ;
      RECT  1142400.0 379800.0 1143600.0 2149200.0 ;
      RECT  1145400.0 378600.0 1146600.0 2148000.0 ;
      RECT  1152600.0 379800.0 1153800.0 2149200.0 ;
      RECT  1155600.0 378600.0 1156800.0 2148000.0 ;
      RECT  1162800.0 379800.0 1164000.0 2149200.0 ;
      RECT  1165800.0 378600.0 1167000.0 2148000.0 ;
      RECT  1173000.0 379800.0 1174200.0 2149200.0 ;
      RECT  1176000.0 378600.0 1177200.0 2148000.0 ;
      RECT  1183200.0 379800.0 1184400.0 2149200.0 ;
      RECT  1186200.0 378600.0 1187400.0 2148000.0 ;
      RECT  1193400.0 379800.0 1194600.0 2149200.0 ;
      RECT  1196400.0 378600.0 1197600.0 2148000.0 ;
      RECT  1203600.0 379800.0 1204800.0 2149200.0 ;
      RECT  1206600.0 378600.0 1207800.0 2148000.0 ;
      RECT  1213800.0 379800.0 1215000.0 2149200.0 ;
      RECT  1216800.0 378600.0 1218000.0 2148000.0 ;
      RECT  1224000.0 379800.0 1225200.0 2149200.0 ;
      RECT  1227000.0 378600.0 1228200.0 2148000.0 ;
      RECT  1234200.0 379800.0 1235400.0 2149200.0 ;
      RECT  1237200.0 378600.0 1238400.0 2148000.0 ;
      RECT  1244400.0 379800.0 1245600.0 2149200.0 ;
      RECT  1247400.0 378600.0 1248600.0 2148000.0 ;
      RECT  1254600.0 379800.0 1255800.0 2149200.0 ;
      RECT  1257600.0 378600.0 1258800.0 2148000.0 ;
      RECT  1264800.0 379800.0 1266000.0 2149200.0 ;
      RECT  1267800.0 378600.0 1269000.0 2148000.0 ;
      RECT  1275000.0 379800.0 1276200.0 2149200.0 ;
      RECT  1278000.0 378600.0 1279200.0 2148000.0 ;
      RECT  1285200.0 379800.0 1286400.0 2149200.0 ;
      RECT  1288200.0 378600.0 1289400.0 2148000.0 ;
      RECT  1295400.0 379800.0 1296600.0 2149200.0 ;
      RECT  1298400.0 378600.0 1299600.0 2148000.0 ;
      RECT  1305600.0 379800.0 1306800.0 2149200.0 ;
      RECT  1308600.0 378600.0 1309800.0 2148000.0 ;
      RECT  1315800.0 379800.0 1317000.0 2149200.0 ;
      RECT  1318800.0 378600.0 1320000.0 2148000.0 ;
      RECT  1326000.0 379800.0 1327200.0 2149200.0 ;
      RECT  1329000.0 378600.0 1330200.0 2148000.0 ;
      RECT  1336200.0 379800.0 1337400.0 2149200.0 ;
      RECT  1339200.0 378600.0 1340400.0 2148000.0 ;
      RECT  1346400.0 379800.0 1347600.0 2149200.0 ;
      RECT  1349400.0 378600.0 1350600.0 2148000.0 ;
      RECT  1356600.0 379800.0 1357800.0 2149200.0 ;
      RECT  1359600.0 378600.0 1360800.0 2148000.0 ;
      RECT  1366800.0 379800.0 1368000.0 2149200.0 ;
      RECT  1369800.0 378600.0 1371000.0 2148000.0 ;
      RECT  1377000.0 379800.0 1378200.0 2149200.0 ;
      RECT  1380000.0 378600.0 1381200.0 2148000.0 ;
      RECT  1387200.0 379800.0 1388400.0 2149200.0 ;
      RECT  1390200.0 378600.0 1391400.0 2148000.0 ;
      RECT  1397400.0 379800.0 1398600.0 2149200.0 ;
      RECT  1400400.0 378600.0 1401600.0 2148000.0 ;
      RECT  1407600.0 379800.0 1408800.0 2149200.0 ;
      RECT  1410600.0 378600.0 1411800.0 2148000.0 ;
      RECT  1417800.0 379800.0 1419000.0 2149200.0 ;
      RECT  1420800.0 378600.0 1422000.0 2148000.0 ;
      RECT  1428000.0 379800.0 1429200.0 2149200.0 ;
      RECT  1431000.0 378600.0 1432200.0 2148000.0 ;
      RECT  1438200.0 379800.0 1439400.0 2149200.0 ;
      RECT  1441200.0 378600.0 1442400.0 2148000.0 ;
      RECT  1448400.0 379800.0 1449600.0 2149200.0 ;
      RECT  1451400.0 378600.0 1452600.0 2148000.0 ;
      RECT  1458600.0 379800.0 1459800.0 2149200.0 ;
      RECT  1461600.0 378600.0 1462800.0 2148000.0 ;
      RECT  1468800.0 379800.0 1470000.0 2149200.0 ;
      RECT  1471800.0 378600.0 1473000.0 2148000.0 ;
      RECT  1479000.0 379800.0 1480200.0 2149200.0 ;
      RECT  1482000.0 378600.0 1483200.0 2148000.0 ;
      RECT  1489200.0 379800.0 1490400.0 2149200.0 ;
      RECT  1492200.0 378600.0 1493400.0 2148000.0 ;
      RECT  1499400.0 379800.0 1500600.0 2149200.0 ;
      RECT  1502400.0 378600.0 1503600.0 2148000.0 ;
      RECT  1509600.0 379800.0 1510800.0 2149200.0 ;
      RECT  1512600.0 378600.0 1513800.0 2148000.0 ;
      RECT  1519800.0 379800.0 1521000.0 2149200.0 ;
      RECT  1522800.0 378600.0 1524000.0 2148000.0 ;
      RECT  220800.0 378600.0 222000.0 2148000.0 ;
      RECT  231000.0 378600.0 232200.0 2148000.0 ;
      RECT  241200.0 378600.0 242400.0 2148000.0 ;
      RECT  251400.0 378600.0 252600.0 2148000.0 ;
      RECT  261600.0 378600.0 262800.0 2148000.0 ;
      RECT  271800.0 378600.0 273000.0 2148000.0 ;
      RECT  282000.0 378600.0 283200.0 2148000.0 ;
      RECT  292200.0 378600.0 293400.0 2148000.0 ;
      RECT  302400.0 378600.0 303600.0 2148000.0 ;
      RECT  312600.0 378600.0 313800.0 2148000.0 ;
      RECT  322800.0 378600.0 324000.0 2148000.0 ;
      RECT  333000.0 378600.0 334200.0 2148000.0 ;
      RECT  343200.0 378600.0 344400.0 2148000.0 ;
      RECT  353400.0 378600.0 354600.0 2148000.0 ;
      RECT  363600.0 378600.0 364800.0 2148000.0 ;
      RECT  373800.0 378600.0 375000.0 2148000.0 ;
      RECT  384000.0 378600.0 385200.0 2148000.0 ;
      RECT  394200.0 378600.0 395400.0 2148000.0 ;
      RECT  404400.0 378600.0 405600.0 2148000.0 ;
      RECT  414600.0 378600.0 415800.0 2148000.0 ;
      RECT  424800.0 378600.0 426000.0 2148000.0 ;
      RECT  435000.0 378600.0 436200.0 2148000.0 ;
      RECT  445200.0 378600.0 446400.0 2148000.0 ;
      RECT  455400.0 378600.0 456600.0 2148000.0 ;
      RECT  465600.0 378600.0 466800.0 2148000.0 ;
      RECT  475800.0 378600.0 477000.0 2148000.0 ;
      RECT  486000.0 378600.0 487200.0 2148000.0 ;
      RECT  496200.0 378600.0 497400.0 2148000.0 ;
      RECT  506400.0 378600.0 507600.0 2148000.0 ;
      RECT  516600.0 378600.0 517800.0 2148000.0 ;
      RECT  526800.0 378600.0 528000.0 2148000.0 ;
      RECT  537000.0 378600.0 538200.0 2148000.0 ;
      RECT  547200.0 378600.0 548400.0 2148000.0 ;
      RECT  557400.0 378600.0 558600.0 2148000.0 ;
      RECT  567600.0 378600.0 568800.0 2148000.0 ;
      RECT  577800.0 378600.0 579000.0 2148000.0 ;
      RECT  588000.0 378600.0 589200.0 2148000.0 ;
      RECT  598200.0 378600.0 599400.0 2148000.0 ;
      RECT  608400.0 378600.0 609600.0 2148000.0 ;
      RECT  618600.0 378600.0 619800.0 2148000.0 ;
      RECT  628800.0 378600.0 630000.0 2148000.0 ;
      RECT  639000.0 378600.0 640200.0 2148000.0 ;
      RECT  649200.0 378600.0 650400.0 2148000.0 ;
      RECT  659400.0 378600.0 660600.0 2148000.0 ;
      RECT  669600.0 378600.0 670800.0 2148000.0 ;
      RECT  679800.0 378600.0 681000.0 2148000.0 ;
      RECT  690000.0 378600.0 691200.0 2148000.0 ;
      RECT  700200.0 378600.0 701400.0 2148000.0 ;
      RECT  710400.0 378600.0 711600.0 2148000.0 ;
      RECT  720600.0 378600.0 721800.0 2148000.0 ;
      RECT  730800.0 378600.0 732000.0 2148000.0 ;
      RECT  741000.0 378600.0 742200.0 2148000.0 ;
      RECT  751200.0 378600.0 752400.0 2148000.0 ;
      RECT  761400.0 378600.0 762600.0 2148000.0 ;
      RECT  771600.0 378600.0 772800.0 2148000.0 ;
      RECT  781800.0 378600.0 783000.0 2148000.0 ;
      RECT  792000.0 378600.0 793200.0 2148000.0 ;
      RECT  802200.0 378600.0 803400.0 2148000.0 ;
      RECT  812400.0 378600.0 813600.0 2148000.0 ;
      RECT  822600.0 378600.0 823800.0 2148000.0 ;
      RECT  832800.0 378600.0 834000.0 2148000.0 ;
      RECT  843000.0 378600.0 844200.0 2148000.0 ;
      RECT  853200.0 378600.0 854400.0 2148000.0 ;
      RECT  863400.0 378600.0 864600.0 2148000.0 ;
      RECT  873600.0 378600.0 874800.0 2148000.0 ;
      RECT  883800.0 378600.0 885000.0 2148000.0 ;
      RECT  894000.0 378600.0 895200.0 2148000.0 ;
      RECT  904200.0 378600.0 905400.0 2148000.0 ;
      RECT  914400.0 378600.0 915600.0 2148000.0 ;
      RECT  924600.0 378600.0 925800.0 2148000.0 ;
      RECT  934800.0 378600.0 936000.0 2148000.0 ;
      RECT  945000.0 378600.0 946200.0 2148000.0 ;
      RECT  955200.0 378600.0 956400.0 2148000.0 ;
      RECT  965400.0 378600.0 966600.0 2148000.0 ;
      RECT  975600.0 378600.0 976800.0 2148000.0 ;
      RECT  985800.0 378600.0 987000.0 2148000.0 ;
      RECT  996000.0 378600.0 997200.0 2148000.0 ;
      RECT  1006200.0 378600.0 1007400.0 2148000.0 ;
      RECT  1016400.0 378600.0 1017600.0 2148000.0 ;
      RECT  1026600.0 378600.0 1027800.0 2148000.0 ;
      RECT  1036800.0 378600.0 1038000.0 2148000.0 ;
      RECT  1047000.0 378600.0 1048200.0 2148000.0 ;
      RECT  1057200.0 378600.0 1058400.0 2148000.0 ;
      RECT  1067400.0 378600.0 1068600.0 2148000.0 ;
      RECT  1077600.0 378600.0 1078800.0 2148000.0 ;
      RECT  1087800.0 378600.0 1089000.0 2148000.0 ;
      RECT  1098000.0 378600.0 1099200.0 2148000.0 ;
      RECT  1108200.0 378600.0 1109400.0 2148000.0 ;
      RECT  1118400.0 378600.0 1119600.0 2148000.0 ;
      RECT  1128600.0 378600.0 1129800.0 2148000.0 ;
      RECT  1138800.0 378600.0 1140000.0 2148000.0 ;
      RECT  1149000.0 378600.0 1150200.0 2148000.0 ;
      RECT  1159200.0 378600.0 1160400.0 2148000.0 ;
      RECT  1169400.0 378600.0 1170600.0 2148000.0 ;
      RECT  1179600.0 378600.0 1180800.0 2148000.0 ;
      RECT  1189800.0 378600.0 1191000.0 2148000.0 ;
      RECT  1200000.0 378600.0 1201200.0 2148000.0 ;
      RECT  1210200.0 378600.0 1211400.0 2148000.0 ;
      RECT  1220400.0 378600.0 1221600.0 2148000.0 ;
      RECT  1230600.0 378600.0 1231800.0 2148000.0 ;
      RECT  1240800.0 378600.0 1242000.0 2148000.0 ;
      RECT  1251000.0 378600.0 1252200.0 2148000.0 ;
      RECT  1261200.0 378600.0 1262400.0 2148000.0 ;
      RECT  1271400.0 378600.0 1272600.0 2148000.0 ;
      RECT  1281600.0 378600.0 1282800.0 2148000.0 ;
      RECT  1291800.0 378600.0 1293000.0 2148000.0 ;
      RECT  1302000.0 378600.0 1303200.0 2148000.0 ;
      RECT  1312200.0 378600.0 1313400.0 2148000.0 ;
      RECT  1322400.0 378600.0 1323600.0 2148000.0 ;
      RECT  1332600.0 378600.0 1333800.0 2148000.0 ;
      RECT  1342800.0 378600.0 1344000.0 2148000.0 ;
      RECT  1353000.0 378600.0 1354200.0 2148000.0 ;
      RECT  1363200.0 378600.0 1364400.0 2148000.0 ;
      RECT  1373400.0 378600.0 1374600.0 2148000.0 ;
      RECT  1383600.0 378600.0 1384800.0 2148000.0 ;
      RECT  1393800.0 378600.0 1395000.0 2148000.0 ;
      RECT  1404000.0 378600.0 1405200.0 2148000.0 ;
      RECT  1414200.0 378600.0 1415400.0 2148000.0 ;
      RECT  1424400.0 378600.0 1425600.0 2148000.0 ;
      RECT  1434600.0 378600.0 1435800.0 2148000.0 ;
      RECT  1444800.0 378600.0 1446000.0 2148000.0 ;
      RECT  1455000.0 378600.0 1456200.0 2148000.0 ;
      RECT  1465200.0 378600.0 1466400.0 2148000.0 ;
      RECT  1475400.0 378600.0 1476600.0 2148000.0 ;
      RECT  1485600.0 378600.0 1486800.0 2148000.0 ;
      RECT  1495800.0 378600.0 1497000.0 2148000.0 ;
      RECT  1506000.0 378600.0 1507200.0 2148000.0 ;
      RECT  1516200.0 378600.0 1517400.0 2148000.0 ;
      RECT  1526400.0 378600.0 1527600.0 2148000.0 ;
      RECT  224400.0 2151600.0 225600.0 2152800.0 ;
      RECT  226800.0 2151600.0 228450.0 2152800.0 ;
      RECT  224400.0 2158800.0 225600.0 2160000.0 ;
      RECT  227550.0 2158800.0 230400.0 2160000.0 ;
      RECT  224400.0 2151600.0 225600.0 2152800.0 ;
      RECT  226800.0 2151600.0 228000.0 2152800.0 ;
      RECT  224400.0 2158800.0 225600.0 2160000.0 ;
      RECT  229200.0 2158800.0 230400.0 2160000.0 ;
      RECT  224550.0 2149200.0 225450.0 2166000.0 ;
      RECT  227550.0 2149200.0 228450.0 2166000.0 ;
      RECT  234600.0 2151600.0 235800.0 2152800.0 ;
      RECT  237000.0 2151600.0 238650.0 2152800.0 ;
      RECT  234600.0 2158800.0 235800.0 2160000.0 ;
      RECT  237750.0 2158800.0 240600.0 2160000.0 ;
      RECT  234600.0 2151600.0 235800.0 2152800.0 ;
      RECT  237000.0 2151600.0 238200.0 2152800.0 ;
      RECT  234600.0 2158800.0 235800.0 2160000.0 ;
      RECT  239400.0 2158800.0 240600.0 2160000.0 ;
      RECT  234750.0 2149200.0 235650.0 2166000.0 ;
      RECT  237750.0 2149200.0 238650.0 2166000.0 ;
      RECT  244800.0 2151600.0 246000.0 2152800.0 ;
      RECT  247200.0 2151600.0 248850.0 2152800.0 ;
      RECT  244800.0 2158800.0 246000.0 2160000.0 ;
      RECT  247950.0 2158800.0 250800.0 2160000.0 ;
      RECT  244800.0 2151600.0 246000.0 2152800.0 ;
      RECT  247200.0 2151600.0 248400.0 2152800.0 ;
      RECT  244800.0 2158800.0 246000.0 2160000.0 ;
      RECT  249600.0 2158800.0 250800.0 2160000.0 ;
      RECT  244950.0 2149200.0 245850.0 2166000.0 ;
      RECT  247950.0 2149200.0 248850.0 2166000.0 ;
      RECT  255000.0 2151600.0 256200.0 2152800.0 ;
      RECT  257400.0 2151600.0 259050.0 2152800.0 ;
      RECT  255000.0 2158800.0 256200.0 2160000.0 ;
      RECT  258150.0 2158800.0 261000.0 2160000.0 ;
      RECT  255000.0 2151600.0 256200.0 2152800.0 ;
      RECT  257400.0 2151600.0 258600.0 2152800.0 ;
      RECT  255000.0 2158800.0 256200.0 2160000.0 ;
      RECT  259800.0 2158800.0 261000.0 2160000.0 ;
      RECT  255150.0 2149200.0 256050.0 2166000.0 ;
      RECT  258150.0 2149200.0 259050.0 2166000.0 ;
      RECT  265200.0 2151600.0 266400.0 2152800.0 ;
      RECT  267600.0 2151600.0 269250.0 2152800.0 ;
      RECT  265200.0 2158800.0 266400.0 2160000.0 ;
      RECT  268350.0 2158800.0 271200.0 2160000.0 ;
      RECT  265200.0 2151600.0 266400.0 2152800.0 ;
      RECT  267600.0 2151600.0 268800.0 2152800.0 ;
      RECT  265200.0 2158800.0 266400.0 2160000.0 ;
      RECT  270000.0 2158800.0 271200.0 2160000.0 ;
      RECT  265350.0 2149200.0 266250.0 2166000.0 ;
      RECT  268350.0 2149200.0 269250.0 2166000.0 ;
      RECT  275400.0 2151600.0 276600.0 2152800.0 ;
      RECT  277800.0 2151600.0 279450.0 2152800.0 ;
      RECT  275400.0 2158800.0 276600.0 2160000.0 ;
      RECT  278550.0 2158800.0 281400.0 2160000.0 ;
      RECT  275400.0 2151600.0 276600.0 2152800.0 ;
      RECT  277800.0 2151600.0 279000.0 2152800.0 ;
      RECT  275400.0 2158800.0 276600.0 2160000.0 ;
      RECT  280200.0 2158800.0 281400.0 2160000.0 ;
      RECT  275550.0 2149200.0 276450.0 2166000.0 ;
      RECT  278550.0 2149200.0 279450.0 2166000.0 ;
      RECT  285600.0 2151600.0 286800.0 2152800.0 ;
      RECT  288000.0 2151600.0 289650.0 2152800.0 ;
      RECT  285600.0 2158800.0 286800.0 2160000.0 ;
      RECT  288750.0 2158800.0 291600.0 2160000.0 ;
      RECT  285600.0 2151600.0 286800.0 2152800.0 ;
      RECT  288000.0 2151600.0 289200.0 2152800.0 ;
      RECT  285600.0 2158800.0 286800.0 2160000.0 ;
      RECT  290400.0 2158800.0 291600.0 2160000.0 ;
      RECT  285750.0 2149200.0 286650.0 2166000.0 ;
      RECT  288750.0 2149200.0 289650.0 2166000.0 ;
      RECT  295800.0 2151600.0 297000.0 2152800.0 ;
      RECT  298200.0 2151600.0 299850.0 2152800.0 ;
      RECT  295800.0 2158800.0 297000.0 2160000.0 ;
      RECT  298950.0 2158800.0 301800.0 2160000.0 ;
      RECT  295800.0 2151600.0 297000.0 2152800.0 ;
      RECT  298200.0 2151600.0 299400.0 2152800.0 ;
      RECT  295800.0 2158800.0 297000.0 2160000.0 ;
      RECT  300600.0 2158800.0 301800.0 2160000.0 ;
      RECT  295950.0 2149200.0 296850.0 2166000.0 ;
      RECT  298950.0 2149200.0 299850.0 2166000.0 ;
      RECT  306000.0 2151600.0 307200.0 2152800.0 ;
      RECT  308400.0 2151600.0 310050.0 2152800.0 ;
      RECT  306000.0 2158800.0 307200.0 2160000.0 ;
      RECT  309150.0 2158800.0 312000.0 2160000.0 ;
      RECT  306000.0 2151600.0 307200.0 2152800.0 ;
      RECT  308400.0 2151600.0 309600.0 2152800.0 ;
      RECT  306000.0 2158800.0 307200.0 2160000.0 ;
      RECT  310800.0 2158800.0 312000.0 2160000.0 ;
      RECT  306150.0 2149200.0 307050.0 2166000.0 ;
      RECT  309150.0 2149200.0 310050.0 2166000.0 ;
      RECT  316200.0 2151600.0 317400.0 2152800.0 ;
      RECT  318600.0 2151600.0 320250.0 2152800.0 ;
      RECT  316200.0 2158800.0 317400.0 2160000.0 ;
      RECT  319350.0 2158800.0 322200.0 2160000.0 ;
      RECT  316200.0 2151600.0 317400.0 2152800.0 ;
      RECT  318600.0 2151600.0 319800.0 2152800.0 ;
      RECT  316200.0 2158800.0 317400.0 2160000.0 ;
      RECT  321000.0 2158800.0 322200.0 2160000.0 ;
      RECT  316350.0 2149200.0 317250.0 2166000.0 ;
      RECT  319350.0 2149200.0 320250.0 2166000.0 ;
      RECT  326400.0 2151600.0 327600.0 2152800.0 ;
      RECT  328800.0 2151600.0 330450.0 2152800.0 ;
      RECT  326400.0 2158800.0 327600.0 2160000.0 ;
      RECT  329550.0 2158800.0 332400.0 2160000.0 ;
      RECT  326400.0 2151600.0 327600.0 2152800.0 ;
      RECT  328800.0 2151600.0 330000.0 2152800.0 ;
      RECT  326400.0 2158800.0 327600.0 2160000.0 ;
      RECT  331200.0 2158800.0 332400.0 2160000.0 ;
      RECT  326550.0 2149200.0 327450.0 2166000.0 ;
      RECT  329550.0 2149200.0 330450.0 2166000.0 ;
      RECT  336600.0 2151600.0 337800.0 2152800.0 ;
      RECT  339000.0 2151600.0 340650.0 2152800.0 ;
      RECT  336600.0 2158800.0 337800.0 2160000.0 ;
      RECT  339750.0 2158800.0 342600.0 2160000.0 ;
      RECT  336600.0 2151600.0 337800.0 2152800.0 ;
      RECT  339000.0 2151600.0 340200.0 2152800.0 ;
      RECT  336600.0 2158800.0 337800.0 2160000.0 ;
      RECT  341400.0 2158800.0 342600.0 2160000.0 ;
      RECT  336750.0 2149200.0 337650.0 2166000.0 ;
      RECT  339750.0 2149200.0 340650.0 2166000.0 ;
      RECT  346800.0 2151600.0 348000.0 2152800.0 ;
      RECT  349200.0 2151600.0 350850.0 2152800.0 ;
      RECT  346800.0 2158800.0 348000.0 2160000.0 ;
      RECT  349950.0 2158800.0 352800.0 2160000.0 ;
      RECT  346800.0 2151600.0 348000.0 2152800.0 ;
      RECT  349200.0 2151600.0 350400.0 2152800.0 ;
      RECT  346800.0 2158800.0 348000.0 2160000.0 ;
      RECT  351600.0 2158800.0 352800.0 2160000.0 ;
      RECT  346950.0 2149200.0 347850.0 2166000.0 ;
      RECT  349950.0 2149200.0 350850.0 2166000.0 ;
      RECT  357000.0 2151600.0 358200.0 2152800.0 ;
      RECT  359400.0 2151600.0 361050.0 2152800.0 ;
      RECT  357000.0 2158800.0 358200.0 2160000.0 ;
      RECT  360150.0 2158800.0 363000.0 2160000.0 ;
      RECT  357000.0 2151600.0 358200.0 2152800.0 ;
      RECT  359400.0 2151600.0 360600.0 2152800.0 ;
      RECT  357000.0 2158800.0 358200.0 2160000.0 ;
      RECT  361800.0 2158800.0 363000.0 2160000.0 ;
      RECT  357150.0 2149200.0 358050.0 2166000.0 ;
      RECT  360150.0 2149200.0 361050.0 2166000.0 ;
      RECT  367200.0 2151600.0 368400.0 2152800.0 ;
      RECT  369600.0 2151600.0 371250.0 2152800.0 ;
      RECT  367200.0 2158800.0 368400.0 2160000.0 ;
      RECT  370350.0 2158800.0 373200.0 2160000.0 ;
      RECT  367200.0 2151600.0 368400.0 2152800.0 ;
      RECT  369600.0 2151600.0 370800.0 2152800.0 ;
      RECT  367200.0 2158800.0 368400.0 2160000.0 ;
      RECT  372000.0 2158800.0 373200.0 2160000.0 ;
      RECT  367350.0 2149200.0 368250.0 2166000.0 ;
      RECT  370350.0 2149200.0 371250.0 2166000.0 ;
      RECT  377400.0 2151600.0 378600.0 2152800.0 ;
      RECT  379800.0 2151600.0 381450.0 2152800.0 ;
      RECT  377400.0 2158800.0 378600.0 2160000.0 ;
      RECT  380550.0 2158800.0 383400.0 2160000.0 ;
      RECT  377400.0 2151600.0 378600.0 2152800.0 ;
      RECT  379800.0 2151600.0 381000.0 2152800.0 ;
      RECT  377400.0 2158800.0 378600.0 2160000.0 ;
      RECT  382200.0 2158800.0 383400.0 2160000.0 ;
      RECT  377550.0 2149200.0 378450.0 2166000.0 ;
      RECT  380550.0 2149200.0 381450.0 2166000.0 ;
      RECT  387600.0 2151600.0 388800.0 2152800.0 ;
      RECT  390000.0 2151600.0 391650.0 2152800.0 ;
      RECT  387600.0 2158800.0 388800.0 2160000.0 ;
      RECT  390750.0 2158800.0 393600.0 2160000.0 ;
      RECT  387600.0 2151600.0 388800.0 2152800.0 ;
      RECT  390000.0 2151600.0 391200.0 2152800.0 ;
      RECT  387600.0 2158800.0 388800.0 2160000.0 ;
      RECT  392400.0 2158800.0 393600.0 2160000.0 ;
      RECT  387750.0 2149200.0 388650.0 2166000.0 ;
      RECT  390750.0 2149200.0 391650.0 2166000.0 ;
      RECT  397800.0 2151600.0 399000.0 2152800.0 ;
      RECT  400200.0 2151600.0 401850.0 2152800.0 ;
      RECT  397800.0 2158800.0 399000.0 2160000.0 ;
      RECT  400950.0 2158800.0 403800.0 2160000.0 ;
      RECT  397800.0 2151600.0 399000.0 2152800.0 ;
      RECT  400200.0 2151600.0 401400.0 2152800.0 ;
      RECT  397800.0 2158800.0 399000.0 2160000.0 ;
      RECT  402600.0 2158800.0 403800.0 2160000.0 ;
      RECT  397950.0 2149200.0 398850.0 2166000.0 ;
      RECT  400950.0 2149200.0 401850.0 2166000.0 ;
      RECT  408000.0 2151600.0 409200.0 2152800.0 ;
      RECT  410400.0 2151600.0 412050.0 2152800.0 ;
      RECT  408000.0 2158800.0 409200.0 2160000.0 ;
      RECT  411150.0 2158800.0 414000.0 2160000.0 ;
      RECT  408000.0 2151600.0 409200.0 2152800.0 ;
      RECT  410400.0 2151600.0 411600.0 2152800.0 ;
      RECT  408000.0 2158800.0 409200.0 2160000.0 ;
      RECT  412800.0 2158800.0 414000.0 2160000.0 ;
      RECT  408150.0 2149200.0 409050.0 2166000.0 ;
      RECT  411150.0 2149200.0 412050.0 2166000.0 ;
      RECT  418200.0 2151600.0 419400.0 2152800.0 ;
      RECT  420600.0 2151600.0 422250.0 2152800.0 ;
      RECT  418200.0 2158800.0 419400.0 2160000.0 ;
      RECT  421350.0 2158800.0 424200.0 2160000.0 ;
      RECT  418200.0 2151600.0 419400.0 2152800.0 ;
      RECT  420600.0 2151600.0 421800.0 2152800.0 ;
      RECT  418200.0 2158800.0 419400.0 2160000.0 ;
      RECT  423000.0 2158800.0 424200.0 2160000.0 ;
      RECT  418350.0 2149200.0 419250.0 2166000.0 ;
      RECT  421350.0 2149200.0 422250.0 2166000.0 ;
      RECT  428400.0 2151600.0 429600.0 2152800.0 ;
      RECT  430800.0 2151600.0 432450.0 2152800.0 ;
      RECT  428400.0 2158800.0 429600.0 2160000.0 ;
      RECT  431550.0 2158800.0 434400.0 2160000.0 ;
      RECT  428400.0 2151600.0 429600.0 2152800.0 ;
      RECT  430800.0 2151600.0 432000.0 2152800.0 ;
      RECT  428400.0 2158800.0 429600.0 2160000.0 ;
      RECT  433200.0 2158800.0 434400.0 2160000.0 ;
      RECT  428550.0 2149200.0 429450.0 2166000.0 ;
      RECT  431550.0 2149200.0 432450.0 2166000.0 ;
      RECT  438600.0 2151600.0 439800.0 2152800.0 ;
      RECT  441000.0 2151600.0 442650.0 2152800.0 ;
      RECT  438600.0 2158800.0 439800.0 2160000.0 ;
      RECT  441750.0 2158800.0 444600.0 2160000.0 ;
      RECT  438600.0 2151600.0 439800.0 2152800.0 ;
      RECT  441000.0 2151600.0 442200.0 2152800.0 ;
      RECT  438600.0 2158800.0 439800.0 2160000.0 ;
      RECT  443400.0 2158800.0 444600.0 2160000.0 ;
      RECT  438750.0 2149200.0 439650.0 2166000.0 ;
      RECT  441750.0 2149200.0 442650.0 2166000.0 ;
      RECT  448800.0 2151600.0 450000.0 2152800.0 ;
      RECT  451200.0 2151600.0 452850.0 2152800.0 ;
      RECT  448800.0 2158800.0 450000.0 2160000.0 ;
      RECT  451950.0 2158800.0 454800.0 2160000.0 ;
      RECT  448800.0 2151600.0 450000.0 2152800.0 ;
      RECT  451200.0 2151600.0 452400.0 2152800.0 ;
      RECT  448800.0 2158800.0 450000.0 2160000.0 ;
      RECT  453600.0 2158800.0 454800.0 2160000.0 ;
      RECT  448950.0 2149200.0 449850.0 2166000.0 ;
      RECT  451950.0 2149200.0 452850.0 2166000.0 ;
      RECT  459000.0 2151600.0 460200.0 2152800.0 ;
      RECT  461400.0 2151600.0 463050.0 2152800.0 ;
      RECT  459000.0 2158800.0 460200.0 2160000.0 ;
      RECT  462150.0 2158800.0 465000.0 2160000.0 ;
      RECT  459000.0 2151600.0 460200.0 2152800.0 ;
      RECT  461400.0 2151600.0 462600.0 2152800.0 ;
      RECT  459000.0 2158800.0 460200.0 2160000.0 ;
      RECT  463800.0 2158800.0 465000.0 2160000.0 ;
      RECT  459150.0 2149200.0 460050.0 2166000.0 ;
      RECT  462150.0 2149200.0 463050.0 2166000.0 ;
      RECT  469200.0 2151600.0 470400.0 2152800.0 ;
      RECT  471600.0 2151600.0 473250.0 2152800.0 ;
      RECT  469200.0 2158800.0 470400.0 2160000.0 ;
      RECT  472350.0 2158800.0 475200.0 2160000.0 ;
      RECT  469200.0 2151600.0 470400.0 2152800.0 ;
      RECT  471600.0 2151600.0 472800.0 2152800.0 ;
      RECT  469200.0 2158800.0 470400.0 2160000.0 ;
      RECT  474000.0 2158800.0 475200.0 2160000.0 ;
      RECT  469350.0 2149200.0 470250.0 2166000.0 ;
      RECT  472350.0 2149200.0 473250.0 2166000.0 ;
      RECT  479400.0 2151600.0 480600.0 2152800.0 ;
      RECT  481800.0 2151600.0 483450.0 2152800.0 ;
      RECT  479400.0 2158800.0 480600.0 2160000.0 ;
      RECT  482550.0 2158800.0 485400.0 2160000.0 ;
      RECT  479400.0 2151600.0 480600.0 2152800.0 ;
      RECT  481800.0 2151600.0 483000.0 2152800.0 ;
      RECT  479400.0 2158800.0 480600.0 2160000.0 ;
      RECT  484200.0 2158800.0 485400.0 2160000.0 ;
      RECT  479550.0 2149200.0 480450.0 2166000.0 ;
      RECT  482550.0 2149200.0 483450.0 2166000.0 ;
      RECT  489600.0 2151600.0 490800.0 2152800.0 ;
      RECT  492000.0 2151600.0 493650.0 2152800.0 ;
      RECT  489600.0 2158800.0 490800.0 2160000.0 ;
      RECT  492750.0 2158800.0 495600.0 2160000.0 ;
      RECT  489600.0 2151600.0 490800.0 2152800.0 ;
      RECT  492000.0 2151600.0 493200.0 2152800.0 ;
      RECT  489600.0 2158800.0 490800.0 2160000.0 ;
      RECT  494400.0 2158800.0 495600.0 2160000.0 ;
      RECT  489750.0 2149200.0 490650.0 2166000.0 ;
      RECT  492750.0 2149200.0 493650.0 2166000.0 ;
      RECT  499800.0 2151600.0 501000.0 2152800.0 ;
      RECT  502200.0 2151600.0 503850.0 2152800.0 ;
      RECT  499800.0 2158800.0 501000.0 2160000.0 ;
      RECT  502950.0 2158800.0 505800.0 2160000.0 ;
      RECT  499800.0 2151600.0 501000.0 2152800.0 ;
      RECT  502200.0 2151600.0 503400.0 2152800.0 ;
      RECT  499800.0 2158800.0 501000.0 2160000.0 ;
      RECT  504600.0 2158800.0 505800.0 2160000.0 ;
      RECT  499950.0 2149200.0 500850.0 2166000.0 ;
      RECT  502950.0 2149200.0 503850.0 2166000.0 ;
      RECT  510000.0 2151600.0 511200.0 2152800.0 ;
      RECT  512400.0 2151600.0 514050.0 2152800.0 ;
      RECT  510000.0 2158800.0 511200.0 2160000.0 ;
      RECT  513150.0 2158800.0 516000.0 2160000.0 ;
      RECT  510000.0 2151600.0 511200.0 2152800.0 ;
      RECT  512400.0 2151600.0 513600.0 2152800.0 ;
      RECT  510000.0 2158800.0 511200.0 2160000.0 ;
      RECT  514800.0 2158800.0 516000.0 2160000.0 ;
      RECT  510150.0 2149200.0 511050.0 2166000.0 ;
      RECT  513150.0 2149200.0 514050.0 2166000.0 ;
      RECT  520200.0 2151600.0 521400.0 2152800.0 ;
      RECT  522600.0 2151600.0 524250.0 2152800.0 ;
      RECT  520200.0 2158800.0 521400.0 2160000.0 ;
      RECT  523350.0 2158800.0 526200.0 2160000.0 ;
      RECT  520200.0 2151600.0 521400.0 2152800.0 ;
      RECT  522600.0 2151600.0 523800.0 2152800.0 ;
      RECT  520200.0 2158800.0 521400.0 2160000.0 ;
      RECT  525000.0 2158800.0 526200.0 2160000.0 ;
      RECT  520350.0 2149200.0 521250.0 2166000.0 ;
      RECT  523350.0 2149200.0 524250.0 2166000.0 ;
      RECT  530400.0 2151600.0 531600.0 2152800.0 ;
      RECT  532800.0 2151600.0 534450.0 2152800.0 ;
      RECT  530400.0 2158800.0 531600.0 2160000.0 ;
      RECT  533550.0 2158800.0 536400.0 2160000.0 ;
      RECT  530400.0 2151600.0 531600.0 2152800.0 ;
      RECT  532800.0 2151600.0 534000.0 2152800.0 ;
      RECT  530400.0 2158800.0 531600.0 2160000.0 ;
      RECT  535200.0 2158800.0 536400.0 2160000.0 ;
      RECT  530550.0 2149200.0 531450.0 2166000.0 ;
      RECT  533550.0 2149200.0 534450.0 2166000.0 ;
      RECT  540600.0 2151600.0 541800.0 2152800.0 ;
      RECT  543000.0 2151600.0 544650.0 2152800.0 ;
      RECT  540600.0 2158800.0 541800.0 2160000.0 ;
      RECT  543750.0 2158800.0 546600.0 2160000.0 ;
      RECT  540600.0 2151600.0 541800.0 2152800.0 ;
      RECT  543000.0 2151600.0 544200.0 2152800.0 ;
      RECT  540600.0 2158800.0 541800.0 2160000.0 ;
      RECT  545400.0 2158800.0 546600.0 2160000.0 ;
      RECT  540750.0 2149200.0 541650.0 2166000.0 ;
      RECT  543750.0 2149200.0 544650.0 2166000.0 ;
      RECT  550800.0 2151600.0 552000.0 2152800.0 ;
      RECT  553200.0 2151600.0 554850.0 2152800.0 ;
      RECT  550800.0 2158800.0 552000.0 2160000.0 ;
      RECT  553950.0 2158800.0 556800.0 2160000.0 ;
      RECT  550800.0 2151600.0 552000.0 2152800.0 ;
      RECT  553200.0 2151600.0 554400.0 2152800.0 ;
      RECT  550800.0 2158800.0 552000.0 2160000.0 ;
      RECT  555600.0 2158800.0 556800.0 2160000.0 ;
      RECT  550950.0 2149200.0 551850.0 2166000.0 ;
      RECT  553950.0 2149200.0 554850.0 2166000.0 ;
      RECT  561000.0 2151600.0 562200.0 2152800.0 ;
      RECT  563400.0 2151600.0 565050.0 2152800.0 ;
      RECT  561000.0 2158800.0 562200.0 2160000.0 ;
      RECT  564150.0 2158800.0 567000.0 2160000.0 ;
      RECT  561000.0 2151600.0 562200.0 2152800.0 ;
      RECT  563400.0 2151600.0 564600.0 2152800.0 ;
      RECT  561000.0 2158800.0 562200.0 2160000.0 ;
      RECT  565800.0 2158800.0 567000.0 2160000.0 ;
      RECT  561150.0 2149200.0 562050.0 2166000.0 ;
      RECT  564150.0 2149200.0 565050.0 2166000.0 ;
      RECT  571200.0 2151600.0 572400.0 2152800.0 ;
      RECT  573600.0 2151600.0 575250.0 2152800.0 ;
      RECT  571200.0 2158800.0 572400.0 2160000.0 ;
      RECT  574350.0 2158800.0 577200.0 2160000.0 ;
      RECT  571200.0 2151600.0 572400.0 2152800.0 ;
      RECT  573600.0 2151600.0 574800.0 2152800.0 ;
      RECT  571200.0 2158800.0 572400.0 2160000.0 ;
      RECT  576000.0 2158800.0 577200.0 2160000.0 ;
      RECT  571350.0 2149200.0 572250.0 2166000.0 ;
      RECT  574350.0 2149200.0 575250.0 2166000.0 ;
      RECT  581400.0 2151600.0 582600.0 2152800.0 ;
      RECT  583800.0 2151600.0 585450.0 2152800.0 ;
      RECT  581400.0 2158800.0 582600.0 2160000.0 ;
      RECT  584550.0 2158800.0 587400.0 2160000.0 ;
      RECT  581400.0 2151600.0 582600.0 2152800.0 ;
      RECT  583800.0 2151600.0 585000.0 2152800.0 ;
      RECT  581400.0 2158800.0 582600.0 2160000.0 ;
      RECT  586200.0 2158800.0 587400.0 2160000.0 ;
      RECT  581550.0 2149200.0 582450.0 2166000.0 ;
      RECT  584550.0 2149200.0 585450.0 2166000.0 ;
      RECT  591600.0 2151600.0 592800.0 2152800.0 ;
      RECT  594000.0 2151600.0 595650.0 2152800.0 ;
      RECT  591600.0 2158800.0 592800.0 2160000.0 ;
      RECT  594750.0 2158800.0 597600.0 2160000.0 ;
      RECT  591600.0 2151600.0 592800.0 2152800.0 ;
      RECT  594000.0 2151600.0 595200.0 2152800.0 ;
      RECT  591600.0 2158800.0 592800.0 2160000.0 ;
      RECT  596400.0 2158800.0 597600.0 2160000.0 ;
      RECT  591750.0 2149200.0 592650.0 2166000.0 ;
      RECT  594750.0 2149200.0 595650.0 2166000.0 ;
      RECT  601800.0 2151600.0 603000.0 2152800.0 ;
      RECT  604200.0 2151600.0 605850.0 2152800.0 ;
      RECT  601800.0 2158800.0 603000.0 2160000.0 ;
      RECT  604950.0 2158800.0 607800.0 2160000.0 ;
      RECT  601800.0 2151600.0 603000.0 2152800.0 ;
      RECT  604200.0 2151600.0 605400.0 2152800.0 ;
      RECT  601800.0 2158800.0 603000.0 2160000.0 ;
      RECT  606600.0 2158800.0 607800.0 2160000.0 ;
      RECT  601950.0 2149200.0 602850.0 2166000.0 ;
      RECT  604950.0 2149200.0 605850.0 2166000.0 ;
      RECT  612000.0 2151600.0 613200.0 2152800.0 ;
      RECT  614400.0 2151600.0 616050.0 2152800.0 ;
      RECT  612000.0 2158800.0 613200.0 2160000.0 ;
      RECT  615150.0 2158800.0 618000.0 2160000.0 ;
      RECT  612000.0 2151600.0 613200.0 2152800.0 ;
      RECT  614400.0 2151600.0 615600.0 2152800.0 ;
      RECT  612000.0 2158800.0 613200.0 2160000.0 ;
      RECT  616800.0 2158800.0 618000.0 2160000.0 ;
      RECT  612150.0 2149200.0 613050.0 2166000.0 ;
      RECT  615150.0 2149200.0 616050.0 2166000.0 ;
      RECT  622200.0 2151600.0 623400.0 2152800.0 ;
      RECT  624600.0 2151600.0 626250.0 2152800.0 ;
      RECT  622200.0 2158800.0 623400.0 2160000.0 ;
      RECT  625350.0 2158800.0 628200.0 2160000.0 ;
      RECT  622200.0 2151600.0 623400.0 2152800.0 ;
      RECT  624600.0 2151600.0 625800.0 2152800.0 ;
      RECT  622200.0 2158800.0 623400.0 2160000.0 ;
      RECT  627000.0 2158800.0 628200.0 2160000.0 ;
      RECT  622350.0 2149200.0 623250.0 2166000.0 ;
      RECT  625350.0 2149200.0 626250.0 2166000.0 ;
      RECT  632400.0 2151600.0 633600.0 2152800.0 ;
      RECT  634800.0 2151600.0 636450.0 2152800.0 ;
      RECT  632400.0 2158800.0 633600.0 2160000.0 ;
      RECT  635550.0 2158800.0 638400.0 2160000.0 ;
      RECT  632400.0 2151600.0 633600.0 2152800.0 ;
      RECT  634800.0 2151600.0 636000.0 2152800.0 ;
      RECT  632400.0 2158800.0 633600.0 2160000.0 ;
      RECT  637200.0 2158800.0 638400.0 2160000.0 ;
      RECT  632550.0 2149200.0 633450.0 2166000.0 ;
      RECT  635550.0 2149200.0 636450.0 2166000.0 ;
      RECT  642600.0 2151600.0 643800.0 2152800.0 ;
      RECT  645000.0 2151600.0 646650.0 2152800.0 ;
      RECT  642600.0 2158800.0 643800.0 2160000.0 ;
      RECT  645750.0 2158800.0 648600.0 2160000.0 ;
      RECT  642600.0 2151600.0 643800.0 2152800.0 ;
      RECT  645000.0 2151600.0 646200.0 2152800.0 ;
      RECT  642600.0 2158800.0 643800.0 2160000.0 ;
      RECT  647400.0 2158800.0 648600.0 2160000.0 ;
      RECT  642750.0 2149200.0 643650.0 2166000.0 ;
      RECT  645750.0 2149200.0 646650.0 2166000.0 ;
      RECT  652800.0 2151600.0 654000.0 2152800.0 ;
      RECT  655200.0 2151600.0 656850.0 2152800.0 ;
      RECT  652800.0 2158800.0 654000.0 2160000.0 ;
      RECT  655950.0 2158800.0 658800.0 2160000.0 ;
      RECT  652800.0 2151600.0 654000.0 2152800.0 ;
      RECT  655200.0 2151600.0 656400.0 2152800.0 ;
      RECT  652800.0 2158800.0 654000.0 2160000.0 ;
      RECT  657600.0 2158800.0 658800.0 2160000.0 ;
      RECT  652950.0 2149200.0 653850.0 2166000.0 ;
      RECT  655950.0 2149200.0 656850.0 2166000.0 ;
      RECT  663000.0 2151600.0 664200.0 2152800.0 ;
      RECT  665400.0 2151600.0 667050.0 2152800.0 ;
      RECT  663000.0 2158800.0 664200.0 2160000.0 ;
      RECT  666150.0 2158800.0 669000.0 2160000.0 ;
      RECT  663000.0 2151600.0 664200.0 2152800.0 ;
      RECT  665400.0 2151600.0 666600.0 2152800.0 ;
      RECT  663000.0 2158800.0 664200.0 2160000.0 ;
      RECT  667800.0 2158800.0 669000.0 2160000.0 ;
      RECT  663150.0 2149200.0 664050.0 2166000.0 ;
      RECT  666150.0 2149200.0 667050.0 2166000.0 ;
      RECT  673200.0 2151600.0 674400.0 2152800.0 ;
      RECT  675600.0 2151600.0 677250.0 2152800.0 ;
      RECT  673200.0 2158800.0 674400.0 2160000.0 ;
      RECT  676350.0 2158800.0 679200.0 2160000.0 ;
      RECT  673200.0 2151600.0 674400.0 2152800.0 ;
      RECT  675600.0 2151600.0 676800.0 2152800.0 ;
      RECT  673200.0 2158800.0 674400.0 2160000.0 ;
      RECT  678000.0 2158800.0 679200.0 2160000.0 ;
      RECT  673350.0 2149200.0 674250.0 2166000.0 ;
      RECT  676350.0 2149200.0 677250.0 2166000.0 ;
      RECT  683400.0 2151600.0 684600.0 2152800.0 ;
      RECT  685800.0 2151600.0 687450.0 2152800.0 ;
      RECT  683400.0 2158800.0 684600.0 2160000.0 ;
      RECT  686550.0 2158800.0 689400.0 2160000.0 ;
      RECT  683400.0 2151600.0 684600.0 2152800.0 ;
      RECT  685800.0 2151600.0 687000.0 2152800.0 ;
      RECT  683400.0 2158800.0 684600.0 2160000.0 ;
      RECT  688200.0 2158800.0 689400.0 2160000.0 ;
      RECT  683550.0 2149200.0 684450.0 2166000.0 ;
      RECT  686550.0 2149200.0 687450.0 2166000.0 ;
      RECT  693600.0 2151600.0 694800.0 2152800.0 ;
      RECT  696000.0 2151600.0 697650.0 2152800.0 ;
      RECT  693600.0 2158800.0 694800.0 2160000.0 ;
      RECT  696750.0 2158800.0 699600.0 2160000.0 ;
      RECT  693600.0 2151600.0 694800.0 2152800.0 ;
      RECT  696000.0 2151600.0 697200.0 2152800.0 ;
      RECT  693600.0 2158800.0 694800.0 2160000.0 ;
      RECT  698400.0 2158800.0 699600.0 2160000.0 ;
      RECT  693750.0 2149200.0 694650.0 2166000.0 ;
      RECT  696750.0 2149200.0 697650.0 2166000.0 ;
      RECT  703800.0 2151600.0 705000.0 2152800.0 ;
      RECT  706200.0 2151600.0 707850.0 2152800.0 ;
      RECT  703800.0 2158800.0 705000.0 2160000.0 ;
      RECT  706950.0 2158800.0 709800.0 2160000.0 ;
      RECT  703800.0 2151600.0 705000.0 2152800.0 ;
      RECT  706200.0 2151600.0 707400.0 2152800.0 ;
      RECT  703800.0 2158800.0 705000.0 2160000.0 ;
      RECT  708600.0 2158800.0 709800.0 2160000.0 ;
      RECT  703950.0 2149200.0 704850.0 2166000.0 ;
      RECT  706950.0 2149200.0 707850.0 2166000.0 ;
      RECT  714000.0 2151600.0 715200.0 2152800.0 ;
      RECT  716400.0 2151600.0 718050.0 2152800.0 ;
      RECT  714000.0 2158800.0 715200.0 2160000.0 ;
      RECT  717150.0 2158800.0 720000.0 2160000.0 ;
      RECT  714000.0 2151600.0 715200.0 2152800.0 ;
      RECT  716400.0 2151600.0 717600.0 2152800.0 ;
      RECT  714000.0 2158800.0 715200.0 2160000.0 ;
      RECT  718800.0 2158800.0 720000.0 2160000.0 ;
      RECT  714150.0 2149200.0 715050.0 2166000.0 ;
      RECT  717150.0 2149200.0 718050.0 2166000.0 ;
      RECT  724200.0 2151600.0 725400.0 2152800.0 ;
      RECT  726600.0 2151600.0 728250.0 2152800.0 ;
      RECT  724200.0 2158800.0 725400.0 2160000.0 ;
      RECT  727350.0 2158800.0 730200.0 2160000.0 ;
      RECT  724200.0 2151600.0 725400.0 2152800.0 ;
      RECT  726600.0 2151600.0 727800.0 2152800.0 ;
      RECT  724200.0 2158800.0 725400.0 2160000.0 ;
      RECT  729000.0 2158800.0 730200.0 2160000.0 ;
      RECT  724350.0 2149200.0 725250.0 2166000.0 ;
      RECT  727350.0 2149200.0 728250.0 2166000.0 ;
      RECT  734400.0 2151600.0 735600.0 2152800.0 ;
      RECT  736800.0 2151600.0 738450.0 2152800.0 ;
      RECT  734400.0 2158800.0 735600.0 2160000.0 ;
      RECT  737550.0 2158800.0 740400.0 2160000.0 ;
      RECT  734400.0 2151600.0 735600.0 2152800.0 ;
      RECT  736800.0 2151600.0 738000.0 2152800.0 ;
      RECT  734400.0 2158800.0 735600.0 2160000.0 ;
      RECT  739200.0 2158800.0 740400.0 2160000.0 ;
      RECT  734550.0 2149200.0 735450.0 2166000.0 ;
      RECT  737550.0 2149200.0 738450.0 2166000.0 ;
      RECT  744600.0 2151600.0 745800.0 2152800.0 ;
      RECT  747000.0 2151600.0 748650.0 2152800.0 ;
      RECT  744600.0 2158800.0 745800.0 2160000.0 ;
      RECT  747750.0 2158800.0 750600.0 2160000.0 ;
      RECT  744600.0 2151600.0 745800.0 2152800.0 ;
      RECT  747000.0 2151600.0 748200.0 2152800.0 ;
      RECT  744600.0 2158800.0 745800.0 2160000.0 ;
      RECT  749400.0 2158800.0 750600.0 2160000.0 ;
      RECT  744750.0 2149200.0 745650.0 2166000.0 ;
      RECT  747750.0 2149200.0 748650.0 2166000.0 ;
      RECT  754800.0 2151600.0 756000.0 2152800.0 ;
      RECT  757200.0 2151600.0 758850.0 2152800.0 ;
      RECT  754800.0 2158800.0 756000.0 2160000.0 ;
      RECT  757950.0 2158800.0 760800.0 2160000.0 ;
      RECT  754800.0 2151600.0 756000.0 2152800.0 ;
      RECT  757200.0 2151600.0 758400.0 2152800.0 ;
      RECT  754800.0 2158800.0 756000.0 2160000.0 ;
      RECT  759600.0 2158800.0 760800.0 2160000.0 ;
      RECT  754950.0 2149200.0 755850.0 2166000.0 ;
      RECT  757950.0 2149200.0 758850.0 2166000.0 ;
      RECT  765000.0 2151600.0 766200.0 2152800.0 ;
      RECT  767400.0 2151600.0 769050.0 2152800.0 ;
      RECT  765000.0 2158800.0 766200.0 2160000.0 ;
      RECT  768150.0 2158800.0 771000.0 2160000.0 ;
      RECT  765000.0 2151600.0 766200.0 2152800.0 ;
      RECT  767400.0 2151600.0 768600.0 2152800.0 ;
      RECT  765000.0 2158800.0 766200.0 2160000.0 ;
      RECT  769800.0 2158800.0 771000.0 2160000.0 ;
      RECT  765150.0 2149200.0 766050.0 2166000.0 ;
      RECT  768150.0 2149200.0 769050.0 2166000.0 ;
      RECT  775200.0 2151600.0 776400.0 2152800.0 ;
      RECT  777600.0 2151600.0 779250.0 2152800.0 ;
      RECT  775200.0 2158800.0 776400.0 2160000.0 ;
      RECT  778350.0 2158800.0 781200.0 2160000.0 ;
      RECT  775200.0 2151600.0 776400.0 2152800.0 ;
      RECT  777600.0 2151600.0 778800.0 2152800.0 ;
      RECT  775200.0 2158800.0 776400.0 2160000.0 ;
      RECT  780000.0 2158800.0 781200.0 2160000.0 ;
      RECT  775350.0 2149200.0 776250.0 2166000.0 ;
      RECT  778350.0 2149200.0 779250.0 2166000.0 ;
      RECT  785400.0 2151600.0 786600.0 2152800.0 ;
      RECT  787800.0 2151600.0 789450.0 2152800.0 ;
      RECT  785400.0 2158800.0 786600.0 2160000.0 ;
      RECT  788550.0 2158800.0 791400.0 2160000.0 ;
      RECT  785400.0 2151600.0 786600.0 2152800.0 ;
      RECT  787800.0 2151600.0 789000.0 2152800.0 ;
      RECT  785400.0 2158800.0 786600.0 2160000.0 ;
      RECT  790200.0 2158800.0 791400.0 2160000.0 ;
      RECT  785550.0 2149200.0 786450.0 2166000.0 ;
      RECT  788550.0 2149200.0 789450.0 2166000.0 ;
      RECT  795600.0 2151600.0 796800.0 2152800.0 ;
      RECT  798000.0 2151600.0 799650.0 2152800.0 ;
      RECT  795600.0 2158800.0 796800.0 2160000.0 ;
      RECT  798750.0 2158800.0 801600.0 2160000.0 ;
      RECT  795600.0 2151600.0 796800.0 2152800.0 ;
      RECT  798000.0 2151600.0 799200.0 2152800.0 ;
      RECT  795600.0 2158800.0 796800.0 2160000.0 ;
      RECT  800400.0 2158800.0 801600.0 2160000.0 ;
      RECT  795750.0 2149200.0 796650.0 2166000.0 ;
      RECT  798750.0 2149200.0 799650.0 2166000.0 ;
      RECT  805800.0 2151600.0 807000.0 2152800.0 ;
      RECT  808200.0 2151600.0 809850.0 2152800.0 ;
      RECT  805800.0 2158800.0 807000.0 2160000.0 ;
      RECT  808950.0 2158800.0 811800.0 2160000.0 ;
      RECT  805800.0 2151600.0 807000.0 2152800.0 ;
      RECT  808200.0 2151600.0 809400.0 2152800.0 ;
      RECT  805800.0 2158800.0 807000.0 2160000.0 ;
      RECT  810600.0 2158800.0 811800.0 2160000.0 ;
      RECT  805950.0 2149200.0 806850.0 2166000.0 ;
      RECT  808950.0 2149200.0 809850.0 2166000.0 ;
      RECT  816000.0 2151600.0 817200.0 2152800.0 ;
      RECT  818400.0 2151600.0 820050.0 2152800.0 ;
      RECT  816000.0 2158800.0 817200.0 2160000.0 ;
      RECT  819150.0 2158800.0 822000.0 2160000.0 ;
      RECT  816000.0 2151600.0 817200.0 2152800.0 ;
      RECT  818400.0 2151600.0 819600.0 2152800.0 ;
      RECT  816000.0 2158800.0 817200.0 2160000.0 ;
      RECT  820800.0 2158800.0 822000.0 2160000.0 ;
      RECT  816150.0 2149200.0 817050.0 2166000.0 ;
      RECT  819150.0 2149200.0 820050.0 2166000.0 ;
      RECT  826200.0 2151600.0 827400.0 2152800.0 ;
      RECT  828600.0 2151600.0 830250.0 2152800.0 ;
      RECT  826200.0 2158800.0 827400.0 2160000.0 ;
      RECT  829350.0 2158800.0 832200.0 2160000.0 ;
      RECT  826200.0 2151600.0 827400.0 2152800.0 ;
      RECT  828600.0 2151600.0 829800.0 2152800.0 ;
      RECT  826200.0 2158800.0 827400.0 2160000.0 ;
      RECT  831000.0 2158800.0 832200.0 2160000.0 ;
      RECT  826350.0 2149200.0 827250.0 2166000.0 ;
      RECT  829350.0 2149200.0 830250.0 2166000.0 ;
      RECT  836400.0 2151600.0 837600.0 2152800.0 ;
      RECT  838800.0 2151600.0 840450.0 2152800.0 ;
      RECT  836400.0 2158800.0 837600.0 2160000.0 ;
      RECT  839550.0 2158800.0 842400.0 2160000.0 ;
      RECT  836400.0 2151600.0 837600.0 2152800.0 ;
      RECT  838800.0 2151600.0 840000.0 2152800.0 ;
      RECT  836400.0 2158800.0 837600.0 2160000.0 ;
      RECT  841200.0 2158800.0 842400.0 2160000.0 ;
      RECT  836550.0 2149200.0 837450.0 2166000.0 ;
      RECT  839550.0 2149200.0 840450.0 2166000.0 ;
      RECT  846600.0 2151600.0 847800.0 2152800.0 ;
      RECT  849000.0 2151600.0 850650.0 2152800.0 ;
      RECT  846600.0 2158800.0 847800.0 2160000.0 ;
      RECT  849750.0 2158800.0 852600.0 2160000.0 ;
      RECT  846600.0 2151600.0 847800.0 2152800.0 ;
      RECT  849000.0 2151600.0 850200.0 2152800.0 ;
      RECT  846600.0 2158800.0 847800.0 2160000.0 ;
      RECT  851400.0 2158800.0 852600.0 2160000.0 ;
      RECT  846750.0 2149200.0 847650.0 2166000.0 ;
      RECT  849750.0 2149200.0 850650.0 2166000.0 ;
      RECT  856800.0 2151600.0 858000.0 2152800.0 ;
      RECT  859200.0 2151600.0 860850.0 2152800.0 ;
      RECT  856800.0 2158800.0 858000.0 2160000.0 ;
      RECT  859950.0 2158800.0 862800.0 2160000.0 ;
      RECT  856800.0 2151600.0 858000.0 2152800.0 ;
      RECT  859200.0 2151600.0 860400.0 2152800.0 ;
      RECT  856800.0 2158800.0 858000.0 2160000.0 ;
      RECT  861600.0 2158800.0 862800.0 2160000.0 ;
      RECT  856950.0 2149200.0 857850.0 2166000.0 ;
      RECT  859950.0 2149200.0 860850.0 2166000.0 ;
      RECT  867000.0 2151600.0 868200.0 2152800.0 ;
      RECT  869400.0 2151600.0 871050.0 2152800.0 ;
      RECT  867000.0 2158800.0 868200.0 2160000.0 ;
      RECT  870150.0 2158800.0 873000.0 2160000.0 ;
      RECT  867000.0 2151600.0 868200.0 2152800.0 ;
      RECT  869400.0 2151600.0 870600.0 2152800.0 ;
      RECT  867000.0 2158800.0 868200.0 2160000.0 ;
      RECT  871800.0 2158800.0 873000.0 2160000.0 ;
      RECT  867150.0 2149200.0 868050.0 2166000.0 ;
      RECT  870150.0 2149200.0 871050.0 2166000.0 ;
      RECT  877200.0 2151600.0 878400.0 2152800.0 ;
      RECT  879600.0 2151600.0 881250.0 2152800.0 ;
      RECT  877200.0 2158800.0 878400.0 2160000.0 ;
      RECT  880350.0 2158800.0 883200.0 2160000.0 ;
      RECT  877200.0 2151600.0 878400.0 2152800.0 ;
      RECT  879600.0 2151600.0 880800.0 2152800.0 ;
      RECT  877200.0 2158800.0 878400.0 2160000.0 ;
      RECT  882000.0 2158800.0 883200.0 2160000.0 ;
      RECT  877350.0 2149200.0 878250.0 2166000.0 ;
      RECT  880350.0 2149200.0 881250.0 2166000.0 ;
      RECT  887400.0 2151600.0 888600.0 2152800.0 ;
      RECT  889800.0 2151600.0 891450.0 2152800.0 ;
      RECT  887400.0 2158800.0 888600.0 2160000.0 ;
      RECT  890550.0 2158800.0 893400.0 2160000.0 ;
      RECT  887400.0 2151600.0 888600.0 2152800.0 ;
      RECT  889800.0 2151600.0 891000.0 2152800.0 ;
      RECT  887400.0 2158800.0 888600.0 2160000.0 ;
      RECT  892200.0 2158800.0 893400.0 2160000.0 ;
      RECT  887550.0 2149200.0 888450.0 2166000.0 ;
      RECT  890550.0 2149200.0 891450.0 2166000.0 ;
      RECT  897600.0 2151600.0 898800.0 2152800.0 ;
      RECT  900000.0 2151600.0 901650.0 2152800.0 ;
      RECT  897600.0 2158800.0 898800.0 2160000.0 ;
      RECT  900750.0 2158800.0 903600.0 2160000.0 ;
      RECT  897600.0 2151600.0 898800.0 2152800.0 ;
      RECT  900000.0 2151600.0 901200.0 2152800.0 ;
      RECT  897600.0 2158800.0 898800.0 2160000.0 ;
      RECT  902400.0 2158800.0 903600.0 2160000.0 ;
      RECT  897750.0 2149200.0 898650.0 2166000.0 ;
      RECT  900750.0 2149200.0 901650.0 2166000.0 ;
      RECT  907800.0 2151600.0 909000.0 2152800.0 ;
      RECT  910200.0 2151600.0 911850.0 2152800.0 ;
      RECT  907800.0 2158800.0 909000.0 2160000.0 ;
      RECT  910950.0 2158800.0 913800.0 2160000.0 ;
      RECT  907800.0 2151600.0 909000.0 2152800.0 ;
      RECT  910200.0 2151600.0 911400.0 2152800.0 ;
      RECT  907800.0 2158800.0 909000.0 2160000.0 ;
      RECT  912600.0 2158800.0 913800.0 2160000.0 ;
      RECT  907950.0 2149200.0 908850.0 2166000.0 ;
      RECT  910950.0 2149200.0 911850.0 2166000.0 ;
      RECT  918000.0 2151600.0 919200.0 2152800.0 ;
      RECT  920400.0 2151600.0 922050.0 2152800.0 ;
      RECT  918000.0 2158800.0 919200.0 2160000.0 ;
      RECT  921150.0 2158800.0 924000.0 2160000.0 ;
      RECT  918000.0 2151600.0 919200.0 2152800.0 ;
      RECT  920400.0 2151600.0 921600.0 2152800.0 ;
      RECT  918000.0 2158800.0 919200.0 2160000.0 ;
      RECT  922800.0 2158800.0 924000.0 2160000.0 ;
      RECT  918150.0 2149200.0 919050.0 2166000.0 ;
      RECT  921150.0 2149200.0 922050.0 2166000.0 ;
      RECT  928200.0 2151600.0 929400.0 2152800.0 ;
      RECT  930600.0 2151600.0 932250.0 2152800.0 ;
      RECT  928200.0 2158800.0 929400.0 2160000.0 ;
      RECT  931350.0 2158800.0 934200.0 2160000.0 ;
      RECT  928200.0 2151600.0 929400.0 2152800.0 ;
      RECT  930600.0 2151600.0 931800.0 2152800.0 ;
      RECT  928200.0 2158800.0 929400.0 2160000.0 ;
      RECT  933000.0 2158800.0 934200.0 2160000.0 ;
      RECT  928350.0 2149200.0 929250.0 2166000.0 ;
      RECT  931350.0 2149200.0 932250.0 2166000.0 ;
      RECT  938400.0 2151600.0 939600.0 2152800.0 ;
      RECT  940800.0 2151600.0 942450.0 2152800.0 ;
      RECT  938400.0 2158800.0 939600.0 2160000.0 ;
      RECT  941550.0 2158800.0 944400.0 2160000.0 ;
      RECT  938400.0 2151600.0 939600.0 2152800.0 ;
      RECT  940800.0 2151600.0 942000.0 2152800.0 ;
      RECT  938400.0 2158800.0 939600.0 2160000.0 ;
      RECT  943200.0 2158800.0 944400.0 2160000.0 ;
      RECT  938550.0 2149200.0 939450.0 2166000.0 ;
      RECT  941550.0 2149200.0 942450.0 2166000.0 ;
      RECT  948600.0 2151600.0 949800.0 2152800.0 ;
      RECT  951000.0 2151600.0 952650.0 2152800.0 ;
      RECT  948600.0 2158800.0 949800.0 2160000.0 ;
      RECT  951750.0 2158800.0 954600.0 2160000.0 ;
      RECT  948600.0 2151600.0 949800.0 2152800.0 ;
      RECT  951000.0 2151600.0 952200.0 2152800.0 ;
      RECT  948600.0 2158800.0 949800.0 2160000.0 ;
      RECT  953400.0 2158800.0 954600.0 2160000.0 ;
      RECT  948750.0 2149200.0 949650.0 2166000.0 ;
      RECT  951750.0 2149200.0 952650.0 2166000.0 ;
      RECT  958800.0 2151600.0 960000.0 2152800.0 ;
      RECT  961200.0 2151600.0 962850.0 2152800.0 ;
      RECT  958800.0 2158800.0 960000.0 2160000.0 ;
      RECT  961950.0 2158800.0 964800.0 2160000.0 ;
      RECT  958800.0 2151600.0 960000.0 2152800.0 ;
      RECT  961200.0 2151600.0 962400.0 2152800.0 ;
      RECT  958800.0 2158800.0 960000.0 2160000.0 ;
      RECT  963600.0 2158800.0 964800.0 2160000.0 ;
      RECT  958950.0 2149200.0 959850.0 2166000.0 ;
      RECT  961950.0 2149200.0 962850.0 2166000.0 ;
      RECT  969000.0 2151600.0 970200.0 2152800.0 ;
      RECT  971400.0 2151600.0 973050.0 2152800.0 ;
      RECT  969000.0 2158800.0 970200.0 2160000.0 ;
      RECT  972150.0 2158800.0 975000.0 2160000.0 ;
      RECT  969000.0 2151600.0 970200.0 2152800.0 ;
      RECT  971400.0 2151600.0 972600.0 2152800.0 ;
      RECT  969000.0 2158800.0 970200.0 2160000.0 ;
      RECT  973800.0 2158800.0 975000.0 2160000.0 ;
      RECT  969150.0 2149200.0 970050.0 2166000.0 ;
      RECT  972150.0 2149200.0 973050.0 2166000.0 ;
      RECT  979200.0 2151600.0 980400.0 2152800.0 ;
      RECT  981600.0 2151600.0 983250.0 2152800.0 ;
      RECT  979200.0 2158800.0 980400.0 2160000.0 ;
      RECT  982350.0 2158800.0 985200.0 2160000.0 ;
      RECT  979200.0 2151600.0 980400.0 2152800.0 ;
      RECT  981600.0 2151600.0 982800.0 2152800.0 ;
      RECT  979200.0 2158800.0 980400.0 2160000.0 ;
      RECT  984000.0 2158800.0 985200.0 2160000.0 ;
      RECT  979350.0 2149200.0 980250.0 2166000.0 ;
      RECT  982350.0 2149200.0 983250.0 2166000.0 ;
      RECT  989400.0 2151600.0 990600.0 2152800.0 ;
      RECT  991800.0 2151600.0 993450.0 2152800.0 ;
      RECT  989400.0 2158800.0 990600.0 2160000.0 ;
      RECT  992550.0 2158800.0 995400.0 2160000.0 ;
      RECT  989400.0 2151600.0 990600.0 2152800.0 ;
      RECT  991800.0 2151600.0 993000.0 2152800.0 ;
      RECT  989400.0 2158800.0 990600.0 2160000.0 ;
      RECT  994200.0 2158800.0 995400.0 2160000.0 ;
      RECT  989550.0 2149200.0 990450.0 2166000.0 ;
      RECT  992550.0 2149200.0 993450.0 2166000.0 ;
      RECT  999600.0 2151600.0 1000800.0 2152800.0 ;
      RECT  1002000.0 2151600.0 1003650.0 2152800.0 ;
      RECT  999600.0 2158800.0 1000800.0 2160000.0 ;
      RECT  1002750.0 2158800.0 1005600.0 2160000.0 ;
      RECT  999600.0 2151600.0 1000800.0 2152800.0 ;
      RECT  1002000.0 2151600.0 1003200.0 2152800.0 ;
      RECT  999600.0 2158800.0 1000800.0 2160000.0 ;
      RECT  1004400.0 2158800.0 1005600.0 2160000.0 ;
      RECT  999750.0 2149200.0 1000650.0 2166000.0 ;
      RECT  1002750.0 2149200.0 1003650.0 2166000.0 ;
      RECT  1009800.0 2151600.0 1011000.0 2152800.0 ;
      RECT  1012200.0 2151600.0 1013850.0 2152800.0 ;
      RECT  1009800.0 2158800.0 1011000.0 2160000.0 ;
      RECT  1012950.0 2158800.0 1015800.0 2160000.0 ;
      RECT  1009800.0 2151600.0 1011000.0 2152800.0 ;
      RECT  1012200.0 2151600.0 1013400.0 2152800.0 ;
      RECT  1009800.0 2158800.0 1011000.0 2160000.0 ;
      RECT  1014600.0 2158800.0 1015800.0 2160000.0 ;
      RECT  1009950.0 2149200.0 1010850.0 2166000.0 ;
      RECT  1012950.0 2149200.0 1013850.0 2166000.0 ;
      RECT  1020000.0 2151600.0 1021200.0 2152800.0 ;
      RECT  1022400.0 2151600.0 1024050.0 2152800.0 ;
      RECT  1020000.0 2158800.0 1021200.0 2160000.0 ;
      RECT  1023150.0 2158800.0 1026000.0 2160000.0 ;
      RECT  1020000.0 2151600.0 1021200.0 2152800.0 ;
      RECT  1022400.0 2151600.0 1023600.0 2152800.0 ;
      RECT  1020000.0 2158800.0 1021200.0 2160000.0 ;
      RECT  1024800.0 2158800.0 1026000.0 2160000.0 ;
      RECT  1020150.0 2149200.0 1021050.0 2166000.0 ;
      RECT  1023150.0 2149200.0 1024050.0 2166000.0 ;
      RECT  1030200.0 2151600.0 1031400.0 2152800.0 ;
      RECT  1032600.0 2151600.0 1034250.0 2152800.0 ;
      RECT  1030200.0 2158800.0 1031400.0 2160000.0 ;
      RECT  1033350.0 2158800.0 1036200.0 2160000.0 ;
      RECT  1030200.0 2151600.0 1031400.0 2152800.0 ;
      RECT  1032600.0 2151600.0 1033800.0 2152800.0 ;
      RECT  1030200.0 2158800.0 1031400.0 2160000.0 ;
      RECT  1035000.0 2158800.0 1036200.0 2160000.0 ;
      RECT  1030350.0 2149200.0 1031250.0 2166000.0 ;
      RECT  1033350.0 2149200.0 1034250.0 2166000.0 ;
      RECT  1040400.0 2151600.0 1041600.0 2152800.0 ;
      RECT  1042800.0 2151600.0 1044450.0 2152800.0 ;
      RECT  1040400.0 2158800.0 1041600.0 2160000.0 ;
      RECT  1043550.0 2158800.0 1046400.0 2160000.0 ;
      RECT  1040400.0 2151600.0 1041600.0 2152800.0 ;
      RECT  1042800.0 2151600.0 1044000.0 2152800.0 ;
      RECT  1040400.0 2158800.0 1041600.0 2160000.0 ;
      RECT  1045200.0 2158800.0 1046400.0 2160000.0 ;
      RECT  1040550.0 2149200.0 1041450.0 2166000.0 ;
      RECT  1043550.0 2149200.0 1044450.0 2166000.0 ;
      RECT  1050600.0 2151600.0 1051800.0 2152800.0 ;
      RECT  1053000.0 2151600.0 1054650.0 2152800.0 ;
      RECT  1050600.0 2158800.0 1051800.0 2160000.0 ;
      RECT  1053750.0 2158800.0 1056600.0 2160000.0 ;
      RECT  1050600.0 2151600.0 1051800.0 2152800.0 ;
      RECT  1053000.0 2151600.0 1054200.0 2152800.0 ;
      RECT  1050600.0 2158800.0 1051800.0 2160000.0 ;
      RECT  1055400.0 2158800.0 1056600.0 2160000.0 ;
      RECT  1050750.0 2149200.0 1051650.0 2166000.0 ;
      RECT  1053750.0 2149200.0 1054650.0 2166000.0 ;
      RECT  1060800.0 2151600.0 1062000.0 2152800.0 ;
      RECT  1063200.0 2151600.0 1064850.0 2152800.0 ;
      RECT  1060800.0 2158800.0 1062000.0 2160000.0 ;
      RECT  1063950.0 2158800.0 1066800.0 2160000.0 ;
      RECT  1060800.0 2151600.0 1062000.0 2152800.0 ;
      RECT  1063200.0 2151600.0 1064400.0 2152800.0 ;
      RECT  1060800.0 2158800.0 1062000.0 2160000.0 ;
      RECT  1065600.0 2158800.0 1066800.0 2160000.0 ;
      RECT  1060950.0 2149200.0 1061850.0 2166000.0 ;
      RECT  1063950.0 2149200.0 1064850.0 2166000.0 ;
      RECT  1071000.0 2151600.0 1072200.0 2152800.0 ;
      RECT  1073400.0 2151600.0 1075050.0 2152800.0 ;
      RECT  1071000.0 2158800.0 1072200.0 2160000.0 ;
      RECT  1074150.0 2158800.0 1077000.0 2160000.0 ;
      RECT  1071000.0 2151600.0 1072200.0 2152800.0 ;
      RECT  1073400.0 2151600.0 1074600.0 2152800.0 ;
      RECT  1071000.0 2158800.0 1072200.0 2160000.0 ;
      RECT  1075800.0 2158800.0 1077000.0 2160000.0 ;
      RECT  1071150.0 2149200.0 1072050.0 2166000.0 ;
      RECT  1074150.0 2149200.0 1075050.0 2166000.0 ;
      RECT  1081200.0 2151600.0 1082400.0 2152800.0 ;
      RECT  1083600.0 2151600.0 1085250.0 2152800.0 ;
      RECT  1081200.0 2158800.0 1082400.0 2160000.0 ;
      RECT  1084350.0 2158800.0 1087200.0 2160000.0 ;
      RECT  1081200.0 2151600.0 1082400.0 2152800.0 ;
      RECT  1083600.0 2151600.0 1084800.0 2152800.0 ;
      RECT  1081200.0 2158800.0 1082400.0 2160000.0 ;
      RECT  1086000.0 2158800.0 1087200.0 2160000.0 ;
      RECT  1081350.0 2149200.0 1082250.0 2166000.0 ;
      RECT  1084350.0 2149200.0 1085250.0 2166000.0 ;
      RECT  1091400.0 2151600.0 1092600.0 2152800.0 ;
      RECT  1093800.0 2151600.0 1095450.0 2152800.0 ;
      RECT  1091400.0 2158800.0 1092600.0 2160000.0 ;
      RECT  1094550.0 2158800.0 1097400.0 2160000.0 ;
      RECT  1091400.0 2151600.0 1092600.0 2152800.0 ;
      RECT  1093800.0 2151600.0 1095000.0 2152800.0 ;
      RECT  1091400.0 2158800.0 1092600.0 2160000.0 ;
      RECT  1096200.0 2158800.0 1097400.0 2160000.0 ;
      RECT  1091550.0 2149200.0 1092450.0 2166000.0 ;
      RECT  1094550.0 2149200.0 1095450.0 2166000.0 ;
      RECT  1101600.0 2151600.0 1102800.0 2152800.0 ;
      RECT  1104000.0 2151600.0 1105650.0 2152800.0 ;
      RECT  1101600.0 2158800.0 1102800.0 2160000.0 ;
      RECT  1104750.0 2158800.0 1107600.0 2160000.0 ;
      RECT  1101600.0 2151600.0 1102800.0 2152800.0 ;
      RECT  1104000.0 2151600.0 1105200.0 2152800.0 ;
      RECT  1101600.0 2158800.0 1102800.0 2160000.0 ;
      RECT  1106400.0 2158800.0 1107600.0 2160000.0 ;
      RECT  1101750.0 2149200.0 1102650.0 2166000.0 ;
      RECT  1104750.0 2149200.0 1105650.0 2166000.0 ;
      RECT  1111800.0 2151600.0 1113000.0 2152800.0 ;
      RECT  1114200.0 2151600.0 1115850.0 2152800.0 ;
      RECT  1111800.0 2158800.0 1113000.0 2160000.0 ;
      RECT  1114950.0 2158800.0 1117800.0 2160000.0 ;
      RECT  1111800.0 2151600.0 1113000.0 2152800.0 ;
      RECT  1114200.0 2151600.0 1115400.0 2152800.0 ;
      RECT  1111800.0 2158800.0 1113000.0 2160000.0 ;
      RECT  1116600.0 2158800.0 1117800.0 2160000.0 ;
      RECT  1111950.0 2149200.0 1112850.0 2166000.0 ;
      RECT  1114950.0 2149200.0 1115850.0 2166000.0 ;
      RECT  1122000.0 2151600.0 1123200.0 2152800.0 ;
      RECT  1124400.0 2151600.0 1126050.0 2152800.0 ;
      RECT  1122000.0 2158800.0 1123200.0 2160000.0 ;
      RECT  1125150.0 2158800.0 1128000.0 2160000.0 ;
      RECT  1122000.0 2151600.0 1123200.0 2152800.0 ;
      RECT  1124400.0 2151600.0 1125600.0 2152800.0 ;
      RECT  1122000.0 2158800.0 1123200.0 2160000.0 ;
      RECT  1126800.0 2158800.0 1128000.0 2160000.0 ;
      RECT  1122150.0 2149200.0 1123050.0 2166000.0 ;
      RECT  1125150.0 2149200.0 1126050.0 2166000.0 ;
      RECT  1132200.0 2151600.0 1133400.0 2152800.0 ;
      RECT  1134600.0 2151600.0 1136250.0 2152800.0 ;
      RECT  1132200.0 2158800.0 1133400.0 2160000.0 ;
      RECT  1135350.0 2158800.0 1138200.0 2160000.0 ;
      RECT  1132200.0 2151600.0 1133400.0 2152800.0 ;
      RECT  1134600.0 2151600.0 1135800.0 2152800.0 ;
      RECT  1132200.0 2158800.0 1133400.0 2160000.0 ;
      RECT  1137000.0 2158800.0 1138200.0 2160000.0 ;
      RECT  1132350.0 2149200.0 1133250.0 2166000.0 ;
      RECT  1135350.0 2149200.0 1136250.0 2166000.0 ;
      RECT  1142400.0 2151600.0 1143600.0 2152800.0 ;
      RECT  1144800.0 2151600.0 1146450.0 2152800.0 ;
      RECT  1142400.0 2158800.0 1143600.0 2160000.0 ;
      RECT  1145550.0 2158800.0 1148400.0 2160000.0 ;
      RECT  1142400.0 2151600.0 1143600.0 2152800.0 ;
      RECT  1144800.0 2151600.0 1146000.0 2152800.0 ;
      RECT  1142400.0 2158800.0 1143600.0 2160000.0 ;
      RECT  1147200.0 2158800.0 1148400.0 2160000.0 ;
      RECT  1142550.0 2149200.0 1143450.0 2166000.0 ;
      RECT  1145550.0 2149200.0 1146450.0 2166000.0 ;
      RECT  1152600.0 2151600.0 1153800.0 2152800.0 ;
      RECT  1155000.0 2151600.0 1156650.0 2152800.0 ;
      RECT  1152600.0 2158800.0 1153800.0 2160000.0 ;
      RECT  1155750.0 2158800.0 1158600.0 2160000.0 ;
      RECT  1152600.0 2151600.0 1153800.0 2152800.0 ;
      RECT  1155000.0 2151600.0 1156200.0 2152800.0 ;
      RECT  1152600.0 2158800.0 1153800.0 2160000.0 ;
      RECT  1157400.0 2158800.0 1158600.0 2160000.0 ;
      RECT  1152750.0 2149200.0 1153650.0 2166000.0 ;
      RECT  1155750.0 2149200.0 1156650.0 2166000.0 ;
      RECT  1162800.0 2151600.0 1164000.0 2152800.0 ;
      RECT  1165200.0 2151600.0 1166850.0 2152800.0 ;
      RECT  1162800.0 2158800.0 1164000.0 2160000.0 ;
      RECT  1165950.0 2158800.0 1168800.0 2160000.0 ;
      RECT  1162800.0 2151600.0 1164000.0 2152800.0 ;
      RECT  1165200.0 2151600.0 1166400.0 2152800.0 ;
      RECT  1162800.0 2158800.0 1164000.0 2160000.0 ;
      RECT  1167600.0 2158800.0 1168800.0 2160000.0 ;
      RECT  1162950.0 2149200.0 1163850.0 2166000.0 ;
      RECT  1165950.0 2149200.0 1166850.0 2166000.0 ;
      RECT  1173000.0 2151600.0 1174200.0 2152800.0 ;
      RECT  1175400.0 2151600.0 1177050.0 2152800.0 ;
      RECT  1173000.0 2158800.0 1174200.0 2160000.0 ;
      RECT  1176150.0 2158800.0 1179000.0 2160000.0 ;
      RECT  1173000.0 2151600.0 1174200.0 2152800.0 ;
      RECT  1175400.0 2151600.0 1176600.0 2152800.0 ;
      RECT  1173000.0 2158800.0 1174200.0 2160000.0 ;
      RECT  1177800.0 2158800.0 1179000.0 2160000.0 ;
      RECT  1173150.0 2149200.0 1174050.0 2166000.0 ;
      RECT  1176150.0 2149200.0 1177050.0 2166000.0 ;
      RECT  1183200.0 2151600.0 1184400.0 2152800.0 ;
      RECT  1185600.0 2151600.0 1187250.0 2152800.0 ;
      RECT  1183200.0 2158800.0 1184400.0 2160000.0 ;
      RECT  1186350.0 2158800.0 1189200.0 2160000.0 ;
      RECT  1183200.0 2151600.0 1184400.0 2152800.0 ;
      RECT  1185600.0 2151600.0 1186800.0 2152800.0 ;
      RECT  1183200.0 2158800.0 1184400.0 2160000.0 ;
      RECT  1188000.0 2158800.0 1189200.0 2160000.0 ;
      RECT  1183350.0 2149200.0 1184250.0 2166000.0 ;
      RECT  1186350.0 2149200.0 1187250.0 2166000.0 ;
      RECT  1193400.0 2151600.0 1194600.0 2152800.0 ;
      RECT  1195800.0 2151600.0 1197450.0 2152800.0 ;
      RECT  1193400.0 2158800.0 1194600.0 2160000.0 ;
      RECT  1196550.0 2158800.0 1199400.0 2160000.0 ;
      RECT  1193400.0 2151600.0 1194600.0 2152800.0 ;
      RECT  1195800.0 2151600.0 1197000.0 2152800.0 ;
      RECT  1193400.0 2158800.0 1194600.0 2160000.0 ;
      RECT  1198200.0 2158800.0 1199400.0 2160000.0 ;
      RECT  1193550.0 2149200.0 1194450.0 2166000.0 ;
      RECT  1196550.0 2149200.0 1197450.0 2166000.0 ;
      RECT  1203600.0 2151600.0 1204800.0 2152800.0 ;
      RECT  1206000.0 2151600.0 1207650.0 2152800.0 ;
      RECT  1203600.0 2158800.0 1204800.0 2160000.0 ;
      RECT  1206750.0 2158800.0 1209600.0 2160000.0 ;
      RECT  1203600.0 2151600.0 1204800.0 2152800.0 ;
      RECT  1206000.0 2151600.0 1207200.0 2152800.0 ;
      RECT  1203600.0 2158800.0 1204800.0 2160000.0 ;
      RECT  1208400.0 2158800.0 1209600.0 2160000.0 ;
      RECT  1203750.0 2149200.0 1204650.0 2166000.0 ;
      RECT  1206750.0 2149200.0 1207650.0 2166000.0 ;
      RECT  1213800.0 2151600.0 1215000.0 2152800.0 ;
      RECT  1216200.0 2151600.0 1217850.0 2152800.0 ;
      RECT  1213800.0 2158800.0 1215000.0 2160000.0 ;
      RECT  1216950.0 2158800.0 1219800.0 2160000.0 ;
      RECT  1213800.0 2151600.0 1215000.0 2152800.0 ;
      RECT  1216200.0 2151600.0 1217400.0 2152800.0 ;
      RECT  1213800.0 2158800.0 1215000.0 2160000.0 ;
      RECT  1218600.0 2158800.0 1219800.0 2160000.0 ;
      RECT  1213950.0 2149200.0 1214850.0 2166000.0 ;
      RECT  1216950.0 2149200.0 1217850.0 2166000.0 ;
      RECT  1224000.0 2151600.0 1225200.0 2152800.0 ;
      RECT  1226400.0 2151600.0 1228050.0 2152800.0 ;
      RECT  1224000.0 2158800.0 1225200.0 2160000.0 ;
      RECT  1227150.0 2158800.0 1230000.0 2160000.0 ;
      RECT  1224000.0 2151600.0 1225200.0 2152800.0 ;
      RECT  1226400.0 2151600.0 1227600.0 2152800.0 ;
      RECT  1224000.0 2158800.0 1225200.0 2160000.0 ;
      RECT  1228800.0 2158800.0 1230000.0 2160000.0 ;
      RECT  1224150.0 2149200.0 1225050.0 2166000.0 ;
      RECT  1227150.0 2149200.0 1228050.0 2166000.0 ;
      RECT  1234200.0 2151600.0 1235400.0 2152800.0 ;
      RECT  1236600.0 2151600.0 1238250.0 2152800.0 ;
      RECT  1234200.0 2158800.0 1235400.0 2160000.0 ;
      RECT  1237350.0 2158800.0 1240200.0 2160000.0 ;
      RECT  1234200.0 2151600.0 1235400.0 2152800.0 ;
      RECT  1236600.0 2151600.0 1237800.0 2152800.0 ;
      RECT  1234200.0 2158800.0 1235400.0 2160000.0 ;
      RECT  1239000.0 2158800.0 1240200.0 2160000.0 ;
      RECT  1234350.0 2149200.0 1235250.0 2166000.0 ;
      RECT  1237350.0 2149200.0 1238250.0 2166000.0 ;
      RECT  1244400.0 2151600.0 1245600.0 2152800.0 ;
      RECT  1246800.0 2151600.0 1248450.0 2152800.0 ;
      RECT  1244400.0 2158800.0 1245600.0 2160000.0 ;
      RECT  1247550.0 2158800.0 1250400.0 2160000.0 ;
      RECT  1244400.0 2151600.0 1245600.0 2152800.0 ;
      RECT  1246800.0 2151600.0 1248000.0 2152800.0 ;
      RECT  1244400.0 2158800.0 1245600.0 2160000.0 ;
      RECT  1249200.0 2158800.0 1250400.0 2160000.0 ;
      RECT  1244550.0 2149200.0 1245450.0 2166000.0 ;
      RECT  1247550.0 2149200.0 1248450.0 2166000.0 ;
      RECT  1254600.0 2151600.0 1255800.0 2152800.0 ;
      RECT  1257000.0 2151600.0 1258650.0 2152800.0 ;
      RECT  1254600.0 2158800.0 1255800.0 2160000.0 ;
      RECT  1257750.0 2158800.0 1260600.0 2160000.0 ;
      RECT  1254600.0 2151600.0 1255800.0 2152800.0 ;
      RECT  1257000.0 2151600.0 1258200.0 2152800.0 ;
      RECT  1254600.0 2158800.0 1255800.0 2160000.0 ;
      RECT  1259400.0 2158800.0 1260600.0 2160000.0 ;
      RECT  1254750.0 2149200.0 1255650.0 2166000.0 ;
      RECT  1257750.0 2149200.0 1258650.0 2166000.0 ;
      RECT  1264800.0 2151600.0 1266000.0 2152800.0 ;
      RECT  1267200.0 2151600.0 1268850.0 2152800.0 ;
      RECT  1264800.0 2158800.0 1266000.0 2160000.0 ;
      RECT  1267950.0 2158800.0 1270800.0 2160000.0 ;
      RECT  1264800.0 2151600.0 1266000.0 2152800.0 ;
      RECT  1267200.0 2151600.0 1268400.0 2152800.0 ;
      RECT  1264800.0 2158800.0 1266000.0 2160000.0 ;
      RECT  1269600.0 2158800.0 1270800.0 2160000.0 ;
      RECT  1264950.0 2149200.0 1265850.0 2166000.0 ;
      RECT  1267950.0 2149200.0 1268850.0 2166000.0 ;
      RECT  1275000.0 2151600.0 1276200.0 2152800.0 ;
      RECT  1277400.0 2151600.0 1279050.0 2152800.0 ;
      RECT  1275000.0 2158800.0 1276200.0 2160000.0 ;
      RECT  1278150.0 2158800.0 1281000.0 2160000.0 ;
      RECT  1275000.0 2151600.0 1276200.0 2152800.0 ;
      RECT  1277400.0 2151600.0 1278600.0 2152800.0 ;
      RECT  1275000.0 2158800.0 1276200.0 2160000.0 ;
      RECT  1279800.0 2158800.0 1281000.0 2160000.0 ;
      RECT  1275150.0 2149200.0 1276050.0 2166000.0 ;
      RECT  1278150.0 2149200.0 1279050.0 2166000.0 ;
      RECT  1285200.0 2151600.0 1286400.0 2152800.0 ;
      RECT  1287600.0 2151600.0 1289250.0 2152800.0 ;
      RECT  1285200.0 2158800.0 1286400.0 2160000.0 ;
      RECT  1288350.0 2158800.0 1291200.0 2160000.0 ;
      RECT  1285200.0 2151600.0 1286400.0 2152800.0 ;
      RECT  1287600.0 2151600.0 1288800.0 2152800.0 ;
      RECT  1285200.0 2158800.0 1286400.0 2160000.0 ;
      RECT  1290000.0 2158800.0 1291200.0 2160000.0 ;
      RECT  1285350.0 2149200.0 1286250.0 2166000.0 ;
      RECT  1288350.0 2149200.0 1289250.0 2166000.0 ;
      RECT  1295400.0 2151600.0 1296600.0 2152800.0 ;
      RECT  1297800.0 2151600.0 1299450.0 2152800.0 ;
      RECT  1295400.0 2158800.0 1296600.0 2160000.0 ;
      RECT  1298550.0 2158800.0 1301400.0 2160000.0 ;
      RECT  1295400.0 2151600.0 1296600.0 2152800.0 ;
      RECT  1297800.0 2151600.0 1299000.0 2152800.0 ;
      RECT  1295400.0 2158800.0 1296600.0 2160000.0 ;
      RECT  1300200.0 2158800.0 1301400.0 2160000.0 ;
      RECT  1295550.0 2149200.0 1296450.0 2166000.0 ;
      RECT  1298550.0 2149200.0 1299450.0 2166000.0 ;
      RECT  1305600.0 2151600.0 1306800.0 2152800.0 ;
      RECT  1308000.0 2151600.0 1309650.0 2152800.0 ;
      RECT  1305600.0 2158800.0 1306800.0 2160000.0 ;
      RECT  1308750.0 2158800.0 1311600.0 2160000.0 ;
      RECT  1305600.0 2151600.0 1306800.0 2152800.0 ;
      RECT  1308000.0 2151600.0 1309200.0 2152800.0 ;
      RECT  1305600.0 2158800.0 1306800.0 2160000.0 ;
      RECT  1310400.0 2158800.0 1311600.0 2160000.0 ;
      RECT  1305750.0 2149200.0 1306650.0 2166000.0 ;
      RECT  1308750.0 2149200.0 1309650.0 2166000.0 ;
      RECT  1315800.0 2151600.0 1317000.0 2152800.0 ;
      RECT  1318200.0 2151600.0 1319850.0 2152800.0 ;
      RECT  1315800.0 2158800.0 1317000.0 2160000.0 ;
      RECT  1318950.0 2158800.0 1321800.0 2160000.0 ;
      RECT  1315800.0 2151600.0 1317000.0 2152800.0 ;
      RECT  1318200.0 2151600.0 1319400.0 2152800.0 ;
      RECT  1315800.0 2158800.0 1317000.0 2160000.0 ;
      RECT  1320600.0 2158800.0 1321800.0 2160000.0 ;
      RECT  1315950.0 2149200.0 1316850.0 2166000.0 ;
      RECT  1318950.0 2149200.0 1319850.0 2166000.0 ;
      RECT  1326000.0 2151600.0 1327200.0 2152800.0 ;
      RECT  1328400.0 2151600.0 1330050.0 2152800.0 ;
      RECT  1326000.0 2158800.0 1327200.0 2160000.0 ;
      RECT  1329150.0 2158800.0 1332000.0 2160000.0 ;
      RECT  1326000.0 2151600.0 1327200.0 2152800.0 ;
      RECT  1328400.0 2151600.0 1329600.0 2152800.0 ;
      RECT  1326000.0 2158800.0 1327200.0 2160000.0 ;
      RECT  1330800.0 2158800.0 1332000.0 2160000.0 ;
      RECT  1326150.0 2149200.0 1327050.0 2166000.0 ;
      RECT  1329150.0 2149200.0 1330050.0 2166000.0 ;
      RECT  1336200.0 2151600.0 1337400.0 2152800.0 ;
      RECT  1338600.0 2151600.0 1340250.0 2152800.0 ;
      RECT  1336200.0 2158800.0 1337400.0 2160000.0 ;
      RECT  1339350.0 2158800.0 1342200.0 2160000.0 ;
      RECT  1336200.0 2151600.0 1337400.0 2152800.0 ;
      RECT  1338600.0 2151600.0 1339800.0 2152800.0 ;
      RECT  1336200.0 2158800.0 1337400.0 2160000.0 ;
      RECT  1341000.0 2158800.0 1342200.0 2160000.0 ;
      RECT  1336350.0 2149200.0 1337250.0 2166000.0 ;
      RECT  1339350.0 2149200.0 1340250.0 2166000.0 ;
      RECT  1346400.0 2151600.0 1347600.0 2152800.0 ;
      RECT  1348800.0 2151600.0 1350450.0 2152800.0 ;
      RECT  1346400.0 2158800.0 1347600.0 2160000.0 ;
      RECT  1349550.0 2158800.0 1352400.0 2160000.0 ;
      RECT  1346400.0 2151600.0 1347600.0 2152800.0 ;
      RECT  1348800.0 2151600.0 1350000.0 2152800.0 ;
      RECT  1346400.0 2158800.0 1347600.0 2160000.0 ;
      RECT  1351200.0 2158800.0 1352400.0 2160000.0 ;
      RECT  1346550.0 2149200.0 1347450.0 2166000.0 ;
      RECT  1349550.0 2149200.0 1350450.0 2166000.0 ;
      RECT  1356600.0 2151600.0 1357800.0 2152800.0 ;
      RECT  1359000.0 2151600.0 1360650.0 2152800.0 ;
      RECT  1356600.0 2158800.0 1357800.0 2160000.0 ;
      RECT  1359750.0 2158800.0 1362600.0 2160000.0 ;
      RECT  1356600.0 2151600.0 1357800.0 2152800.0 ;
      RECT  1359000.0 2151600.0 1360200.0 2152800.0 ;
      RECT  1356600.0 2158800.0 1357800.0 2160000.0 ;
      RECT  1361400.0 2158800.0 1362600.0 2160000.0 ;
      RECT  1356750.0 2149200.0 1357650.0 2166000.0 ;
      RECT  1359750.0 2149200.0 1360650.0 2166000.0 ;
      RECT  1366800.0 2151600.0 1368000.0 2152800.0 ;
      RECT  1369200.0 2151600.0 1370850.0 2152800.0 ;
      RECT  1366800.0 2158800.0 1368000.0 2160000.0 ;
      RECT  1369950.0 2158800.0 1372800.0 2160000.0 ;
      RECT  1366800.0 2151600.0 1368000.0 2152800.0 ;
      RECT  1369200.0 2151600.0 1370400.0 2152800.0 ;
      RECT  1366800.0 2158800.0 1368000.0 2160000.0 ;
      RECT  1371600.0 2158800.0 1372800.0 2160000.0 ;
      RECT  1366950.0 2149200.0 1367850.0 2166000.0 ;
      RECT  1369950.0 2149200.0 1370850.0 2166000.0 ;
      RECT  1377000.0 2151600.0 1378200.0 2152800.0 ;
      RECT  1379400.0 2151600.0 1381050.0 2152800.0 ;
      RECT  1377000.0 2158800.0 1378200.0 2160000.0 ;
      RECT  1380150.0 2158800.0 1383000.0 2160000.0 ;
      RECT  1377000.0 2151600.0 1378200.0 2152800.0 ;
      RECT  1379400.0 2151600.0 1380600.0 2152800.0 ;
      RECT  1377000.0 2158800.0 1378200.0 2160000.0 ;
      RECT  1381800.0 2158800.0 1383000.0 2160000.0 ;
      RECT  1377150.0 2149200.0 1378050.0 2166000.0 ;
      RECT  1380150.0 2149200.0 1381050.0 2166000.0 ;
      RECT  1387200.0 2151600.0 1388400.0 2152800.0 ;
      RECT  1389600.0 2151600.0 1391250.0 2152800.0 ;
      RECT  1387200.0 2158800.0 1388400.0 2160000.0 ;
      RECT  1390350.0 2158800.0 1393200.0 2160000.0 ;
      RECT  1387200.0 2151600.0 1388400.0 2152800.0 ;
      RECT  1389600.0 2151600.0 1390800.0 2152800.0 ;
      RECT  1387200.0 2158800.0 1388400.0 2160000.0 ;
      RECT  1392000.0 2158800.0 1393200.0 2160000.0 ;
      RECT  1387350.0 2149200.0 1388250.0 2166000.0 ;
      RECT  1390350.0 2149200.0 1391250.0 2166000.0 ;
      RECT  1397400.0 2151600.0 1398600.0 2152800.0 ;
      RECT  1399800.0 2151600.0 1401450.0 2152800.0 ;
      RECT  1397400.0 2158800.0 1398600.0 2160000.0 ;
      RECT  1400550.0 2158800.0 1403400.0 2160000.0 ;
      RECT  1397400.0 2151600.0 1398600.0 2152800.0 ;
      RECT  1399800.0 2151600.0 1401000.0 2152800.0 ;
      RECT  1397400.0 2158800.0 1398600.0 2160000.0 ;
      RECT  1402200.0 2158800.0 1403400.0 2160000.0 ;
      RECT  1397550.0 2149200.0 1398450.0 2166000.0 ;
      RECT  1400550.0 2149200.0 1401450.0 2166000.0 ;
      RECT  1407600.0 2151600.0 1408800.0 2152800.0 ;
      RECT  1410000.0 2151600.0 1411650.0 2152800.0 ;
      RECT  1407600.0 2158800.0 1408800.0 2160000.0 ;
      RECT  1410750.0 2158800.0 1413600.0 2160000.0 ;
      RECT  1407600.0 2151600.0 1408800.0 2152800.0 ;
      RECT  1410000.0 2151600.0 1411200.0 2152800.0 ;
      RECT  1407600.0 2158800.0 1408800.0 2160000.0 ;
      RECT  1412400.0 2158800.0 1413600.0 2160000.0 ;
      RECT  1407750.0 2149200.0 1408650.0 2166000.0 ;
      RECT  1410750.0 2149200.0 1411650.0 2166000.0 ;
      RECT  1417800.0 2151600.0 1419000.0 2152800.0 ;
      RECT  1420200.0 2151600.0 1421850.0 2152800.0 ;
      RECT  1417800.0 2158800.0 1419000.0 2160000.0 ;
      RECT  1420950.0 2158800.0 1423800.0 2160000.0 ;
      RECT  1417800.0 2151600.0 1419000.0 2152800.0 ;
      RECT  1420200.0 2151600.0 1421400.0 2152800.0 ;
      RECT  1417800.0 2158800.0 1419000.0 2160000.0 ;
      RECT  1422600.0 2158800.0 1423800.0 2160000.0 ;
      RECT  1417950.0 2149200.0 1418850.0 2166000.0 ;
      RECT  1420950.0 2149200.0 1421850.0 2166000.0 ;
      RECT  1428000.0 2151600.0 1429200.0 2152800.0 ;
      RECT  1430400.0 2151600.0 1432050.0 2152800.0 ;
      RECT  1428000.0 2158800.0 1429200.0 2160000.0 ;
      RECT  1431150.0 2158800.0 1434000.0 2160000.0 ;
      RECT  1428000.0 2151600.0 1429200.0 2152800.0 ;
      RECT  1430400.0 2151600.0 1431600.0 2152800.0 ;
      RECT  1428000.0 2158800.0 1429200.0 2160000.0 ;
      RECT  1432800.0 2158800.0 1434000.0 2160000.0 ;
      RECT  1428150.0 2149200.0 1429050.0 2166000.0 ;
      RECT  1431150.0 2149200.0 1432050.0 2166000.0 ;
      RECT  1438200.0 2151600.0 1439400.0 2152800.0 ;
      RECT  1440600.0 2151600.0 1442250.0 2152800.0 ;
      RECT  1438200.0 2158800.0 1439400.0 2160000.0 ;
      RECT  1441350.0 2158800.0 1444200.0 2160000.0 ;
      RECT  1438200.0 2151600.0 1439400.0 2152800.0 ;
      RECT  1440600.0 2151600.0 1441800.0 2152800.0 ;
      RECT  1438200.0 2158800.0 1439400.0 2160000.0 ;
      RECT  1443000.0 2158800.0 1444200.0 2160000.0 ;
      RECT  1438350.0 2149200.0 1439250.0 2166000.0 ;
      RECT  1441350.0 2149200.0 1442250.0 2166000.0 ;
      RECT  1448400.0 2151600.0 1449600.0 2152800.0 ;
      RECT  1450800.0 2151600.0 1452450.0 2152800.0 ;
      RECT  1448400.0 2158800.0 1449600.0 2160000.0 ;
      RECT  1451550.0 2158800.0 1454400.0 2160000.0 ;
      RECT  1448400.0 2151600.0 1449600.0 2152800.0 ;
      RECT  1450800.0 2151600.0 1452000.0 2152800.0 ;
      RECT  1448400.0 2158800.0 1449600.0 2160000.0 ;
      RECT  1453200.0 2158800.0 1454400.0 2160000.0 ;
      RECT  1448550.0 2149200.0 1449450.0 2166000.0 ;
      RECT  1451550.0 2149200.0 1452450.0 2166000.0 ;
      RECT  1458600.0 2151600.0 1459800.0 2152800.0 ;
      RECT  1461000.0 2151600.0 1462650.0 2152800.0 ;
      RECT  1458600.0 2158800.0 1459800.0 2160000.0 ;
      RECT  1461750.0 2158800.0 1464600.0 2160000.0 ;
      RECT  1458600.0 2151600.0 1459800.0 2152800.0 ;
      RECT  1461000.0 2151600.0 1462200.0 2152800.0 ;
      RECT  1458600.0 2158800.0 1459800.0 2160000.0 ;
      RECT  1463400.0 2158800.0 1464600.0 2160000.0 ;
      RECT  1458750.0 2149200.0 1459650.0 2166000.0 ;
      RECT  1461750.0 2149200.0 1462650.0 2166000.0 ;
      RECT  1468800.0 2151600.0 1470000.0 2152800.0 ;
      RECT  1471200.0 2151600.0 1472850.0 2152800.0 ;
      RECT  1468800.0 2158800.0 1470000.0 2160000.0 ;
      RECT  1471950.0 2158800.0 1474800.0 2160000.0 ;
      RECT  1468800.0 2151600.0 1470000.0 2152800.0 ;
      RECT  1471200.0 2151600.0 1472400.0 2152800.0 ;
      RECT  1468800.0 2158800.0 1470000.0 2160000.0 ;
      RECT  1473600.0 2158800.0 1474800.0 2160000.0 ;
      RECT  1468950.0 2149200.0 1469850.0 2166000.0 ;
      RECT  1471950.0 2149200.0 1472850.0 2166000.0 ;
      RECT  1479000.0 2151600.0 1480200.0 2152800.0 ;
      RECT  1481400.0 2151600.0 1483050.0 2152800.0 ;
      RECT  1479000.0 2158800.0 1480200.0 2160000.0 ;
      RECT  1482150.0 2158800.0 1485000.0 2160000.0 ;
      RECT  1479000.0 2151600.0 1480200.0 2152800.0 ;
      RECT  1481400.0 2151600.0 1482600.0 2152800.0 ;
      RECT  1479000.0 2158800.0 1480200.0 2160000.0 ;
      RECT  1483800.0 2158800.0 1485000.0 2160000.0 ;
      RECT  1479150.0 2149200.0 1480050.0 2166000.0 ;
      RECT  1482150.0 2149200.0 1483050.0 2166000.0 ;
      RECT  1489200.0 2151600.0 1490400.0 2152800.0 ;
      RECT  1491600.0 2151600.0 1493250.0 2152800.0 ;
      RECT  1489200.0 2158800.0 1490400.0 2160000.0 ;
      RECT  1492350.0 2158800.0 1495200.0 2160000.0 ;
      RECT  1489200.0 2151600.0 1490400.0 2152800.0 ;
      RECT  1491600.0 2151600.0 1492800.0 2152800.0 ;
      RECT  1489200.0 2158800.0 1490400.0 2160000.0 ;
      RECT  1494000.0 2158800.0 1495200.0 2160000.0 ;
      RECT  1489350.0 2149200.0 1490250.0 2166000.0 ;
      RECT  1492350.0 2149200.0 1493250.0 2166000.0 ;
      RECT  1499400.0 2151600.0 1500600.0 2152800.0 ;
      RECT  1501800.0 2151600.0 1503450.0 2152800.0 ;
      RECT  1499400.0 2158800.0 1500600.0 2160000.0 ;
      RECT  1502550.0 2158800.0 1505400.0 2160000.0 ;
      RECT  1499400.0 2151600.0 1500600.0 2152800.0 ;
      RECT  1501800.0 2151600.0 1503000.0 2152800.0 ;
      RECT  1499400.0 2158800.0 1500600.0 2160000.0 ;
      RECT  1504200.0 2158800.0 1505400.0 2160000.0 ;
      RECT  1499550.0 2149200.0 1500450.0 2166000.0 ;
      RECT  1502550.0 2149200.0 1503450.0 2166000.0 ;
      RECT  1509600.0 2151600.0 1510800.0 2152800.0 ;
      RECT  1512000.0 2151600.0 1513650.0 2152800.0 ;
      RECT  1509600.0 2158800.0 1510800.0 2160000.0 ;
      RECT  1512750.0 2158800.0 1515600.0 2160000.0 ;
      RECT  1509600.0 2151600.0 1510800.0 2152800.0 ;
      RECT  1512000.0 2151600.0 1513200.0 2152800.0 ;
      RECT  1509600.0 2158800.0 1510800.0 2160000.0 ;
      RECT  1514400.0 2158800.0 1515600.0 2160000.0 ;
      RECT  1509750.0 2149200.0 1510650.0 2166000.0 ;
      RECT  1512750.0 2149200.0 1513650.0 2166000.0 ;
      RECT  1519800.0 2151600.0 1521000.0 2152800.0 ;
      RECT  1522200.0 2151600.0 1523850.0 2152800.0 ;
      RECT  1519800.0 2158800.0 1521000.0 2160000.0 ;
      RECT  1522950.0 2158800.0 1525800.0 2160000.0 ;
      RECT  1519800.0 2151600.0 1521000.0 2152800.0 ;
      RECT  1522200.0 2151600.0 1523400.0 2152800.0 ;
      RECT  1519800.0 2158800.0 1521000.0 2160000.0 ;
      RECT  1524600.0 2158800.0 1525800.0 2160000.0 ;
      RECT  1519950.0 2149200.0 1520850.0 2166000.0 ;
      RECT  1522950.0 2149200.0 1523850.0 2166000.0 ;
      RECT  224550.0 2149200.0 225450.0 2166000.0 ;
      RECT  227550.0 2149200.0 228450.0 2166000.0 ;
      RECT  234750.0 2149200.0 235650.0 2166000.0 ;
      RECT  237750.0 2149200.0 238650.0 2166000.0 ;
      RECT  244950.0 2149200.0 245850.0 2166000.0 ;
      RECT  247950.0 2149200.0 248850.0 2166000.0 ;
      RECT  255150.0 2149200.0 256050.0 2166000.0 ;
      RECT  258150.0 2149200.0 259050.0 2166000.0 ;
      RECT  265350.0 2149200.0 266250.0 2166000.0 ;
      RECT  268350.0 2149200.0 269250.0 2166000.0 ;
      RECT  275550.0 2149200.0 276450.0 2166000.0 ;
      RECT  278550.0 2149200.0 279450.0 2166000.0 ;
      RECT  285750.0 2149200.0 286650.0 2166000.0 ;
      RECT  288750.0 2149200.0 289650.0 2166000.0 ;
      RECT  295950.0 2149200.0 296850.0 2166000.0 ;
      RECT  298950.0 2149200.0 299850.0 2166000.0 ;
      RECT  306150.0 2149200.0 307050.0 2166000.0 ;
      RECT  309150.0 2149200.0 310050.0 2166000.0 ;
      RECT  316350.0 2149200.0 317250.0 2166000.0 ;
      RECT  319350.0 2149200.0 320250.0 2166000.0 ;
      RECT  326550.0 2149200.0 327450.0 2166000.0 ;
      RECT  329550.0 2149200.0 330450.0 2166000.0 ;
      RECT  336750.0 2149200.0 337650.0 2166000.0 ;
      RECT  339750.0 2149200.0 340650.0 2166000.0 ;
      RECT  346950.0 2149200.0 347850.0 2166000.0 ;
      RECT  349950.0 2149200.0 350850.0 2166000.0 ;
      RECT  357150.0 2149200.0 358050.0 2166000.0 ;
      RECT  360150.0 2149200.0 361050.0 2166000.0 ;
      RECT  367350.0 2149200.0 368250.0 2166000.0 ;
      RECT  370350.0 2149200.0 371250.0 2166000.0 ;
      RECT  377550.0 2149200.0 378450.0 2166000.0 ;
      RECT  380550.0 2149200.0 381450.0 2166000.0 ;
      RECT  387750.0 2149200.0 388650.0 2166000.0 ;
      RECT  390750.0 2149200.0 391650.0 2166000.0 ;
      RECT  397950.0 2149200.0 398850.0 2166000.0 ;
      RECT  400950.0 2149200.0 401850.0 2166000.0 ;
      RECT  408150.0 2149200.0 409050.0 2166000.0 ;
      RECT  411150.0 2149200.0 412050.0 2166000.0 ;
      RECT  418350.0 2149200.0 419250.0 2166000.0 ;
      RECT  421350.0 2149200.0 422250.0 2166000.0 ;
      RECT  428550.0 2149200.0 429450.0 2166000.0 ;
      RECT  431550.0 2149200.0 432450.0 2166000.0 ;
      RECT  438750.0 2149200.0 439650.0 2166000.0 ;
      RECT  441750.0 2149200.0 442650.0 2166000.0 ;
      RECT  448950.0 2149200.0 449850.0 2166000.0 ;
      RECT  451950.0 2149200.0 452850.0 2166000.0 ;
      RECT  459150.0 2149200.0 460050.0 2166000.0 ;
      RECT  462150.0 2149200.0 463050.0 2166000.0 ;
      RECT  469350.0 2149200.0 470250.0 2166000.0 ;
      RECT  472350.0 2149200.0 473250.0 2166000.0 ;
      RECT  479550.0 2149200.0 480450.0 2166000.0 ;
      RECT  482550.0 2149200.0 483450.0 2166000.0 ;
      RECT  489750.0 2149200.0 490650.0 2166000.0 ;
      RECT  492750.0 2149200.0 493650.0 2166000.0 ;
      RECT  499950.0 2149200.0 500850.0 2166000.0 ;
      RECT  502950.0 2149200.0 503850.0 2166000.0 ;
      RECT  510150.0 2149200.0 511050.0 2166000.0 ;
      RECT  513150.0 2149200.0 514050.0 2166000.0 ;
      RECT  520350.0 2149200.0 521250.0 2166000.0 ;
      RECT  523350.0 2149200.0 524250.0 2166000.0 ;
      RECT  530550.0 2149200.0 531450.0 2166000.0 ;
      RECT  533550.0 2149200.0 534450.0 2166000.0 ;
      RECT  540750.0 2149200.0 541650.0 2166000.0 ;
      RECT  543750.0 2149200.0 544650.0 2166000.0 ;
      RECT  550950.0 2149200.0 551850.0 2166000.0 ;
      RECT  553950.0 2149200.0 554850.0 2166000.0 ;
      RECT  561150.0 2149200.0 562050.0 2166000.0 ;
      RECT  564150.0 2149200.0 565050.0 2166000.0 ;
      RECT  571350.0 2149200.0 572250.0 2166000.0 ;
      RECT  574350.0 2149200.0 575250.0 2166000.0 ;
      RECT  581550.0 2149200.0 582450.0 2166000.0 ;
      RECT  584550.0 2149200.0 585450.0 2166000.0 ;
      RECT  591750.0 2149200.0 592650.0 2166000.0 ;
      RECT  594750.0 2149200.0 595650.0 2166000.0 ;
      RECT  601950.0 2149200.0 602850.0 2166000.0 ;
      RECT  604950.0 2149200.0 605850.0 2166000.0 ;
      RECT  612150.0 2149200.0 613050.0 2166000.0 ;
      RECT  615150.0 2149200.0 616050.0 2166000.0 ;
      RECT  622350.0 2149200.0 623250.0 2166000.0 ;
      RECT  625350.0 2149200.0 626250.0 2166000.0 ;
      RECT  632550.0 2149200.0 633450.0 2166000.0 ;
      RECT  635550.0 2149200.0 636450.0 2166000.0 ;
      RECT  642750.0 2149200.0 643650.0 2166000.0 ;
      RECT  645750.0 2149200.0 646650.0 2166000.0 ;
      RECT  652950.0 2149200.0 653850.0 2166000.0 ;
      RECT  655950.0 2149200.0 656850.0 2166000.0 ;
      RECT  663150.0 2149200.0 664050.0 2166000.0 ;
      RECT  666150.0 2149200.0 667050.0 2166000.0 ;
      RECT  673350.0 2149200.0 674250.0 2166000.0 ;
      RECT  676350.0 2149200.0 677250.0 2166000.0 ;
      RECT  683550.0 2149200.0 684450.0 2166000.0 ;
      RECT  686550.0 2149200.0 687450.0 2166000.0 ;
      RECT  693750.0 2149200.0 694650.0 2166000.0 ;
      RECT  696750.0 2149200.0 697650.0 2166000.0 ;
      RECT  703950.0 2149200.0 704850.0 2166000.0 ;
      RECT  706950.0 2149200.0 707850.0 2166000.0 ;
      RECT  714150.0 2149200.0 715050.0 2166000.0 ;
      RECT  717150.0 2149200.0 718050.0 2166000.0 ;
      RECT  724350.0 2149200.0 725250.0 2166000.0 ;
      RECT  727350.0 2149200.0 728250.0 2166000.0 ;
      RECT  734550.0 2149200.0 735450.0 2166000.0 ;
      RECT  737550.0 2149200.0 738450.0 2166000.0 ;
      RECT  744750.0 2149200.0 745650.0 2166000.0 ;
      RECT  747750.0 2149200.0 748650.0 2166000.0 ;
      RECT  754950.0 2149200.0 755850.0 2166000.0 ;
      RECT  757950.0 2149200.0 758850.0 2166000.0 ;
      RECT  765150.0 2149200.0 766050.0 2166000.0 ;
      RECT  768150.0 2149200.0 769050.0 2166000.0 ;
      RECT  775350.0 2149200.0 776250.0 2166000.0 ;
      RECT  778350.0 2149200.0 779250.0 2166000.0 ;
      RECT  785550.0 2149200.0 786450.0 2166000.0 ;
      RECT  788550.0 2149200.0 789450.0 2166000.0 ;
      RECT  795750.0 2149200.0 796650.0 2166000.0 ;
      RECT  798750.0 2149200.0 799650.0 2166000.0 ;
      RECT  805950.0 2149200.0 806850.0 2166000.0 ;
      RECT  808950.0 2149200.0 809850.0 2166000.0 ;
      RECT  816150.0 2149200.0 817050.0 2166000.0 ;
      RECT  819150.0 2149200.0 820050.0 2166000.0 ;
      RECT  826350.0 2149200.0 827250.0 2166000.0 ;
      RECT  829350.0 2149200.0 830250.0 2166000.0 ;
      RECT  836550.0 2149200.0 837450.0 2166000.0 ;
      RECT  839550.0 2149200.0 840450.0 2166000.0 ;
      RECT  846750.0 2149200.0 847650.0 2166000.0 ;
      RECT  849750.0 2149200.0 850650.0 2166000.0 ;
      RECT  856950.0 2149200.0 857850.0 2166000.0 ;
      RECT  859950.0 2149200.0 860850.0 2166000.0 ;
      RECT  867150.0 2149200.0 868050.0 2166000.0 ;
      RECT  870150.0 2149200.0 871050.0 2166000.0 ;
      RECT  877350.0 2149200.0 878250.0 2166000.0 ;
      RECT  880350.0 2149200.0 881250.0 2166000.0 ;
      RECT  887550.0 2149200.0 888450.0 2166000.0 ;
      RECT  890550.0 2149200.0 891450.0 2166000.0 ;
      RECT  897750.0 2149200.0 898650.0 2166000.0 ;
      RECT  900750.0 2149200.0 901650.0 2166000.0 ;
      RECT  907950.0 2149200.0 908850.0 2166000.0 ;
      RECT  910950.0 2149200.0 911850.0 2166000.0 ;
      RECT  918150.0 2149200.0 919050.0 2166000.0 ;
      RECT  921150.0 2149200.0 922050.0 2166000.0 ;
      RECT  928350.0 2149200.0 929250.0 2166000.0 ;
      RECT  931350.0 2149200.0 932250.0 2166000.0 ;
      RECT  938550.0 2149200.0 939450.0 2166000.0 ;
      RECT  941550.0 2149200.0 942450.0 2166000.0 ;
      RECT  948750.0 2149200.0 949650.0 2166000.0 ;
      RECT  951750.0 2149200.0 952650.0 2166000.0 ;
      RECT  958950.0 2149200.0 959850.0 2166000.0 ;
      RECT  961950.0 2149200.0 962850.0 2166000.0 ;
      RECT  969150.0 2149200.0 970050.0 2166000.0 ;
      RECT  972150.0 2149200.0 973050.0 2166000.0 ;
      RECT  979350.0 2149200.0 980250.0 2166000.0 ;
      RECT  982350.0 2149200.0 983250.0 2166000.0 ;
      RECT  989550.0 2149200.0 990450.0 2166000.0 ;
      RECT  992550.0 2149200.0 993450.0 2166000.0 ;
      RECT  999750.0 2149200.0 1000650.0 2166000.0 ;
      RECT  1002750.0 2149200.0 1003650.0 2166000.0 ;
      RECT  1009950.0 2149200.0 1010850.0 2166000.0 ;
      RECT  1012950.0 2149200.0 1013850.0 2166000.0 ;
      RECT  1020150.0 2149200.0 1021050.0 2166000.0 ;
      RECT  1023150.0 2149200.0 1024050.0 2166000.0 ;
      RECT  1030350.0 2149200.0 1031250.0 2166000.0 ;
      RECT  1033350.0 2149200.0 1034250.0 2166000.0 ;
      RECT  1040550.0 2149200.0 1041450.0 2166000.0 ;
      RECT  1043550.0 2149200.0 1044450.0 2166000.0 ;
      RECT  1050750.0 2149200.0 1051650.0 2166000.0 ;
      RECT  1053750.0 2149200.0 1054650.0 2166000.0 ;
      RECT  1060950.0 2149200.0 1061850.0 2166000.0 ;
      RECT  1063950.0 2149200.0 1064850.0 2166000.0 ;
      RECT  1071150.0 2149200.0 1072050.0 2166000.0 ;
      RECT  1074150.0 2149200.0 1075050.0 2166000.0 ;
      RECT  1081350.0 2149200.0 1082250.0 2166000.0 ;
      RECT  1084350.0 2149200.0 1085250.0 2166000.0 ;
      RECT  1091550.0 2149200.0 1092450.0 2166000.0 ;
      RECT  1094550.0 2149200.0 1095450.0 2166000.0 ;
      RECT  1101750.0 2149200.0 1102650.0 2166000.0 ;
      RECT  1104750.0 2149200.0 1105650.0 2166000.0 ;
      RECT  1111950.0 2149200.0 1112850.0 2166000.0 ;
      RECT  1114950.0 2149200.0 1115850.0 2166000.0 ;
      RECT  1122150.0 2149200.0 1123050.0 2166000.0 ;
      RECT  1125150.0 2149200.0 1126050.0 2166000.0 ;
      RECT  1132350.0 2149200.0 1133250.0 2166000.0 ;
      RECT  1135350.0 2149200.0 1136250.0 2166000.0 ;
      RECT  1142550.0 2149200.0 1143450.0 2166000.0 ;
      RECT  1145550.0 2149200.0 1146450.0 2166000.0 ;
      RECT  1152750.0 2149200.0 1153650.0 2166000.0 ;
      RECT  1155750.0 2149200.0 1156650.0 2166000.0 ;
      RECT  1162950.0 2149200.0 1163850.0 2166000.0 ;
      RECT  1165950.0 2149200.0 1166850.0 2166000.0 ;
      RECT  1173150.0 2149200.0 1174050.0 2166000.0 ;
      RECT  1176150.0 2149200.0 1177050.0 2166000.0 ;
      RECT  1183350.0 2149200.0 1184250.0 2166000.0 ;
      RECT  1186350.0 2149200.0 1187250.0 2166000.0 ;
      RECT  1193550.0 2149200.0 1194450.0 2166000.0 ;
      RECT  1196550.0 2149200.0 1197450.0 2166000.0 ;
      RECT  1203750.0 2149200.0 1204650.0 2166000.0 ;
      RECT  1206750.0 2149200.0 1207650.0 2166000.0 ;
      RECT  1213950.0 2149200.0 1214850.0 2166000.0 ;
      RECT  1216950.0 2149200.0 1217850.0 2166000.0 ;
      RECT  1224150.0 2149200.0 1225050.0 2166000.0 ;
      RECT  1227150.0 2149200.0 1228050.0 2166000.0 ;
      RECT  1234350.0 2149200.0 1235250.0 2166000.0 ;
      RECT  1237350.0 2149200.0 1238250.0 2166000.0 ;
      RECT  1244550.0 2149200.0 1245450.0 2166000.0 ;
      RECT  1247550.0 2149200.0 1248450.0 2166000.0 ;
      RECT  1254750.0 2149200.0 1255650.0 2166000.0 ;
      RECT  1257750.0 2149200.0 1258650.0 2166000.0 ;
      RECT  1264950.0 2149200.0 1265850.0 2166000.0 ;
      RECT  1267950.0 2149200.0 1268850.0 2166000.0 ;
      RECT  1275150.0 2149200.0 1276050.0 2166000.0 ;
      RECT  1278150.0 2149200.0 1279050.0 2166000.0 ;
      RECT  1285350.0 2149200.0 1286250.0 2166000.0 ;
      RECT  1288350.0 2149200.0 1289250.0 2166000.0 ;
      RECT  1295550.0 2149200.0 1296450.0 2166000.0 ;
      RECT  1298550.0 2149200.0 1299450.0 2166000.0 ;
      RECT  1305750.0 2149200.0 1306650.0 2166000.0 ;
      RECT  1308750.0 2149200.0 1309650.0 2166000.0 ;
      RECT  1315950.0 2149200.0 1316850.0 2166000.0 ;
      RECT  1318950.0 2149200.0 1319850.0 2166000.0 ;
      RECT  1326150.0 2149200.0 1327050.0 2166000.0 ;
      RECT  1329150.0 2149200.0 1330050.0 2166000.0 ;
      RECT  1336350.0 2149200.0 1337250.0 2166000.0 ;
      RECT  1339350.0 2149200.0 1340250.0 2166000.0 ;
      RECT  1346550.0 2149200.0 1347450.0 2166000.0 ;
      RECT  1349550.0 2149200.0 1350450.0 2166000.0 ;
      RECT  1356750.0 2149200.0 1357650.0 2166000.0 ;
      RECT  1359750.0 2149200.0 1360650.0 2166000.0 ;
      RECT  1366950.0 2149200.0 1367850.0 2166000.0 ;
      RECT  1369950.0 2149200.0 1370850.0 2166000.0 ;
      RECT  1377150.0 2149200.0 1378050.0 2166000.0 ;
      RECT  1380150.0 2149200.0 1381050.0 2166000.0 ;
      RECT  1387350.0 2149200.0 1388250.0 2166000.0 ;
      RECT  1390350.0 2149200.0 1391250.0 2166000.0 ;
      RECT  1397550.0 2149200.0 1398450.0 2166000.0 ;
      RECT  1400550.0 2149200.0 1401450.0 2166000.0 ;
      RECT  1407750.0 2149200.0 1408650.0 2166000.0 ;
      RECT  1410750.0 2149200.0 1411650.0 2166000.0 ;
      RECT  1417950.0 2149200.0 1418850.0 2166000.0 ;
      RECT  1420950.0 2149200.0 1421850.0 2166000.0 ;
      RECT  1428150.0 2149200.0 1429050.0 2166000.0 ;
      RECT  1431150.0 2149200.0 1432050.0 2166000.0 ;
      RECT  1438350.0 2149200.0 1439250.0 2166000.0 ;
      RECT  1441350.0 2149200.0 1442250.0 2166000.0 ;
      RECT  1448550.0 2149200.0 1449450.0 2166000.0 ;
      RECT  1451550.0 2149200.0 1452450.0 2166000.0 ;
      RECT  1458750.0 2149200.0 1459650.0 2166000.0 ;
      RECT  1461750.0 2149200.0 1462650.0 2166000.0 ;
      RECT  1468950.0 2149200.0 1469850.0 2166000.0 ;
      RECT  1471950.0 2149200.0 1472850.0 2166000.0 ;
      RECT  1479150.0 2149200.0 1480050.0 2166000.0 ;
      RECT  1482150.0 2149200.0 1483050.0 2166000.0 ;
      RECT  1489350.0 2149200.0 1490250.0 2166000.0 ;
      RECT  1492350.0 2149200.0 1493250.0 2166000.0 ;
      RECT  1499550.0 2149200.0 1500450.0 2166000.0 ;
      RECT  1502550.0 2149200.0 1503450.0 2166000.0 ;
      RECT  1509750.0 2149200.0 1510650.0 2166000.0 ;
      RECT  1512750.0 2149200.0 1513650.0 2166000.0 ;
      RECT  1519950.0 2149200.0 1520850.0 2166000.0 ;
      RECT  1522950.0 2149200.0 1523850.0 2166000.0 ;
      RECT  234600.0 342750.0 235500.0 353250.0 ;
      RECT  237600.0 340650.0 238500.0 353250.0 ;
      RECT  244800.0 342750.0 245700.0 353250.0 ;
      RECT  247800.0 340650.0 248700.0 353250.0 ;
      RECT  255000.0 342750.0 255900.0 353250.0 ;
      RECT  258000.0 340650.0 258900.0 353250.0 ;
      RECT  275400.0 342750.0 276300.0 353250.0 ;
      RECT  278400.0 340650.0 279300.0 353250.0 ;
      RECT  285600.0 342750.0 286500.0 353250.0 ;
      RECT  288600.0 340650.0 289500.0 353250.0 ;
      RECT  295800.0 342750.0 296700.0 353250.0 ;
      RECT  298800.0 340650.0 299700.0 353250.0 ;
      RECT  316200.0 342750.0 317100.0 353250.0 ;
      RECT  319200.0 340650.0 320100.0 353250.0 ;
      RECT  326400.0 342750.0 327300.0 353250.0 ;
      RECT  329400.0 340650.0 330300.0 353250.0 ;
      RECT  336600.0 342750.0 337500.0 353250.0 ;
      RECT  339600.0 340650.0 340500.0 353250.0 ;
      RECT  357000.0 342750.0 357900.0 353250.0 ;
      RECT  360000.0 340650.0 360900.0 353250.0 ;
      RECT  367200.0 342750.0 368100.0 353250.0 ;
      RECT  370200.0 340650.0 371100.0 353250.0 ;
      RECT  377400.0 342750.0 378300.0 353250.0 ;
      RECT  380400.0 340650.0 381300.0 353250.0 ;
      RECT  397800.0 342750.0 398700.0 353250.0 ;
      RECT  400800.0 340650.0 401700.0 353250.0 ;
      RECT  408000.0 342750.0 408900.0 353250.0 ;
      RECT  411000.0 340650.0 411900.0 353250.0 ;
      RECT  418200.0 342750.0 419100.0 353250.0 ;
      RECT  421200.0 340650.0 422100.0 353250.0 ;
      RECT  438600.0 342750.0 439500.0 353250.0 ;
      RECT  441600.0 340650.0 442500.0 353250.0 ;
      RECT  448800.0 342750.0 449700.0 353250.0 ;
      RECT  451800.0 340650.0 452700.0 353250.0 ;
      RECT  459000.0 342750.0 459900.0 353250.0 ;
      RECT  462000.0 340650.0 462900.0 353250.0 ;
      RECT  479400.0 342750.0 480300.0 353250.0 ;
      RECT  482400.0 340650.0 483300.0 353250.0 ;
      RECT  489600.0 342750.0 490500.0 353250.0 ;
      RECT  492600.0 340650.0 493500.0 353250.0 ;
      RECT  499800.0 342750.0 500700.0 353250.0 ;
      RECT  502800.0 340650.0 503700.0 353250.0 ;
      RECT  520200.0 342750.0 521100.0 353250.0 ;
      RECT  523200.0 340650.0 524100.0 353250.0 ;
      RECT  530400.0 342750.0 531300.0 353250.0 ;
      RECT  533400.0 340650.0 534300.0 353250.0 ;
      RECT  540600.0 342750.0 541500.0 353250.0 ;
      RECT  543600.0 340650.0 544500.0 353250.0 ;
      RECT  561000.0 342750.0 561900.0 353250.0 ;
      RECT  564000.0 340650.0 564900.0 353250.0 ;
      RECT  571200.0 342750.0 572100.0 353250.0 ;
      RECT  574200.0 340650.0 575100.0 353250.0 ;
      RECT  581400.0 342750.0 582300.0 353250.0 ;
      RECT  584400.0 340650.0 585300.0 353250.0 ;
      RECT  601800.0 342750.0 602700.0 353250.0 ;
      RECT  604800.0 340650.0 605700.0 353250.0 ;
      RECT  612000.0 342750.0 612900.0 353250.0 ;
      RECT  615000.0 340650.0 615900.0 353250.0 ;
      RECT  622200.0 342750.0 623100.0 353250.0 ;
      RECT  625200.0 340650.0 626100.0 353250.0 ;
      RECT  642600.0 342750.0 643500.0 353250.0 ;
      RECT  645600.0 340650.0 646500.0 353250.0 ;
      RECT  652800.0 342750.0 653700.0 353250.0 ;
      RECT  655800.0 340650.0 656700.0 353250.0 ;
      RECT  663000.0 342750.0 663900.0 353250.0 ;
      RECT  666000.0 340650.0 666900.0 353250.0 ;
      RECT  683400.0 342750.0 684300.0 353250.0 ;
      RECT  686400.0 340650.0 687300.0 353250.0 ;
      RECT  693600.0 342750.0 694500.0 353250.0 ;
      RECT  696600.0 340650.0 697500.0 353250.0 ;
      RECT  703800.0 342750.0 704700.0 353250.0 ;
      RECT  706800.0 340650.0 707700.0 353250.0 ;
      RECT  724200.0 342750.0 725100.0 353250.0 ;
      RECT  727200.0 340650.0 728100.0 353250.0 ;
      RECT  734400.0 342750.0 735300.0 353250.0 ;
      RECT  737400.0 340650.0 738300.0 353250.0 ;
      RECT  744600.0 342750.0 745500.0 353250.0 ;
      RECT  747600.0 340650.0 748500.0 353250.0 ;
      RECT  765000.0 342750.0 765900.0 353250.0 ;
      RECT  768000.0 340650.0 768900.0 353250.0 ;
      RECT  775200.0 342750.0 776100.0 353250.0 ;
      RECT  778200.0 340650.0 779100.0 353250.0 ;
      RECT  785400.0 342750.0 786300.0 353250.0 ;
      RECT  788400.0 340650.0 789300.0 353250.0 ;
      RECT  805800.0 342750.0 806700.0 353250.0 ;
      RECT  808800.0 340650.0 809700.0 353250.0 ;
      RECT  816000.0 342750.0 816900.0 353250.0 ;
      RECT  819000.0 340650.0 819900.0 353250.0 ;
      RECT  826200.0 342750.0 827100.0 353250.0 ;
      RECT  829200.0 340650.0 830100.0 353250.0 ;
      RECT  846600.0 342750.0 847500.0 353250.0 ;
      RECT  849600.0 340650.0 850500.0 353250.0 ;
      RECT  856800.0 342750.0 857700.0 353250.0 ;
      RECT  859800.0 340650.0 860700.0 353250.0 ;
      RECT  867000.0 342750.0 867900.0 353250.0 ;
      RECT  870000.0 340650.0 870900.0 353250.0 ;
      RECT  887400.0 342750.0 888300.0 353250.0 ;
      RECT  890400.0 340650.0 891300.0 353250.0 ;
      RECT  897600.0 342750.0 898500.0 353250.0 ;
      RECT  900600.0 340650.0 901500.0 353250.0 ;
      RECT  907800.0 342750.0 908700.0 353250.0 ;
      RECT  910800.0 340650.0 911700.0 353250.0 ;
      RECT  928200.0 342750.0 929100.0 353250.0 ;
      RECT  931200.0 340650.0 932100.0 353250.0 ;
      RECT  938400.0 342750.0 939300.0 353250.0 ;
      RECT  941400.0 340650.0 942300.0 353250.0 ;
      RECT  948600.0 342750.0 949500.0 353250.0 ;
      RECT  951600.0 340650.0 952500.0 353250.0 ;
      RECT  969000.0 342750.0 969900.0 353250.0 ;
      RECT  972000.0 340650.0 972900.0 353250.0 ;
      RECT  979200.0 342750.0 980100.0 353250.0 ;
      RECT  982200.0 340650.0 983100.0 353250.0 ;
      RECT  989400.0 342750.0 990300.0 353250.0 ;
      RECT  992400.0 340650.0 993300.0 353250.0 ;
      RECT  1009800.0 342750.0 1010700.0 353250.0 ;
      RECT  1012800.0 340650.0 1013700.0 353250.0 ;
      RECT  1020000.0 342750.0 1020900.0 353250.0 ;
      RECT  1023000.0 340650.0 1023900.0 353250.0 ;
      RECT  1030200.0 342750.0 1031100.0 353250.0 ;
      RECT  1033200.0 340650.0 1034100.0 353250.0 ;
      RECT  1050600.0 342750.0 1051500.0 353250.0 ;
      RECT  1053600.0 340650.0 1054500.0 353250.0 ;
      RECT  1060800.0 342750.0 1061700.0 353250.0 ;
      RECT  1063800.0 340650.0 1064700.0 353250.0 ;
      RECT  1071000.0 342750.0 1071900.0 353250.0 ;
      RECT  1074000.0 340650.0 1074900.0 353250.0 ;
      RECT  1091400.0 342750.0 1092300.0 353250.0 ;
      RECT  1094400.0 340650.0 1095300.0 353250.0 ;
      RECT  1101600.0 342750.0 1102500.0 353250.0 ;
      RECT  1104600.0 340650.0 1105500.0 353250.0 ;
      RECT  1111800.0 342750.0 1112700.0 353250.0 ;
      RECT  1114800.0 340650.0 1115700.0 353250.0 ;
      RECT  1132200.0 342750.0 1133100.0 353250.0 ;
      RECT  1135200.0 340650.0 1136100.0 353250.0 ;
      RECT  1142400.0 342750.0 1143300.0 353250.0 ;
      RECT  1145400.0 340650.0 1146300.0 353250.0 ;
      RECT  1152600.0 342750.0 1153500.0 353250.0 ;
      RECT  1155600.0 340650.0 1156500.0 353250.0 ;
      RECT  1173000.0 342750.0 1173900.0 353250.0 ;
      RECT  1176000.0 340650.0 1176900.0 353250.0 ;
      RECT  1183200.0 342750.0 1184100.0 353250.0 ;
      RECT  1186200.0 340650.0 1187100.0 353250.0 ;
      RECT  1193400.0 342750.0 1194300.0 353250.0 ;
      RECT  1196400.0 340650.0 1197300.0 353250.0 ;
      RECT  1213800.0 342750.0 1214700.0 353250.0 ;
      RECT  1216800.0 340650.0 1217700.0 353250.0 ;
      RECT  1224000.0 342750.0 1224900.0 353250.0 ;
      RECT  1227000.0 340650.0 1227900.0 353250.0 ;
      RECT  1234200.0 342750.0 1235100.0 353250.0 ;
      RECT  1237200.0 340650.0 1238100.0 353250.0 ;
      RECT  1254600.0 342750.0 1255500.0 353250.0 ;
      RECT  1257600.0 340650.0 1258500.0 353250.0 ;
      RECT  1264800.0 342750.0 1265700.0 353250.0 ;
      RECT  1267800.0 340650.0 1268700.0 353250.0 ;
      RECT  1275000.0 342750.0 1275900.0 353250.0 ;
      RECT  1278000.0 340650.0 1278900.0 353250.0 ;
      RECT  1295400.0 342750.0 1296300.0 353250.0 ;
      RECT  1298400.0 340650.0 1299300.0 353250.0 ;
      RECT  1305600.0 342750.0 1306500.0 353250.0 ;
      RECT  1308600.0 340650.0 1309500.0 353250.0 ;
      RECT  1315800.0 342750.0 1316700.0 353250.0 ;
      RECT  1318800.0 340650.0 1319700.0 353250.0 ;
      RECT  1336200.0 342750.0 1337100.0 353250.0 ;
      RECT  1339200.0 340650.0 1340100.0 353250.0 ;
      RECT  1346400.0 342750.0 1347300.0 353250.0 ;
      RECT  1349400.0 340650.0 1350300.0 353250.0 ;
      RECT  1356600.0 342750.0 1357500.0 353250.0 ;
      RECT  1359600.0 340650.0 1360500.0 353250.0 ;
      RECT  1377000.0 342750.0 1377900.0 353250.0 ;
      RECT  1380000.0 340650.0 1380900.0 353250.0 ;
      RECT  1387200.0 342750.0 1388100.0 353250.0 ;
      RECT  1390200.0 340650.0 1391100.0 353250.0 ;
      RECT  1397400.0 342750.0 1398300.0 353250.0 ;
      RECT  1400400.0 340650.0 1401300.0 353250.0 ;
      RECT  1417800.0 342750.0 1418700.0 353250.0 ;
      RECT  1420800.0 340650.0 1421700.0 353250.0 ;
      RECT  1428000.0 342750.0 1428900.0 353250.0 ;
      RECT  1431000.0 340650.0 1431900.0 353250.0 ;
      RECT  1438200.0 342750.0 1439100.0 353250.0 ;
      RECT  1441200.0 340650.0 1442100.0 353250.0 ;
      RECT  1458600.0 342750.0 1459500.0 353250.0 ;
      RECT  1461600.0 340650.0 1462500.0 353250.0 ;
      RECT  1468800.0 342750.0 1469700.0 353250.0 ;
      RECT  1471800.0 340650.0 1472700.0 353250.0 ;
      RECT  1479000.0 342750.0 1479900.0 353250.0 ;
      RECT  1482000.0 340650.0 1482900.0 353250.0 ;
      RECT  1499400.0 342750.0 1500300.0 353250.0 ;
      RECT  1502400.0 340650.0 1503300.0 353250.0 ;
      RECT  1509600.0 342750.0 1510500.0 353250.0 ;
      RECT  1512600.0 340650.0 1513500.0 353250.0 ;
      RECT  1519800.0 342750.0 1520700.0 353250.0 ;
      RECT  1522800.0 340650.0 1523700.0 353250.0 ;
      RECT  224400.0 361950.0 225300.0 362850.0 ;
      RECT  224850.0 361950.0 225750.0 362850.0 ;
      RECT  224400.0 355050.0 225300.0 362400.0 ;
      RECT  224850.0 361950.0 225300.0 362850.0 ;
      RECT  224850.0 362400.0 225750.0 369750.0 ;
      RECT  227400.0 368250.0 228300.0 369150.0 ;
      RECT  227250.0 368250.0 228150.0 369150.0 ;
      RECT  227400.0 368700.0 228300.0 376950.0 ;
      RECT  227700.0 368250.0 227850.0 369150.0 ;
      RECT  227250.0 360450.0 228150.0 368700.0 ;
      RECT  224250.0 376350.0 225450.0 377550.0 ;
      RECT  227250.0 354450.0 228450.0 355650.0 ;
      RECT  224700.0 369750.0 225900.0 370950.0 ;
      RECT  227100.0 359250.0 228300.0 360450.0 ;
      RECT  231000.0 357450.0 232200.0 358650.0 ;
      RECT  224400.0 376950.0 225300.0 378750.0 ;
      RECT  227400.0 376950.0 228300.0 378750.0 ;
      RECT  224400.0 353250.0 225300.0 355050.0 ;
      RECT  227400.0 353250.0 228300.0 355050.0 ;
      RECT  220800.0 353250.0 221700.0 378750.0 ;
      RECT  231000.0 353250.0 231900.0 378750.0 ;
      RECT  234600.0 361950.0 235500.0 362850.0 ;
      RECT  235050.0 361950.0 235950.0 362850.0 ;
      RECT  234600.0 355050.0 235500.0 362400.0 ;
      RECT  235050.0 361950.0 235500.0 362850.0 ;
      RECT  235050.0 362400.0 235950.0 369750.0 ;
      RECT  237600.0 368250.0 238500.0 369150.0 ;
      RECT  237450.0 368250.0 238350.0 369150.0 ;
      RECT  237600.0 368700.0 238500.0 376950.0 ;
      RECT  237900.0 368250.0 238050.0 369150.0 ;
      RECT  237450.0 360450.0 238350.0 368700.0 ;
      RECT  234450.0 376350.0 235650.0 377550.0 ;
      RECT  237450.0 354450.0 238650.0 355650.0 ;
      RECT  234900.0 369750.0 236100.0 370950.0 ;
      RECT  237300.0 359250.0 238500.0 360450.0 ;
      RECT  241200.0 357450.0 242400.0 358650.0 ;
      RECT  234600.0 376950.0 235500.0 378750.0 ;
      RECT  237600.0 376950.0 238500.0 378750.0 ;
      RECT  234600.0 353250.0 235500.0 355050.0 ;
      RECT  237600.0 353250.0 238500.0 355050.0 ;
      RECT  231000.0 353250.0 231900.0 378750.0 ;
      RECT  241200.0 353250.0 242100.0 378750.0 ;
      RECT  244800.0 361950.0 245700.0 362850.0 ;
      RECT  245250.0 361950.0 246150.0 362850.0 ;
      RECT  244800.0 355050.0 245700.0 362400.0 ;
      RECT  245250.0 361950.0 245700.0 362850.0 ;
      RECT  245250.0 362400.0 246150.0 369750.0 ;
      RECT  247800.0 368250.0 248700.0 369150.0 ;
      RECT  247650.0 368250.0 248550.0 369150.0 ;
      RECT  247800.0 368700.0 248700.0 376950.0 ;
      RECT  248100.0 368250.0 248250.0 369150.0 ;
      RECT  247650.0 360450.0 248550.0 368700.0 ;
      RECT  244650.0 376350.0 245850.0 377550.0 ;
      RECT  247650.0 354450.0 248850.0 355650.0 ;
      RECT  245100.0 369750.0 246300.0 370950.0 ;
      RECT  247500.0 359250.0 248700.0 360450.0 ;
      RECT  251400.0 357450.0 252600.0 358650.0 ;
      RECT  244800.0 376950.0 245700.0 378750.0 ;
      RECT  247800.0 376950.0 248700.0 378750.0 ;
      RECT  244800.0 353250.0 245700.0 355050.0 ;
      RECT  247800.0 353250.0 248700.0 355050.0 ;
      RECT  241200.0 353250.0 242100.0 378750.0 ;
      RECT  251400.0 353250.0 252300.0 378750.0 ;
      RECT  255000.0 361950.0 255900.0 362850.0 ;
      RECT  255450.0 361950.0 256350.0 362850.0 ;
      RECT  255000.0 355050.0 255900.0 362400.0 ;
      RECT  255450.0 361950.0 255900.0 362850.0 ;
      RECT  255450.0 362400.0 256350.0 369750.0 ;
      RECT  258000.0 368250.0 258900.0 369150.0 ;
      RECT  257850.0 368250.0 258750.0 369150.0 ;
      RECT  258000.0 368700.0 258900.0 376950.0 ;
      RECT  258300.0 368250.0 258450.0 369150.0 ;
      RECT  257850.0 360450.0 258750.0 368700.0 ;
      RECT  254850.0 376350.0 256050.0 377550.0 ;
      RECT  257850.0 354450.0 259050.0 355650.0 ;
      RECT  255300.0 369750.0 256500.0 370950.0 ;
      RECT  257700.0 359250.0 258900.0 360450.0 ;
      RECT  261600.0 357450.0 262800.0 358650.0 ;
      RECT  255000.0 376950.0 255900.0 378750.0 ;
      RECT  258000.0 376950.0 258900.0 378750.0 ;
      RECT  255000.0 353250.0 255900.0 355050.0 ;
      RECT  258000.0 353250.0 258900.0 355050.0 ;
      RECT  251400.0 353250.0 252300.0 378750.0 ;
      RECT  261600.0 353250.0 262500.0 378750.0 ;
      RECT  265200.0 361950.0 266100.0 362850.0 ;
      RECT  265650.0 361950.0 266550.0 362850.0 ;
      RECT  265200.0 355050.0 266100.0 362400.0 ;
      RECT  265650.0 361950.0 266100.0 362850.0 ;
      RECT  265650.0 362400.0 266550.0 369750.0 ;
      RECT  268200.0 368250.0 269100.0 369150.0 ;
      RECT  268050.0 368250.0 268950.0 369150.0 ;
      RECT  268200.0 368700.0 269100.0 376950.0 ;
      RECT  268500.0 368250.0 268650.0 369150.0 ;
      RECT  268050.0 360450.0 268950.0 368700.0 ;
      RECT  265050.0 376350.0 266250.0 377550.0 ;
      RECT  268050.0 354450.0 269250.0 355650.0 ;
      RECT  265500.0 369750.0 266700.0 370950.0 ;
      RECT  267900.0 359250.0 269100.0 360450.0 ;
      RECT  271800.0 357450.0 273000.0 358650.0 ;
      RECT  265200.0 376950.0 266100.0 378750.0 ;
      RECT  268200.0 376950.0 269100.0 378750.0 ;
      RECT  265200.0 353250.0 266100.0 355050.0 ;
      RECT  268200.0 353250.0 269100.0 355050.0 ;
      RECT  261600.0 353250.0 262500.0 378750.0 ;
      RECT  271800.0 353250.0 272700.0 378750.0 ;
      RECT  275400.0 361950.0 276300.0 362850.0 ;
      RECT  275850.0 361950.0 276750.0 362850.0 ;
      RECT  275400.0 355050.0 276300.0 362400.0 ;
      RECT  275850.0 361950.0 276300.0 362850.0 ;
      RECT  275850.0 362400.0 276750.0 369750.0 ;
      RECT  278400.0 368250.0 279300.0 369150.0 ;
      RECT  278250.0 368250.0 279150.0 369150.0 ;
      RECT  278400.0 368700.0 279300.0 376950.0 ;
      RECT  278700.0 368250.0 278850.0 369150.0 ;
      RECT  278250.0 360450.0 279150.0 368700.0 ;
      RECT  275250.0 376350.0 276450.0 377550.0 ;
      RECT  278250.0 354450.0 279450.0 355650.0 ;
      RECT  275700.0 369750.0 276900.0 370950.0 ;
      RECT  278100.0 359250.0 279300.0 360450.0 ;
      RECT  282000.0 357450.0 283200.0 358650.0 ;
      RECT  275400.0 376950.0 276300.0 378750.0 ;
      RECT  278400.0 376950.0 279300.0 378750.0 ;
      RECT  275400.0 353250.0 276300.0 355050.0 ;
      RECT  278400.0 353250.0 279300.0 355050.0 ;
      RECT  271800.0 353250.0 272700.0 378750.0 ;
      RECT  282000.0 353250.0 282900.0 378750.0 ;
      RECT  285600.0 361950.0 286500.0 362850.0 ;
      RECT  286050.0 361950.0 286950.0 362850.0 ;
      RECT  285600.0 355050.0 286500.0 362400.0 ;
      RECT  286050.0 361950.0 286500.0 362850.0 ;
      RECT  286050.0 362400.0 286950.0 369750.0 ;
      RECT  288600.0 368250.0 289500.0 369150.0 ;
      RECT  288450.0 368250.0 289350.0 369150.0 ;
      RECT  288600.0 368700.0 289500.0 376950.0 ;
      RECT  288900.0 368250.0 289050.0 369150.0 ;
      RECT  288450.0 360450.0 289350.0 368700.0 ;
      RECT  285450.0 376350.0 286650.0 377550.0 ;
      RECT  288450.0 354450.0 289650.0 355650.0 ;
      RECT  285900.0 369750.0 287100.0 370950.0 ;
      RECT  288300.0 359250.0 289500.0 360450.0 ;
      RECT  292200.0 357450.0 293400.0 358650.0 ;
      RECT  285600.0 376950.0 286500.0 378750.0 ;
      RECT  288600.0 376950.0 289500.0 378750.0 ;
      RECT  285600.0 353250.0 286500.0 355050.0 ;
      RECT  288600.0 353250.0 289500.0 355050.0 ;
      RECT  282000.0 353250.0 282900.0 378750.0 ;
      RECT  292200.0 353250.0 293100.0 378750.0 ;
      RECT  295800.0 361950.0 296700.0 362850.0 ;
      RECT  296250.0 361950.0 297150.0 362850.0 ;
      RECT  295800.0 355050.0 296700.0 362400.0 ;
      RECT  296250.0 361950.0 296700.0 362850.0 ;
      RECT  296250.0 362400.0 297150.0 369750.0 ;
      RECT  298800.0 368250.0 299700.0 369150.0 ;
      RECT  298650.0 368250.0 299550.0 369150.0 ;
      RECT  298800.0 368700.0 299700.0 376950.0 ;
      RECT  299100.0 368250.0 299250.0 369150.0 ;
      RECT  298650.0 360450.0 299550.0 368700.0 ;
      RECT  295650.0 376350.0 296850.0 377550.0 ;
      RECT  298650.0 354450.0 299850.0 355650.0 ;
      RECT  296100.0 369750.0 297300.0 370950.0 ;
      RECT  298500.0 359250.0 299700.0 360450.0 ;
      RECT  302400.0 357450.0 303600.0 358650.0 ;
      RECT  295800.0 376950.0 296700.0 378750.0 ;
      RECT  298800.0 376950.0 299700.0 378750.0 ;
      RECT  295800.0 353250.0 296700.0 355050.0 ;
      RECT  298800.0 353250.0 299700.0 355050.0 ;
      RECT  292200.0 353250.0 293100.0 378750.0 ;
      RECT  302400.0 353250.0 303300.0 378750.0 ;
      RECT  306000.0 361950.0 306900.0 362850.0 ;
      RECT  306450.0 361950.0 307350.0 362850.0 ;
      RECT  306000.0 355050.0 306900.0 362400.0 ;
      RECT  306450.0 361950.0 306900.0 362850.0 ;
      RECT  306450.0 362400.0 307350.0 369750.0 ;
      RECT  309000.0 368250.0 309900.0 369150.0 ;
      RECT  308850.0 368250.0 309750.0 369150.0 ;
      RECT  309000.0 368700.0 309900.0 376950.0 ;
      RECT  309300.0 368250.0 309450.0 369150.0 ;
      RECT  308850.0 360450.0 309750.0 368700.0 ;
      RECT  305850.0 376350.0 307050.0 377550.0 ;
      RECT  308850.0 354450.0 310050.0 355650.0 ;
      RECT  306300.0 369750.0 307500.0 370950.0 ;
      RECT  308700.0 359250.0 309900.0 360450.0 ;
      RECT  312600.0 357450.0 313800.0 358650.0 ;
      RECT  306000.0 376950.0 306900.0 378750.0 ;
      RECT  309000.0 376950.0 309900.0 378750.0 ;
      RECT  306000.0 353250.0 306900.0 355050.0 ;
      RECT  309000.0 353250.0 309900.0 355050.0 ;
      RECT  302400.0 353250.0 303300.0 378750.0 ;
      RECT  312600.0 353250.0 313500.0 378750.0 ;
      RECT  316200.0 361950.0 317100.0 362850.0 ;
      RECT  316650.0 361950.0 317550.0 362850.0 ;
      RECT  316200.0 355050.0 317100.0 362400.0 ;
      RECT  316650.0 361950.0 317100.0 362850.0 ;
      RECT  316650.0 362400.0 317550.0 369750.0 ;
      RECT  319200.0 368250.0 320100.0 369150.0 ;
      RECT  319050.0 368250.0 319950.0 369150.0 ;
      RECT  319200.0 368700.0 320100.0 376950.0 ;
      RECT  319500.0 368250.0 319650.0 369150.0 ;
      RECT  319050.0 360450.0 319950.0 368700.0 ;
      RECT  316050.0 376350.0 317250.0 377550.0 ;
      RECT  319050.0 354450.0 320250.0 355650.0 ;
      RECT  316500.0 369750.0 317700.0 370950.0 ;
      RECT  318900.0 359250.0 320100.0 360450.0 ;
      RECT  322800.0 357450.0 324000.0 358650.0 ;
      RECT  316200.0 376950.0 317100.0 378750.0 ;
      RECT  319200.0 376950.0 320100.0 378750.0 ;
      RECT  316200.0 353250.0 317100.0 355050.0 ;
      RECT  319200.0 353250.0 320100.0 355050.0 ;
      RECT  312600.0 353250.0 313500.0 378750.0 ;
      RECT  322800.0 353250.0 323700.0 378750.0 ;
      RECT  326400.0 361950.0 327300.0 362850.0 ;
      RECT  326850.0 361950.0 327750.0 362850.0 ;
      RECT  326400.0 355050.0 327300.0 362400.0 ;
      RECT  326850.0 361950.0 327300.0 362850.0 ;
      RECT  326850.0 362400.0 327750.0 369750.0 ;
      RECT  329400.0 368250.0 330300.0 369150.0 ;
      RECT  329250.0 368250.0 330150.0 369150.0 ;
      RECT  329400.0 368700.0 330300.0 376950.0 ;
      RECT  329700.0 368250.0 329850.0 369150.0 ;
      RECT  329250.0 360450.0 330150.0 368700.0 ;
      RECT  326250.0 376350.0 327450.0 377550.0 ;
      RECT  329250.0 354450.0 330450.0 355650.0 ;
      RECT  326700.0 369750.0 327900.0 370950.0 ;
      RECT  329100.0 359250.0 330300.0 360450.0 ;
      RECT  333000.0 357450.0 334200.0 358650.0 ;
      RECT  326400.0 376950.0 327300.0 378750.0 ;
      RECT  329400.0 376950.0 330300.0 378750.0 ;
      RECT  326400.0 353250.0 327300.0 355050.0 ;
      RECT  329400.0 353250.0 330300.0 355050.0 ;
      RECT  322800.0 353250.0 323700.0 378750.0 ;
      RECT  333000.0 353250.0 333900.0 378750.0 ;
      RECT  336600.0 361950.0 337500.0 362850.0 ;
      RECT  337050.0 361950.0 337950.0 362850.0 ;
      RECT  336600.0 355050.0 337500.0 362400.0 ;
      RECT  337050.0 361950.0 337500.0 362850.0 ;
      RECT  337050.0 362400.0 337950.0 369750.0 ;
      RECT  339600.0 368250.0 340500.0 369150.0 ;
      RECT  339450.0 368250.0 340350.0 369150.0 ;
      RECT  339600.0 368700.0 340500.0 376950.0 ;
      RECT  339900.0 368250.0 340050.0 369150.0 ;
      RECT  339450.0 360450.0 340350.0 368700.0 ;
      RECT  336450.0 376350.0 337650.0 377550.0 ;
      RECT  339450.0 354450.0 340650.0 355650.0 ;
      RECT  336900.0 369750.0 338100.0 370950.0 ;
      RECT  339300.0 359250.0 340500.0 360450.0 ;
      RECT  343200.0 357450.0 344400.0 358650.0 ;
      RECT  336600.0 376950.0 337500.0 378750.0 ;
      RECT  339600.0 376950.0 340500.0 378750.0 ;
      RECT  336600.0 353250.0 337500.0 355050.0 ;
      RECT  339600.0 353250.0 340500.0 355050.0 ;
      RECT  333000.0 353250.0 333900.0 378750.0 ;
      RECT  343200.0 353250.0 344100.0 378750.0 ;
      RECT  346800.0 361950.0 347700.0 362850.0 ;
      RECT  347250.0 361950.0 348150.0 362850.0 ;
      RECT  346800.0 355050.0 347700.0 362400.0 ;
      RECT  347250.0 361950.0 347700.0 362850.0 ;
      RECT  347250.0 362400.0 348150.0 369750.0 ;
      RECT  349800.0 368250.0 350700.0 369150.0 ;
      RECT  349650.0 368250.0 350550.0 369150.0 ;
      RECT  349800.0 368700.0 350700.0 376950.0 ;
      RECT  350100.0 368250.0 350250.0 369150.0 ;
      RECT  349650.0 360450.0 350550.0 368700.0 ;
      RECT  346650.0 376350.0 347850.0 377550.0 ;
      RECT  349650.0 354450.0 350850.0 355650.0 ;
      RECT  347100.0 369750.0 348300.0 370950.0 ;
      RECT  349500.0 359250.0 350700.0 360450.0 ;
      RECT  353400.0 357450.0 354600.0 358650.0 ;
      RECT  346800.0 376950.0 347700.0 378750.0 ;
      RECT  349800.0 376950.0 350700.0 378750.0 ;
      RECT  346800.0 353250.0 347700.0 355050.0 ;
      RECT  349800.0 353250.0 350700.0 355050.0 ;
      RECT  343200.0 353250.0 344100.0 378750.0 ;
      RECT  353400.0 353250.0 354300.0 378750.0 ;
      RECT  357000.0 361950.0 357900.0 362850.0 ;
      RECT  357450.0 361950.0 358350.0 362850.0 ;
      RECT  357000.0 355050.0 357900.0 362400.0 ;
      RECT  357450.0 361950.0 357900.0 362850.0 ;
      RECT  357450.0 362400.0 358350.0 369750.0 ;
      RECT  360000.0 368250.0 360900.0 369150.0 ;
      RECT  359850.0 368250.0 360750.0 369150.0 ;
      RECT  360000.0 368700.0 360900.0 376950.0 ;
      RECT  360300.0 368250.0 360450.0 369150.0 ;
      RECT  359850.0 360450.0 360750.0 368700.0 ;
      RECT  356850.0 376350.0 358050.0 377550.0 ;
      RECT  359850.0 354450.0 361050.0 355650.0 ;
      RECT  357300.0 369750.0 358500.0 370950.0 ;
      RECT  359700.0 359250.0 360900.0 360450.0 ;
      RECT  363600.0 357450.0 364800.0 358650.0 ;
      RECT  357000.0 376950.0 357900.0 378750.0 ;
      RECT  360000.0 376950.0 360900.0 378750.0 ;
      RECT  357000.0 353250.0 357900.0 355050.0 ;
      RECT  360000.0 353250.0 360900.0 355050.0 ;
      RECT  353400.0 353250.0 354300.0 378750.0 ;
      RECT  363600.0 353250.0 364500.0 378750.0 ;
      RECT  367200.0 361950.0 368100.0 362850.0 ;
      RECT  367650.0 361950.0 368550.0 362850.0 ;
      RECT  367200.0 355050.0 368100.0 362400.0 ;
      RECT  367650.0 361950.0 368100.0 362850.0 ;
      RECT  367650.0 362400.0 368550.0 369750.0 ;
      RECT  370200.0 368250.0 371100.0 369150.0 ;
      RECT  370050.0 368250.0 370950.0 369150.0 ;
      RECT  370200.0 368700.0 371100.0 376950.0 ;
      RECT  370500.0 368250.0 370650.0 369150.0 ;
      RECT  370050.0 360450.0 370950.0 368700.0 ;
      RECT  367050.0 376350.0 368250.0 377550.0 ;
      RECT  370050.0 354450.0 371250.0 355650.0 ;
      RECT  367500.0 369750.0 368700.0 370950.0 ;
      RECT  369900.0 359250.0 371100.0 360450.0 ;
      RECT  373800.0 357450.0 375000.0 358650.0 ;
      RECT  367200.0 376950.0 368100.0 378750.0 ;
      RECT  370200.0 376950.0 371100.0 378750.0 ;
      RECT  367200.0 353250.0 368100.0 355050.0 ;
      RECT  370200.0 353250.0 371100.0 355050.0 ;
      RECT  363600.0 353250.0 364500.0 378750.0 ;
      RECT  373800.0 353250.0 374700.0 378750.0 ;
      RECT  377400.0 361950.0 378300.0 362850.0 ;
      RECT  377850.0 361950.0 378750.0 362850.0 ;
      RECT  377400.0 355050.0 378300.0 362400.0 ;
      RECT  377850.0 361950.0 378300.0 362850.0 ;
      RECT  377850.0 362400.0 378750.0 369750.0 ;
      RECT  380400.0 368250.0 381300.0 369150.0 ;
      RECT  380250.0 368250.0 381150.0 369150.0 ;
      RECT  380400.0 368700.0 381300.0 376950.0 ;
      RECT  380700.0 368250.0 380850.0 369150.0 ;
      RECT  380250.0 360450.0 381150.0 368700.0 ;
      RECT  377250.0 376350.0 378450.0 377550.0 ;
      RECT  380250.0 354450.0 381450.0 355650.0 ;
      RECT  377700.0 369750.0 378900.0 370950.0 ;
      RECT  380100.0 359250.0 381300.0 360450.0 ;
      RECT  384000.0 357450.0 385200.0 358650.0 ;
      RECT  377400.0 376950.0 378300.0 378750.0 ;
      RECT  380400.0 376950.0 381300.0 378750.0 ;
      RECT  377400.0 353250.0 378300.0 355050.0 ;
      RECT  380400.0 353250.0 381300.0 355050.0 ;
      RECT  373800.0 353250.0 374700.0 378750.0 ;
      RECT  384000.0 353250.0 384900.0 378750.0 ;
      RECT  387600.0 361950.0 388500.0 362850.0 ;
      RECT  388050.0 361950.0 388950.0 362850.0 ;
      RECT  387600.0 355050.0 388500.0 362400.0 ;
      RECT  388050.0 361950.0 388500.0 362850.0 ;
      RECT  388050.0 362400.0 388950.0 369750.0 ;
      RECT  390600.0 368250.0 391500.0 369150.0 ;
      RECT  390450.0 368250.0 391350.0 369150.0 ;
      RECT  390600.0 368700.0 391500.0 376950.0 ;
      RECT  390900.0 368250.0 391050.0 369150.0 ;
      RECT  390450.0 360450.0 391350.0 368700.0 ;
      RECT  387450.0 376350.0 388650.0 377550.0 ;
      RECT  390450.0 354450.0 391650.0 355650.0 ;
      RECT  387900.0 369750.0 389100.0 370950.0 ;
      RECT  390300.0 359250.0 391500.0 360450.0 ;
      RECT  394200.0 357450.0 395400.0 358650.0 ;
      RECT  387600.0 376950.0 388500.0 378750.0 ;
      RECT  390600.0 376950.0 391500.0 378750.0 ;
      RECT  387600.0 353250.0 388500.0 355050.0 ;
      RECT  390600.0 353250.0 391500.0 355050.0 ;
      RECT  384000.0 353250.0 384900.0 378750.0 ;
      RECT  394200.0 353250.0 395100.0 378750.0 ;
      RECT  397800.0 361950.0 398700.0 362850.0 ;
      RECT  398250.0 361950.0 399150.0 362850.0 ;
      RECT  397800.0 355050.0 398700.0 362400.0 ;
      RECT  398250.0 361950.0 398700.0 362850.0 ;
      RECT  398250.0 362400.0 399150.0 369750.0 ;
      RECT  400800.0 368250.0 401700.0 369150.0 ;
      RECT  400650.0 368250.0 401550.0 369150.0 ;
      RECT  400800.0 368700.0 401700.0 376950.0 ;
      RECT  401100.0 368250.0 401250.0 369150.0 ;
      RECT  400650.0 360450.0 401550.0 368700.0 ;
      RECT  397650.0 376350.0 398850.0 377550.0 ;
      RECT  400650.0 354450.0 401850.0 355650.0 ;
      RECT  398100.0 369750.0 399300.0 370950.0 ;
      RECT  400500.0 359250.0 401700.0 360450.0 ;
      RECT  404400.0 357450.0 405600.0 358650.0 ;
      RECT  397800.0 376950.0 398700.0 378750.0 ;
      RECT  400800.0 376950.0 401700.0 378750.0 ;
      RECT  397800.0 353250.0 398700.0 355050.0 ;
      RECT  400800.0 353250.0 401700.0 355050.0 ;
      RECT  394200.0 353250.0 395100.0 378750.0 ;
      RECT  404400.0 353250.0 405300.0 378750.0 ;
      RECT  408000.0 361950.0 408900.0 362850.0 ;
      RECT  408450.0 361950.0 409350.0 362850.0 ;
      RECT  408000.0 355050.0 408900.0 362400.0 ;
      RECT  408450.0 361950.0 408900.0 362850.0 ;
      RECT  408450.0 362400.0 409350.0 369750.0 ;
      RECT  411000.0 368250.0 411900.0 369150.0 ;
      RECT  410850.0 368250.0 411750.0 369150.0 ;
      RECT  411000.0 368700.0 411900.0 376950.0 ;
      RECT  411300.0 368250.0 411450.0 369150.0 ;
      RECT  410850.0 360450.0 411750.0 368700.0 ;
      RECT  407850.0 376350.0 409050.0 377550.0 ;
      RECT  410850.0 354450.0 412050.0 355650.0 ;
      RECT  408300.0 369750.0 409500.0 370950.0 ;
      RECT  410700.0 359250.0 411900.0 360450.0 ;
      RECT  414600.0 357450.0 415800.0 358650.0 ;
      RECT  408000.0 376950.0 408900.0 378750.0 ;
      RECT  411000.0 376950.0 411900.0 378750.0 ;
      RECT  408000.0 353250.0 408900.0 355050.0 ;
      RECT  411000.0 353250.0 411900.0 355050.0 ;
      RECT  404400.0 353250.0 405300.0 378750.0 ;
      RECT  414600.0 353250.0 415500.0 378750.0 ;
      RECT  418200.0 361950.0 419100.0 362850.0 ;
      RECT  418650.0 361950.0 419550.0 362850.0 ;
      RECT  418200.0 355050.0 419100.0 362400.0 ;
      RECT  418650.0 361950.0 419100.0 362850.0 ;
      RECT  418650.0 362400.0 419550.0 369750.0 ;
      RECT  421200.0 368250.0 422100.0 369150.0 ;
      RECT  421050.0 368250.0 421950.0 369150.0 ;
      RECT  421200.0 368700.0 422100.0 376950.0 ;
      RECT  421500.0 368250.0 421650.0 369150.0 ;
      RECT  421050.0 360450.0 421950.0 368700.0 ;
      RECT  418050.0 376350.0 419250.0 377550.0 ;
      RECT  421050.0 354450.0 422250.0 355650.0 ;
      RECT  418500.0 369750.0 419700.0 370950.0 ;
      RECT  420900.0 359250.0 422100.0 360450.0 ;
      RECT  424800.0 357450.0 426000.0 358650.0 ;
      RECT  418200.0 376950.0 419100.0 378750.0 ;
      RECT  421200.0 376950.0 422100.0 378750.0 ;
      RECT  418200.0 353250.0 419100.0 355050.0 ;
      RECT  421200.0 353250.0 422100.0 355050.0 ;
      RECT  414600.0 353250.0 415500.0 378750.0 ;
      RECT  424800.0 353250.0 425700.0 378750.0 ;
      RECT  428400.0 361950.0 429300.0 362850.0 ;
      RECT  428850.0 361950.0 429750.0 362850.0 ;
      RECT  428400.0 355050.0 429300.0 362400.0 ;
      RECT  428850.0 361950.0 429300.0 362850.0 ;
      RECT  428850.0 362400.0 429750.0 369750.0 ;
      RECT  431400.0 368250.0 432300.0 369150.0 ;
      RECT  431250.0 368250.0 432150.0 369150.0 ;
      RECT  431400.0 368700.0 432300.0 376950.0 ;
      RECT  431700.0 368250.0 431850.0 369150.0 ;
      RECT  431250.0 360450.0 432150.0 368700.0 ;
      RECT  428250.0 376350.0 429450.0 377550.0 ;
      RECT  431250.0 354450.0 432450.0 355650.0 ;
      RECT  428700.0 369750.0 429900.0 370950.0 ;
      RECT  431100.0 359250.0 432300.0 360450.0 ;
      RECT  435000.0 357450.0 436200.0 358650.0 ;
      RECT  428400.0 376950.0 429300.0 378750.0 ;
      RECT  431400.0 376950.0 432300.0 378750.0 ;
      RECT  428400.0 353250.0 429300.0 355050.0 ;
      RECT  431400.0 353250.0 432300.0 355050.0 ;
      RECT  424800.0 353250.0 425700.0 378750.0 ;
      RECT  435000.0 353250.0 435900.0 378750.0 ;
      RECT  438600.0 361950.0 439500.0 362850.0 ;
      RECT  439050.0 361950.0 439950.0 362850.0 ;
      RECT  438600.0 355050.0 439500.0 362400.0 ;
      RECT  439050.0 361950.0 439500.0 362850.0 ;
      RECT  439050.0 362400.0 439950.0 369750.0 ;
      RECT  441600.0 368250.0 442500.0 369150.0 ;
      RECT  441450.0 368250.0 442350.0 369150.0 ;
      RECT  441600.0 368700.0 442500.0 376950.0 ;
      RECT  441900.0 368250.0 442050.0 369150.0 ;
      RECT  441450.0 360450.0 442350.0 368700.0 ;
      RECT  438450.0 376350.0 439650.0 377550.0 ;
      RECT  441450.0 354450.0 442650.0 355650.0 ;
      RECT  438900.0 369750.0 440100.0 370950.0 ;
      RECT  441300.0 359250.0 442500.0 360450.0 ;
      RECT  445200.0 357450.0 446400.0 358650.0 ;
      RECT  438600.0 376950.0 439500.0 378750.0 ;
      RECT  441600.0 376950.0 442500.0 378750.0 ;
      RECT  438600.0 353250.0 439500.0 355050.0 ;
      RECT  441600.0 353250.0 442500.0 355050.0 ;
      RECT  435000.0 353250.0 435900.0 378750.0 ;
      RECT  445200.0 353250.0 446100.0 378750.0 ;
      RECT  448800.0 361950.0 449700.0 362850.0 ;
      RECT  449250.0 361950.0 450150.0 362850.0 ;
      RECT  448800.0 355050.0 449700.0 362400.0 ;
      RECT  449250.0 361950.0 449700.0 362850.0 ;
      RECT  449250.0 362400.0 450150.0 369750.0 ;
      RECT  451800.0 368250.0 452700.0 369150.0 ;
      RECT  451650.0 368250.0 452550.0 369150.0 ;
      RECT  451800.0 368700.0 452700.0 376950.0 ;
      RECT  452100.0 368250.0 452250.0 369150.0 ;
      RECT  451650.0 360450.0 452550.0 368700.0 ;
      RECT  448650.0 376350.0 449850.0 377550.0 ;
      RECT  451650.0 354450.0 452850.0 355650.0 ;
      RECT  449100.0 369750.0 450300.0 370950.0 ;
      RECT  451500.0 359250.0 452700.0 360450.0 ;
      RECT  455400.0 357450.0 456600.0 358650.0 ;
      RECT  448800.0 376950.0 449700.0 378750.0 ;
      RECT  451800.0 376950.0 452700.0 378750.0 ;
      RECT  448800.0 353250.0 449700.0 355050.0 ;
      RECT  451800.0 353250.0 452700.0 355050.0 ;
      RECT  445200.0 353250.0 446100.0 378750.0 ;
      RECT  455400.0 353250.0 456300.0 378750.0 ;
      RECT  459000.0 361950.0 459900.0 362850.0 ;
      RECT  459450.0 361950.0 460350.0 362850.0 ;
      RECT  459000.0 355050.0 459900.0 362400.0 ;
      RECT  459450.0 361950.0 459900.0 362850.0 ;
      RECT  459450.0 362400.0 460350.0 369750.0 ;
      RECT  462000.0 368250.0 462900.0 369150.0 ;
      RECT  461850.0 368250.0 462750.0 369150.0 ;
      RECT  462000.0 368700.0 462900.0 376950.0 ;
      RECT  462300.0 368250.0 462450.0 369150.0 ;
      RECT  461850.0 360450.0 462750.0 368700.0 ;
      RECT  458850.0 376350.0 460050.0 377550.0 ;
      RECT  461850.0 354450.0 463050.0 355650.0 ;
      RECT  459300.0 369750.0 460500.0 370950.0 ;
      RECT  461700.0 359250.0 462900.0 360450.0 ;
      RECT  465600.0 357450.0 466800.0 358650.0 ;
      RECT  459000.0 376950.0 459900.0 378750.0 ;
      RECT  462000.0 376950.0 462900.0 378750.0 ;
      RECT  459000.0 353250.0 459900.0 355050.0 ;
      RECT  462000.0 353250.0 462900.0 355050.0 ;
      RECT  455400.0 353250.0 456300.0 378750.0 ;
      RECT  465600.0 353250.0 466500.0 378750.0 ;
      RECT  469200.0 361950.0 470100.0 362850.0 ;
      RECT  469650.0 361950.0 470550.0 362850.0 ;
      RECT  469200.0 355050.0 470100.0 362400.0 ;
      RECT  469650.0 361950.0 470100.0 362850.0 ;
      RECT  469650.0 362400.0 470550.0 369750.0 ;
      RECT  472200.0 368250.0 473100.0 369150.0 ;
      RECT  472050.0 368250.0 472950.0 369150.0 ;
      RECT  472200.0 368700.0 473100.0 376950.0 ;
      RECT  472500.0 368250.0 472650.0 369150.0 ;
      RECT  472050.0 360450.0 472950.0 368700.0 ;
      RECT  469050.0 376350.0 470250.0 377550.0 ;
      RECT  472050.0 354450.0 473250.0 355650.0 ;
      RECT  469500.0 369750.0 470700.0 370950.0 ;
      RECT  471900.0 359250.0 473100.0 360450.0 ;
      RECT  475800.0 357450.0 477000.0 358650.0 ;
      RECT  469200.0 376950.0 470100.0 378750.0 ;
      RECT  472200.0 376950.0 473100.0 378750.0 ;
      RECT  469200.0 353250.0 470100.0 355050.0 ;
      RECT  472200.0 353250.0 473100.0 355050.0 ;
      RECT  465600.0 353250.0 466500.0 378750.0 ;
      RECT  475800.0 353250.0 476700.0 378750.0 ;
      RECT  479400.0 361950.0 480300.0 362850.0 ;
      RECT  479850.0 361950.0 480750.0 362850.0 ;
      RECT  479400.0 355050.0 480300.0 362400.0 ;
      RECT  479850.0 361950.0 480300.0 362850.0 ;
      RECT  479850.0 362400.0 480750.0 369750.0 ;
      RECT  482400.0 368250.0 483300.0 369150.0 ;
      RECT  482250.0 368250.0 483150.0 369150.0 ;
      RECT  482400.0 368700.0 483300.0 376950.0 ;
      RECT  482700.0 368250.0 482850.0 369150.0 ;
      RECT  482250.0 360450.0 483150.0 368700.0 ;
      RECT  479250.0 376350.0 480450.0 377550.0 ;
      RECT  482250.0 354450.0 483450.0 355650.0 ;
      RECT  479700.0 369750.0 480900.0 370950.0 ;
      RECT  482100.0 359250.0 483300.0 360450.0 ;
      RECT  486000.0 357450.0 487200.0 358650.0 ;
      RECT  479400.0 376950.0 480300.0 378750.0 ;
      RECT  482400.0 376950.0 483300.0 378750.0 ;
      RECT  479400.0 353250.0 480300.0 355050.0 ;
      RECT  482400.0 353250.0 483300.0 355050.0 ;
      RECT  475800.0 353250.0 476700.0 378750.0 ;
      RECT  486000.0 353250.0 486900.0 378750.0 ;
      RECT  489600.0 361950.0 490500.0 362850.0 ;
      RECT  490050.0 361950.0 490950.0 362850.0 ;
      RECT  489600.0 355050.0 490500.0 362400.0 ;
      RECT  490050.0 361950.0 490500.0 362850.0 ;
      RECT  490050.0 362400.0 490950.0 369750.0 ;
      RECT  492600.0 368250.0 493500.0 369150.0 ;
      RECT  492450.0 368250.0 493350.0 369150.0 ;
      RECT  492600.0 368700.0 493500.0 376950.0 ;
      RECT  492900.0 368250.0 493050.0 369150.0 ;
      RECT  492450.0 360450.0 493350.0 368700.0 ;
      RECT  489450.0 376350.0 490650.0 377550.0 ;
      RECT  492450.0 354450.0 493650.0 355650.0 ;
      RECT  489900.0 369750.0 491100.0 370950.0 ;
      RECT  492300.0 359250.0 493500.0 360450.0 ;
      RECT  496200.0 357450.0 497400.0 358650.0 ;
      RECT  489600.0 376950.0 490500.0 378750.0 ;
      RECT  492600.0 376950.0 493500.0 378750.0 ;
      RECT  489600.0 353250.0 490500.0 355050.0 ;
      RECT  492600.0 353250.0 493500.0 355050.0 ;
      RECT  486000.0 353250.0 486900.0 378750.0 ;
      RECT  496200.0 353250.0 497100.0 378750.0 ;
      RECT  499800.0 361950.0 500700.0 362850.0 ;
      RECT  500250.0 361950.0 501150.0 362850.0 ;
      RECT  499800.0 355050.0 500700.0 362400.0 ;
      RECT  500250.0 361950.0 500700.0 362850.0 ;
      RECT  500250.0 362400.0 501150.0 369750.0 ;
      RECT  502800.0 368250.0 503700.0 369150.0 ;
      RECT  502650.0 368250.0 503550.0 369150.0 ;
      RECT  502800.0 368700.0 503700.0 376950.0 ;
      RECT  503100.0 368250.0 503250.0 369150.0 ;
      RECT  502650.0 360450.0 503550.0 368700.0 ;
      RECT  499650.0 376350.0 500850.0 377550.0 ;
      RECT  502650.0 354450.0 503850.0 355650.0 ;
      RECT  500100.0 369750.0 501300.0 370950.0 ;
      RECT  502500.0 359250.0 503700.0 360450.0 ;
      RECT  506400.0 357450.0 507600.0 358650.0 ;
      RECT  499800.0 376950.0 500700.0 378750.0 ;
      RECT  502800.0 376950.0 503700.0 378750.0 ;
      RECT  499800.0 353250.0 500700.0 355050.0 ;
      RECT  502800.0 353250.0 503700.0 355050.0 ;
      RECT  496200.0 353250.0 497100.0 378750.0 ;
      RECT  506400.0 353250.0 507300.0 378750.0 ;
      RECT  510000.0 361950.0 510900.0 362850.0 ;
      RECT  510450.0 361950.0 511350.0 362850.0 ;
      RECT  510000.0 355050.0 510900.0 362400.0 ;
      RECT  510450.0 361950.0 510900.0 362850.0 ;
      RECT  510450.0 362400.0 511350.0 369750.0 ;
      RECT  513000.0 368250.0 513900.0 369150.0 ;
      RECT  512850.0 368250.0 513750.0 369150.0 ;
      RECT  513000.0 368700.0 513900.0 376950.0 ;
      RECT  513300.0 368250.0 513450.0 369150.0 ;
      RECT  512850.0 360450.0 513750.0 368700.0 ;
      RECT  509850.0 376350.0 511050.0 377550.0 ;
      RECT  512850.0 354450.0 514050.0 355650.0 ;
      RECT  510300.0 369750.0 511500.0 370950.0 ;
      RECT  512700.0 359250.0 513900.0 360450.0 ;
      RECT  516600.0 357450.0 517800.0 358650.0 ;
      RECT  510000.0 376950.0 510900.0 378750.0 ;
      RECT  513000.0 376950.0 513900.0 378750.0 ;
      RECT  510000.0 353250.0 510900.0 355050.0 ;
      RECT  513000.0 353250.0 513900.0 355050.0 ;
      RECT  506400.0 353250.0 507300.0 378750.0 ;
      RECT  516600.0 353250.0 517500.0 378750.0 ;
      RECT  520200.0 361950.0 521100.0 362850.0 ;
      RECT  520650.0 361950.0 521550.0 362850.0 ;
      RECT  520200.0 355050.0 521100.0 362400.0 ;
      RECT  520650.0 361950.0 521100.0 362850.0 ;
      RECT  520650.0 362400.0 521550.0 369750.0 ;
      RECT  523200.0 368250.0 524100.0 369150.0 ;
      RECT  523050.0 368250.0 523950.0 369150.0 ;
      RECT  523200.0 368700.0 524100.0 376950.0 ;
      RECT  523500.0 368250.0 523650.0 369150.0 ;
      RECT  523050.0 360450.0 523950.0 368700.0 ;
      RECT  520050.0 376350.0 521250.0 377550.0 ;
      RECT  523050.0 354450.0 524250.0 355650.0 ;
      RECT  520500.0 369750.0 521700.0 370950.0 ;
      RECT  522900.0 359250.0 524100.0 360450.0 ;
      RECT  526800.0 357450.0 528000.0 358650.0 ;
      RECT  520200.0 376950.0 521100.0 378750.0 ;
      RECT  523200.0 376950.0 524100.0 378750.0 ;
      RECT  520200.0 353250.0 521100.0 355050.0 ;
      RECT  523200.0 353250.0 524100.0 355050.0 ;
      RECT  516600.0 353250.0 517500.0 378750.0 ;
      RECT  526800.0 353250.0 527700.0 378750.0 ;
      RECT  530400.0 361950.0 531300.0 362850.0 ;
      RECT  530850.0 361950.0 531750.0 362850.0 ;
      RECT  530400.0 355050.0 531300.0 362400.0 ;
      RECT  530850.0 361950.0 531300.0 362850.0 ;
      RECT  530850.0 362400.0 531750.0 369750.0 ;
      RECT  533400.0 368250.0 534300.0 369150.0 ;
      RECT  533250.0 368250.0 534150.0 369150.0 ;
      RECT  533400.0 368700.0 534300.0 376950.0 ;
      RECT  533700.0 368250.0 533850.0 369150.0 ;
      RECT  533250.0 360450.0 534150.0 368700.0 ;
      RECT  530250.0 376350.0 531450.0 377550.0 ;
      RECT  533250.0 354450.0 534450.0 355650.0 ;
      RECT  530700.0 369750.0 531900.0 370950.0 ;
      RECT  533100.0 359250.0 534300.0 360450.0 ;
      RECT  537000.0 357450.0 538200.0 358650.0 ;
      RECT  530400.0 376950.0 531300.0 378750.0 ;
      RECT  533400.0 376950.0 534300.0 378750.0 ;
      RECT  530400.0 353250.0 531300.0 355050.0 ;
      RECT  533400.0 353250.0 534300.0 355050.0 ;
      RECT  526800.0 353250.0 527700.0 378750.0 ;
      RECT  537000.0 353250.0 537900.0 378750.0 ;
      RECT  540600.0 361950.0 541500.0 362850.0 ;
      RECT  541050.0 361950.0 541950.0 362850.0 ;
      RECT  540600.0 355050.0 541500.0 362400.0 ;
      RECT  541050.0 361950.0 541500.0 362850.0 ;
      RECT  541050.0 362400.0 541950.0 369750.0 ;
      RECT  543600.0 368250.0 544500.0 369150.0 ;
      RECT  543450.0 368250.0 544350.0 369150.0 ;
      RECT  543600.0 368700.0 544500.0 376950.0 ;
      RECT  543900.0 368250.0 544050.0 369150.0 ;
      RECT  543450.0 360450.0 544350.0 368700.0 ;
      RECT  540450.0 376350.0 541650.0 377550.0 ;
      RECT  543450.0 354450.0 544650.0 355650.0 ;
      RECT  540900.0 369750.0 542100.0 370950.0 ;
      RECT  543300.0 359250.0 544500.0 360450.0 ;
      RECT  547200.0 357450.0 548400.0 358650.0 ;
      RECT  540600.0 376950.0 541500.0 378750.0 ;
      RECT  543600.0 376950.0 544500.0 378750.0 ;
      RECT  540600.0 353250.0 541500.0 355050.0 ;
      RECT  543600.0 353250.0 544500.0 355050.0 ;
      RECT  537000.0 353250.0 537900.0 378750.0 ;
      RECT  547200.0 353250.0 548100.0 378750.0 ;
      RECT  550800.0 361950.0 551700.0 362850.0 ;
      RECT  551250.0 361950.0 552150.0 362850.0 ;
      RECT  550800.0 355050.0 551700.0 362400.0 ;
      RECT  551250.0 361950.0 551700.0 362850.0 ;
      RECT  551250.0 362400.0 552150.0 369750.0 ;
      RECT  553800.0 368250.0 554700.0 369150.0 ;
      RECT  553650.0 368250.0 554550.0 369150.0 ;
      RECT  553800.0 368700.0 554700.0 376950.0 ;
      RECT  554100.0 368250.0 554250.0 369150.0 ;
      RECT  553650.0 360450.0 554550.0 368700.0 ;
      RECT  550650.0 376350.0 551850.0 377550.0 ;
      RECT  553650.0 354450.0 554850.0 355650.0 ;
      RECT  551100.0 369750.0 552300.0 370950.0 ;
      RECT  553500.0 359250.0 554700.0 360450.0 ;
      RECT  557400.0 357450.0 558600.0 358650.0 ;
      RECT  550800.0 376950.0 551700.0 378750.0 ;
      RECT  553800.0 376950.0 554700.0 378750.0 ;
      RECT  550800.0 353250.0 551700.0 355050.0 ;
      RECT  553800.0 353250.0 554700.0 355050.0 ;
      RECT  547200.0 353250.0 548100.0 378750.0 ;
      RECT  557400.0 353250.0 558300.0 378750.0 ;
      RECT  561000.0 361950.0 561900.0 362850.0 ;
      RECT  561450.0 361950.0 562350.0 362850.0 ;
      RECT  561000.0 355050.0 561900.0 362400.0 ;
      RECT  561450.0 361950.0 561900.0 362850.0 ;
      RECT  561450.0 362400.0 562350.0 369750.0 ;
      RECT  564000.0 368250.0 564900.0 369150.0 ;
      RECT  563850.0 368250.0 564750.0 369150.0 ;
      RECT  564000.0 368700.0 564900.0 376950.0 ;
      RECT  564300.0 368250.0 564450.0 369150.0 ;
      RECT  563850.0 360450.0 564750.0 368700.0 ;
      RECT  560850.0 376350.0 562050.0 377550.0 ;
      RECT  563850.0 354450.0 565050.0 355650.0 ;
      RECT  561300.0 369750.0 562500.0 370950.0 ;
      RECT  563700.0 359250.0 564900.0 360450.0 ;
      RECT  567600.0 357450.0 568800.0 358650.0 ;
      RECT  561000.0 376950.0 561900.0 378750.0 ;
      RECT  564000.0 376950.0 564900.0 378750.0 ;
      RECT  561000.0 353250.0 561900.0 355050.0 ;
      RECT  564000.0 353250.0 564900.0 355050.0 ;
      RECT  557400.0 353250.0 558300.0 378750.0 ;
      RECT  567600.0 353250.0 568500.0 378750.0 ;
      RECT  571200.0 361950.0 572100.0 362850.0 ;
      RECT  571650.0 361950.0 572550.0 362850.0 ;
      RECT  571200.0 355050.0 572100.0 362400.0 ;
      RECT  571650.0 361950.0 572100.0 362850.0 ;
      RECT  571650.0 362400.0 572550.0 369750.0 ;
      RECT  574200.0 368250.0 575100.0 369150.0 ;
      RECT  574050.0 368250.0 574950.0 369150.0 ;
      RECT  574200.0 368700.0 575100.0 376950.0 ;
      RECT  574500.0 368250.0 574650.0 369150.0 ;
      RECT  574050.0 360450.0 574950.0 368700.0 ;
      RECT  571050.0 376350.0 572250.0 377550.0 ;
      RECT  574050.0 354450.0 575250.0 355650.0 ;
      RECT  571500.0 369750.0 572700.0 370950.0 ;
      RECT  573900.0 359250.0 575100.0 360450.0 ;
      RECT  577800.0 357450.0 579000.0 358650.0 ;
      RECT  571200.0 376950.0 572100.0 378750.0 ;
      RECT  574200.0 376950.0 575100.0 378750.0 ;
      RECT  571200.0 353250.0 572100.0 355050.0 ;
      RECT  574200.0 353250.0 575100.0 355050.0 ;
      RECT  567600.0 353250.0 568500.0 378750.0 ;
      RECT  577800.0 353250.0 578700.0 378750.0 ;
      RECT  581400.0 361950.0 582300.0 362850.0 ;
      RECT  581850.0 361950.0 582750.0 362850.0 ;
      RECT  581400.0 355050.0 582300.0 362400.0 ;
      RECT  581850.0 361950.0 582300.0 362850.0 ;
      RECT  581850.0 362400.0 582750.0 369750.0 ;
      RECT  584400.0 368250.0 585300.0 369150.0 ;
      RECT  584250.0 368250.0 585150.0 369150.0 ;
      RECT  584400.0 368700.0 585300.0 376950.0 ;
      RECT  584700.0 368250.0 584850.0 369150.0 ;
      RECT  584250.0 360450.0 585150.0 368700.0 ;
      RECT  581250.0 376350.0 582450.0 377550.0 ;
      RECT  584250.0 354450.0 585450.0 355650.0 ;
      RECT  581700.0 369750.0 582900.0 370950.0 ;
      RECT  584100.0 359250.0 585300.0 360450.0 ;
      RECT  588000.0 357450.0 589200.0 358650.0 ;
      RECT  581400.0 376950.0 582300.0 378750.0 ;
      RECT  584400.0 376950.0 585300.0 378750.0 ;
      RECT  581400.0 353250.0 582300.0 355050.0 ;
      RECT  584400.0 353250.0 585300.0 355050.0 ;
      RECT  577800.0 353250.0 578700.0 378750.0 ;
      RECT  588000.0 353250.0 588900.0 378750.0 ;
      RECT  591600.0 361950.0 592500.0 362850.0 ;
      RECT  592050.0 361950.0 592950.0 362850.0 ;
      RECT  591600.0 355050.0 592500.0 362400.0 ;
      RECT  592050.0 361950.0 592500.0 362850.0 ;
      RECT  592050.0 362400.0 592950.0 369750.0 ;
      RECT  594600.0 368250.0 595500.0 369150.0 ;
      RECT  594450.0 368250.0 595350.0 369150.0 ;
      RECT  594600.0 368700.0 595500.0 376950.0 ;
      RECT  594900.0 368250.0 595050.0 369150.0 ;
      RECT  594450.0 360450.0 595350.0 368700.0 ;
      RECT  591450.0 376350.0 592650.0 377550.0 ;
      RECT  594450.0 354450.0 595650.0 355650.0 ;
      RECT  591900.0 369750.0 593100.0 370950.0 ;
      RECT  594300.0 359250.0 595500.0 360450.0 ;
      RECT  598200.0 357450.0 599400.0 358650.0 ;
      RECT  591600.0 376950.0 592500.0 378750.0 ;
      RECT  594600.0 376950.0 595500.0 378750.0 ;
      RECT  591600.0 353250.0 592500.0 355050.0 ;
      RECT  594600.0 353250.0 595500.0 355050.0 ;
      RECT  588000.0 353250.0 588900.0 378750.0 ;
      RECT  598200.0 353250.0 599100.0 378750.0 ;
      RECT  601800.0 361950.0 602700.0 362850.0 ;
      RECT  602250.0 361950.0 603150.0 362850.0 ;
      RECT  601800.0 355050.0 602700.0 362400.0 ;
      RECT  602250.0 361950.0 602700.0 362850.0 ;
      RECT  602250.0 362400.0 603150.0 369750.0 ;
      RECT  604800.0 368250.0 605700.0 369150.0 ;
      RECT  604650.0 368250.0 605550.0 369150.0 ;
      RECT  604800.0 368700.0 605700.0 376950.0 ;
      RECT  605100.0 368250.0 605250.0 369150.0 ;
      RECT  604650.0 360450.0 605550.0 368700.0 ;
      RECT  601650.0 376350.0 602850.0 377550.0 ;
      RECT  604650.0 354450.0 605850.0 355650.0 ;
      RECT  602100.0 369750.0 603300.0 370950.0 ;
      RECT  604500.0 359250.0 605700.0 360450.0 ;
      RECT  608400.0 357450.0 609600.0 358650.0 ;
      RECT  601800.0 376950.0 602700.0 378750.0 ;
      RECT  604800.0 376950.0 605700.0 378750.0 ;
      RECT  601800.0 353250.0 602700.0 355050.0 ;
      RECT  604800.0 353250.0 605700.0 355050.0 ;
      RECT  598200.0 353250.0 599100.0 378750.0 ;
      RECT  608400.0 353250.0 609300.0 378750.0 ;
      RECT  612000.0 361950.0 612900.0 362850.0 ;
      RECT  612450.0 361950.0 613350.0 362850.0 ;
      RECT  612000.0 355050.0 612900.0 362400.0 ;
      RECT  612450.0 361950.0 612900.0 362850.0 ;
      RECT  612450.0 362400.0 613350.0 369750.0 ;
      RECT  615000.0 368250.0 615900.0 369150.0 ;
      RECT  614850.0 368250.0 615750.0 369150.0 ;
      RECT  615000.0 368700.0 615900.0 376950.0 ;
      RECT  615300.0 368250.0 615450.0 369150.0 ;
      RECT  614850.0 360450.0 615750.0 368700.0 ;
      RECT  611850.0 376350.0 613050.0 377550.0 ;
      RECT  614850.0 354450.0 616050.0 355650.0 ;
      RECT  612300.0 369750.0 613500.0 370950.0 ;
      RECT  614700.0 359250.0 615900.0 360450.0 ;
      RECT  618600.0 357450.0 619800.0 358650.0 ;
      RECT  612000.0 376950.0 612900.0 378750.0 ;
      RECT  615000.0 376950.0 615900.0 378750.0 ;
      RECT  612000.0 353250.0 612900.0 355050.0 ;
      RECT  615000.0 353250.0 615900.0 355050.0 ;
      RECT  608400.0 353250.0 609300.0 378750.0 ;
      RECT  618600.0 353250.0 619500.0 378750.0 ;
      RECT  622200.0 361950.0 623100.0 362850.0 ;
      RECT  622650.0 361950.0 623550.0 362850.0 ;
      RECT  622200.0 355050.0 623100.0 362400.0 ;
      RECT  622650.0 361950.0 623100.0 362850.0 ;
      RECT  622650.0 362400.0 623550.0 369750.0 ;
      RECT  625200.0 368250.0 626100.0 369150.0 ;
      RECT  625050.0 368250.0 625950.0 369150.0 ;
      RECT  625200.0 368700.0 626100.0 376950.0 ;
      RECT  625500.0 368250.0 625650.0 369150.0 ;
      RECT  625050.0 360450.0 625950.0 368700.0 ;
      RECT  622050.0 376350.0 623250.0 377550.0 ;
      RECT  625050.0 354450.0 626250.0 355650.0 ;
      RECT  622500.0 369750.0 623700.0 370950.0 ;
      RECT  624900.0 359250.0 626100.0 360450.0 ;
      RECT  628800.0 357450.0 630000.0 358650.0 ;
      RECT  622200.0 376950.0 623100.0 378750.0 ;
      RECT  625200.0 376950.0 626100.0 378750.0 ;
      RECT  622200.0 353250.0 623100.0 355050.0 ;
      RECT  625200.0 353250.0 626100.0 355050.0 ;
      RECT  618600.0 353250.0 619500.0 378750.0 ;
      RECT  628800.0 353250.0 629700.0 378750.0 ;
      RECT  632400.0 361950.0 633300.0 362850.0 ;
      RECT  632850.0 361950.0 633750.0 362850.0 ;
      RECT  632400.0 355050.0 633300.0 362400.0 ;
      RECT  632850.0 361950.0 633300.0 362850.0 ;
      RECT  632850.0 362400.0 633750.0 369750.0 ;
      RECT  635400.0 368250.0 636300.0 369150.0 ;
      RECT  635250.0 368250.0 636150.0 369150.0 ;
      RECT  635400.0 368700.0 636300.0 376950.0 ;
      RECT  635700.0 368250.0 635850.0 369150.0 ;
      RECT  635250.0 360450.0 636150.0 368700.0 ;
      RECT  632250.0 376350.0 633450.0 377550.0 ;
      RECT  635250.0 354450.0 636450.0 355650.0 ;
      RECT  632700.0 369750.0 633900.0 370950.0 ;
      RECT  635100.0 359250.0 636300.0 360450.0 ;
      RECT  639000.0 357450.0 640200.0 358650.0 ;
      RECT  632400.0 376950.0 633300.0 378750.0 ;
      RECT  635400.0 376950.0 636300.0 378750.0 ;
      RECT  632400.0 353250.0 633300.0 355050.0 ;
      RECT  635400.0 353250.0 636300.0 355050.0 ;
      RECT  628800.0 353250.0 629700.0 378750.0 ;
      RECT  639000.0 353250.0 639900.0 378750.0 ;
      RECT  642600.0 361950.0 643500.0 362850.0 ;
      RECT  643050.0 361950.0 643950.0 362850.0 ;
      RECT  642600.0 355050.0 643500.0 362400.0 ;
      RECT  643050.0 361950.0 643500.0 362850.0 ;
      RECT  643050.0 362400.0 643950.0 369750.0 ;
      RECT  645600.0 368250.0 646500.0 369150.0 ;
      RECT  645450.0 368250.0 646350.0 369150.0 ;
      RECT  645600.0 368700.0 646500.0 376950.0 ;
      RECT  645900.0 368250.0 646050.0 369150.0 ;
      RECT  645450.0 360450.0 646350.0 368700.0 ;
      RECT  642450.0 376350.0 643650.0 377550.0 ;
      RECT  645450.0 354450.0 646650.0 355650.0 ;
      RECT  642900.0 369750.0 644100.0 370950.0 ;
      RECT  645300.0 359250.0 646500.0 360450.0 ;
      RECT  649200.0 357450.0 650400.0 358650.0 ;
      RECT  642600.0 376950.0 643500.0 378750.0 ;
      RECT  645600.0 376950.0 646500.0 378750.0 ;
      RECT  642600.0 353250.0 643500.0 355050.0 ;
      RECT  645600.0 353250.0 646500.0 355050.0 ;
      RECT  639000.0 353250.0 639900.0 378750.0 ;
      RECT  649200.0 353250.0 650100.0 378750.0 ;
      RECT  652800.0 361950.0 653700.0 362850.0 ;
      RECT  653250.0 361950.0 654150.0 362850.0 ;
      RECT  652800.0 355050.0 653700.0 362400.0 ;
      RECT  653250.0 361950.0 653700.0 362850.0 ;
      RECT  653250.0 362400.0 654150.0 369750.0 ;
      RECT  655800.0 368250.0 656700.0 369150.0 ;
      RECT  655650.0 368250.0 656550.0 369150.0 ;
      RECT  655800.0 368700.0 656700.0 376950.0 ;
      RECT  656100.0 368250.0 656250.0 369150.0 ;
      RECT  655650.0 360450.0 656550.0 368700.0 ;
      RECT  652650.0 376350.0 653850.0 377550.0 ;
      RECT  655650.0 354450.0 656850.0 355650.0 ;
      RECT  653100.0 369750.0 654300.0 370950.0 ;
      RECT  655500.0 359250.0 656700.0 360450.0 ;
      RECT  659400.0 357450.0 660600.0 358650.0 ;
      RECT  652800.0 376950.0 653700.0 378750.0 ;
      RECT  655800.0 376950.0 656700.0 378750.0 ;
      RECT  652800.0 353250.0 653700.0 355050.0 ;
      RECT  655800.0 353250.0 656700.0 355050.0 ;
      RECT  649200.0 353250.0 650100.0 378750.0 ;
      RECT  659400.0 353250.0 660300.0 378750.0 ;
      RECT  663000.0 361950.0 663900.0 362850.0 ;
      RECT  663450.0 361950.0 664350.0 362850.0 ;
      RECT  663000.0 355050.0 663900.0 362400.0 ;
      RECT  663450.0 361950.0 663900.0 362850.0 ;
      RECT  663450.0 362400.0 664350.0 369750.0 ;
      RECT  666000.0 368250.0 666900.0 369150.0 ;
      RECT  665850.0 368250.0 666750.0 369150.0 ;
      RECT  666000.0 368700.0 666900.0 376950.0 ;
      RECT  666300.0 368250.0 666450.0 369150.0 ;
      RECT  665850.0 360450.0 666750.0 368700.0 ;
      RECT  662850.0 376350.0 664050.0 377550.0 ;
      RECT  665850.0 354450.0 667050.0 355650.0 ;
      RECT  663300.0 369750.0 664500.0 370950.0 ;
      RECT  665700.0 359250.0 666900.0 360450.0 ;
      RECT  669600.0 357450.0 670800.0 358650.0 ;
      RECT  663000.0 376950.0 663900.0 378750.0 ;
      RECT  666000.0 376950.0 666900.0 378750.0 ;
      RECT  663000.0 353250.0 663900.0 355050.0 ;
      RECT  666000.0 353250.0 666900.0 355050.0 ;
      RECT  659400.0 353250.0 660300.0 378750.0 ;
      RECT  669600.0 353250.0 670500.0 378750.0 ;
      RECT  673200.0 361950.0 674100.0 362850.0 ;
      RECT  673650.0 361950.0 674550.0 362850.0 ;
      RECT  673200.0 355050.0 674100.0 362400.0 ;
      RECT  673650.0 361950.0 674100.0 362850.0 ;
      RECT  673650.0 362400.0 674550.0 369750.0 ;
      RECT  676200.0 368250.0 677100.0 369150.0 ;
      RECT  676050.0 368250.0 676950.0 369150.0 ;
      RECT  676200.0 368700.0 677100.0 376950.0 ;
      RECT  676500.0 368250.0 676650.0 369150.0 ;
      RECT  676050.0 360450.0 676950.0 368700.0 ;
      RECT  673050.0 376350.0 674250.0 377550.0 ;
      RECT  676050.0 354450.0 677250.0 355650.0 ;
      RECT  673500.0 369750.0 674700.0 370950.0 ;
      RECT  675900.0 359250.0 677100.0 360450.0 ;
      RECT  679800.0 357450.0 681000.0 358650.0 ;
      RECT  673200.0 376950.0 674100.0 378750.0 ;
      RECT  676200.0 376950.0 677100.0 378750.0 ;
      RECT  673200.0 353250.0 674100.0 355050.0 ;
      RECT  676200.0 353250.0 677100.0 355050.0 ;
      RECT  669600.0 353250.0 670500.0 378750.0 ;
      RECT  679800.0 353250.0 680700.0 378750.0 ;
      RECT  683400.0 361950.0 684300.0 362850.0 ;
      RECT  683850.0 361950.0 684750.0 362850.0 ;
      RECT  683400.0 355050.0 684300.0 362400.0 ;
      RECT  683850.0 361950.0 684300.0 362850.0 ;
      RECT  683850.0 362400.0 684750.0 369750.0 ;
      RECT  686400.0 368250.0 687300.0 369150.0 ;
      RECT  686250.0 368250.0 687150.0 369150.0 ;
      RECT  686400.0 368700.0 687300.0 376950.0 ;
      RECT  686700.0 368250.0 686850.0 369150.0 ;
      RECT  686250.0 360450.0 687150.0 368700.0 ;
      RECT  683250.0 376350.0 684450.0 377550.0 ;
      RECT  686250.0 354450.0 687450.0 355650.0 ;
      RECT  683700.0 369750.0 684900.0 370950.0 ;
      RECT  686100.0 359250.0 687300.0 360450.0 ;
      RECT  690000.0 357450.0 691200.0 358650.0 ;
      RECT  683400.0 376950.0 684300.0 378750.0 ;
      RECT  686400.0 376950.0 687300.0 378750.0 ;
      RECT  683400.0 353250.0 684300.0 355050.0 ;
      RECT  686400.0 353250.0 687300.0 355050.0 ;
      RECT  679800.0 353250.0 680700.0 378750.0 ;
      RECT  690000.0 353250.0 690900.0 378750.0 ;
      RECT  693600.0 361950.0 694500.0 362850.0 ;
      RECT  694050.0 361950.0 694950.0 362850.0 ;
      RECT  693600.0 355050.0 694500.0 362400.0 ;
      RECT  694050.0 361950.0 694500.0 362850.0 ;
      RECT  694050.0 362400.0 694950.0 369750.0 ;
      RECT  696600.0 368250.0 697500.0 369150.0 ;
      RECT  696450.0 368250.0 697350.0 369150.0 ;
      RECT  696600.0 368700.0 697500.0 376950.0 ;
      RECT  696900.0 368250.0 697050.0 369150.0 ;
      RECT  696450.0 360450.0 697350.0 368700.0 ;
      RECT  693450.0 376350.0 694650.0 377550.0 ;
      RECT  696450.0 354450.0 697650.0 355650.0 ;
      RECT  693900.0 369750.0 695100.0 370950.0 ;
      RECT  696300.0 359250.0 697500.0 360450.0 ;
      RECT  700200.0 357450.0 701400.0 358650.0 ;
      RECT  693600.0 376950.0 694500.0 378750.0 ;
      RECT  696600.0 376950.0 697500.0 378750.0 ;
      RECT  693600.0 353250.0 694500.0 355050.0 ;
      RECT  696600.0 353250.0 697500.0 355050.0 ;
      RECT  690000.0 353250.0 690900.0 378750.0 ;
      RECT  700200.0 353250.0 701100.0 378750.0 ;
      RECT  703800.0 361950.0 704700.0 362850.0 ;
      RECT  704250.0 361950.0 705150.0 362850.0 ;
      RECT  703800.0 355050.0 704700.0 362400.0 ;
      RECT  704250.0 361950.0 704700.0 362850.0 ;
      RECT  704250.0 362400.0 705150.0 369750.0 ;
      RECT  706800.0 368250.0 707700.0 369150.0 ;
      RECT  706650.0 368250.0 707550.0 369150.0 ;
      RECT  706800.0 368700.0 707700.0 376950.0 ;
      RECT  707100.0 368250.0 707250.0 369150.0 ;
      RECT  706650.0 360450.0 707550.0 368700.0 ;
      RECT  703650.0 376350.0 704850.0 377550.0 ;
      RECT  706650.0 354450.0 707850.0 355650.0 ;
      RECT  704100.0 369750.0 705300.0 370950.0 ;
      RECT  706500.0 359250.0 707700.0 360450.0 ;
      RECT  710400.0 357450.0 711600.0 358650.0 ;
      RECT  703800.0 376950.0 704700.0 378750.0 ;
      RECT  706800.0 376950.0 707700.0 378750.0 ;
      RECT  703800.0 353250.0 704700.0 355050.0 ;
      RECT  706800.0 353250.0 707700.0 355050.0 ;
      RECT  700200.0 353250.0 701100.0 378750.0 ;
      RECT  710400.0 353250.0 711300.0 378750.0 ;
      RECT  714000.0 361950.0 714900.0 362850.0 ;
      RECT  714450.0 361950.0 715350.0 362850.0 ;
      RECT  714000.0 355050.0 714900.0 362400.0 ;
      RECT  714450.0 361950.0 714900.0 362850.0 ;
      RECT  714450.0 362400.0 715350.0 369750.0 ;
      RECT  717000.0 368250.0 717900.0 369150.0 ;
      RECT  716850.0 368250.0 717750.0 369150.0 ;
      RECT  717000.0 368700.0 717900.0 376950.0 ;
      RECT  717300.0 368250.0 717450.0 369150.0 ;
      RECT  716850.0 360450.0 717750.0 368700.0 ;
      RECT  713850.0 376350.0 715050.0 377550.0 ;
      RECT  716850.0 354450.0 718050.0 355650.0 ;
      RECT  714300.0 369750.0 715500.0 370950.0 ;
      RECT  716700.0 359250.0 717900.0 360450.0 ;
      RECT  720600.0 357450.0 721800.0 358650.0 ;
      RECT  714000.0 376950.0 714900.0 378750.0 ;
      RECT  717000.0 376950.0 717900.0 378750.0 ;
      RECT  714000.0 353250.0 714900.0 355050.0 ;
      RECT  717000.0 353250.0 717900.0 355050.0 ;
      RECT  710400.0 353250.0 711300.0 378750.0 ;
      RECT  720600.0 353250.0 721500.0 378750.0 ;
      RECT  724200.0 361950.0 725100.0 362850.0 ;
      RECT  724650.0 361950.0 725550.0 362850.0 ;
      RECT  724200.0 355050.0 725100.0 362400.0 ;
      RECT  724650.0 361950.0 725100.0 362850.0 ;
      RECT  724650.0 362400.0 725550.0 369750.0 ;
      RECT  727200.0 368250.0 728100.0 369150.0 ;
      RECT  727050.0 368250.0 727950.0 369150.0 ;
      RECT  727200.0 368700.0 728100.0 376950.0 ;
      RECT  727500.0 368250.0 727650.0 369150.0 ;
      RECT  727050.0 360450.0 727950.0 368700.0 ;
      RECT  724050.0 376350.0 725250.0 377550.0 ;
      RECT  727050.0 354450.0 728250.0 355650.0 ;
      RECT  724500.0 369750.0 725700.0 370950.0 ;
      RECT  726900.0 359250.0 728100.0 360450.0 ;
      RECT  730800.0 357450.0 732000.0 358650.0 ;
      RECT  724200.0 376950.0 725100.0 378750.0 ;
      RECT  727200.0 376950.0 728100.0 378750.0 ;
      RECT  724200.0 353250.0 725100.0 355050.0 ;
      RECT  727200.0 353250.0 728100.0 355050.0 ;
      RECT  720600.0 353250.0 721500.0 378750.0 ;
      RECT  730800.0 353250.0 731700.0 378750.0 ;
      RECT  734400.0 361950.0 735300.0 362850.0 ;
      RECT  734850.0 361950.0 735750.0 362850.0 ;
      RECT  734400.0 355050.0 735300.0 362400.0 ;
      RECT  734850.0 361950.0 735300.0 362850.0 ;
      RECT  734850.0 362400.0 735750.0 369750.0 ;
      RECT  737400.0 368250.0 738300.0 369150.0 ;
      RECT  737250.0 368250.0 738150.0 369150.0 ;
      RECT  737400.0 368700.0 738300.0 376950.0 ;
      RECT  737700.0 368250.0 737850.0 369150.0 ;
      RECT  737250.0 360450.0 738150.0 368700.0 ;
      RECT  734250.0 376350.0 735450.0 377550.0 ;
      RECT  737250.0 354450.0 738450.0 355650.0 ;
      RECT  734700.0 369750.0 735900.0 370950.0 ;
      RECT  737100.0 359250.0 738300.0 360450.0 ;
      RECT  741000.0 357450.0 742200.0 358650.0 ;
      RECT  734400.0 376950.0 735300.0 378750.0 ;
      RECT  737400.0 376950.0 738300.0 378750.0 ;
      RECT  734400.0 353250.0 735300.0 355050.0 ;
      RECT  737400.0 353250.0 738300.0 355050.0 ;
      RECT  730800.0 353250.0 731700.0 378750.0 ;
      RECT  741000.0 353250.0 741900.0 378750.0 ;
      RECT  744600.0 361950.0 745500.0 362850.0 ;
      RECT  745050.0 361950.0 745950.0 362850.0 ;
      RECT  744600.0 355050.0 745500.0 362400.0 ;
      RECT  745050.0 361950.0 745500.0 362850.0 ;
      RECT  745050.0 362400.0 745950.0 369750.0 ;
      RECT  747600.0 368250.0 748500.0 369150.0 ;
      RECT  747450.0 368250.0 748350.0 369150.0 ;
      RECT  747600.0 368700.0 748500.0 376950.0 ;
      RECT  747900.0 368250.0 748050.0 369150.0 ;
      RECT  747450.0 360450.0 748350.0 368700.0 ;
      RECT  744450.0 376350.0 745650.0 377550.0 ;
      RECT  747450.0 354450.0 748650.0 355650.0 ;
      RECT  744900.0 369750.0 746100.0 370950.0 ;
      RECT  747300.0 359250.0 748500.0 360450.0 ;
      RECT  751200.0 357450.0 752400.0 358650.0 ;
      RECT  744600.0 376950.0 745500.0 378750.0 ;
      RECT  747600.0 376950.0 748500.0 378750.0 ;
      RECT  744600.0 353250.0 745500.0 355050.0 ;
      RECT  747600.0 353250.0 748500.0 355050.0 ;
      RECT  741000.0 353250.0 741900.0 378750.0 ;
      RECT  751200.0 353250.0 752100.0 378750.0 ;
      RECT  754800.0 361950.0 755700.0 362850.0 ;
      RECT  755250.0 361950.0 756150.0 362850.0 ;
      RECT  754800.0 355050.0 755700.0 362400.0 ;
      RECT  755250.0 361950.0 755700.0 362850.0 ;
      RECT  755250.0 362400.0 756150.0 369750.0 ;
      RECT  757800.0 368250.0 758700.0 369150.0 ;
      RECT  757650.0 368250.0 758550.0 369150.0 ;
      RECT  757800.0 368700.0 758700.0 376950.0 ;
      RECT  758100.0 368250.0 758250.0 369150.0 ;
      RECT  757650.0 360450.0 758550.0 368700.0 ;
      RECT  754650.0 376350.0 755850.0 377550.0 ;
      RECT  757650.0 354450.0 758850.0 355650.0 ;
      RECT  755100.0 369750.0 756300.0 370950.0 ;
      RECT  757500.0 359250.0 758700.0 360450.0 ;
      RECT  761400.0 357450.0 762600.0 358650.0 ;
      RECT  754800.0 376950.0 755700.0 378750.0 ;
      RECT  757800.0 376950.0 758700.0 378750.0 ;
      RECT  754800.0 353250.0 755700.0 355050.0 ;
      RECT  757800.0 353250.0 758700.0 355050.0 ;
      RECT  751200.0 353250.0 752100.0 378750.0 ;
      RECT  761400.0 353250.0 762300.0 378750.0 ;
      RECT  765000.0 361950.0 765900.0 362850.0 ;
      RECT  765450.0 361950.0 766350.0 362850.0 ;
      RECT  765000.0 355050.0 765900.0 362400.0 ;
      RECT  765450.0 361950.0 765900.0 362850.0 ;
      RECT  765450.0 362400.0 766350.0 369750.0 ;
      RECT  768000.0 368250.0 768900.0 369150.0 ;
      RECT  767850.0 368250.0 768750.0 369150.0 ;
      RECT  768000.0 368700.0 768900.0 376950.0 ;
      RECT  768300.0 368250.0 768450.0 369150.0 ;
      RECT  767850.0 360450.0 768750.0 368700.0 ;
      RECT  764850.0 376350.0 766050.0 377550.0 ;
      RECT  767850.0 354450.0 769050.0 355650.0 ;
      RECT  765300.0 369750.0 766500.0 370950.0 ;
      RECT  767700.0 359250.0 768900.0 360450.0 ;
      RECT  771600.0 357450.0 772800.0 358650.0 ;
      RECT  765000.0 376950.0 765900.0 378750.0 ;
      RECT  768000.0 376950.0 768900.0 378750.0 ;
      RECT  765000.0 353250.0 765900.0 355050.0 ;
      RECT  768000.0 353250.0 768900.0 355050.0 ;
      RECT  761400.0 353250.0 762300.0 378750.0 ;
      RECT  771600.0 353250.0 772500.0 378750.0 ;
      RECT  775200.0 361950.0 776100.0 362850.0 ;
      RECT  775650.0 361950.0 776550.0 362850.0 ;
      RECT  775200.0 355050.0 776100.0 362400.0 ;
      RECT  775650.0 361950.0 776100.0 362850.0 ;
      RECT  775650.0 362400.0 776550.0 369750.0 ;
      RECT  778200.0 368250.0 779100.0 369150.0 ;
      RECT  778050.0 368250.0 778950.0 369150.0 ;
      RECT  778200.0 368700.0 779100.0 376950.0 ;
      RECT  778500.0 368250.0 778650.0 369150.0 ;
      RECT  778050.0 360450.0 778950.0 368700.0 ;
      RECT  775050.0 376350.0 776250.0 377550.0 ;
      RECT  778050.0 354450.0 779250.0 355650.0 ;
      RECT  775500.0 369750.0 776700.0 370950.0 ;
      RECT  777900.0 359250.0 779100.0 360450.0 ;
      RECT  781800.0 357450.0 783000.0 358650.0 ;
      RECT  775200.0 376950.0 776100.0 378750.0 ;
      RECT  778200.0 376950.0 779100.0 378750.0 ;
      RECT  775200.0 353250.0 776100.0 355050.0 ;
      RECT  778200.0 353250.0 779100.0 355050.0 ;
      RECT  771600.0 353250.0 772500.0 378750.0 ;
      RECT  781800.0 353250.0 782700.0 378750.0 ;
      RECT  785400.0 361950.0 786300.0 362850.0 ;
      RECT  785850.0 361950.0 786750.0 362850.0 ;
      RECT  785400.0 355050.0 786300.0 362400.0 ;
      RECT  785850.0 361950.0 786300.0 362850.0 ;
      RECT  785850.0 362400.0 786750.0 369750.0 ;
      RECT  788400.0 368250.0 789300.0 369150.0 ;
      RECT  788250.0 368250.0 789150.0 369150.0 ;
      RECT  788400.0 368700.0 789300.0 376950.0 ;
      RECT  788700.0 368250.0 788850.0 369150.0 ;
      RECT  788250.0 360450.0 789150.0 368700.0 ;
      RECT  785250.0 376350.0 786450.0 377550.0 ;
      RECT  788250.0 354450.0 789450.0 355650.0 ;
      RECT  785700.0 369750.0 786900.0 370950.0 ;
      RECT  788100.0 359250.0 789300.0 360450.0 ;
      RECT  792000.0 357450.0 793200.0 358650.0 ;
      RECT  785400.0 376950.0 786300.0 378750.0 ;
      RECT  788400.0 376950.0 789300.0 378750.0 ;
      RECT  785400.0 353250.0 786300.0 355050.0 ;
      RECT  788400.0 353250.0 789300.0 355050.0 ;
      RECT  781800.0 353250.0 782700.0 378750.0 ;
      RECT  792000.0 353250.0 792900.0 378750.0 ;
      RECT  795600.0 361950.0 796500.0 362850.0 ;
      RECT  796050.0 361950.0 796950.0 362850.0 ;
      RECT  795600.0 355050.0 796500.0 362400.0 ;
      RECT  796050.0 361950.0 796500.0 362850.0 ;
      RECT  796050.0 362400.0 796950.0 369750.0 ;
      RECT  798600.0 368250.0 799500.0 369150.0 ;
      RECT  798450.0 368250.0 799350.0 369150.0 ;
      RECT  798600.0 368700.0 799500.0 376950.0 ;
      RECT  798900.0 368250.0 799050.0 369150.0 ;
      RECT  798450.0 360450.0 799350.0 368700.0 ;
      RECT  795450.0 376350.0 796650.0 377550.0 ;
      RECT  798450.0 354450.0 799650.0 355650.0 ;
      RECT  795900.0 369750.0 797100.0 370950.0 ;
      RECT  798300.0 359250.0 799500.0 360450.0 ;
      RECT  802200.0 357450.0 803400.0 358650.0 ;
      RECT  795600.0 376950.0 796500.0 378750.0 ;
      RECT  798600.0 376950.0 799500.0 378750.0 ;
      RECT  795600.0 353250.0 796500.0 355050.0 ;
      RECT  798600.0 353250.0 799500.0 355050.0 ;
      RECT  792000.0 353250.0 792900.0 378750.0 ;
      RECT  802200.0 353250.0 803100.0 378750.0 ;
      RECT  805800.0 361950.0 806700.0 362850.0 ;
      RECT  806250.0 361950.0 807150.0 362850.0 ;
      RECT  805800.0 355050.0 806700.0 362400.0 ;
      RECT  806250.0 361950.0 806700.0 362850.0 ;
      RECT  806250.0 362400.0 807150.0 369750.0 ;
      RECT  808800.0 368250.0 809700.0 369150.0 ;
      RECT  808650.0 368250.0 809550.0 369150.0 ;
      RECT  808800.0 368700.0 809700.0 376950.0 ;
      RECT  809100.0 368250.0 809250.0 369150.0 ;
      RECT  808650.0 360450.0 809550.0 368700.0 ;
      RECT  805650.0 376350.0 806850.0 377550.0 ;
      RECT  808650.0 354450.0 809850.0 355650.0 ;
      RECT  806100.0 369750.0 807300.0 370950.0 ;
      RECT  808500.0 359250.0 809700.0 360450.0 ;
      RECT  812400.0 357450.0 813600.0 358650.0 ;
      RECT  805800.0 376950.0 806700.0 378750.0 ;
      RECT  808800.0 376950.0 809700.0 378750.0 ;
      RECT  805800.0 353250.0 806700.0 355050.0 ;
      RECT  808800.0 353250.0 809700.0 355050.0 ;
      RECT  802200.0 353250.0 803100.0 378750.0 ;
      RECT  812400.0 353250.0 813300.0 378750.0 ;
      RECT  816000.0 361950.0 816900.0 362850.0 ;
      RECT  816450.0 361950.0 817350.0 362850.0 ;
      RECT  816000.0 355050.0 816900.0 362400.0 ;
      RECT  816450.0 361950.0 816900.0 362850.0 ;
      RECT  816450.0 362400.0 817350.0 369750.0 ;
      RECT  819000.0 368250.0 819900.0 369150.0 ;
      RECT  818850.0 368250.0 819750.0 369150.0 ;
      RECT  819000.0 368700.0 819900.0 376950.0 ;
      RECT  819300.0 368250.0 819450.0 369150.0 ;
      RECT  818850.0 360450.0 819750.0 368700.0 ;
      RECT  815850.0 376350.0 817050.0 377550.0 ;
      RECT  818850.0 354450.0 820050.0 355650.0 ;
      RECT  816300.0 369750.0 817500.0 370950.0 ;
      RECT  818700.0 359250.0 819900.0 360450.0 ;
      RECT  822600.0 357450.0 823800.0 358650.0 ;
      RECT  816000.0 376950.0 816900.0 378750.0 ;
      RECT  819000.0 376950.0 819900.0 378750.0 ;
      RECT  816000.0 353250.0 816900.0 355050.0 ;
      RECT  819000.0 353250.0 819900.0 355050.0 ;
      RECT  812400.0 353250.0 813300.0 378750.0 ;
      RECT  822600.0 353250.0 823500.0 378750.0 ;
      RECT  826200.0 361950.0 827100.0 362850.0 ;
      RECT  826650.0 361950.0 827550.0 362850.0 ;
      RECT  826200.0 355050.0 827100.0 362400.0 ;
      RECT  826650.0 361950.0 827100.0 362850.0 ;
      RECT  826650.0 362400.0 827550.0 369750.0 ;
      RECT  829200.0 368250.0 830100.0 369150.0 ;
      RECT  829050.0 368250.0 829950.0 369150.0 ;
      RECT  829200.0 368700.0 830100.0 376950.0 ;
      RECT  829500.0 368250.0 829650.0 369150.0 ;
      RECT  829050.0 360450.0 829950.0 368700.0 ;
      RECT  826050.0 376350.0 827250.0 377550.0 ;
      RECT  829050.0 354450.0 830250.0 355650.0 ;
      RECT  826500.0 369750.0 827700.0 370950.0 ;
      RECT  828900.0 359250.0 830100.0 360450.0 ;
      RECT  832800.0 357450.0 834000.0 358650.0 ;
      RECT  826200.0 376950.0 827100.0 378750.0 ;
      RECT  829200.0 376950.0 830100.0 378750.0 ;
      RECT  826200.0 353250.0 827100.0 355050.0 ;
      RECT  829200.0 353250.0 830100.0 355050.0 ;
      RECT  822600.0 353250.0 823500.0 378750.0 ;
      RECT  832800.0 353250.0 833700.0 378750.0 ;
      RECT  836400.0 361950.0 837300.0 362850.0 ;
      RECT  836850.0 361950.0 837750.0 362850.0 ;
      RECT  836400.0 355050.0 837300.0 362400.0 ;
      RECT  836850.0 361950.0 837300.0 362850.0 ;
      RECT  836850.0 362400.0 837750.0 369750.0 ;
      RECT  839400.0 368250.0 840300.0 369150.0 ;
      RECT  839250.0 368250.0 840150.0 369150.0 ;
      RECT  839400.0 368700.0 840300.0 376950.0 ;
      RECT  839700.0 368250.0 839850.0 369150.0 ;
      RECT  839250.0 360450.0 840150.0 368700.0 ;
      RECT  836250.0 376350.0 837450.0 377550.0 ;
      RECT  839250.0 354450.0 840450.0 355650.0 ;
      RECT  836700.0 369750.0 837900.0 370950.0 ;
      RECT  839100.0 359250.0 840300.0 360450.0 ;
      RECT  843000.0 357450.0 844200.0 358650.0 ;
      RECT  836400.0 376950.0 837300.0 378750.0 ;
      RECT  839400.0 376950.0 840300.0 378750.0 ;
      RECT  836400.0 353250.0 837300.0 355050.0 ;
      RECT  839400.0 353250.0 840300.0 355050.0 ;
      RECT  832800.0 353250.0 833700.0 378750.0 ;
      RECT  843000.0 353250.0 843900.0 378750.0 ;
      RECT  846600.0 361950.0 847500.0 362850.0 ;
      RECT  847050.0 361950.0 847950.0 362850.0 ;
      RECT  846600.0 355050.0 847500.0 362400.0 ;
      RECT  847050.0 361950.0 847500.0 362850.0 ;
      RECT  847050.0 362400.0 847950.0 369750.0 ;
      RECT  849600.0 368250.0 850500.0 369150.0 ;
      RECT  849450.0 368250.0 850350.0 369150.0 ;
      RECT  849600.0 368700.0 850500.0 376950.0 ;
      RECT  849900.0 368250.0 850050.0 369150.0 ;
      RECT  849450.0 360450.0 850350.0 368700.0 ;
      RECT  846450.0 376350.0 847650.0 377550.0 ;
      RECT  849450.0 354450.0 850650.0 355650.0 ;
      RECT  846900.0 369750.0 848100.0 370950.0 ;
      RECT  849300.0 359250.0 850500.0 360450.0 ;
      RECT  853200.0 357450.0 854400.0 358650.0 ;
      RECT  846600.0 376950.0 847500.0 378750.0 ;
      RECT  849600.0 376950.0 850500.0 378750.0 ;
      RECT  846600.0 353250.0 847500.0 355050.0 ;
      RECT  849600.0 353250.0 850500.0 355050.0 ;
      RECT  843000.0 353250.0 843900.0 378750.0 ;
      RECT  853200.0 353250.0 854100.0 378750.0 ;
      RECT  856800.0 361950.0 857700.0 362850.0 ;
      RECT  857250.0 361950.0 858150.0 362850.0 ;
      RECT  856800.0 355050.0 857700.0 362400.0 ;
      RECT  857250.0 361950.0 857700.0 362850.0 ;
      RECT  857250.0 362400.0 858150.0 369750.0 ;
      RECT  859800.0 368250.0 860700.0 369150.0 ;
      RECT  859650.0 368250.0 860550.0 369150.0 ;
      RECT  859800.0 368700.0 860700.0 376950.0 ;
      RECT  860100.0 368250.0 860250.0 369150.0 ;
      RECT  859650.0 360450.0 860550.0 368700.0 ;
      RECT  856650.0 376350.0 857850.0 377550.0 ;
      RECT  859650.0 354450.0 860850.0 355650.0 ;
      RECT  857100.0 369750.0 858300.0 370950.0 ;
      RECT  859500.0 359250.0 860700.0 360450.0 ;
      RECT  863400.0 357450.0 864600.0 358650.0 ;
      RECT  856800.0 376950.0 857700.0 378750.0 ;
      RECT  859800.0 376950.0 860700.0 378750.0 ;
      RECT  856800.0 353250.0 857700.0 355050.0 ;
      RECT  859800.0 353250.0 860700.0 355050.0 ;
      RECT  853200.0 353250.0 854100.0 378750.0 ;
      RECT  863400.0 353250.0 864300.0 378750.0 ;
      RECT  867000.0 361950.0 867900.0 362850.0 ;
      RECT  867450.0 361950.0 868350.0 362850.0 ;
      RECT  867000.0 355050.0 867900.0 362400.0 ;
      RECT  867450.0 361950.0 867900.0 362850.0 ;
      RECT  867450.0 362400.0 868350.0 369750.0 ;
      RECT  870000.0 368250.0 870900.0 369150.0 ;
      RECT  869850.0 368250.0 870750.0 369150.0 ;
      RECT  870000.0 368700.0 870900.0 376950.0 ;
      RECT  870300.0 368250.0 870450.0 369150.0 ;
      RECT  869850.0 360450.0 870750.0 368700.0 ;
      RECT  866850.0 376350.0 868050.0 377550.0 ;
      RECT  869850.0 354450.0 871050.0 355650.0 ;
      RECT  867300.0 369750.0 868500.0 370950.0 ;
      RECT  869700.0 359250.0 870900.0 360450.0 ;
      RECT  873600.0 357450.0 874800.0 358650.0 ;
      RECT  867000.0 376950.0 867900.0 378750.0 ;
      RECT  870000.0 376950.0 870900.0 378750.0 ;
      RECT  867000.0 353250.0 867900.0 355050.0 ;
      RECT  870000.0 353250.0 870900.0 355050.0 ;
      RECT  863400.0 353250.0 864300.0 378750.0 ;
      RECT  873600.0 353250.0 874500.0 378750.0 ;
      RECT  877200.0 361950.0 878100.0 362850.0 ;
      RECT  877650.0 361950.0 878550.0 362850.0 ;
      RECT  877200.0 355050.0 878100.0 362400.0 ;
      RECT  877650.0 361950.0 878100.0 362850.0 ;
      RECT  877650.0 362400.0 878550.0 369750.0 ;
      RECT  880200.0 368250.0 881100.0 369150.0 ;
      RECT  880050.0 368250.0 880950.0 369150.0 ;
      RECT  880200.0 368700.0 881100.0 376950.0 ;
      RECT  880500.0 368250.0 880650.0 369150.0 ;
      RECT  880050.0 360450.0 880950.0 368700.0 ;
      RECT  877050.0 376350.0 878250.0 377550.0 ;
      RECT  880050.0 354450.0 881250.0 355650.0 ;
      RECT  877500.0 369750.0 878700.0 370950.0 ;
      RECT  879900.0 359250.0 881100.0 360450.0 ;
      RECT  883800.0 357450.0 885000.0 358650.0 ;
      RECT  877200.0 376950.0 878100.0 378750.0 ;
      RECT  880200.0 376950.0 881100.0 378750.0 ;
      RECT  877200.0 353250.0 878100.0 355050.0 ;
      RECT  880200.0 353250.0 881100.0 355050.0 ;
      RECT  873600.0 353250.0 874500.0 378750.0 ;
      RECT  883800.0 353250.0 884700.0 378750.0 ;
      RECT  887400.0 361950.0 888300.0 362850.0 ;
      RECT  887850.0 361950.0 888750.0 362850.0 ;
      RECT  887400.0 355050.0 888300.0 362400.0 ;
      RECT  887850.0 361950.0 888300.0 362850.0 ;
      RECT  887850.0 362400.0 888750.0 369750.0 ;
      RECT  890400.0 368250.0 891300.0 369150.0 ;
      RECT  890250.0 368250.0 891150.0 369150.0 ;
      RECT  890400.0 368700.0 891300.0 376950.0 ;
      RECT  890700.0 368250.0 890850.0 369150.0 ;
      RECT  890250.0 360450.0 891150.0 368700.0 ;
      RECT  887250.0 376350.0 888450.0 377550.0 ;
      RECT  890250.0 354450.0 891450.0 355650.0 ;
      RECT  887700.0 369750.0 888900.0 370950.0 ;
      RECT  890100.0 359250.0 891300.0 360450.0 ;
      RECT  894000.0 357450.0 895200.0 358650.0 ;
      RECT  887400.0 376950.0 888300.0 378750.0 ;
      RECT  890400.0 376950.0 891300.0 378750.0 ;
      RECT  887400.0 353250.0 888300.0 355050.0 ;
      RECT  890400.0 353250.0 891300.0 355050.0 ;
      RECT  883800.0 353250.0 884700.0 378750.0 ;
      RECT  894000.0 353250.0 894900.0 378750.0 ;
      RECT  897600.0 361950.0 898500.0 362850.0 ;
      RECT  898050.0 361950.0 898950.0 362850.0 ;
      RECT  897600.0 355050.0 898500.0 362400.0 ;
      RECT  898050.0 361950.0 898500.0 362850.0 ;
      RECT  898050.0 362400.0 898950.0 369750.0 ;
      RECT  900600.0 368250.0 901500.0 369150.0 ;
      RECT  900450.0 368250.0 901350.0 369150.0 ;
      RECT  900600.0 368700.0 901500.0 376950.0 ;
      RECT  900900.0 368250.0 901050.0 369150.0 ;
      RECT  900450.0 360450.0 901350.0 368700.0 ;
      RECT  897450.0 376350.0 898650.0 377550.0 ;
      RECT  900450.0 354450.0 901650.0 355650.0 ;
      RECT  897900.0 369750.0 899100.0 370950.0 ;
      RECT  900300.0 359250.0 901500.0 360450.0 ;
      RECT  904200.0 357450.0 905400.0 358650.0 ;
      RECT  897600.0 376950.0 898500.0 378750.0 ;
      RECT  900600.0 376950.0 901500.0 378750.0 ;
      RECT  897600.0 353250.0 898500.0 355050.0 ;
      RECT  900600.0 353250.0 901500.0 355050.0 ;
      RECT  894000.0 353250.0 894900.0 378750.0 ;
      RECT  904200.0 353250.0 905100.0 378750.0 ;
      RECT  907800.0 361950.0 908700.0 362850.0 ;
      RECT  908250.0 361950.0 909150.0 362850.0 ;
      RECT  907800.0 355050.0 908700.0 362400.0 ;
      RECT  908250.0 361950.0 908700.0 362850.0 ;
      RECT  908250.0 362400.0 909150.0 369750.0 ;
      RECT  910800.0 368250.0 911700.0 369150.0 ;
      RECT  910650.0 368250.0 911550.0 369150.0 ;
      RECT  910800.0 368700.0 911700.0 376950.0 ;
      RECT  911100.0 368250.0 911250.0 369150.0 ;
      RECT  910650.0 360450.0 911550.0 368700.0 ;
      RECT  907650.0 376350.0 908850.0 377550.0 ;
      RECT  910650.0 354450.0 911850.0 355650.0 ;
      RECT  908100.0 369750.0 909300.0 370950.0 ;
      RECT  910500.0 359250.0 911700.0 360450.0 ;
      RECT  914400.0 357450.0 915600.0 358650.0 ;
      RECT  907800.0 376950.0 908700.0 378750.0 ;
      RECT  910800.0 376950.0 911700.0 378750.0 ;
      RECT  907800.0 353250.0 908700.0 355050.0 ;
      RECT  910800.0 353250.0 911700.0 355050.0 ;
      RECT  904200.0 353250.0 905100.0 378750.0 ;
      RECT  914400.0 353250.0 915300.0 378750.0 ;
      RECT  918000.0 361950.0 918900.0 362850.0 ;
      RECT  918450.0 361950.0 919350.0 362850.0 ;
      RECT  918000.0 355050.0 918900.0 362400.0 ;
      RECT  918450.0 361950.0 918900.0 362850.0 ;
      RECT  918450.0 362400.0 919350.0 369750.0 ;
      RECT  921000.0 368250.0 921900.0 369150.0 ;
      RECT  920850.0 368250.0 921750.0 369150.0 ;
      RECT  921000.0 368700.0 921900.0 376950.0 ;
      RECT  921300.0 368250.0 921450.0 369150.0 ;
      RECT  920850.0 360450.0 921750.0 368700.0 ;
      RECT  917850.0 376350.0 919050.0 377550.0 ;
      RECT  920850.0 354450.0 922050.0 355650.0 ;
      RECT  918300.0 369750.0 919500.0 370950.0 ;
      RECT  920700.0 359250.0 921900.0 360450.0 ;
      RECT  924600.0 357450.0 925800.0 358650.0 ;
      RECT  918000.0 376950.0 918900.0 378750.0 ;
      RECT  921000.0 376950.0 921900.0 378750.0 ;
      RECT  918000.0 353250.0 918900.0 355050.0 ;
      RECT  921000.0 353250.0 921900.0 355050.0 ;
      RECT  914400.0 353250.0 915300.0 378750.0 ;
      RECT  924600.0 353250.0 925500.0 378750.0 ;
      RECT  928200.0 361950.0 929100.0 362850.0 ;
      RECT  928650.0 361950.0 929550.0 362850.0 ;
      RECT  928200.0 355050.0 929100.0 362400.0 ;
      RECT  928650.0 361950.0 929100.0 362850.0 ;
      RECT  928650.0 362400.0 929550.0 369750.0 ;
      RECT  931200.0 368250.0 932100.0 369150.0 ;
      RECT  931050.0 368250.0 931950.0 369150.0 ;
      RECT  931200.0 368700.0 932100.0 376950.0 ;
      RECT  931500.0 368250.0 931650.0 369150.0 ;
      RECT  931050.0 360450.0 931950.0 368700.0 ;
      RECT  928050.0 376350.0 929250.0 377550.0 ;
      RECT  931050.0 354450.0 932250.0 355650.0 ;
      RECT  928500.0 369750.0 929700.0 370950.0 ;
      RECT  930900.0 359250.0 932100.0 360450.0 ;
      RECT  934800.0 357450.0 936000.0 358650.0 ;
      RECT  928200.0 376950.0 929100.0 378750.0 ;
      RECT  931200.0 376950.0 932100.0 378750.0 ;
      RECT  928200.0 353250.0 929100.0 355050.0 ;
      RECT  931200.0 353250.0 932100.0 355050.0 ;
      RECT  924600.0 353250.0 925500.0 378750.0 ;
      RECT  934800.0 353250.0 935700.0 378750.0 ;
      RECT  938400.0 361950.0 939300.0 362850.0 ;
      RECT  938850.0 361950.0 939750.0 362850.0 ;
      RECT  938400.0 355050.0 939300.0 362400.0 ;
      RECT  938850.0 361950.0 939300.0 362850.0 ;
      RECT  938850.0 362400.0 939750.0 369750.0 ;
      RECT  941400.0 368250.0 942300.0 369150.0 ;
      RECT  941250.0 368250.0 942150.0 369150.0 ;
      RECT  941400.0 368700.0 942300.0 376950.0 ;
      RECT  941700.0 368250.0 941850.0 369150.0 ;
      RECT  941250.0 360450.0 942150.0 368700.0 ;
      RECT  938250.0 376350.0 939450.0 377550.0 ;
      RECT  941250.0 354450.0 942450.0 355650.0 ;
      RECT  938700.0 369750.0 939900.0 370950.0 ;
      RECT  941100.0 359250.0 942300.0 360450.0 ;
      RECT  945000.0 357450.0 946200.0 358650.0 ;
      RECT  938400.0 376950.0 939300.0 378750.0 ;
      RECT  941400.0 376950.0 942300.0 378750.0 ;
      RECT  938400.0 353250.0 939300.0 355050.0 ;
      RECT  941400.0 353250.0 942300.0 355050.0 ;
      RECT  934800.0 353250.0 935700.0 378750.0 ;
      RECT  945000.0 353250.0 945900.0 378750.0 ;
      RECT  948600.0 361950.0 949500.0 362850.0 ;
      RECT  949050.0 361950.0 949950.0 362850.0 ;
      RECT  948600.0 355050.0 949500.0 362400.0 ;
      RECT  949050.0 361950.0 949500.0 362850.0 ;
      RECT  949050.0 362400.0 949950.0 369750.0 ;
      RECT  951600.0 368250.0 952500.0 369150.0 ;
      RECT  951450.0 368250.0 952350.0 369150.0 ;
      RECT  951600.0 368700.0 952500.0 376950.0 ;
      RECT  951900.0 368250.0 952050.0 369150.0 ;
      RECT  951450.0 360450.0 952350.0 368700.0 ;
      RECT  948450.0 376350.0 949650.0 377550.0 ;
      RECT  951450.0 354450.0 952650.0 355650.0 ;
      RECT  948900.0 369750.0 950100.0 370950.0 ;
      RECT  951300.0 359250.0 952500.0 360450.0 ;
      RECT  955200.0 357450.0 956400.0 358650.0 ;
      RECT  948600.0 376950.0 949500.0 378750.0 ;
      RECT  951600.0 376950.0 952500.0 378750.0 ;
      RECT  948600.0 353250.0 949500.0 355050.0 ;
      RECT  951600.0 353250.0 952500.0 355050.0 ;
      RECT  945000.0 353250.0 945900.0 378750.0 ;
      RECT  955200.0 353250.0 956100.0 378750.0 ;
      RECT  958800.0 361950.0 959700.0 362850.0 ;
      RECT  959250.0 361950.0 960150.0 362850.0 ;
      RECT  958800.0 355050.0 959700.0 362400.0 ;
      RECT  959250.0 361950.0 959700.0 362850.0 ;
      RECT  959250.0 362400.0 960150.0 369750.0 ;
      RECT  961800.0 368250.0 962700.0 369150.0 ;
      RECT  961650.0 368250.0 962550.0 369150.0 ;
      RECT  961800.0 368700.0 962700.0 376950.0 ;
      RECT  962100.0 368250.0 962250.0 369150.0 ;
      RECT  961650.0 360450.0 962550.0 368700.0 ;
      RECT  958650.0 376350.0 959850.0 377550.0 ;
      RECT  961650.0 354450.0 962850.0 355650.0 ;
      RECT  959100.0 369750.0 960300.0 370950.0 ;
      RECT  961500.0 359250.0 962700.0 360450.0 ;
      RECT  965400.0 357450.0 966600.0 358650.0 ;
      RECT  958800.0 376950.0 959700.0 378750.0 ;
      RECT  961800.0 376950.0 962700.0 378750.0 ;
      RECT  958800.0 353250.0 959700.0 355050.0 ;
      RECT  961800.0 353250.0 962700.0 355050.0 ;
      RECT  955200.0 353250.0 956100.0 378750.0 ;
      RECT  965400.0 353250.0 966300.0 378750.0 ;
      RECT  969000.0 361950.0 969900.0 362850.0 ;
      RECT  969450.0 361950.0 970350.0 362850.0 ;
      RECT  969000.0 355050.0 969900.0 362400.0 ;
      RECT  969450.0 361950.0 969900.0 362850.0 ;
      RECT  969450.0 362400.0 970350.0 369750.0 ;
      RECT  972000.0 368250.0 972900.0 369150.0 ;
      RECT  971850.0 368250.0 972750.0 369150.0 ;
      RECT  972000.0 368700.0 972900.0 376950.0 ;
      RECT  972300.0 368250.0 972450.0 369150.0 ;
      RECT  971850.0 360450.0 972750.0 368700.0 ;
      RECT  968850.0 376350.0 970050.0 377550.0 ;
      RECT  971850.0 354450.0 973050.0 355650.0 ;
      RECT  969300.0 369750.0 970500.0 370950.0 ;
      RECT  971700.0 359250.0 972900.0 360450.0 ;
      RECT  975600.0 357450.0 976800.0 358650.0 ;
      RECT  969000.0 376950.0 969900.0 378750.0 ;
      RECT  972000.0 376950.0 972900.0 378750.0 ;
      RECT  969000.0 353250.0 969900.0 355050.0 ;
      RECT  972000.0 353250.0 972900.0 355050.0 ;
      RECT  965400.0 353250.0 966300.0 378750.0 ;
      RECT  975600.0 353250.0 976500.0 378750.0 ;
      RECT  979200.0 361950.0 980100.0 362850.0 ;
      RECT  979650.0 361950.0 980550.0 362850.0 ;
      RECT  979200.0 355050.0 980100.0 362400.0 ;
      RECT  979650.0 361950.0 980100.0 362850.0 ;
      RECT  979650.0 362400.0 980550.0 369750.0 ;
      RECT  982200.0 368250.0 983100.0 369150.0 ;
      RECT  982050.0 368250.0 982950.0 369150.0 ;
      RECT  982200.0 368700.0 983100.0 376950.0 ;
      RECT  982500.0 368250.0 982650.0 369150.0 ;
      RECT  982050.0 360450.0 982950.0 368700.0 ;
      RECT  979050.0 376350.0 980250.0 377550.0 ;
      RECT  982050.0 354450.0 983250.0 355650.0 ;
      RECT  979500.0 369750.0 980700.0 370950.0 ;
      RECT  981900.0 359250.0 983100.0 360450.0 ;
      RECT  985800.0 357450.0 987000.0 358650.0 ;
      RECT  979200.0 376950.0 980100.0 378750.0 ;
      RECT  982200.0 376950.0 983100.0 378750.0 ;
      RECT  979200.0 353250.0 980100.0 355050.0 ;
      RECT  982200.0 353250.0 983100.0 355050.0 ;
      RECT  975600.0 353250.0 976500.0 378750.0 ;
      RECT  985800.0 353250.0 986700.0 378750.0 ;
      RECT  989400.0 361950.0 990300.0 362850.0 ;
      RECT  989850.0 361950.0 990750.0 362850.0 ;
      RECT  989400.0 355050.0 990300.0 362400.0 ;
      RECT  989850.0 361950.0 990300.0 362850.0 ;
      RECT  989850.0 362400.0 990750.0 369750.0 ;
      RECT  992400.0 368250.0 993300.0 369150.0 ;
      RECT  992250.0 368250.0 993150.0 369150.0 ;
      RECT  992400.0 368700.0 993300.0 376950.0 ;
      RECT  992700.0 368250.0 992850.0 369150.0 ;
      RECT  992250.0 360450.0 993150.0 368700.0 ;
      RECT  989250.0 376350.0 990450.0 377550.0 ;
      RECT  992250.0 354450.0 993450.0 355650.0 ;
      RECT  989700.0 369750.0 990900.0 370950.0 ;
      RECT  992100.0 359250.0 993300.0 360450.0 ;
      RECT  996000.0 357450.0 997200.0 358650.0 ;
      RECT  989400.0 376950.0 990300.0 378750.0 ;
      RECT  992400.0 376950.0 993300.0 378750.0 ;
      RECT  989400.0 353250.0 990300.0 355050.0 ;
      RECT  992400.0 353250.0 993300.0 355050.0 ;
      RECT  985800.0 353250.0 986700.0 378750.0 ;
      RECT  996000.0 353250.0 996900.0 378750.0 ;
      RECT  999600.0 361950.0 1000500.0 362850.0 ;
      RECT  1000050.0 361950.0 1000950.0 362850.0 ;
      RECT  999600.0 355050.0 1000500.0 362400.0 ;
      RECT  1000050.0 361950.0 1000500.0 362850.0 ;
      RECT  1000050.0 362400.0 1000950.0 369750.0 ;
      RECT  1002600.0 368250.0 1003500.0 369150.0 ;
      RECT  1002450.0 368250.0 1003350.0 369150.0 ;
      RECT  1002600.0 368700.0 1003500.0 376950.0 ;
      RECT  1002900.0 368250.0 1003050.0 369150.0 ;
      RECT  1002450.0 360450.0 1003350.0 368700.0 ;
      RECT  999450.0 376350.0 1000650.0 377550.0 ;
      RECT  1002450.0 354450.0 1003650.0 355650.0 ;
      RECT  999900.0 369750.0 1001100.0 370950.0 ;
      RECT  1002300.0 359250.0 1003500.0 360450.0 ;
      RECT  1006200.0 357450.0 1007400.0 358650.0 ;
      RECT  999600.0 376950.0 1000500.0 378750.0 ;
      RECT  1002600.0 376950.0 1003500.0 378750.0 ;
      RECT  999600.0 353250.0 1000500.0 355050.0 ;
      RECT  1002600.0 353250.0 1003500.0 355050.0 ;
      RECT  996000.0 353250.0 996900.0 378750.0 ;
      RECT  1006200.0 353250.0 1007100.0 378750.0 ;
      RECT  1009800.0 361950.0 1010700.0 362850.0 ;
      RECT  1010250.0 361950.0 1011150.0 362850.0 ;
      RECT  1009800.0 355050.0 1010700.0 362400.0 ;
      RECT  1010250.0 361950.0 1010700.0 362850.0 ;
      RECT  1010250.0 362400.0 1011150.0 369750.0 ;
      RECT  1012800.0 368250.0 1013700.0 369150.0 ;
      RECT  1012650.0 368250.0 1013550.0 369150.0 ;
      RECT  1012800.0 368700.0 1013700.0 376950.0 ;
      RECT  1013100.0 368250.0 1013250.0 369150.0 ;
      RECT  1012650.0 360450.0 1013550.0 368700.0 ;
      RECT  1009650.0 376350.0 1010850.0 377550.0 ;
      RECT  1012650.0 354450.0 1013850.0 355650.0 ;
      RECT  1010100.0 369750.0 1011300.0 370950.0 ;
      RECT  1012500.0 359250.0 1013700.0 360450.0 ;
      RECT  1016400.0 357450.0 1017600.0 358650.0 ;
      RECT  1009800.0 376950.0 1010700.0 378750.0 ;
      RECT  1012800.0 376950.0 1013700.0 378750.0 ;
      RECT  1009800.0 353250.0 1010700.0 355050.0 ;
      RECT  1012800.0 353250.0 1013700.0 355050.0 ;
      RECT  1006200.0 353250.0 1007100.0 378750.0 ;
      RECT  1016400.0 353250.0 1017300.0 378750.0 ;
      RECT  1020000.0 361950.0 1020900.0 362850.0 ;
      RECT  1020450.0 361950.0 1021350.0 362850.0 ;
      RECT  1020000.0 355050.0 1020900.0 362400.0 ;
      RECT  1020450.0 361950.0 1020900.0 362850.0 ;
      RECT  1020450.0 362400.0 1021350.0 369750.0 ;
      RECT  1023000.0 368250.0 1023900.0 369150.0 ;
      RECT  1022850.0 368250.0 1023750.0 369150.0 ;
      RECT  1023000.0 368700.0 1023900.0 376950.0 ;
      RECT  1023300.0 368250.0 1023450.0 369150.0 ;
      RECT  1022850.0 360450.0 1023750.0 368700.0 ;
      RECT  1019850.0 376350.0 1021050.0 377550.0 ;
      RECT  1022850.0 354450.0 1024050.0 355650.0 ;
      RECT  1020300.0 369750.0 1021500.0 370950.0 ;
      RECT  1022700.0 359250.0 1023900.0 360450.0 ;
      RECT  1026600.0 357450.0 1027800.0 358650.0 ;
      RECT  1020000.0 376950.0 1020900.0 378750.0 ;
      RECT  1023000.0 376950.0 1023900.0 378750.0 ;
      RECT  1020000.0 353250.0 1020900.0 355050.0 ;
      RECT  1023000.0 353250.0 1023900.0 355050.0 ;
      RECT  1016400.0 353250.0 1017300.0 378750.0 ;
      RECT  1026600.0 353250.0 1027500.0 378750.0 ;
      RECT  1030200.0 361950.0 1031100.0 362850.0 ;
      RECT  1030650.0 361950.0 1031550.0 362850.0 ;
      RECT  1030200.0 355050.0 1031100.0 362400.0 ;
      RECT  1030650.0 361950.0 1031100.0 362850.0 ;
      RECT  1030650.0 362400.0 1031550.0 369750.0 ;
      RECT  1033200.0 368250.0 1034100.0 369150.0 ;
      RECT  1033050.0 368250.0 1033950.0 369150.0 ;
      RECT  1033200.0 368700.0 1034100.0 376950.0 ;
      RECT  1033500.0 368250.0 1033650.0 369150.0 ;
      RECT  1033050.0 360450.0 1033950.0 368700.0 ;
      RECT  1030050.0 376350.0 1031250.0 377550.0 ;
      RECT  1033050.0 354450.0 1034250.0 355650.0 ;
      RECT  1030500.0 369750.0 1031700.0 370950.0 ;
      RECT  1032900.0 359250.0 1034100.0 360450.0 ;
      RECT  1036800.0 357450.0 1038000.0 358650.0 ;
      RECT  1030200.0 376950.0 1031100.0 378750.0 ;
      RECT  1033200.0 376950.0 1034100.0 378750.0 ;
      RECT  1030200.0 353250.0 1031100.0 355050.0 ;
      RECT  1033200.0 353250.0 1034100.0 355050.0 ;
      RECT  1026600.0 353250.0 1027500.0 378750.0 ;
      RECT  1036800.0 353250.0 1037700.0 378750.0 ;
      RECT  1040400.0 361950.0 1041300.0 362850.0 ;
      RECT  1040850.0 361950.0 1041750.0 362850.0 ;
      RECT  1040400.0 355050.0 1041300.0 362400.0 ;
      RECT  1040850.0 361950.0 1041300.0 362850.0 ;
      RECT  1040850.0 362400.0 1041750.0 369750.0 ;
      RECT  1043400.0 368250.0 1044300.0 369150.0 ;
      RECT  1043250.0 368250.0 1044150.0 369150.0 ;
      RECT  1043400.0 368700.0 1044300.0 376950.0 ;
      RECT  1043700.0 368250.0 1043850.0 369150.0 ;
      RECT  1043250.0 360450.0 1044150.0 368700.0 ;
      RECT  1040250.0 376350.0 1041450.0 377550.0 ;
      RECT  1043250.0 354450.0 1044450.0 355650.0 ;
      RECT  1040700.0 369750.0 1041900.0 370950.0 ;
      RECT  1043100.0 359250.0 1044300.0 360450.0 ;
      RECT  1047000.0 357450.0 1048200.0 358650.0 ;
      RECT  1040400.0 376950.0 1041300.0 378750.0 ;
      RECT  1043400.0 376950.0 1044300.0 378750.0 ;
      RECT  1040400.0 353250.0 1041300.0 355050.0 ;
      RECT  1043400.0 353250.0 1044300.0 355050.0 ;
      RECT  1036800.0 353250.0 1037700.0 378750.0 ;
      RECT  1047000.0 353250.0 1047900.0 378750.0 ;
      RECT  1050600.0 361950.0 1051500.0 362850.0 ;
      RECT  1051050.0 361950.0 1051950.0 362850.0 ;
      RECT  1050600.0 355050.0 1051500.0 362400.0 ;
      RECT  1051050.0 361950.0 1051500.0 362850.0 ;
      RECT  1051050.0 362400.0 1051950.0 369750.0 ;
      RECT  1053600.0 368250.0 1054500.0 369150.0 ;
      RECT  1053450.0 368250.0 1054350.0 369150.0 ;
      RECT  1053600.0 368700.0 1054500.0 376950.0 ;
      RECT  1053900.0 368250.0 1054050.0 369150.0 ;
      RECT  1053450.0 360450.0 1054350.0 368700.0 ;
      RECT  1050450.0 376350.0 1051650.0 377550.0 ;
      RECT  1053450.0 354450.0 1054650.0 355650.0 ;
      RECT  1050900.0 369750.0 1052100.0 370950.0 ;
      RECT  1053300.0 359250.0 1054500.0 360450.0 ;
      RECT  1057200.0 357450.0 1058400.0 358650.0 ;
      RECT  1050600.0 376950.0 1051500.0 378750.0 ;
      RECT  1053600.0 376950.0 1054500.0 378750.0 ;
      RECT  1050600.0 353250.0 1051500.0 355050.0 ;
      RECT  1053600.0 353250.0 1054500.0 355050.0 ;
      RECT  1047000.0 353250.0 1047900.0 378750.0 ;
      RECT  1057200.0 353250.0 1058100.0 378750.0 ;
      RECT  1060800.0 361950.0 1061700.0 362850.0 ;
      RECT  1061250.0 361950.0 1062150.0 362850.0 ;
      RECT  1060800.0 355050.0 1061700.0 362400.0 ;
      RECT  1061250.0 361950.0 1061700.0 362850.0 ;
      RECT  1061250.0 362400.0 1062150.0 369750.0 ;
      RECT  1063800.0 368250.0 1064700.0 369150.0 ;
      RECT  1063650.0 368250.0 1064550.0 369150.0 ;
      RECT  1063800.0 368700.0 1064700.0 376950.0 ;
      RECT  1064100.0 368250.0 1064250.0 369150.0 ;
      RECT  1063650.0 360450.0 1064550.0 368700.0 ;
      RECT  1060650.0 376350.0 1061850.0 377550.0 ;
      RECT  1063650.0 354450.0 1064850.0 355650.0 ;
      RECT  1061100.0 369750.0 1062300.0 370950.0 ;
      RECT  1063500.0 359250.0 1064700.0 360450.0 ;
      RECT  1067400.0 357450.0 1068600.0 358650.0 ;
      RECT  1060800.0 376950.0 1061700.0 378750.0 ;
      RECT  1063800.0 376950.0 1064700.0 378750.0 ;
      RECT  1060800.0 353250.0 1061700.0 355050.0 ;
      RECT  1063800.0 353250.0 1064700.0 355050.0 ;
      RECT  1057200.0 353250.0 1058100.0 378750.0 ;
      RECT  1067400.0 353250.0 1068300.0 378750.0 ;
      RECT  1071000.0 361950.0 1071900.0 362850.0 ;
      RECT  1071450.0 361950.0 1072350.0 362850.0 ;
      RECT  1071000.0 355050.0 1071900.0 362400.0 ;
      RECT  1071450.0 361950.0 1071900.0 362850.0 ;
      RECT  1071450.0 362400.0 1072350.0 369750.0 ;
      RECT  1074000.0 368250.0 1074900.0 369150.0 ;
      RECT  1073850.0 368250.0 1074750.0 369150.0 ;
      RECT  1074000.0 368700.0 1074900.0 376950.0 ;
      RECT  1074300.0 368250.0 1074450.0 369150.0 ;
      RECT  1073850.0 360450.0 1074750.0 368700.0 ;
      RECT  1070850.0 376350.0 1072050.0 377550.0 ;
      RECT  1073850.0 354450.0 1075050.0 355650.0 ;
      RECT  1071300.0 369750.0 1072500.0 370950.0 ;
      RECT  1073700.0 359250.0 1074900.0 360450.0 ;
      RECT  1077600.0 357450.0 1078800.0 358650.0 ;
      RECT  1071000.0 376950.0 1071900.0 378750.0 ;
      RECT  1074000.0 376950.0 1074900.0 378750.0 ;
      RECT  1071000.0 353250.0 1071900.0 355050.0 ;
      RECT  1074000.0 353250.0 1074900.0 355050.0 ;
      RECT  1067400.0 353250.0 1068300.0 378750.0 ;
      RECT  1077600.0 353250.0 1078500.0 378750.0 ;
      RECT  1081200.0 361950.0 1082100.0 362850.0 ;
      RECT  1081650.0 361950.0 1082550.0 362850.0 ;
      RECT  1081200.0 355050.0 1082100.0 362400.0 ;
      RECT  1081650.0 361950.0 1082100.0 362850.0 ;
      RECT  1081650.0 362400.0 1082550.0 369750.0 ;
      RECT  1084200.0 368250.0 1085100.0 369150.0 ;
      RECT  1084050.0 368250.0 1084950.0 369150.0 ;
      RECT  1084200.0 368700.0 1085100.0 376950.0 ;
      RECT  1084500.0 368250.0 1084650.0 369150.0 ;
      RECT  1084050.0 360450.0 1084950.0 368700.0 ;
      RECT  1081050.0 376350.0 1082250.0 377550.0 ;
      RECT  1084050.0 354450.0 1085250.0 355650.0 ;
      RECT  1081500.0 369750.0 1082700.0 370950.0 ;
      RECT  1083900.0 359250.0 1085100.0 360450.0 ;
      RECT  1087800.0 357450.0 1089000.0 358650.0 ;
      RECT  1081200.0 376950.0 1082100.0 378750.0 ;
      RECT  1084200.0 376950.0 1085100.0 378750.0 ;
      RECT  1081200.0 353250.0 1082100.0 355050.0 ;
      RECT  1084200.0 353250.0 1085100.0 355050.0 ;
      RECT  1077600.0 353250.0 1078500.0 378750.0 ;
      RECT  1087800.0 353250.0 1088700.0 378750.0 ;
      RECT  1091400.0 361950.0 1092300.0 362850.0 ;
      RECT  1091850.0 361950.0 1092750.0 362850.0 ;
      RECT  1091400.0 355050.0 1092300.0 362400.0 ;
      RECT  1091850.0 361950.0 1092300.0 362850.0 ;
      RECT  1091850.0 362400.0 1092750.0 369750.0 ;
      RECT  1094400.0 368250.0 1095300.0 369150.0 ;
      RECT  1094250.0 368250.0 1095150.0 369150.0 ;
      RECT  1094400.0 368700.0 1095300.0 376950.0 ;
      RECT  1094700.0 368250.0 1094850.0 369150.0 ;
      RECT  1094250.0 360450.0 1095150.0 368700.0 ;
      RECT  1091250.0 376350.0 1092450.0 377550.0 ;
      RECT  1094250.0 354450.0 1095450.0 355650.0 ;
      RECT  1091700.0 369750.0 1092900.0 370950.0 ;
      RECT  1094100.0 359250.0 1095300.0 360450.0 ;
      RECT  1098000.0 357450.0 1099200.0 358650.0 ;
      RECT  1091400.0 376950.0 1092300.0 378750.0 ;
      RECT  1094400.0 376950.0 1095300.0 378750.0 ;
      RECT  1091400.0 353250.0 1092300.0 355050.0 ;
      RECT  1094400.0 353250.0 1095300.0 355050.0 ;
      RECT  1087800.0 353250.0 1088700.0 378750.0 ;
      RECT  1098000.0 353250.0 1098900.0 378750.0 ;
      RECT  1101600.0 361950.0 1102500.0 362850.0 ;
      RECT  1102050.0 361950.0 1102950.0 362850.0 ;
      RECT  1101600.0 355050.0 1102500.0 362400.0 ;
      RECT  1102050.0 361950.0 1102500.0 362850.0 ;
      RECT  1102050.0 362400.0 1102950.0 369750.0 ;
      RECT  1104600.0 368250.0 1105500.0 369150.0 ;
      RECT  1104450.0 368250.0 1105350.0 369150.0 ;
      RECT  1104600.0 368700.0 1105500.0 376950.0 ;
      RECT  1104900.0 368250.0 1105050.0 369150.0 ;
      RECT  1104450.0 360450.0 1105350.0 368700.0 ;
      RECT  1101450.0 376350.0 1102650.0 377550.0 ;
      RECT  1104450.0 354450.0 1105650.0 355650.0 ;
      RECT  1101900.0 369750.0 1103100.0 370950.0 ;
      RECT  1104300.0 359250.0 1105500.0 360450.0 ;
      RECT  1108200.0 357450.0 1109400.0 358650.0 ;
      RECT  1101600.0 376950.0 1102500.0 378750.0 ;
      RECT  1104600.0 376950.0 1105500.0 378750.0 ;
      RECT  1101600.0 353250.0 1102500.0 355050.0 ;
      RECT  1104600.0 353250.0 1105500.0 355050.0 ;
      RECT  1098000.0 353250.0 1098900.0 378750.0 ;
      RECT  1108200.0 353250.0 1109100.0 378750.0 ;
      RECT  1111800.0 361950.0 1112700.0 362850.0 ;
      RECT  1112250.0 361950.0 1113150.0 362850.0 ;
      RECT  1111800.0 355050.0 1112700.0 362400.0 ;
      RECT  1112250.0 361950.0 1112700.0 362850.0 ;
      RECT  1112250.0 362400.0 1113150.0 369750.0 ;
      RECT  1114800.0 368250.0 1115700.0 369150.0 ;
      RECT  1114650.0 368250.0 1115550.0 369150.0 ;
      RECT  1114800.0 368700.0 1115700.0 376950.0 ;
      RECT  1115100.0 368250.0 1115250.0 369150.0 ;
      RECT  1114650.0 360450.0 1115550.0 368700.0 ;
      RECT  1111650.0 376350.0 1112850.0 377550.0 ;
      RECT  1114650.0 354450.0 1115850.0 355650.0 ;
      RECT  1112100.0 369750.0 1113300.0 370950.0 ;
      RECT  1114500.0 359250.0 1115700.0 360450.0 ;
      RECT  1118400.0 357450.0 1119600.0 358650.0 ;
      RECT  1111800.0 376950.0 1112700.0 378750.0 ;
      RECT  1114800.0 376950.0 1115700.0 378750.0 ;
      RECT  1111800.0 353250.0 1112700.0 355050.0 ;
      RECT  1114800.0 353250.0 1115700.0 355050.0 ;
      RECT  1108200.0 353250.0 1109100.0 378750.0 ;
      RECT  1118400.0 353250.0 1119300.0 378750.0 ;
      RECT  1122000.0 361950.0 1122900.0 362850.0 ;
      RECT  1122450.0 361950.0 1123350.0 362850.0 ;
      RECT  1122000.0 355050.0 1122900.0 362400.0 ;
      RECT  1122450.0 361950.0 1122900.0 362850.0 ;
      RECT  1122450.0 362400.0 1123350.0 369750.0 ;
      RECT  1125000.0 368250.0 1125900.0 369150.0 ;
      RECT  1124850.0 368250.0 1125750.0 369150.0 ;
      RECT  1125000.0 368700.0 1125900.0 376950.0 ;
      RECT  1125300.0 368250.0 1125450.0 369150.0 ;
      RECT  1124850.0 360450.0 1125750.0 368700.0 ;
      RECT  1121850.0 376350.0 1123050.0 377550.0 ;
      RECT  1124850.0 354450.0 1126050.0 355650.0 ;
      RECT  1122300.0 369750.0 1123500.0 370950.0 ;
      RECT  1124700.0 359250.0 1125900.0 360450.0 ;
      RECT  1128600.0 357450.0 1129800.0 358650.0 ;
      RECT  1122000.0 376950.0 1122900.0 378750.0 ;
      RECT  1125000.0 376950.0 1125900.0 378750.0 ;
      RECT  1122000.0 353250.0 1122900.0 355050.0 ;
      RECT  1125000.0 353250.0 1125900.0 355050.0 ;
      RECT  1118400.0 353250.0 1119300.0 378750.0 ;
      RECT  1128600.0 353250.0 1129500.0 378750.0 ;
      RECT  1132200.0 361950.0 1133100.0 362850.0 ;
      RECT  1132650.0 361950.0 1133550.0 362850.0 ;
      RECT  1132200.0 355050.0 1133100.0 362400.0 ;
      RECT  1132650.0 361950.0 1133100.0 362850.0 ;
      RECT  1132650.0 362400.0 1133550.0 369750.0 ;
      RECT  1135200.0 368250.0 1136100.0 369150.0 ;
      RECT  1135050.0 368250.0 1135950.0 369150.0 ;
      RECT  1135200.0 368700.0 1136100.0 376950.0 ;
      RECT  1135500.0 368250.0 1135650.0 369150.0 ;
      RECT  1135050.0 360450.0 1135950.0 368700.0 ;
      RECT  1132050.0 376350.0 1133250.0 377550.0 ;
      RECT  1135050.0 354450.0 1136250.0 355650.0 ;
      RECT  1132500.0 369750.0 1133700.0 370950.0 ;
      RECT  1134900.0 359250.0 1136100.0 360450.0 ;
      RECT  1138800.0 357450.0 1140000.0 358650.0 ;
      RECT  1132200.0 376950.0 1133100.0 378750.0 ;
      RECT  1135200.0 376950.0 1136100.0 378750.0 ;
      RECT  1132200.0 353250.0 1133100.0 355050.0 ;
      RECT  1135200.0 353250.0 1136100.0 355050.0 ;
      RECT  1128600.0 353250.0 1129500.0 378750.0 ;
      RECT  1138800.0 353250.0 1139700.0 378750.0 ;
      RECT  1142400.0 361950.0 1143300.0 362850.0 ;
      RECT  1142850.0 361950.0 1143750.0 362850.0 ;
      RECT  1142400.0 355050.0 1143300.0 362400.0 ;
      RECT  1142850.0 361950.0 1143300.0 362850.0 ;
      RECT  1142850.0 362400.0 1143750.0 369750.0 ;
      RECT  1145400.0 368250.0 1146300.0 369150.0 ;
      RECT  1145250.0 368250.0 1146150.0 369150.0 ;
      RECT  1145400.0 368700.0 1146300.0 376950.0 ;
      RECT  1145700.0 368250.0 1145850.0 369150.0 ;
      RECT  1145250.0 360450.0 1146150.0 368700.0 ;
      RECT  1142250.0 376350.0 1143450.0 377550.0 ;
      RECT  1145250.0 354450.0 1146450.0 355650.0 ;
      RECT  1142700.0 369750.0 1143900.0 370950.0 ;
      RECT  1145100.0 359250.0 1146300.0 360450.0 ;
      RECT  1149000.0 357450.0 1150200.0 358650.0 ;
      RECT  1142400.0 376950.0 1143300.0 378750.0 ;
      RECT  1145400.0 376950.0 1146300.0 378750.0 ;
      RECT  1142400.0 353250.0 1143300.0 355050.0 ;
      RECT  1145400.0 353250.0 1146300.0 355050.0 ;
      RECT  1138800.0 353250.0 1139700.0 378750.0 ;
      RECT  1149000.0 353250.0 1149900.0 378750.0 ;
      RECT  1152600.0 361950.0 1153500.0 362850.0 ;
      RECT  1153050.0 361950.0 1153950.0 362850.0 ;
      RECT  1152600.0 355050.0 1153500.0 362400.0 ;
      RECT  1153050.0 361950.0 1153500.0 362850.0 ;
      RECT  1153050.0 362400.0 1153950.0 369750.0 ;
      RECT  1155600.0 368250.0 1156500.0 369150.0 ;
      RECT  1155450.0 368250.0 1156350.0 369150.0 ;
      RECT  1155600.0 368700.0 1156500.0 376950.0 ;
      RECT  1155900.0 368250.0 1156050.0 369150.0 ;
      RECT  1155450.0 360450.0 1156350.0 368700.0 ;
      RECT  1152450.0 376350.0 1153650.0 377550.0 ;
      RECT  1155450.0 354450.0 1156650.0 355650.0 ;
      RECT  1152900.0 369750.0 1154100.0 370950.0 ;
      RECT  1155300.0 359250.0 1156500.0 360450.0 ;
      RECT  1159200.0 357450.0 1160400.0 358650.0 ;
      RECT  1152600.0 376950.0 1153500.0 378750.0 ;
      RECT  1155600.0 376950.0 1156500.0 378750.0 ;
      RECT  1152600.0 353250.0 1153500.0 355050.0 ;
      RECT  1155600.0 353250.0 1156500.0 355050.0 ;
      RECT  1149000.0 353250.0 1149900.0 378750.0 ;
      RECT  1159200.0 353250.0 1160100.0 378750.0 ;
      RECT  1162800.0 361950.0 1163700.0 362850.0 ;
      RECT  1163250.0 361950.0 1164150.0 362850.0 ;
      RECT  1162800.0 355050.0 1163700.0 362400.0 ;
      RECT  1163250.0 361950.0 1163700.0 362850.0 ;
      RECT  1163250.0 362400.0 1164150.0 369750.0 ;
      RECT  1165800.0 368250.0 1166700.0 369150.0 ;
      RECT  1165650.0 368250.0 1166550.0 369150.0 ;
      RECT  1165800.0 368700.0 1166700.0 376950.0 ;
      RECT  1166100.0 368250.0 1166250.0 369150.0 ;
      RECT  1165650.0 360450.0 1166550.0 368700.0 ;
      RECT  1162650.0 376350.0 1163850.0 377550.0 ;
      RECT  1165650.0 354450.0 1166850.0 355650.0 ;
      RECT  1163100.0 369750.0 1164300.0 370950.0 ;
      RECT  1165500.0 359250.0 1166700.0 360450.0 ;
      RECT  1169400.0 357450.0 1170600.0 358650.0 ;
      RECT  1162800.0 376950.0 1163700.0 378750.0 ;
      RECT  1165800.0 376950.0 1166700.0 378750.0 ;
      RECT  1162800.0 353250.0 1163700.0 355050.0 ;
      RECT  1165800.0 353250.0 1166700.0 355050.0 ;
      RECT  1159200.0 353250.0 1160100.0 378750.0 ;
      RECT  1169400.0 353250.0 1170300.0 378750.0 ;
      RECT  1173000.0 361950.0 1173900.0 362850.0 ;
      RECT  1173450.0 361950.0 1174350.0 362850.0 ;
      RECT  1173000.0 355050.0 1173900.0 362400.0 ;
      RECT  1173450.0 361950.0 1173900.0 362850.0 ;
      RECT  1173450.0 362400.0 1174350.0 369750.0 ;
      RECT  1176000.0 368250.0 1176900.0 369150.0 ;
      RECT  1175850.0 368250.0 1176750.0 369150.0 ;
      RECT  1176000.0 368700.0 1176900.0 376950.0 ;
      RECT  1176300.0 368250.0 1176450.0 369150.0 ;
      RECT  1175850.0 360450.0 1176750.0 368700.0 ;
      RECT  1172850.0 376350.0 1174050.0 377550.0 ;
      RECT  1175850.0 354450.0 1177050.0 355650.0 ;
      RECT  1173300.0 369750.0 1174500.0 370950.0 ;
      RECT  1175700.0 359250.0 1176900.0 360450.0 ;
      RECT  1179600.0 357450.0 1180800.0 358650.0 ;
      RECT  1173000.0 376950.0 1173900.0 378750.0 ;
      RECT  1176000.0 376950.0 1176900.0 378750.0 ;
      RECT  1173000.0 353250.0 1173900.0 355050.0 ;
      RECT  1176000.0 353250.0 1176900.0 355050.0 ;
      RECT  1169400.0 353250.0 1170300.0 378750.0 ;
      RECT  1179600.0 353250.0 1180500.0 378750.0 ;
      RECT  1183200.0 361950.0 1184100.0 362850.0 ;
      RECT  1183650.0 361950.0 1184550.0 362850.0 ;
      RECT  1183200.0 355050.0 1184100.0 362400.0 ;
      RECT  1183650.0 361950.0 1184100.0 362850.0 ;
      RECT  1183650.0 362400.0 1184550.0 369750.0 ;
      RECT  1186200.0 368250.0 1187100.0 369150.0 ;
      RECT  1186050.0 368250.0 1186950.0 369150.0 ;
      RECT  1186200.0 368700.0 1187100.0 376950.0 ;
      RECT  1186500.0 368250.0 1186650.0 369150.0 ;
      RECT  1186050.0 360450.0 1186950.0 368700.0 ;
      RECT  1183050.0 376350.0 1184250.0 377550.0 ;
      RECT  1186050.0 354450.0 1187250.0 355650.0 ;
      RECT  1183500.0 369750.0 1184700.0 370950.0 ;
      RECT  1185900.0 359250.0 1187100.0 360450.0 ;
      RECT  1189800.0 357450.0 1191000.0 358650.0 ;
      RECT  1183200.0 376950.0 1184100.0 378750.0 ;
      RECT  1186200.0 376950.0 1187100.0 378750.0 ;
      RECT  1183200.0 353250.0 1184100.0 355050.0 ;
      RECT  1186200.0 353250.0 1187100.0 355050.0 ;
      RECT  1179600.0 353250.0 1180500.0 378750.0 ;
      RECT  1189800.0 353250.0 1190700.0 378750.0 ;
      RECT  1193400.0 361950.0 1194300.0 362850.0 ;
      RECT  1193850.0 361950.0 1194750.0 362850.0 ;
      RECT  1193400.0 355050.0 1194300.0 362400.0 ;
      RECT  1193850.0 361950.0 1194300.0 362850.0 ;
      RECT  1193850.0 362400.0 1194750.0 369750.0 ;
      RECT  1196400.0 368250.0 1197300.0 369150.0 ;
      RECT  1196250.0 368250.0 1197150.0 369150.0 ;
      RECT  1196400.0 368700.0 1197300.0 376950.0 ;
      RECT  1196700.0 368250.0 1196850.0 369150.0 ;
      RECT  1196250.0 360450.0 1197150.0 368700.0 ;
      RECT  1193250.0 376350.0 1194450.0 377550.0 ;
      RECT  1196250.0 354450.0 1197450.0 355650.0 ;
      RECT  1193700.0 369750.0 1194900.0 370950.0 ;
      RECT  1196100.0 359250.0 1197300.0 360450.0 ;
      RECT  1200000.0 357450.0 1201200.0 358650.0 ;
      RECT  1193400.0 376950.0 1194300.0 378750.0 ;
      RECT  1196400.0 376950.0 1197300.0 378750.0 ;
      RECT  1193400.0 353250.0 1194300.0 355050.0 ;
      RECT  1196400.0 353250.0 1197300.0 355050.0 ;
      RECT  1189800.0 353250.0 1190700.0 378750.0 ;
      RECT  1200000.0 353250.0 1200900.0 378750.0 ;
      RECT  1203600.0 361950.0 1204500.0 362850.0 ;
      RECT  1204050.0 361950.0 1204950.0 362850.0 ;
      RECT  1203600.0 355050.0 1204500.0 362400.0 ;
      RECT  1204050.0 361950.0 1204500.0 362850.0 ;
      RECT  1204050.0 362400.0 1204950.0 369750.0 ;
      RECT  1206600.0 368250.0 1207500.0 369150.0 ;
      RECT  1206450.0 368250.0 1207350.0 369150.0 ;
      RECT  1206600.0 368700.0 1207500.0 376950.0 ;
      RECT  1206900.0 368250.0 1207050.0 369150.0 ;
      RECT  1206450.0 360450.0 1207350.0 368700.0 ;
      RECT  1203450.0 376350.0 1204650.0 377550.0 ;
      RECT  1206450.0 354450.0 1207650.0 355650.0 ;
      RECT  1203900.0 369750.0 1205100.0 370950.0 ;
      RECT  1206300.0 359250.0 1207500.0 360450.0 ;
      RECT  1210200.0 357450.0 1211400.0 358650.0 ;
      RECT  1203600.0 376950.0 1204500.0 378750.0 ;
      RECT  1206600.0 376950.0 1207500.0 378750.0 ;
      RECT  1203600.0 353250.0 1204500.0 355050.0 ;
      RECT  1206600.0 353250.0 1207500.0 355050.0 ;
      RECT  1200000.0 353250.0 1200900.0 378750.0 ;
      RECT  1210200.0 353250.0 1211100.0 378750.0 ;
      RECT  1213800.0 361950.0 1214700.0 362850.0 ;
      RECT  1214250.0 361950.0 1215150.0 362850.0 ;
      RECT  1213800.0 355050.0 1214700.0 362400.0 ;
      RECT  1214250.0 361950.0 1214700.0 362850.0 ;
      RECT  1214250.0 362400.0 1215150.0 369750.0 ;
      RECT  1216800.0 368250.0 1217700.0 369150.0 ;
      RECT  1216650.0 368250.0 1217550.0 369150.0 ;
      RECT  1216800.0 368700.0 1217700.0 376950.0 ;
      RECT  1217100.0 368250.0 1217250.0 369150.0 ;
      RECT  1216650.0 360450.0 1217550.0 368700.0 ;
      RECT  1213650.0 376350.0 1214850.0 377550.0 ;
      RECT  1216650.0 354450.0 1217850.0 355650.0 ;
      RECT  1214100.0 369750.0 1215300.0 370950.0 ;
      RECT  1216500.0 359250.0 1217700.0 360450.0 ;
      RECT  1220400.0 357450.0 1221600.0 358650.0 ;
      RECT  1213800.0 376950.0 1214700.0 378750.0 ;
      RECT  1216800.0 376950.0 1217700.0 378750.0 ;
      RECT  1213800.0 353250.0 1214700.0 355050.0 ;
      RECT  1216800.0 353250.0 1217700.0 355050.0 ;
      RECT  1210200.0 353250.0 1211100.0 378750.0 ;
      RECT  1220400.0 353250.0 1221300.0 378750.0 ;
      RECT  1224000.0 361950.0 1224900.0 362850.0 ;
      RECT  1224450.0 361950.0 1225350.0 362850.0 ;
      RECT  1224000.0 355050.0 1224900.0 362400.0 ;
      RECT  1224450.0 361950.0 1224900.0 362850.0 ;
      RECT  1224450.0 362400.0 1225350.0 369750.0 ;
      RECT  1227000.0 368250.0 1227900.0 369150.0 ;
      RECT  1226850.0 368250.0 1227750.0 369150.0 ;
      RECT  1227000.0 368700.0 1227900.0 376950.0 ;
      RECT  1227300.0 368250.0 1227450.0 369150.0 ;
      RECT  1226850.0 360450.0 1227750.0 368700.0 ;
      RECT  1223850.0 376350.0 1225050.0 377550.0 ;
      RECT  1226850.0 354450.0 1228050.0 355650.0 ;
      RECT  1224300.0 369750.0 1225500.0 370950.0 ;
      RECT  1226700.0 359250.0 1227900.0 360450.0 ;
      RECT  1230600.0 357450.0 1231800.0 358650.0 ;
      RECT  1224000.0 376950.0 1224900.0 378750.0 ;
      RECT  1227000.0 376950.0 1227900.0 378750.0 ;
      RECT  1224000.0 353250.0 1224900.0 355050.0 ;
      RECT  1227000.0 353250.0 1227900.0 355050.0 ;
      RECT  1220400.0 353250.0 1221300.0 378750.0 ;
      RECT  1230600.0 353250.0 1231500.0 378750.0 ;
      RECT  1234200.0 361950.0 1235100.0 362850.0 ;
      RECT  1234650.0 361950.0 1235550.0 362850.0 ;
      RECT  1234200.0 355050.0 1235100.0 362400.0 ;
      RECT  1234650.0 361950.0 1235100.0 362850.0 ;
      RECT  1234650.0 362400.0 1235550.0 369750.0 ;
      RECT  1237200.0 368250.0 1238100.0 369150.0 ;
      RECT  1237050.0 368250.0 1237950.0 369150.0 ;
      RECT  1237200.0 368700.0 1238100.0 376950.0 ;
      RECT  1237500.0 368250.0 1237650.0 369150.0 ;
      RECT  1237050.0 360450.0 1237950.0 368700.0 ;
      RECT  1234050.0 376350.0 1235250.0 377550.0 ;
      RECT  1237050.0 354450.0 1238250.0 355650.0 ;
      RECT  1234500.0 369750.0 1235700.0 370950.0 ;
      RECT  1236900.0 359250.0 1238100.0 360450.0 ;
      RECT  1240800.0 357450.0 1242000.0 358650.0 ;
      RECT  1234200.0 376950.0 1235100.0 378750.0 ;
      RECT  1237200.0 376950.0 1238100.0 378750.0 ;
      RECT  1234200.0 353250.0 1235100.0 355050.0 ;
      RECT  1237200.0 353250.0 1238100.0 355050.0 ;
      RECT  1230600.0 353250.0 1231500.0 378750.0 ;
      RECT  1240800.0 353250.0 1241700.0 378750.0 ;
      RECT  1244400.0 361950.0 1245300.0 362850.0 ;
      RECT  1244850.0 361950.0 1245750.0 362850.0 ;
      RECT  1244400.0 355050.0 1245300.0 362400.0 ;
      RECT  1244850.0 361950.0 1245300.0 362850.0 ;
      RECT  1244850.0 362400.0 1245750.0 369750.0 ;
      RECT  1247400.0 368250.0 1248300.0 369150.0 ;
      RECT  1247250.0 368250.0 1248150.0 369150.0 ;
      RECT  1247400.0 368700.0 1248300.0 376950.0 ;
      RECT  1247700.0 368250.0 1247850.0 369150.0 ;
      RECT  1247250.0 360450.0 1248150.0 368700.0 ;
      RECT  1244250.0 376350.0 1245450.0 377550.0 ;
      RECT  1247250.0 354450.0 1248450.0 355650.0 ;
      RECT  1244700.0 369750.0 1245900.0 370950.0 ;
      RECT  1247100.0 359250.0 1248300.0 360450.0 ;
      RECT  1251000.0 357450.0 1252200.0 358650.0 ;
      RECT  1244400.0 376950.0 1245300.0 378750.0 ;
      RECT  1247400.0 376950.0 1248300.0 378750.0 ;
      RECT  1244400.0 353250.0 1245300.0 355050.0 ;
      RECT  1247400.0 353250.0 1248300.0 355050.0 ;
      RECT  1240800.0 353250.0 1241700.0 378750.0 ;
      RECT  1251000.0 353250.0 1251900.0 378750.0 ;
      RECT  1254600.0 361950.0 1255500.0 362850.0 ;
      RECT  1255050.0 361950.0 1255950.0 362850.0 ;
      RECT  1254600.0 355050.0 1255500.0 362400.0 ;
      RECT  1255050.0 361950.0 1255500.0 362850.0 ;
      RECT  1255050.0 362400.0 1255950.0 369750.0 ;
      RECT  1257600.0 368250.0 1258500.0 369150.0 ;
      RECT  1257450.0 368250.0 1258350.0 369150.0 ;
      RECT  1257600.0 368700.0 1258500.0 376950.0 ;
      RECT  1257900.0 368250.0 1258050.0 369150.0 ;
      RECT  1257450.0 360450.0 1258350.0 368700.0 ;
      RECT  1254450.0 376350.0 1255650.0 377550.0 ;
      RECT  1257450.0 354450.0 1258650.0 355650.0 ;
      RECT  1254900.0 369750.0 1256100.0 370950.0 ;
      RECT  1257300.0 359250.0 1258500.0 360450.0 ;
      RECT  1261200.0 357450.0 1262400.0 358650.0 ;
      RECT  1254600.0 376950.0 1255500.0 378750.0 ;
      RECT  1257600.0 376950.0 1258500.0 378750.0 ;
      RECT  1254600.0 353250.0 1255500.0 355050.0 ;
      RECT  1257600.0 353250.0 1258500.0 355050.0 ;
      RECT  1251000.0 353250.0 1251900.0 378750.0 ;
      RECT  1261200.0 353250.0 1262100.0 378750.0 ;
      RECT  1264800.0 361950.0 1265700.0 362850.0 ;
      RECT  1265250.0 361950.0 1266150.0 362850.0 ;
      RECT  1264800.0 355050.0 1265700.0 362400.0 ;
      RECT  1265250.0 361950.0 1265700.0 362850.0 ;
      RECT  1265250.0 362400.0 1266150.0 369750.0 ;
      RECT  1267800.0 368250.0 1268700.0 369150.0 ;
      RECT  1267650.0 368250.0 1268550.0 369150.0 ;
      RECT  1267800.0 368700.0 1268700.0 376950.0 ;
      RECT  1268100.0 368250.0 1268250.0 369150.0 ;
      RECT  1267650.0 360450.0 1268550.0 368700.0 ;
      RECT  1264650.0 376350.0 1265850.0 377550.0 ;
      RECT  1267650.0 354450.0 1268850.0 355650.0 ;
      RECT  1265100.0 369750.0 1266300.0 370950.0 ;
      RECT  1267500.0 359250.0 1268700.0 360450.0 ;
      RECT  1271400.0 357450.0 1272600.0 358650.0 ;
      RECT  1264800.0 376950.0 1265700.0 378750.0 ;
      RECT  1267800.0 376950.0 1268700.0 378750.0 ;
      RECT  1264800.0 353250.0 1265700.0 355050.0 ;
      RECT  1267800.0 353250.0 1268700.0 355050.0 ;
      RECT  1261200.0 353250.0 1262100.0 378750.0 ;
      RECT  1271400.0 353250.0 1272300.0 378750.0 ;
      RECT  1275000.0 361950.0 1275900.0 362850.0 ;
      RECT  1275450.0 361950.0 1276350.0 362850.0 ;
      RECT  1275000.0 355050.0 1275900.0 362400.0 ;
      RECT  1275450.0 361950.0 1275900.0 362850.0 ;
      RECT  1275450.0 362400.0 1276350.0 369750.0 ;
      RECT  1278000.0 368250.0 1278900.0 369150.0 ;
      RECT  1277850.0 368250.0 1278750.0 369150.0 ;
      RECT  1278000.0 368700.0 1278900.0 376950.0 ;
      RECT  1278300.0 368250.0 1278450.0 369150.0 ;
      RECT  1277850.0 360450.0 1278750.0 368700.0 ;
      RECT  1274850.0 376350.0 1276050.0 377550.0 ;
      RECT  1277850.0 354450.0 1279050.0 355650.0 ;
      RECT  1275300.0 369750.0 1276500.0 370950.0 ;
      RECT  1277700.0 359250.0 1278900.0 360450.0 ;
      RECT  1281600.0 357450.0 1282800.0 358650.0 ;
      RECT  1275000.0 376950.0 1275900.0 378750.0 ;
      RECT  1278000.0 376950.0 1278900.0 378750.0 ;
      RECT  1275000.0 353250.0 1275900.0 355050.0 ;
      RECT  1278000.0 353250.0 1278900.0 355050.0 ;
      RECT  1271400.0 353250.0 1272300.0 378750.0 ;
      RECT  1281600.0 353250.0 1282500.0 378750.0 ;
      RECT  1285200.0 361950.0 1286100.0 362850.0 ;
      RECT  1285650.0 361950.0 1286550.0 362850.0 ;
      RECT  1285200.0 355050.0 1286100.0 362400.0 ;
      RECT  1285650.0 361950.0 1286100.0 362850.0 ;
      RECT  1285650.0 362400.0 1286550.0 369750.0 ;
      RECT  1288200.0 368250.0 1289100.0 369150.0 ;
      RECT  1288050.0 368250.0 1288950.0 369150.0 ;
      RECT  1288200.0 368700.0 1289100.0 376950.0 ;
      RECT  1288500.0 368250.0 1288650.0 369150.0 ;
      RECT  1288050.0 360450.0 1288950.0 368700.0 ;
      RECT  1285050.0 376350.0 1286250.0 377550.0 ;
      RECT  1288050.0 354450.0 1289250.0 355650.0 ;
      RECT  1285500.0 369750.0 1286700.0 370950.0 ;
      RECT  1287900.0 359250.0 1289100.0 360450.0 ;
      RECT  1291800.0 357450.0 1293000.0 358650.0 ;
      RECT  1285200.0 376950.0 1286100.0 378750.0 ;
      RECT  1288200.0 376950.0 1289100.0 378750.0 ;
      RECT  1285200.0 353250.0 1286100.0 355050.0 ;
      RECT  1288200.0 353250.0 1289100.0 355050.0 ;
      RECT  1281600.0 353250.0 1282500.0 378750.0 ;
      RECT  1291800.0 353250.0 1292700.0 378750.0 ;
      RECT  1295400.0 361950.0 1296300.0 362850.0 ;
      RECT  1295850.0 361950.0 1296750.0 362850.0 ;
      RECT  1295400.0 355050.0 1296300.0 362400.0 ;
      RECT  1295850.0 361950.0 1296300.0 362850.0 ;
      RECT  1295850.0 362400.0 1296750.0 369750.0 ;
      RECT  1298400.0 368250.0 1299300.0 369150.0 ;
      RECT  1298250.0 368250.0 1299150.0 369150.0 ;
      RECT  1298400.0 368700.0 1299300.0 376950.0 ;
      RECT  1298700.0 368250.0 1298850.0 369150.0 ;
      RECT  1298250.0 360450.0 1299150.0 368700.0 ;
      RECT  1295250.0 376350.0 1296450.0 377550.0 ;
      RECT  1298250.0 354450.0 1299450.0 355650.0 ;
      RECT  1295700.0 369750.0 1296900.0 370950.0 ;
      RECT  1298100.0 359250.0 1299300.0 360450.0 ;
      RECT  1302000.0 357450.0 1303200.0 358650.0 ;
      RECT  1295400.0 376950.0 1296300.0 378750.0 ;
      RECT  1298400.0 376950.0 1299300.0 378750.0 ;
      RECT  1295400.0 353250.0 1296300.0 355050.0 ;
      RECT  1298400.0 353250.0 1299300.0 355050.0 ;
      RECT  1291800.0 353250.0 1292700.0 378750.0 ;
      RECT  1302000.0 353250.0 1302900.0 378750.0 ;
      RECT  1305600.0 361950.0 1306500.0 362850.0 ;
      RECT  1306050.0 361950.0 1306950.0 362850.0 ;
      RECT  1305600.0 355050.0 1306500.0 362400.0 ;
      RECT  1306050.0 361950.0 1306500.0 362850.0 ;
      RECT  1306050.0 362400.0 1306950.0 369750.0 ;
      RECT  1308600.0 368250.0 1309500.0 369150.0 ;
      RECT  1308450.0 368250.0 1309350.0 369150.0 ;
      RECT  1308600.0 368700.0 1309500.0 376950.0 ;
      RECT  1308900.0 368250.0 1309050.0 369150.0 ;
      RECT  1308450.0 360450.0 1309350.0 368700.0 ;
      RECT  1305450.0 376350.0 1306650.0 377550.0 ;
      RECT  1308450.0 354450.0 1309650.0 355650.0 ;
      RECT  1305900.0 369750.0 1307100.0 370950.0 ;
      RECT  1308300.0 359250.0 1309500.0 360450.0 ;
      RECT  1312200.0 357450.0 1313400.0 358650.0 ;
      RECT  1305600.0 376950.0 1306500.0 378750.0 ;
      RECT  1308600.0 376950.0 1309500.0 378750.0 ;
      RECT  1305600.0 353250.0 1306500.0 355050.0 ;
      RECT  1308600.0 353250.0 1309500.0 355050.0 ;
      RECT  1302000.0 353250.0 1302900.0 378750.0 ;
      RECT  1312200.0 353250.0 1313100.0 378750.0 ;
      RECT  1315800.0 361950.0 1316700.0 362850.0 ;
      RECT  1316250.0 361950.0 1317150.0 362850.0 ;
      RECT  1315800.0 355050.0 1316700.0 362400.0 ;
      RECT  1316250.0 361950.0 1316700.0 362850.0 ;
      RECT  1316250.0 362400.0 1317150.0 369750.0 ;
      RECT  1318800.0 368250.0 1319700.0 369150.0 ;
      RECT  1318650.0 368250.0 1319550.0 369150.0 ;
      RECT  1318800.0 368700.0 1319700.0 376950.0 ;
      RECT  1319100.0 368250.0 1319250.0 369150.0 ;
      RECT  1318650.0 360450.0 1319550.0 368700.0 ;
      RECT  1315650.0 376350.0 1316850.0 377550.0 ;
      RECT  1318650.0 354450.0 1319850.0 355650.0 ;
      RECT  1316100.0 369750.0 1317300.0 370950.0 ;
      RECT  1318500.0 359250.0 1319700.0 360450.0 ;
      RECT  1322400.0 357450.0 1323600.0 358650.0 ;
      RECT  1315800.0 376950.0 1316700.0 378750.0 ;
      RECT  1318800.0 376950.0 1319700.0 378750.0 ;
      RECT  1315800.0 353250.0 1316700.0 355050.0 ;
      RECT  1318800.0 353250.0 1319700.0 355050.0 ;
      RECT  1312200.0 353250.0 1313100.0 378750.0 ;
      RECT  1322400.0 353250.0 1323300.0 378750.0 ;
      RECT  1326000.0 361950.0 1326900.0 362850.0 ;
      RECT  1326450.0 361950.0 1327350.0 362850.0 ;
      RECT  1326000.0 355050.0 1326900.0 362400.0 ;
      RECT  1326450.0 361950.0 1326900.0 362850.0 ;
      RECT  1326450.0 362400.0 1327350.0 369750.0 ;
      RECT  1329000.0 368250.0 1329900.0 369150.0 ;
      RECT  1328850.0 368250.0 1329750.0 369150.0 ;
      RECT  1329000.0 368700.0 1329900.0 376950.0 ;
      RECT  1329300.0 368250.0 1329450.0 369150.0 ;
      RECT  1328850.0 360450.0 1329750.0 368700.0 ;
      RECT  1325850.0 376350.0 1327050.0 377550.0 ;
      RECT  1328850.0 354450.0 1330050.0 355650.0 ;
      RECT  1326300.0 369750.0 1327500.0 370950.0 ;
      RECT  1328700.0 359250.0 1329900.0 360450.0 ;
      RECT  1332600.0 357450.0 1333800.0 358650.0 ;
      RECT  1326000.0 376950.0 1326900.0 378750.0 ;
      RECT  1329000.0 376950.0 1329900.0 378750.0 ;
      RECT  1326000.0 353250.0 1326900.0 355050.0 ;
      RECT  1329000.0 353250.0 1329900.0 355050.0 ;
      RECT  1322400.0 353250.0 1323300.0 378750.0 ;
      RECT  1332600.0 353250.0 1333500.0 378750.0 ;
      RECT  1336200.0 361950.0 1337100.0 362850.0 ;
      RECT  1336650.0 361950.0 1337550.0 362850.0 ;
      RECT  1336200.0 355050.0 1337100.0 362400.0 ;
      RECT  1336650.0 361950.0 1337100.0 362850.0 ;
      RECT  1336650.0 362400.0 1337550.0 369750.0 ;
      RECT  1339200.0 368250.0 1340100.0 369150.0 ;
      RECT  1339050.0 368250.0 1339950.0 369150.0 ;
      RECT  1339200.0 368700.0 1340100.0 376950.0 ;
      RECT  1339500.0 368250.0 1339650.0 369150.0 ;
      RECT  1339050.0 360450.0 1339950.0 368700.0 ;
      RECT  1336050.0 376350.0 1337250.0 377550.0 ;
      RECT  1339050.0 354450.0 1340250.0 355650.0 ;
      RECT  1336500.0 369750.0 1337700.0 370950.0 ;
      RECT  1338900.0 359250.0 1340100.0 360450.0 ;
      RECT  1342800.0 357450.0 1344000.0 358650.0 ;
      RECT  1336200.0 376950.0 1337100.0 378750.0 ;
      RECT  1339200.0 376950.0 1340100.0 378750.0 ;
      RECT  1336200.0 353250.0 1337100.0 355050.0 ;
      RECT  1339200.0 353250.0 1340100.0 355050.0 ;
      RECT  1332600.0 353250.0 1333500.0 378750.0 ;
      RECT  1342800.0 353250.0 1343700.0 378750.0 ;
      RECT  1346400.0 361950.0 1347300.0 362850.0 ;
      RECT  1346850.0 361950.0 1347750.0 362850.0 ;
      RECT  1346400.0 355050.0 1347300.0 362400.0 ;
      RECT  1346850.0 361950.0 1347300.0 362850.0 ;
      RECT  1346850.0 362400.0 1347750.0 369750.0 ;
      RECT  1349400.0 368250.0 1350300.0 369150.0 ;
      RECT  1349250.0 368250.0 1350150.0 369150.0 ;
      RECT  1349400.0 368700.0 1350300.0 376950.0 ;
      RECT  1349700.0 368250.0 1349850.0 369150.0 ;
      RECT  1349250.0 360450.0 1350150.0 368700.0 ;
      RECT  1346250.0 376350.0 1347450.0 377550.0 ;
      RECT  1349250.0 354450.0 1350450.0 355650.0 ;
      RECT  1346700.0 369750.0 1347900.0 370950.0 ;
      RECT  1349100.0 359250.0 1350300.0 360450.0 ;
      RECT  1353000.0 357450.0 1354200.0 358650.0 ;
      RECT  1346400.0 376950.0 1347300.0 378750.0 ;
      RECT  1349400.0 376950.0 1350300.0 378750.0 ;
      RECT  1346400.0 353250.0 1347300.0 355050.0 ;
      RECT  1349400.0 353250.0 1350300.0 355050.0 ;
      RECT  1342800.0 353250.0 1343700.0 378750.0 ;
      RECT  1353000.0 353250.0 1353900.0 378750.0 ;
      RECT  1356600.0 361950.0 1357500.0 362850.0 ;
      RECT  1357050.0 361950.0 1357950.0 362850.0 ;
      RECT  1356600.0 355050.0 1357500.0 362400.0 ;
      RECT  1357050.0 361950.0 1357500.0 362850.0 ;
      RECT  1357050.0 362400.0 1357950.0 369750.0 ;
      RECT  1359600.0 368250.0 1360500.0 369150.0 ;
      RECT  1359450.0 368250.0 1360350.0 369150.0 ;
      RECT  1359600.0 368700.0 1360500.0 376950.0 ;
      RECT  1359900.0 368250.0 1360050.0 369150.0 ;
      RECT  1359450.0 360450.0 1360350.0 368700.0 ;
      RECT  1356450.0 376350.0 1357650.0 377550.0 ;
      RECT  1359450.0 354450.0 1360650.0 355650.0 ;
      RECT  1356900.0 369750.0 1358100.0 370950.0 ;
      RECT  1359300.0 359250.0 1360500.0 360450.0 ;
      RECT  1363200.0 357450.0 1364400.0 358650.0 ;
      RECT  1356600.0 376950.0 1357500.0 378750.0 ;
      RECT  1359600.0 376950.0 1360500.0 378750.0 ;
      RECT  1356600.0 353250.0 1357500.0 355050.0 ;
      RECT  1359600.0 353250.0 1360500.0 355050.0 ;
      RECT  1353000.0 353250.0 1353900.0 378750.0 ;
      RECT  1363200.0 353250.0 1364100.0 378750.0 ;
      RECT  1366800.0 361950.0 1367700.0 362850.0 ;
      RECT  1367250.0 361950.0 1368150.0 362850.0 ;
      RECT  1366800.0 355050.0 1367700.0 362400.0 ;
      RECT  1367250.0 361950.0 1367700.0 362850.0 ;
      RECT  1367250.0 362400.0 1368150.0 369750.0 ;
      RECT  1369800.0 368250.0 1370700.0 369150.0 ;
      RECT  1369650.0 368250.0 1370550.0 369150.0 ;
      RECT  1369800.0 368700.0 1370700.0 376950.0 ;
      RECT  1370100.0 368250.0 1370250.0 369150.0 ;
      RECT  1369650.0 360450.0 1370550.0 368700.0 ;
      RECT  1366650.0 376350.0 1367850.0 377550.0 ;
      RECT  1369650.0 354450.0 1370850.0 355650.0 ;
      RECT  1367100.0 369750.0 1368300.0 370950.0 ;
      RECT  1369500.0 359250.0 1370700.0 360450.0 ;
      RECT  1373400.0 357450.0 1374600.0 358650.0 ;
      RECT  1366800.0 376950.0 1367700.0 378750.0 ;
      RECT  1369800.0 376950.0 1370700.0 378750.0 ;
      RECT  1366800.0 353250.0 1367700.0 355050.0 ;
      RECT  1369800.0 353250.0 1370700.0 355050.0 ;
      RECT  1363200.0 353250.0 1364100.0 378750.0 ;
      RECT  1373400.0 353250.0 1374300.0 378750.0 ;
      RECT  1377000.0 361950.0 1377900.0 362850.0 ;
      RECT  1377450.0 361950.0 1378350.0 362850.0 ;
      RECT  1377000.0 355050.0 1377900.0 362400.0 ;
      RECT  1377450.0 361950.0 1377900.0 362850.0 ;
      RECT  1377450.0 362400.0 1378350.0 369750.0 ;
      RECT  1380000.0 368250.0 1380900.0 369150.0 ;
      RECT  1379850.0 368250.0 1380750.0 369150.0 ;
      RECT  1380000.0 368700.0 1380900.0 376950.0 ;
      RECT  1380300.0 368250.0 1380450.0 369150.0 ;
      RECT  1379850.0 360450.0 1380750.0 368700.0 ;
      RECT  1376850.0 376350.0 1378050.0 377550.0 ;
      RECT  1379850.0 354450.0 1381050.0 355650.0 ;
      RECT  1377300.0 369750.0 1378500.0 370950.0 ;
      RECT  1379700.0 359250.0 1380900.0 360450.0 ;
      RECT  1383600.0 357450.0 1384800.0 358650.0 ;
      RECT  1377000.0 376950.0 1377900.0 378750.0 ;
      RECT  1380000.0 376950.0 1380900.0 378750.0 ;
      RECT  1377000.0 353250.0 1377900.0 355050.0 ;
      RECT  1380000.0 353250.0 1380900.0 355050.0 ;
      RECT  1373400.0 353250.0 1374300.0 378750.0 ;
      RECT  1383600.0 353250.0 1384500.0 378750.0 ;
      RECT  1387200.0 361950.0 1388100.0 362850.0 ;
      RECT  1387650.0 361950.0 1388550.0 362850.0 ;
      RECT  1387200.0 355050.0 1388100.0 362400.0 ;
      RECT  1387650.0 361950.0 1388100.0 362850.0 ;
      RECT  1387650.0 362400.0 1388550.0 369750.0 ;
      RECT  1390200.0 368250.0 1391100.0 369150.0 ;
      RECT  1390050.0 368250.0 1390950.0 369150.0 ;
      RECT  1390200.0 368700.0 1391100.0 376950.0 ;
      RECT  1390500.0 368250.0 1390650.0 369150.0 ;
      RECT  1390050.0 360450.0 1390950.0 368700.0 ;
      RECT  1387050.0 376350.0 1388250.0 377550.0 ;
      RECT  1390050.0 354450.0 1391250.0 355650.0 ;
      RECT  1387500.0 369750.0 1388700.0 370950.0 ;
      RECT  1389900.0 359250.0 1391100.0 360450.0 ;
      RECT  1393800.0 357450.0 1395000.0 358650.0 ;
      RECT  1387200.0 376950.0 1388100.0 378750.0 ;
      RECT  1390200.0 376950.0 1391100.0 378750.0 ;
      RECT  1387200.0 353250.0 1388100.0 355050.0 ;
      RECT  1390200.0 353250.0 1391100.0 355050.0 ;
      RECT  1383600.0 353250.0 1384500.0 378750.0 ;
      RECT  1393800.0 353250.0 1394700.0 378750.0 ;
      RECT  1397400.0 361950.0 1398300.0 362850.0 ;
      RECT  1397850.0 361950.0 1398750.0 362850.0 ;
      RECT  1397400.0 355050.0 1398300.0 362400.0 ;
      RECT  1397850.0 361950.0 1398300.0 362850.0 ;
      RECT  1397850.0 362400.0 1398750.0 369750.0 ;
      RECT  1400400.0 368250.0 1401300.0 369150.0 ;
      RECT  1400250.0 368250.0 1401150.0 369150.0 ;
      RECT  1400400.0 368700.0 1401300.0 376950.0 ;
      RECT  1400700.0 368250.0 1400850.0 369150.0 ;
      RECT  1400250.0 360450.0 1401150.0 368700.0 ;
      RECT  1397250.0 376350.0 1398450.0 377550.0 ;
      RECT  1400250.0 354450.0 1401450.0 355650.0 ;
      RECT  1397700.0 369750.0 1398900.0 370950.0 ;
      RECT  1400100.0 359250.0 1401300.0 360450.0 ;
      RECT  1404000.0 357450.0 1405200.0 358650.0 ;
      RECT  1397400.0 376950.0 1398300.0 378750.0 ;
      RECT  1400400.0 376950.0 1401300.0 378750.0 ;
      RECT  1397400.0 353250.0 1398300.0 355050.0 ;
      RECT  1400400.0 353250.0 1401300.0 355050.0 ;
      RECT  1393800.0 353250.0 1394700.0 378750.0 ;
      RECT  1404000.0 353250.0 1404900.0 378750.0 ;
      RECT  1407600.0 361950.0 1408500.0 362850.0 ;
      RECT  1408050.0 361950.0 1408950.0 362850.0 ;
      RECT  1407600.0 355050.0 1408500.0 362400.0 ;
      RECT  1408050.0 361950.0 1408500.0 362850.0 ;
      RECT  1408050.0 362400.0 1408950.0 369750.0 ;
      RECT  1410600.0 368250.0 1411500.0 369150.0 ;
      RECT  1410450.0 368250.0 1411350.0 369150.0 ;
      RECT  1410600.0 368700.0 1411500.0 376950.0 ;
      RECT  1410900.0 368250.0 1411050.0 369150.0 ;
      RECT  1410450.0 360450.0 1411350.0 368700.0 ;
      RECT  1407450.0 376350.0 1408650.0 377550.0 ;
      RECT  1410450.0 354450.0 1411650.0 355650.0 ;
      RECT  1407900.0 369750.0 1409100.0 370950.0 ;
      RECT  1410300.0 359250.0 1411500.0 360450.0 ;
      RECT  1414200.0 357450.0 1415400.0 358650.0 ;
      RECT  1407600.0 376950.0 1408500.0 378750.0 ;
      RECT  1410600.0 376950.0 1411500.0 378750.0 ;
      RECT  1407600.0 353250.0 1408500.0 355050.0 ;
      RECT  1410600.0 353250.0 1411500.0 355050.0 ;
      RECT  1404000.0 353250.0 1404900.0 378750.0 ;
      RECT  1414200.0 353250.0 1415100.0 378750.0 ;
      RECT  1417800.0 361950.0 1418700.0 362850.0 ;
      RECT  1418250.0 361950.0 1419150.0 362850.0 ;
      RECT  1417800.0 355050.0 1418700.0 362400.0 ;
      RECT  1418250.0 361950.0 1418700.0 362850.0 ;
      RECT  1418250.0 362400.0 1419150.0 369750.0 ;
      RECT  1420800.0 368250.0 1421700.0 369150.0 ;
      RECT  1420650.0 368250.0 1421550.0 369150.0 ;
      RECT  1420800.0 368700.0 1421700.0 376950.0 ;
      RECT  1421100.0 368250.0 1421250.0 369150.0 ;
      RECT  1420650.0 360450.0 1421550.0 368700.0 ;
      RECT  1417650.0 376350.0 1418850.0 377550.0 ;
      RECT  1420650.0 354450.0 1421850.0 355650.0 ;
      RECT  1418100.0 369750.0 1419300.0 370950.0 ;
      RECT  1420500.0 359250.0 1421700.0 360450.0 ;
      RECT  1424400.0 357450.0 1425600.0 358650.0 ;
      RECT  1417800.0 376950.0 1418700.0 378750.0 ;
      RECT  1420800.0 376950.0 1421700.0 378750.0 ;
      RECT  1417800.0 353250.0 1418700.0 355050.0 ;
      RECT  1420800.0 353250.0 1421700.0 355050.0 ;
      RECT  1414200.0 353250.0 1415100.0 378750.0 ;
      RECT  1424400.0 353250.0 1425300.0 378750.0 ;
      RECT  1428000.0 361950.0 1428900.0 362850.0 ;
      RECT  1428450.0 361950.0 1429350.0 362850.0 ;
      RECT  1428000.0 355050.0 1428900.0 362400.0 ;
      RECT  1428450.0 361950.0 1428900.0 362850.0 ;
      RECT  1428450.0 362400.0 1429350.0 369750.0 ;
      RECT  1431000.0 368250.0 1431900.0 369150.0 ;
      RECT  1430850.0 368250.0 1431750.0 369150.0 ;
      RECT  1431000.0 368700.0 1431900.0 376950.0 ;
      RECT  1431300.0 368250.0 1431450.0 369150.0 ;
      RECT  1430850.0 360450.0 1431750.0 368700.0 ;
      RECT  1427850.0 376350.0 1429050.0 377550.0 ;
      RECT  1430850.0 354450.0 1432050.0 355650.0 ;
      RECT  1428300.0 369750.0 1429500.0 370950.0 ;
      RECT  1430700.0 359250.0 1431900.0 360450.0 ;
      RECT  1434600.0 357450.0 1435800.0 358650.0 ;
      RECT  1428000.0 376950.0 1428900.0 378750.0 ;
      RECT  1431000.0 376950.0 1431900.0 378750.0 ;
      RECT  1428000.0 353250.0 1428900.0 355050.0 ;
      RECT  1431000.0 353250.0 1431900.0 355050.0 ;
      RECT  1424400.0 353250.0 1425300.0 378750.0 ;
      RECT  1434600.0 353250.0 1435500.0 378750.0 ;
      RECT  1438200.0 361950.0 1439100.0 362850.0 ;
      RECT  1438650.0 361950.0 1439550.0 362850.0 ;
      RECT  1438200.0 355050.0 1439100.0 362400.0 ;
      RECT  1438650.0 361950.0 1439100.0 362850.0 ;
      RECT  1438650.0 362400.0 1439550.0 369750.0 ;
      RECT  1441200.0 368250.0 1442100.0 369150.0 ;
      RECT  1441050.0 368250.0 1441950.0 369150.0 ;
      RECT  1441200.0 368700.0 1442100.0 376950.0 ;
      RECT  1441500.0 368250.0 1441650.0 369150.0 ;
      RECT  1441050.0 360450.0 1441950.0 368700.0 ;
      RECT  1438050.0 376350.0 1439250.0 377550.0 ;
      RECT  1441050.0 354450.0 1442250.0 355650.0 ;
      RECT  1438500.0 369750.0 1439700.0 370950.0 ;
      RECT  1440900.0 359250.0 1442100.0 360450.0 ;
      RECT  1444800.0 357450.0 1446000.0 358650.0 ;
      RECT  1438200.0 376950.0 1439100.0 378750.0 ;
      RECT  1441200.0 376950.0 1442100.0 378750.0 ;
      RECT  1438200.0 353250.0 1439100.0 355050.0 ;
      RECT  1441200.0 353250.0 1442100.0 355050.0 ;
      RECT  1434600.0 353250.0 1435500.0 378750.0 ;
      RECT  1444800.0 353250.0 1445700.0 378750.0 ;
      RECT  1448400.0 361950.0 1449300.0 362850.0 ;
      RECT  1448850.0 361950.0 1449750.0 362850.0 ;
      RECT  1448400.0 355050.0 1449300.0 362400.0 ;
      RECT  1448850.0 361950.0 1449300.0 362850.0 ;
      RECT  1448850.0 362400.0 1449750.0 369750.0 ;
      RECT  1451400.0 368250.0 1452300.0 369150.0 ;
      RECT  1451250.0 368250.0 1452150.0 369150.0 ;
      RECT  1451400.0 368700.0 1452300.0 376950.0 ;
      RECT  1451700.0 368250.0 1451850.0 369150.0 ;
      RECT  1451250.0 360450.0 1452150.0 368700.0 ;
      RECT  1448250.0 376350.0 1449450.0 377550.0 ;
      RECT  1451250.0 354450.0 1452450.0 355650.0 ;
      RECT  1448700.0 369750.0 1449900.0 370950.0 ;
      RECT  1451100.0 359250.0 1452300.0 360450.0 ;
      RECT  1455000.0 357450.0 1456200.0 358650.0 ;
      RECT  1448400.0 376950.0 1449300.0 378750.0 ;
      RECT  1451400.0 376950.0 1452300.0 378750.0 ;
      RECT  1448400.0 353250.0 1449300.0 355050.0 ;
      RECT  1451400.0 353250.0 1452300.0 355050.0 ;
      RECT  1444800.0 353250.0 1445700.0 378750.0 ;
      RECT  1455000.0 353250.0 1455900.0 378750.0 ;
      RECT  1458600.0 361950.0 1459500.0 362850.0 ;
      RECT  1459050.0 361950.0 1459950.0 362850.0 ;
      RECT  1458600.0 355050.0 1459500.0 362400.0 ;
      RECT  1459050.0 361950.0 1459500.0 362850.0 ;
      RECT  1459050.0 362400.0 1459950.0 369750.0 ;
      RECT  1461600.0 368250.0 1462500.0 369150.0 ;
      RECT  1461450.0 368250.0 1462350.0 369150.0 ;
      RECT  1461600.0 368700.0 1462500.0 376950.0 ;
      RECT  1461900.0 368250.0 1462050.0 369150.0 ;
      RECT  1461450.0 360450.0 1462350.0 368700.0 ;
      RECT  1458450.0 376350.0 1459650.0 377550.0 ;
      RECT  1461450.0 354450.0 1462650.0 355650.0 ;
      RECT  1458900.0 369750.0 1460100.0 370950.0 ;
      RECT  1461300.0 359250.0 1462500.0 360450.0 ;
      RECT  1465200.0 357450.0 1466400.0 358650.0 ;
      RECT  1458600.0 376950.0 1459500.0 378750.0 ;
      RECT  1461600.0 376950.0 1462500.0 378750.0 ;
      RECT  1458600.0 353250.0 1459500.0 355050.0 ;
      RECT  1461600.0 353250.0 1462500.0 355050.0 ;
      RECT  1455000.0 353250.0 1455900.0 378750.0 ;
      RECT  1465200.0 353250.0 1466100.0 378750.0 ;
      RECT  1468800.0 361950.0 1469700.0 362850.0 ;
      RECT  1469250.0 361950.0 1470150.0 362850.0 ;
      RECT  1468800.0 355050.0 1469700.0 362400.0 ;
      RECT  1469250.0 361950.0 1469700.0 362850.0 ;
      RECT  1469250.0 362400.0 1470150.0 369750.0 ;
      RECT  1471800.0 368250.0 1472700.0 369150.0 ;
      RECT  1471650.0 368250.0 1472550.0 369150.0 ;
      RECT  1471800.0 368700.0 1472700.0 376950.0 ;
      RECT  1472100.0 368250.0 1472250.0 369150.0 ;
      RECT  1471650.0 360450.0 1472550.0 368700.0 ;
      RECT  1468650.0 376350.0 1469850.0 377550.0 ;
      RECT  1471650.0 354450.0 1472850.0 355650.0 ;
      RECT  1469100.0 369750.0 1470300.0 370950.0 ;
      RECT  1471500.0 359250.0 1472700.0 360450.0 ;
      RECT  1475400.0 357450.0 1476600.0 358650.0 ;
      RECT  1468800.0 376950.0 1469700.0 378750.0 ;
      RECT  1471800.0 376950.0 1472700.0 378750.0 ;
      RECT  1468800.0 353250.0 1469700.0 355050.0 ;
      RECT  1471800.0 353250.0 1472700.0 355050.0 ;
      RECT  1465200.0 353250.0 1466100.0 378750.0 ;
      RECT  1475400.0 353250.0 1476300.0 378750.0 ;
      RECT  1479000.0 361950.0 1479900.0 362850.0 ;
      RECT  1479450.0 361950.0 1480350.0 362850.0 ;
      RECT  1479000.0 355050.0 1479900.0 362400.0 ;
      RECT  1479450.0 361950.0 1479900.0 362850.0 ;
      RECT  1479450.0 362400.0 1480350.0 369750.0 ;
      RECT  1482000.0 368250.0 1482900.0 369150.0 ;
      RECT  1481850.0 368250.0 1482750.0 369150.0 ;
      RECT  1482000.0 368700.0 1482900.0 376950.0 ;
      RECT  1482300.0 368250.0 1482450.0 369150.0 ;
      RECT  1481850.0 360450.0 1482750.0 368700.0 ;
      RECT  1478850.0 376350.0 1480050.0 377550.0 ;
      RECT  1481850.0 354450.0 1483050.0 355650.0 ;
      RECT  1479300.0 369750.0 1480500.0 370950.0 ;
      RECT  1481700.0 359250.0 1482900.0 360450.0 ;
      RECT  1485600.0 357450.0 1486800.0 358650.0 ;
      RECT  1479000.0 376950.0 1479900.0 378750.0 ;
      RECT  1482000.0 376950.0 1482900.0 378750.0 ;
      RECT  1479000.0 353250.0 1479900.0 355050.0 ;
      RECT  1482000.0 353250.0 1482900.0 355050.0 ;
      RECT  1475400.0 353250.0 1476300.0 378750.0 ;
      RECT  1485600.0 353250.0 1486500.0 378750.0 ;
      RECT  1489200.0 361950.0 1490100.0 362850.0 ;
      RECT  1489650.0 361950.0 1490550.0 362850.0 ;
      RECT  1489200.0 355050.0 1490100.0 362400.0 ;
      RECT  1489650.0 361950.0 1490100.0 362850.0 ;
      RECT  1489650.0 362400.0 1490550.0 369750.0 ;
      RECT  1492200.0 368250.0 1493100.0 369150.0 ;
      RECT  1492050.0 368250.0 1492950.0 369150.0 ;
      RECT  1492200.0 368700.0 1493100.0 376950.0 ;
      RECT  1492500.0 368250.0 1492650.0 369150.0 ;
      RECT  1492050.0 360450.0 1492950.0 368700.0 ;
      RECT  1489050.0 376350.0 1490250.0 377550.0 ;
      RECT  1492050.0 354450.0 1493250.0 355650.0 ;
      RECT  1489500.0 369750.0 1490700.0 370950.0 ;
      RECT  1491900.0 359250.0 1493100.0 360450.0 ;
      RECT  1495800.0 357450.0 1497000.0 358650.0 ;
      RECT  1489200.0 376950.0 1490100.0 378750.0 ;
      RECT  1492200.0 376950.0 1493100.0 378750.0 ;
      RECT  1489200.0 353250.0 1490100.0 355050.0 ;
      RECT  1492200.0 353250.0 1493100.0 355050.0 ;
      RECT  1485600.0 353250.0 1486500.0 378750.0 ;
      RECT  1495800.0 353250.0 1496700.0 378750.0 ;
      RECT  1499400.0 361950.0 1500300.0 362850.0 ;
      RECT  1499850.0 361950.0 1500750.0 362850.0 ;
      RECT  1499400.0 355050.0 1500300.0 362400.0 ;
      RECT  1499850.0 361950.0 1500300.0 362850.0 ;
      RECT  1499850.0 362400.0 1500750.0 369750.0 ;
      RECT  1502400.0 368250.0 1503300.0 369150.0 ;
      RECT  1502250.0 368250.0 1503150.0 369150.0 ;
      RECT  1502400.0 368700.0 1503300.0 376950.0 ;
      RECT  1502700.0 368250.0 1502850.0 369150.0 ;
      RECT  1502250.0 360450.0 1503150.0 368700.0 ;
      RECT  1499250.0 376350.0 1500450.0 377550.0 ;
      RECT  1502250.0 354450.0 1503450.0 355650.0 ;
      RECT  1499700.0 369750.0 1500900.0 370950.0 ;
      RECT  1502100.0 359250.0 1503300.0 360450.0 ;
      RECT  1506000.0 357450.0 1507200.0 358650.0 ;
      RECT  1499400.0 376950.0 1500300.0 378750.0 ;
      RECT  1502400.0 376950.0 1503300.0 378750.0 ;
      RECT  1499400.0 353250.0 1500300.0 355050.0 ;
      RECT  1502400.0 353250.0 1503300.0 355050.0 ;
      RECT  1495800.0 353250.0 1496700.0 378750.0 ;
      RECT  1506000.0 353250.0 1506900.0 378750.0 ;
      RECT  1509600.0 361950.0 1510500.0 362850.0 ;
      RECT  1510050.0 361950.0 1510950.0 362850.0 ;
      RECT  1509600.0 355050.0 1510500.0 362400.0 ;
      RECT  1510050.0 361950.0 1510500.0 362850.0 ;
      RECT  1510050.0 362400.0 1510950.0 369750.0 ;
      RECT  1512600.0 368250.0 1513500.0 369150.0 ;
      RECT  1512450.0 368250.0 1513350.0 369150.0 ;
      RECT  1512600.0 368700.0 1513500.0 376950.0 ;
      RECT  1512900.0 368250.0 1513050.0 369150.0 ;
      RECT  1512450.0 360450.0 1513350.0 368700.0 ;
      RECT  1509450.0 376350.0 1510650.0 377550.0 ;
      RECT  1512450.0 354450.0 1513650.0 355650.0 ;
      RECT  1509900.0 369750.0 1511100.0 370950.0 ;
      RECT  1512300.0 359250.0 1513500.0 360450.0 ;
      RECT  1516200.0 357450.0 1517400.0 358650.0 ;
      RECT  1509600.0 376950.0 1510500.0 378750.0 ;
      RECT  1512600.0 376950.0 1513500.0 378750.0 ;
      RECT  1509600.0 353250.0 1510500.0 355050.0 ;
      RECT  1512600.0 353250.0 1513500.0 355050.0 ;
      RECT  1506000.0 353250.0 1506900.0 378750.0 ;
      RECT  1516200.0 353250.0 1517100.0 378750.0 ;
      RECT  1519800.0 361950.0 1520700.0 362850.0 ;
      RECT  1520250.0 361950.0 1521150.0 362850.0 ;
      RECT  1519800.0 355050.0 1520700.0 362400.0 ;
      RECT  1520250.0 361950.0 1520700.0 362850.0 ;
      RECT  1520250.0 362400.0 1521150.0 369750.0 ;
      RECT  1522800.0 368250.0 1523700.0 369150.0 ;
      RECT  1522650.0 368250.0 1523550.0 369150.0 ;
      RECT  1522800.0 368700.0 1523700.0 376950.0 ;
      RECT  1523100.0 368250.0 1523250.0 369150.0 ;
      RECT  1522650.0 360450.0 1523550.0 368700.0 ;
      RECT  1519650.0 376350.0 1520850.0 377550.0 ;
      RECT  1522650.0 354450.0 1523850.0 355650.0 ;
      RECT  1520100.0 369750.0 1521300.0 370950.0 ;
      RECT  1522500.0 359250.0 1523700.0 360450.0 ;
      RECT  1526400.0 357450.0 1527600.0 358650.0 ;
      RECT  1519800.0 376950.0 1520700.0 378750.0 ;
      RECT  1522800.0 376950.0 1523700.0 378750.0 ;
      RECT  1519800.0 353250.0 1520700.0 355050.0 ;
      RECT  1522800.0 353250.0 1523700.0 355050.0 ;
      RECT  1516200.0 353250.0 1517100.0 378750.0 ;
      RECT  1526400.0 353250.0 1527300.0 378750.0 ;
      RECT  225600.0 342750.0 224400.0 343950.0 ;
      RECT  227400.0 340650.0 226200.0 341850.0 ;
      RECT  235800.0 342750.0 234600.0 343950.0 ;
      RECT  237600.0 340650.0 236400.0 341850.0 ;
      RECT  246000.0 342750.0 244800.0 343950.0 ;
      RECT  247800.0 340650.0 246600.0 341850.0 ;
      RECT  256200.0 342750.0 255000.0 343950.0 ;
      RECT  258000.0 340650.0 256800.0 341850.0 ;
      RECT  266400.0 342750.0 265200.0 343950.0 ;
      RECT  268200.0 340650.0 267000.0 341850.0 ;
      RECT  276600.0 342750.0 275400.0 343950.0 ;
      RECT  278400.0 340650.0 277200.0 341850.0 ;
      RECT  286800.0 342750.0 285600.0 343950.0 ;
      RECT  288600.0 340650.0 287400.0 341850.0 ;
      RECT  297000.0 342750.0 295800.0 343950.0 ;
      RECT  298800.0 340650.0 297600.0 341850.0 ;
      RECT  307200.0 342750.0 306000.0 343950.0 ;
      RECT  309000.0 340650.0 307800.0 341850.0 ;
      RECT  317400.0 342750.0 316200.0 343950.0 ;
      RECT  319200.0 340650.0 318000.0 341850.0 ;
      RECT  327600.0 342750.0 326400.0 343950.0 ;
      RECT  329400.0 340650.0 328200.0 341850.0 ;
      RECT  337800.0 342750.0 336600.0 343950.0 ;
      RECT  339600.0 340650.0 338400.0 341850.0 ;
      RECT  348000.0 342750.0 346800.0 343950.0 ;
      RECT  349800.0 340650.0 348600.0 341850.0 ;
      RECT  358200.0 342750.0 357000.0 343950.0 ;
      RECT  360000.0 340650.0 358800.0 341850.0 ;
      RECT  368400.0 342750.0 367200.0 343950.0 ;
      RECT  370200.0 340650.0 369000.0 341850.0 ;
      RECT  378600.0 342750.0 377400.0 343950.0 ;
      RECT  380400.0 340650.0 379200.0 341850.0 ;
      RECT  388800.0 342750.0 387600.0 343950.0 ;
      RECT  390600.0 340650.0 389400.0 341850.0 ;
      RECT  399000.0 342750.0 397800.0 343950.0 ;
      RECT  400800.0 340650.0 399600.0 341850.0 ;
      RECT  409200.0 342750.0 408000.0 343950.0 ;
      RECT  411000.0 340650.0 409800.0 341850.0 ;
      RECT  419400.0 342750.0 418200.0 343950.0 ;
      RECT  421200.0 340650.0 420000.0 341850.0 ;
      RECT  429600.0 342750.0 428400.0 343950.0 ;
      RECT  431400.0 340650.0 430200.0 341850.0 ;
      RECT  439800.0 342750.0 438600.0 343950.0 ;
      RECT  441600.0 340650.0 440400.0 341850.0 ;
      RECT  450000.0 342750.0 448800.0 343950.0 ;
      RECT  451800.0 340650.0 450600.0 341850.0 ;
      RECT  460200.0 342750.0 459000.0 343950.0 ;
      RECT  462000.0 340650.0 460800.0 341850.0 ;
      RECT  470400.0 342750.0 469200.0 343950.0 ;
      RECT  472200.0 340650.0 471000.0 341850.0 ;
      RECT  480600.0 342750.0 479400.0 343950.0 ;
      RECT  482400.0 340650.0 481200.0 341850.0 ;
      RECT  490800.0 342750.0 489600.0 343950.0 ;
      RECT  492600.0 340650.0 491400.0 341850.0 ;
      RECT  501000.0 342750.0 499800.0 343950.0 ;
      RECT  502800.0 340650.0 501600.0 341850.0 ;
      RECT  511200.0 342750.0 510000.0 343950.0 ;
      RECT  513000.0 340650.0 511800.0 341850.0 ;
      RECT  521400.0 342750.0 520200.0 343950.0 ;
      RECT  523200.0 340650.0 522000.0 341850.0 ;
      RECT  531600.0 342750.0 530400.0 343950.0 ;
      RECT  533400.0 340650.0 532200.0 341850.0 ;
      RECT  541800.0 342750.0 540600.0 343950.0 ;
      RECT  543600.0 340650.0 542400.0 341850.0 ;
      RECT  552000.0 342750.0 550800.0 343950.0 ;
      RECT  553800.0 340650.0 552600.0 341850.0 ;
      RECT  562200.0 342750.0 561000.0 343950.0 ;
      RECT  564000.0 340650.0 562800.0 341850.0 ;
      RECT  572400.0 342750.0 571200.0 343950.0 ;
      RECT  574200.0 340650.0 573000.0 341850.0 ;
      RECT  582600.0 342750.0 581400.0 343950.0 ;
      RECT  584400.0 340650.0 583200.0 341850.0 ;
      RECT  592800.0 342750.0 591600.0 343950.0 ;
      RECT  594600.0 340650.0 593400.0 341850.0 ;
      RECT  603000.0 342750.0 601800.0 343950.0 ;
      RECT  604800.0 340650.0 603600.0 341850.0 ;
      RECT  613200.0 342750.0 612000.0 343950.0 ;
      RECT  615000.0 340650.0 613800.0 341850.0 ;
      RECT  623400.0 342750.0 622200.0 343950.0 ;
      RECT  625200.0 340650.0 624000.0 341850.0 ;
      RECT  633600.0 342750.0 632400.0 343950.0 ;
      RECT  635400.0 340650.0 634200.0 341850.0 ;
      RECT  643800.0 342750.0 642600.0 343950.0 ;
      RECT  645600.0 340650.0 644400.0 341850.0 ;
      RECT  654000.0 342750.0 652800.0 343950.0 ;
      RECT  655800.0 340650.0 654600.0 341850.0 ;
      RECT  664200.0 342750.0 663000.0 343950.0 ;
      RECT  666000.0 340650.0 664800.0 341850.0 ;
      RECT  674400.0 342750.0 673200.0 343950.0 ;
      RECT  676200.0 340650.0 675000.0 341850.0 ;
      RECT  684600.0 342750.0 683400.0 343950.0 ;
      RECT  686400.0 340650.0 685200.0 341850.0 ;
      RECT  694800.0 342750.0 693600.0 343950.0 ;
      RECT  696600.0 340650.0 695400.0 341850.0 ;
      RECT  705000.0 342750.0 703800.0 343950.0 ;
      RECT  706800.0 340650.0 705600.0 341850.0 ;
      RECT  715200.0 342750.0 714000.0 343950.0 ;
      RECT  717000.0 340650.0 715800.0 341850.0 ;
      RECT  725400.0 342750.0 724200.0 343950.0 ;
      RECT  727200.0 340650.0 726000.0 341850.0 ;
      RECT  735600.0 342750.0 734400.0 343950.0 ;
      RECT  737400.0 340650.0 736200.0 341850.0 ;
      RECT  745800.0 342750.0 744600.0 343950.0 ;
      RECT  747600.0 340650.0 746400.0 341850.0 ;
      RECT  756000.0 342750.0 754800.0 343950.0 ;
      RECT  757800.0 340650.0 756600.0 341850.0 ;
      RECT  766200.0 342750.0 765000.0 343950.0 ;
      RECT  768000.0 340650.0 766800.0 341850.0 ;
      RECT  776400.0 342750.0 775200.0 343950.0 ;
      RECT  778200.0 340650.0 777000.0 341850.0 ;
      RECT  786600.0 342750.0 785400.0 343950.0 ;
      RECT  788400.0 340650.0 787200.0 341850.0 ;
      RECT  796800.0 342750.0 795600.0 343950.0 ;
      RECT  798600.0 340650.0 797400.0 341850.0 ;
      RECT  807000.0 342750.0 805800.0 343950.0 ;
      RECT  808800.0 340650.0 807600.0 341850.0 ;
      RECT  817200.0 342750.0 816000.0 343950.0 ;
      RECT  819000.0 340650.0 817800.0 341850.0 ;
      RECT  827400.0 342750.0 826200.0 343950.0 ;
      RECT  829200.0 340650.0 828000.0 341850.0 ;
      RECT  837600.0 342750.0 836400.0 343950.0 ;
      RECT  839400.0 340650.0 838200.0 341850.0 ;
      RECT  847800.0 342750.0 846600.0 343950.0 ;
      RECT  849600.0 340650.0 848400.0 341850.0 ;
      RECT  858000.0 342750.0 856800.0 343950.0 ;
      RECT  859800.0 340650.0 858600.0 341850.0 ;
      RECT  868200.0 342750.0 867000.0 343950.0 ;
      RECT  870000.0 340650.0 868800.0 341850.0 ;
      RECT  878400.0 342750.0 877200.0 343950.0 ;
      RECT  880200.0 340650.0 879000.0 341850.0 ;
      RECT  888600.0 342750.0 887400.0 343950.0 ;
      RECT  890400.0 340650.0 889200.0 341850.0 ;
      RECT  898800.0 342750.0 897600.0 343950.0 ;
      RECT  900600.0 340650.0 899400.0 341850.0 ;
      RECT  909000.0 342750.0 907800.0 343950.0 ;
      RECT  910800.0 340650.0 909600.0 341850.0 ;
      RECT  919200.0 342750.0 918000.0 343950.0 ;
      RECT  921000.0 340650.0 919800.0 341850.0 ;
      RECT  929400.0 342750.0 928200.0 343950.0 ;
      RECT  931200.0 340650.0 930000.0 341850.0 ;
      RECT  939600.0 342750.0 938400.0 343950.0 ;
      RECT  941400.0 340650.0 940200.0 341850.0 ;
      RECT  949800.0 342750.0 948600.0 343950.0 ;
      RECT  951600.0 340650.0 950400.0 341850.0 ;
      RECT  960000.0 342750.0 958800.0 343950.0 ;
      RECT  961800.0 340650.0 960600.0 341850.0 ;
      RECT  970200.0 342750.0 969000.0 343950.0 ;
      RECT  972000.0 340650.0 970800.0 341850.0 ;
      RECT  980400.0 342750.0 979200.0 343950.0 ;
      RECT  982200.0 340650.0 981000.0 341850.0 ;
      RECT  990600.0 342750.0 989400.0 343950.0 ;
      RECT  992400.0 340650.0 991200.0 341850.0 ;
      RECT  1000800.0 342750.0 999600.0 343950.0 ;
      RECT  1002600.0 340650.0 1001400.0 341850.0 ;
      RECT  1011000.0 342750.0 1009800.0 343950.0 ;
      RECT  1012800.0 340650.0 1011600.0 341850.0 ;
      RECT  1021200.0 342750.0 1020000.0 343950.0 ;
      RECT  1023000.0 340650.0 1021800.0 341850.0 ;
      RECT  1031400.0 342750.0 1030200.0 343950.0 ;
      RECT  1033200.0 340650.0 1032000.0 341850.0 ;
      RECT  1041600.0 342750.0 1040400.0 343950.0 ;
      RECT  1043400.0 340650.0 1042200.0 341850.0 ;
      RECT  1051800.0 342750.0 1050600.0 343950.0 ;
      RECT  1053600.0 340650.0 1052400.0 341850.0 ;
      RECT  1062000.0 342750.0 1060800.0 343950.0 ;
      RECT  1063800.0 340650.0 1062600.0 341850.0 ;
      RECT  1072200.0 342750.0 1071000.0 343950.0 ;
      RECT  1074000.0 340650.0 1072800.0 341850.0 ;
      RECT  1082400.0 342750.0 1081200.0 343950.0 ;
      RECT  1084200.0 340650.0 1083000.0 341850.0 ;
      RECT  1092600.0 342750.0 1091400.0 343950.0 ;
      RECT  1094400.0 340650.0 1093200.0 341850.0 ;
      RECT  1102800.0 342750.0 1101600.0 343950.0 ;
      RECT  1104600.0 340650.0 1103400.0 341850.0 ;
      RECT  1113000.0 342750.0 1111800.0 343950.0 ;
      RECT  1114800.0 340650.0 1113600.0 341850.0 ;
      RECT  1123200.0 342750.0 1122000.0 343950.0 ;
      RECT  1125000.0 340650.0 1123800.0 341850.0 ;
      RECT  1133400.0 342750.0 1132200.0 343950.0 ;
      RECT  1135200.0 340650.0 1134000.0 341850.0 ;
      RECT  1143600.0 342750.0 1142400.0 343950.0 ;
      RECT  1145400.0 340650.0 1144200.0 341850.0 ;
      RECT  1153800.0 342750.0 1152600.0 343950.0 ;
      RECT  1155600.0 340650.0 1154400.0 341850.0 ;
      RECT  1164000.0 342750.0 1162800.0 343950.0 ;
      RECT  1165800.0 340650.0 1164600.0 341850.0 ;
      RECT  1174200.0 342750.0 1173000.0 343950.0 ;
      RECT  1176000.0 340650.0 1174800.0 341850.0 ;
      RECT  1184400.0 342750.0 1183200.0 343950.0 ;
      RECT  1186200.0 340650.0 1185000.0 341850.0 ;
      RECT  1194600.0 342750.0 1193400.0 343950.0 ;
      RECT  1196400.0 340650.0 1195200.0 341850.0 ;
      RECT  1204800.0 342750.0 1203600.0 343950.0 ;
      RECT  1206600.0 340650.0 1205400.0 341850.0 ;
      RECT  1215000.0 342750.0 1213800.0 343950.0 ;
      RECT  1216800.0 340650.0 1215600.0 341850.0 ;
      RECT  1225200.0 342750.0 1224000.0 343950.0 ;
      RECT  1227000.0 340650.0 1225800.0 341850.0 ;
      RECT  1235400.0 342750.0 1234200.0 343950.0 ;
      RECT  1237200.0 340650.0 1236000.0 341850.0 ;
      RECT  1245600.0 342750.0 1244400.0 343950.0 ;
      RECT  1247400.0 340650.0 1246200.0 341850.0 ;
      RECT  1255800.0 342750.0 1254600.0 343950.0 ;
      RECT  1257600.0 340650.0 1256400.0 341850.0 ;
      RECT  1266000.0 342750.0 1264800.0 343950.0 ;
      RECT  1267800.0 340650.0 1266600.0 341850.0 ;
      RECT  1276200.0 342750.0 1275000.0 343950.0 ;
      RECT  1278000.0 340650.0 1276800.0 341850.0 ;
      RECT  1286400.0 342750.0 1285200.0 343950.0 ;
      RECT  1288200.0 340650.0 1287000.0 341850.0 ;
      RECT  1296600.0 342750.0 1295400.0 343950.0 ;
      RECT  1298400.0 340650.0 1297200.0 341850.0 ;
      RECT  1306800.0 342750.0 1305600.0 343950.0 ;
      RECT  1308600.0 340650.0 1307400.0 341850.0 ;
      RECT  1317000.0 342750.0 1315800.0 343950.0 ;
      RECT  1318800.0 340650.0 1317600.0 341850.0 ;
      RECT  1327200.0 342750.0 1326000.0 343950.0 ;
      RECT  1329000.0 340650.0 1327800.0 341850.0 ;
      RECT  1337400.0 342750.0 1336200.0 343950.0 ;
      RECT  1339200.0 340650.0 1338000.0 341850.0 ;
      RECT  1347600.0 342750.0 1346400.0 343950.0 ;
      RECT  1349400.0 340650.0 1348200.0 341850.0 ;
      RECT  1357800.0 342750.0 1356600.0 343950.0 ;
      RECT  1359600.0 340650.0 1358400.0 341850.0 ;
      RECT  1368000.0 342750.0 1366800.0 343950.0 ;
      RECT  1369800.0 340650.0 1368600.0 341850.0 ;
      RECT  1378200.0 342750.0 1377000.0 343950.0 ;
      RECT  1380000.0 340650.0 1378800.0 341850.0 ;
      RECT  1388400.0 342750.0 1387200.0 343950.0 ;
      RECT  1390200.0 340650.0 1389000.0 341850.0 ;
      RECT  1398600.0 342750.0 1397400.0 343950.0 ;
      RECT  1400400.0 340650.0 1399200.0 341850.0 ;
      RECT  1408800.0 342750.0 1407600.0 343950.0 ;
      RECT  1410600.0 340650.0 1409400.0 341850.0 ;
      RECT  1419000.0 342750.0 1417800.0 343950.0 ;
      RECT  1420800.0 340650.0 1419600.0 341850.0 ;
      RECT  1429200.0 342750.0 1428000.0 343950.0 ;
      RECT  1431000.0 340650.0 1429800.0 341850.0 ;
      RECT  1439400.0 342750.0 1438200.0 343950.0 ;
      RECT  1441200.0 340650.0 1440000.0 341850.0 ;
      RECT  1449600.0 342750.0 1448400.0 343950.0 ;
      RECT  1451400.0 340650.0 1450200.0 341850.0 ;
      RECT  1459800.0 342750.0 1458600.0 343950.0 ;
      RECT  1461600.0 340650.0 1460400.0 341850.0 ;
      RECT  1470000.0 342750.0 1468800.0 343950.0 ;
      RECT  1471800.0 340650.0 1470600.0 341850.0 ;
      RECT  1480200.0 342750.0 1479000.0 343950.0 ;
      RECT  1482000.0 340650.0 1480800.0 341850.0 ;
      RECT  1490400.0 342750.0 1489200.0 343950.0 ;
      RECT  1492200.0 340650.0 1491000.0 341850.0 ;
      RECT  1500600.0 342750.0 1499400.0 343950.0 ;
      RECT  1502400.0 340650.0 1501200.0 341850.0 ;
      RECT  1510800.0 342750.0 1509600.0 343950.0 ;
      RECT  1512600.0 340650.0 1511400.0 341850.0 ;
      RECT  1521000.0 342750.0 1519800.0 343950.0 ;
      RECT  1522800.0 340650.0 1521600.0 341850.0 ;
      RECT  224400.0 376950.0 225300.0 378750.0 ;
      RECT  227400.0 376950.0 228300.0 378750.0 ;
      RECT  234600.0 376950.0 235500.0 378750.0 ;
      RECT  237600.0 376950.0 238500.0 378750.0 ;
      RECT  244800.0 376950.0 245700.0 378750.0 ;
      RECT  247800.0 376950.0 248700.0 378750.0 ;
      RECT  255000.0 376950.0 255900.0 378750.0 ;
      RECT  258000.0 376950.0 258900.0 378750.0 ;
      RECT  265200.0 376950.0 266100.0 378750.0 ;
      RECT  268200.0 376950.0 269100.0 378750.0 ;
      RECT  275400.0 376950.0 276300.0 378750.0 ;
      RECT  278400.0 376950.0 279300.0 378750.0 ;
      RECT  285600.0 376950.0 286500.0 378750.0 ;
      RECT  288600.0 376950.0 289500.0 378750.0 ;
      RECT  295800.0 376950.0 296700.0 378750.0 ;
      RECT  298800.0 376950.0 299700.0 378750.0 ;
      RECT  306000.0 376950.0 306900.0 378750.0 ;
      RECT  309000.0 376950.0 309900.0 378750.0 ;
      RECT  316200.0 376950.0 317100.0 378750.0 ;
      RECT  319200.0 376950.0 320100.0 378750.0 ;
      RECT  326400.0 376950.0 327300.0 378750.0 ;
      RECT  329400.0 376950.0 330300.0 378750.0 ;
      RECT  336600.0 376950.0 337500.0 378750.0 ;
      RECT  339600.0 376950.0 340500.0 378750.0 ;
      RECT  346800.0 376950.0 347700.0 378750.0 ;
      RECT  349800.0 376950.0 350700.0 378750.0 ;
      RECT  357000.0 376950.0 357900.0 378750.0 ;
      RECT  360000.0 376950.0 360900.0 378750.0 ;
      RECT  367200.0 376950.0 368100.0 378750.0 ;
      RECT  370200.0 376950.0 371100.0 378750.0 ;
      RECT  377400.0 376950.0 378300.0 378750.0 ;
      RECT  380400.0 376950.0 381300.0 378750.0 ;
      RECT  387600.0 376950.0 388500.0 378750.0 ;
      RECT  390600.0 376950.0 391500.0 378750.0 ;
      RECT  397800.0 376950.0 398700.0 378750.0 ;
      RECT  400800.0 376950.0 401700.0 378750.0 ;
      RECT  408000.0 376950.0 408900.0 378750.0 ;
      RECT  411000.0 376950.0 411900.0 378750.0 ;
      RECT  418200.0 376950.0 419100.0 378750.0 ;
      RECT  421200.0 376950.0 422100.0 378750.0 ;
      RECT  428400.0 376950.0 429300.0 378750.0 ;
      RECT  431400.0 376950.0 432300.0 378750.0 ;
      RECT  438600.0 376950.0 439500.0 378750.0 ;
      RECT  441600.0 376950.0 442500.0 378750.0 ;
      RECT  448800.0 376950.0 449700.0 378750.0 ;
      RECT  451800.0 376950.0 452700.0 378750.0 ;
      RECT  459000.0 376950.0 459900.0 378750.0 ;
      RECT  462000.0 376950.0 462900.0 378750.0 ;
      RECT  469200.0 376950.0 470100.0 378750.0 ;
      RECT  472200.0 376950.0 473100.0 378750.0 ;
      RECT  479400.0 376950.0 480300.0 378750.0 ;
      RECT  482400.0 376950.0 483300.0 378750.0 ;
      RECT  489600.0 376950.0 490500.0 378750.0 ;
      RECT  492600.0 376950.0 493500.0 378750.0 ;
      RECT  499800.0 376950.0 500700.0 378750.0 ;
      RECT  502800.0 376950.0 503700.0 378750.0 ;
      RECT  510000.0 376950.0 510900.0 378750.0 ;
      RECT  513000.0 376950.0 513900.0 378750.0 ;
      RECT  520200.0 376950.0 521100.0 378750.0 ;
      RECT  523200.0 376950.0 524100.0 378750.0 ;
      RECT  530400.0 376950.0 531300.0 378750.0 ;
      RECT  533400.0 376950.0 534300.0 378750.0 ;
      RECT  540600.0 376950.0 541500.0 378750.0 ;
      RECT  543600.0 376950.0 544500.0 378750.0 ;
      RECT  550800.0 376950.0 551700.0 378750.0 ;
      RECT  553800.0 376950.0 554700.0 378750.0 ;
      RECT  561000.0 376950.0 561900.0 378750.0 ;
      RECT  564000.0 376950.0 564900.0 378750.0 ;
      RECT  571200.0 376950.0 572100.0 378750.0 ;
      RECT  574200.0 376950.0 575100.0 378750.0 ;
      RECT  581400.0 376950.0 582300.0 378750.0 ;
      RECT  584400.0 376950.0 585300.0 378750.0 ;
      RECT  591600.0 376950.0 592500.0 378750.0 ;
      RECT  594600.0 376950.0 595500.0 378750.0 ;
      RECT  601800.0 376950.0 602700.0 378750.0 ;
      RECT  604800.0 376950.0 605700.0 378750.0 ;
      RECT  612000.0 376950.0 612900.0 378750.0 ;
      RECT  615000.0 376950.0 615900.0 378750.0 ;
      RECT  622200.0 376950.0 623100.0 378750.0 ;
      RECT  625200.0 376950.0 626100.0 378750.0 ;
      RECT  632400.0 376950.0 633300.0 378750.0 ;
      RECT  635400.0 376950.0 636300.0 378750.0 ;
      RECT  642600.0 376950.0 643500.0 378750.0 ;
      RECT  645600.0 376950.0 646500.0 378750.0 ;
      RECT  652800.0 376950.0 653700.0 378750.0 ;
      RECT  655800.0 376950.0 656700.0 378750.0 ;
      RECT  663000.0 376950.0 663900.0 378750.0 ;
      RECT  666000.0 376950.0 666900.0 378750.0 ;
      RECT  673200.0 376950.0 674100.0 378750.0 ;
      RECT  676200.0 376950.0 677100.0 378750.0 ;
      RECT  683400.0 376950.0 684300.0 378750.0 ;
      RECT  686400.0 376950.0 687300.0 378750.0 ;
      RECT  693600.0 376950.0 694500.0 378750.0 ;
      RECT  696600.0 376950.0 697500.0 378750.0 ;
      RECT  703800.0 376950.0 704700.0 378750.0 ;
      RECT  706800.0 376950.0 707700.0 378750.0 ;
      RECT  714000.0 376950.0 714900.0 378750.0 ;
      RECT  717000.0 376950.0 717900.0 378750.0 ;
      RECT  724200.0 376950.0 725100.0 378750.0 ;
      RECT  727200.0 376950.0 728100.0 378750.0 ;
      RECT  734400.0 376950.0 735300.0 378750.0 ;
      RECT  737400.0 376950.0 738300.0 378750.0 ;
      RECT  744600.0 376950.0 745500.0 378750.0 ;
      RECT  747600.0 376950.0 748500.0 378750.0 ;
      RECT  754800.0 376950.0 755700.0 378750.0 ;
      RECT  757800.0 376950.0 758700.0 378750.0 ;
      RECT  765000.0 376950.0 765900.0 378750.0 ;
      RECT  768000.0 376950.0 768900.0 378750.0 ;
      RECT  775200.0 376950.0 776100.0 378750.0 ;
      RECT  778200.0 376950.0 779100.0 378750.0 ;
      RECT  785400.0 376950.0 786300.0 378750.0 ;
      RECT  788400.0 376950.0 789300.0 378750.0 ;
      RECT  795600.0 376950.0 796500.0 378750.0 ;
      RECT  798600.0 376950.0 799500.0 378750.0 ;
      RECT  805800.0 376950.0 806700.0 378750.0 ;
      RECT  808800.0 376950.0 809700.0 378750.0 ;
      RECT  816000.0 376950.0 816900.0 378750.0 ;
      RECT  819000.0 376950.0 819900.0 378750.0 ;
      RECT  826200.0 376950.0 827100.0 378750.0 ;
      RECT  829200.0 376950.0 830100.0 378750.0 ;
      RECT  836400.0 376950.0 837300.0 378750.0 ;
      RECT  839400.0 376950.0 840300.0 378750.0 ;
      RECT  846600.0 376950.0 847500.0 378750.0 ;
      RECT  849600.0 376950.0 850500.0 378750.0 ;
      RECT  856800.0 376950.0 857700.0 378750.0 ;
      RECT  859800.0 376950.0 860700.0 378750.0 ;
      RECT  867000.0 376950.0 867900.0 378750.0 ;
      RECT  870000.0 376950.0 870900.0 378750.0 ;
      RECT  877200.0 376950.0 878100.0 378750.0 ;
      RECT  880200.0 376950.0 881100.0 378750.0 ;
      RECT  887400.0 376950.0 888300.0 378750.0 ;
      RECT  890400.0 376950.0 891300.0 378750.0 ;
      RECT  897600.0 376950.0 898500.0 378750.0 ;
      RECT  900600.0 376950.0 901500.0 378750.0 ;
      RECT  907800.0 376950.0 908700.0 378750.0 ;
      RECT  910800.0 376950.0 911700.0 378750.0 ;
      RECT  918000.0 376950.0 918900.0 378750.0 ;
      RECT  921000.0 376950.0 921900.0 378750.0 ;
      RECT  928200.0 376950.0 929100.0 378750.0 ;
      RECT  931200.0 376950.0 932100.0 378750.0 ;
      RECT  938400.0 376950.0 939300.0 378750.0 ;
      RECT  941400.0 376950.0 942300.0 378750.0 ;
      RECT  948600.0 376950.0 949500.0 378750.0 ;
      RECT  951600.0 376950.0 952500.0 378750.0 ;
      RECT  958800.0 376950.0 959700.0 378750.0 ;
      RECT  961800.0 376950.0 962700.0 378750.0 ;
      RECT  969000.0 376950.0 969900.0 378750.0 ;
      RECT  972000.0 376950.0 972900.0 378750.0 ;
      RECT  979200.0 376950.0 980100.0 378750.0 ;
      RECT  982200.0 376950.0 983100.0 378750.0 ;
      RECT  989400.0 376950.0 990300.0 378750.0 ;
      RECT  992400.0 376950.0 993300.0 378750.0 ;
      RECT  999600.0 376950.0 1000500.0 378750.0 ;
      RECT  1002600.0 376950.0 1003500.0 378750.0 ;
      RECT  1009800.0 376950.0 1010700.0 378750.0 ;
      RECT  1012800.0 376950.0 1013700.0 378750.0 ;
      RECT  1020000.0 376950.0 1020900.0 378750.0 ;
      RECT  1023000.0 376950.0 1023900.0 378750.0 ;
      RECT  1030200.0 376950.0 1031100.0 378750.0 ;
      RECT  1033200.0 376950.0 1034100.0 378750.0 ;
      RECT  1040400.0 376950.0 1041300.0 378750.0 ;
      RECT  1043400.0 376950.0 1044300.0 378750.0 ;
      RECT  1050600.0 376950.0 1051500.0 378750.0 ;
      RECT  1053600.0 376950.0 1054500.0 378750.0 ;
      RECT  1060800.0 376950.0 1061700.0 378750.0 ;
      RECT  1063800.0 376950.0 1064700.0 378750.0 ;
      RECT  1071000.0 376950.0 1071900.0 378750.0 ;
      RECT  1074000.0 376950.0 1074900.0 378750.0 ;
      RECT  1081200.0 376950.0 1082100.0 378750.0 ;
      RECT  1084200.0 376950.0 1085100.0 378750.0 ;
      RECT  1091400.0 376950.0 1092300.0 378750.0 ;
      RECT  1094400.0 376950.0 1095300.0 378750.0 ;
      RECT  1101600.0 376950.0 1102500.0 378750.0 ;
      RECT  1104600.0 376950.0 1105500.0 378750.0 ;
      RECT  1111800.0 376950.0 1112700.0 378750.0 ;
      RECT  1114800.0 376950.0 1115700.0 378750.0 ;
      RECT  1122000.0 376950.0 1122900.0 378750.0 ;
      RECT  1125000.0 376950.0 1125900.0 378750.0 ;
      RECT  1132200.0 376950.0 1133100.0 378750.0 ;
      RECT  1135200.0 376950.0 1136100.0 378750.0 ;
      RECT  1142400.0 376950.0 1143300.0 378750.0 ;
      RECT  1145400.0 376950.0 1146300.0 378750.0 ;
      RECT  1152600.0 376950.0 1153500.0 378750.0 ;
      RECT  1155600.0 376950.0 1156500.0 378750.0 ;
      RECT  1162800.0 376950.0 1163700.0 378750.0 ;
      RECT  1165800.0 376950.0 1166700.0 378750.0 ;
      RECT  1173000.0 376950.0 1173900.0 378750.0 ;
      RECT  1176000.0 376950.0 1176900.0 378750.0 ;
      RECT  1183200.0 376950.0 1184100.0 378750.0 ;
      RECT  1186200.0 376950.0 1187100.0 378750.0 ;
      RECT  1193400.0 376950.0 1194300.0 378750.0 ;
      RECT  1196400.0 376950.0 1197300.0 378750.0 ;
      RECT  1203600.0 376950.0 1204500.0 378750.0 ;
      RECT  1206600.0 376950.0 1207500.0 378750.0 ;
      RECT  1213800.0 376950.0 1214700.0 378750.0 ;
      RECT  1216800.0 376950.0 1217700.0 378750.0 ;
      RECT  1224000.0 376950.0 1224900.0 378750.0 ;
      RECT  1227000.0 376950.0 1227900.0 378750.0 ;
      RECT  1234200.0 376950.0 1235100.0 378750.0 ;
      RECT  1237200.0 376950.0 1238100.0 378750.0 ;
      RECT  1244400.0 376950.0 1245300.0 378750.0 ;
      RECT  1247400.0 376950.0 1248300.0 378750.0 ;
      RECT  1254600.0 376950.0 1255500.0 378750.0 ;
      RECT  1257600.0 376950.0 1258500.0 378750.0 ;
      RECT  1264800.0 376950.0 1265700.0 378750.0 ;
      RECT  1267800.0 376950.0 1268700.0 378750.0 ;
      RECT  1275000.0 376950.0 1275900.0 378750.0 ;
      RECT  1278000.0 376950.0 1278900.0 378750.0 ;
      RECT  1285200.0 376950.0 1286100.0 378750.0 ;
      RECT  1288200.0 376950.0 1289100.0 378750.0 ;
      RECT  1295400.0 376950.0 1296300.0 378750.0 ;
      RECT  1298400.0 376950.0 1299300.0 378750.0 ;
      RECT  1305600.0 376950.0 1306500.0 378750.0 ;
      RECT  1308600.0 376950.0 1309500.0 378750.0 ;
      RECT  1315800.0 376950.0 1316700.0 378750.0 ;
      RECT  1318800.0 376950.0 1319700.0 378750.0 ;
      RECT  1326000.0 376950.0 1326900.0 378750.0 ;
      RECT  1329000.0 376950.0 1329900.0 378750.0 ;
      RECT  1336200.0 376950.0 1337100.0 378750.0 ;
      RECT  1339200.0 376950.0 1340100.0 378750.0 ;
      RECT  1346400.0 376950.0 1347300.0 378750.0 ;
      RECT  1349400.0 376950.0 1350300.0 378750.0 ;
      RECT  1356600.0 376950.0 1357500.0 378750.0 ;
      RECT  1359600.0 376950.0 1360500.0 378750.0 ;
      RECT  1366800.0 376950.0 1367700.0 378750.0 ;
      RECT  1369800.0 376950.0 1370700.0 378750.0 ;
      RECT  1377000.0 376950.0 1377900.0 378750.0 ;
      RECT  1380000.0 376950.0 1380900.0 378750.0 ;
      RECT  1387200.0 376950.0 1388100.0 378750.0 ;
      RECT  1390200.0 376950.0 1391100.0 378750.0 ;
      RECT  1397400.0 376950.0 1398300.0 378750.0 ;
      RECT  1400400.0 376950.0 1401300.0 378750.0 ;
      RECT  1407600.0 376950.0 1408500.0 378750.0 ;
      RECT  1410600.0 376950.0 1411500.0 378750.0 ;
      RECT  1417800.0 376950.0 1418700.0 378750.0 ;
      RECT  1420800.0 376950.0 1421700.0 378750.0 ;
      RECT  1428000.0 376950.0 1428900.0 378750.0 ;
      RECT  1431000.0 376950.0 1431900.0 378750.0 ;
      RECT  1438200.0 376950.0 1439100.0 378750.0 ;
      RECT  1441200.0 376950.0 1442100.0 378750.0 ;
      RECT  1448400.0 376950.0 1449300.0 378750.0 ;
      RECT  1451400.0 376950.0 1452300.0 378750.0 ;
      RECT  1458600.0 376950.0 1459500.0 378750.0 ;
      RECT  1461600.0 376950.0 1462500.0 378750.0 ;
      RECT  1468800.0 376950.0 1469700.0 378750.0 ;
      RECT  1471800.0 376950.0 1472700.0 378750.0 ;
      RECT  1479000.0 376950.0 1479900.0 378750.0 ;
      RECT  1482000.0 376950.0 1482900.0 378750.0 ;
      RECT  1489200.0 376950.0 1490100.0 378750.0 ;
      RECT  1492200.0 376950.0 1493100.0 378750.0 ;
      RECT  1499400.0 376950.0 1500300.0 378750.0 ;
      RECT  1502400.0 376950.0 1503300.0 378750.0 ;
      RECT  1509600.0 376950.0 1510500.0 378750.0 ;
      RECT  1512600.0 376950.0 1513500.0 378750.0 ;
      RECT  1519800.0 376950.0 1520700.0 378750.0 ;
      RECT  1522800.0 376950.0 1523700.0 378750.0 ;
      RECT  224400.0 338550.0 225300.0 353250.0 ;
      RECT  227400.0 338550.0 228300.0 353250.0 ;
      RECT  265200.0 338550.0 266100.0 353250.0 ;
      RECT  268200.0 338550.0 269100.0 353250.0 ;
      RECT  306000.0 338550.0 306900.0 353250.0 ;
      RECT  309000.0 338550.0 309900.0 353250.0 ;
      RECT  346800.0 338550.0 347700.0 353250.0 ;
      RECT  349800.0 338550.0 350700.0 353250.0 ;
      RECT  387600.0 338550.0 388500.0 353250.0 ;
      RECT  390600.0 338550.0 391500.0 353250.0 ;
      RECT  428400.0 338550.0 429300.0 353250.0 ;
      RECT  431400.0 338550.0 432300.0 353250.0 ;
      RECT  469200.0 338550.0 470100.0 353250.0 ;
      RECT  472200.0 338550.0 473100.0 353250.0 ;
      RECT  510000.0 338550.0 510900.0 353250.0 ;
      RECT  513000.0 338550.0 513900.0 353250.0 ;
      RECT  550800.0 338550.0 551700.0 353250.0 ;
      RECT  553800.0 338550.0 554700.0 353250.0 ;
      RECT  591600.0 338550.0 592500.0 353250.0 ;
      RECT  594600.0 338550.0 595500.0 353250.0 ;
      RECT  632400.0 338550.0 633300.0 353250.0 ;
      RECT  635400.0 338550.0 636300.0 353250.0 ;
      RECT  673200.0 338550.0 674100.0 353250.0 ;
      RECT  676200.0 338550.0 677100.0 353250.0 ;
      RECT  714000.0 338550.0 714900.0 353250.0 ;
      RECT  717000.0 338550.0 717900.0 353250.0 ;
      RECT  754800.0 338550.0 755700.0 353250.0 ;
      RECT  757800.0 338550.0 758700.0 353250.0 ;
      RECT  795600.0 338550.0 796500.0 353250.0 ;
      RECT  798600.0 338550.0 799500.0 353250.0 ;
      RECT  836400.0 338550.0 837300.0 353250.0 ;
      RECT  839400.0 338550.0 840300.0 353250.0 ;
      RECT  877200.0 338550.0 878100.0 353250.0 ;
      RECT  880200.0 338550.0 881100.0 353250.0 ;
      RECT  918000.0 338550.0 918900.0 353250.0 ;
      RECT  921000.0 338550.0 921900.0 353250.0 ;
      RECT  958800.0 338550.0 959700.0 353250.0 ;
      RECT  961800.0 338550.0 962700.0 353250.0 ;
      RECT  999600.0 338550.0 1000500.0 353250.0 ;
      RECT  1002600.0 338550.0 1003500.0 353250.0 ;
      RECT  1040400.0 338550.0 1041300.0 353250.0 ;
      RECT  1043400.0 338550.0 1044300.0 353250.0 ;
      RECT  1081200.0 338550.0 1082100.0 353250.0 ;
      RECT  1084200.0 338550.0 1085100.0 353250.0 ;
      RECT  1122000.0 338550.0 1122900.0 353250.0 ;
      RECT  1125000.0 338550.0 1125900.0 353250.0 ;
      RECT  1162800.0 338550.0 1163700.0 353250.0 ;
      RECT  1165800.0 338550.0 1166700.0 353250.0 ;
      RECT  1203600.0 338550.0 1204500.0 353250.0 ;
      RECT  1206600.0 338550.0 1207500.0 353250.0 ;
      RECT  1244400.0 338550.0 1245300.0 353250.0 ;
      RECT  1247400.0 338550.0 1248300.0 353250.0 ;
      RECT  1285200.0 338550.0 1286100.0 353250.0 ;
      RECT  1288200.0 338550.0 1289100.0 353250.0 ;
      RECT  1326000.0 338550.0 1326900.0 353250.0 ;
      RECT  1329000.0 338550.0 1329900.0 353250.0 ;
      RECT  1366800.0 338550.0 1367700.0 353250.0 ;
      RECT  1369800.0 338550.0 1370700.0 353250.0 ;
      RECT  1407600.0 338550.0 1408500.0 353250.0 ;
      RECT  1410600.0 338550.0 1411500.0 353250.0 ;
      RECT  1448400.0 338550.0 1449300.0 353250.0 ;
      RECT  1451400.0 338550.0 1452300.0 353250.0 ;
      RECT  1489200.0 338550.0 1490100.0 353250.0 ;
      RECT  1492200.0 338550.0 1493100.0 353250.0 ;
      RECT  220800.0 338550.0 221700.0 378750.0 ;
      RECT  231000.0 338550.0 231900.0 378750.0 ;
      RECT  241200.0 338550.0 242100.0 378750.0 ;
      RECT  251400.0 338550.0 252300.0 378750.0 ;
      RECT  261600.0 338550.0 262500.0 378750.0 ;
      RECT  271800.0 338550.0 272700.0 378750.0 ;
      RECT  282000.0 338550.0 282900.0 378750.0 ;
      RECT  292200.0 338550.0 293100.0 378750.0 ;
      RECT  302400.0 338550.0 303300.0 378750.0 ;
      RECT  312600.0 338550.0 313500.0 378750.0 ;
      RECT  322800.0 338550.0 323700.0 378750.0 ;
      RECT  333000.0 338550.0 333900.0 378750.0 ;
      RECT  343200.0 338550.0 344100.0 378750.0 ;
      RECT  353400.0 338550.0 354300.0 378750.0 ;
      RECT  363600.0 338550.0 364500.0 378750.0 ;
      RECT  373800.0 338550.0 374700.0 378750.0 ;
      RECT  384000.0 338550.0 384900.0 378750.0 ;
      RECT  394200.0 338550.0 395100.0 378750.0 ;
      RECT  404400.0 338550.0 405300.0 378750.0 ;
      RECT  414600.0 338550.0 415500.0 378750.0 ;
      RECT  424800.0 338550.0 425700.0 378750.0 ;
      RECT  435000.0 338550.0 435900.0 378750.0 ;
      RECT  445200.0 338550.0 446100.0 378750.0 ;
      RECT  455400.0 338550.0 456300.0 378750.0 ;
      RECT  465600.0 338550.0 466500.0 378750.0 ;
      RECT  475800.0 338550.0 476700.0 378750.0 ;
      RECT  486000.0 338550.0 486900.0 378750.0 ;
      RECT  496200.0 338550.0 497100.0 378750.0 ;
      RECT  506400.0 338550.0 507300.0 378750.0 ;
      RECT  516600.0 338550.0 517500.0 378750.0 ;
      RECT  526800.0 338550.0 527700.0 378750.0 ;
      RECT  537000.0 338550.0 537900.0 378750.0 ;
      RECT  547200.0 338550.0 548100.0 378750.0 ;
      RECT  557400.0 338550.0 558300.0 378750.0 ;
      RECT  567600.0 338550.0 568500.0 378750.0 ;
      RECT  577800.0 338550.0 578700.0 378750.0 ;
      RECT  588000.0 338550.0 588900.0 378750.0 ;
      RECT  598200.0 338550.0 599100.0 378750.0 ;
      RECT  608400.0 338550.0 609300.0 378750.0 ;
      RECT  618600.0 338550.0 619500.0 378750.0 ;
      RECT  628800.0 338550.0 629700.0 378750.0 ;
      RECT  639000.0 338550.0 639900.0 378750.0 ;
      RECT  649200.0 338550.0 650100.0 378750.0 ;
      RECT  659400.0 338550.0 660300.0 378750.0 ;
      RECT  669600.0 338550.0 670500.0 378750.0 ;
      RECT  679800.0 338550.0 680700.0 378750.0 ;
      RECT  690000.0 338550.0 690900.0 378750.0 ;
      RECT  700200.0 338550.0 701100.0 378750.0 ;
      RECT  710400.0 338550.0 711300.0 378750.0 ;
      RECT  720600.0 338550.0 721500.0 378750.0 ;
      RECT  730800.0 338550.0 731700.0 378750.0 ;
      RECT  741000.0 338550.0 741900.0 378750.0 ;
      RECT  751200.0 338550.0 752100.0 378750.0 ;
      RECT  761400.0 338550.0 762300.0 378750.0 ;
      RECT  771600.0 338550.0 772500.0 378750.0 ;
      RECT  781800.0 338550.0 782700.0 378750.0 ;
      RECT  792000.0 338550.0 792900.0 378750.0 ;
      RECT  802200.0 338550.0 803100.0 378750.0 ;
      RECT  812400.0 338550.0 813300.0 378750.0 ;
      RECT  822600.0 338550.0 823500.0 378750.0 ;
      RECT  832800.0 338550.0 833700.0 378750.0 ;
      RECT  843000.0 338550.0 843900.0 378750.0 ;
      RECT  853200.0 338550.0 854100.0 378750.0 ;
      RECT  863400.0 338550.0 864300.0 378750.0 ;
      RECT  873600.0 338550.0 874500.0 378750.0 ;
      RECT  883800.0 338550.0 884700.0 378750.0 ;
      RECT  894000.0 338550.0 894900.0 378750.0 ;
      RECT  904200.0 338550.0 905100.0 378750.0 ;
      RECT  914400.0 338550.0 915300.0 378750.0 ;
      RECT  924600.0 338550.0 925500.0 378750.0 ;
      RECT  934800.0 338550.0 935700.0 378750.0 ;
      RECT  945000.0 338550.0 945900.0 378750.0 ;
      RECT  955200.0 338550.0 956100.0 378750.0 ;
      RECT  965400.0 338550.0 966300.0 378750.0 ;
      RECT  975600.0 338550.0 976500.0 378750.0 ;
      RECT  985800.0 338550.0 986700.0 378750.0 ;
      RECT  996000.0 338550.0 996900.0 378750.0 ;
      RECT  1006200.0 338550.0 1007100.0 378750.0 ;
      RECT  1016400.0 338550.0 1017300.0 378750.0 ;
      RECT  1026600.0 338550.0 1027500.0 378750.0 ;
      RECT  1036800.0 338550.0 1037700.0 378750.0 ;
      RECT  1047000.0 338550.0 1047900.0 378750.0 ;
      RECT  1057200.0 338550.0 1058100.0 378750.0 ;
      RECT  1067400.0 338550.0 1068300.0 378750.0 ;
      RECT  1077600.0 338550.0 1078500.0 378750.0 ;
      RECT  1087800.0 338550.0 1088700.0 378750.0 ;
      RECT  1098000.0 338550.0 1098900.0 378750.0 ;
      RECT  1108200.0 338550.0 1109100.0 378750.0 ;
      RECT  1118400.0 338550.0 1119300.0 378750.0 ;
      RECT  1128600.0 338550.0 1129500.0 378750.0 ;
      RECT  1138800.0 338550.0 1139700.0 378750.0 ;
      RECT  1149000.0 338550.0 1149900.0 378750.0 ;
      RECT  1159200.0 338550.0 1160100.0 378750.0 ;
      RECT  1169400.0 338550.0 1170300.0 378750.0 ;
      RECT  1179600.0 338550.0 1180500.0 378750.0 ;
      RECT  1189800.0 338550.0 1190700.0 378750.0 ;
      RECT  1200000.0 338550.0 1200900.0 378750.0 ;
      RECT  1210200.0 338550.0 1211100.0 378750.0 ;
      RECT  1220400.0 338550.0 1221300.0 378750.0 ;
      RECT  1230600.0 338550.0 1231500.0 378750.0 ;
      RECT  1240800.0 338550.0 1241700.0 378750.0 ;
      RECT  1251000.0 338550.0 1251900.0 378750.0 ;
      RECT  1261200.0 338550.0 1262100.0 378750.0 ;
      RECT  1271400.0 338550.0 1272300.0 378750.0 ;
      RECT  1281600.0 338550.0 1282500.0 378750.0 ;
      RECT  1291800.0 338550.0 1292700.0 378750.0 ;
      RECT  1302000.0 338550.0 1302900.0 378750.0 ;
      RECT  1312200.0 338550.0 1313100.0 378750.0 ;
      RECT  1322400.0 338550.0 1323300.0 378750.0 ;
      RECT  1332600.0 338550.0 1333500.0 378750.0 ;
      RECT  1342800.0 338550.0 1343700.0 378750.0 ;
      RECT  1353000.0 338550.0 1353900.0 378750.0 ;
      RECT  1363200.0 338550.0 1364100.0 378750.0 ;
      RECT  1373400.0 338550.0 1374300.0 378750.0 ;
      RECT  1383600.0 338550.0 1384500.0 378750.0 ;
      RECT  1393800.0 338550.0 1394700.0 378750.0 ;
      RECT  1404000.0 338550.0 1404900.0 378750.0 ;
      RECT  1414200.0 338550.0 1415100.0 378750.0 ;
      RECT  1424400.0 338550.0 1425300.0 378750.0 ;
      RECT  1434600.0 338550.0 1435500.0 378750.0 ;
      RECT  1444800.0 338550.0 1445700.0 378750.0 ;
      RECT  1455000.0 338550.0 1455900.0 378750.0 ;
      RECT  1465200.0 338550.0 1466100.0 378750.0 ;
      RECT  1475400.0 338550.0 1476300.0 378750.0 ;
      RECT  1485600.0 338550.0 1486500.0 378750.0 ;
      RECT  1495800.0 338550.0 1496700.0 378750.0 ;
      RECT  1506000.0 338550.0 1506900.0 378750.0 ;
      RECT  1516200.0 338550.0 1517100.0 378750.0 ;
      RECT  122100.0 600.0 123000.0 54000.0 ;
      RECT  125100.0 600.0 126000.0 54000.0 ;
      RECT  116100.0 600.0 117000.0 54000.0 ;
      RECT  119100.0 600.0 120000.0 54000.0 ;
      RECT  132450.0 7950.0 133350.0 8850.0 ;
      RECT  134850.0 7950.0 135750.0 8850.0 ;
      RECT  132450.0 8400.0 133350.0 11250.0 ;
      RECT  132900.0 7950.0 135300.0 8850.0 ;
      RECT  134850.0 3750.0 135750.0 8400.0 ;
      RECT  132300.0 11250.0 133500.0 12450.0 ;
      RECT  134700.0 2550.0 135900.0 3750.0 ;
      RECT  135900.0 7800.0 134700.0 9000.0 ;
      RECT  132450.0 20850.0 133350.0 19950.0 ;
      RECT  134850.0 20850.0 135750.0 19950.0 ;
      RECT  132450.0 20400.0 133350.0 17550.0 ;
      RECT  132900.0 20850.0 135300.0 19950.0 ;
      RECT  134850.0 25050.0 135750.0 20400.0 ;
      RECT  132300.0 17550.0 133500.0 16350.0 ;
      RECT  134700.0 26250.0 135900.0 25050.0 ;
      RECT  135900.0 21000.0 134700.0 19800.0 ;
      RECT  132450.0 35550.0 133350.0 36450.0 ;
      RECT  134850.0 35550.0 135750.0 36450.0 ;
      RECT  132450.0 36000.0 133350.0 38850.0 ;
      RECT  132900.0 35550.0 135300.0 36450.0 ;
      RECT  134850.0 31350.0 135750.0 36000.0 ;
      RECT  132300.0 38850.0 133500.0 40050.0 ;
      RECT  134700.0 30150.0 135900.0 31350.0 ;
      RECT  135900.0 35400.0 134700.0 36600.0 ;
      RECT  132450.0 48450.0 133350.0 47550.0 ;
      RECT  134850.0 48450.0 135750.0 47550.0 ;
      RECT  132450.0 48000.0 133350.0 45150.0 ;
      RECT  132900.0 48450.0 135300.0 47550.0 ;
      RECT  134850.0 52650.0 135750.0 48000.0 ;
      RECT  132300.0 45150.0 133500.0 43950.0 ;
      RECT  134700.0 53850.0 135900.0 52650.0 ;
      RECT  135900.0 48600.0 134700.0 47400.0 ;
      RECT  117150.0 11100.0 115950.0 12300.0 ;
      RECT  98550.0 6600.0 97350.0 7800.0 ;
      RECT  120150.0 24900.0 118950.0 26100.0 ;
      RECT  101550.0 21000.0 100350.0 22200.0 ;
      RECT  98550.0 29700.0 97350.0 30900.0 ;
      RECT  123150.0 29700.0 121950.0 30900.0 ;
      RECT  101550.0 43500.0 100350.0 44700.0 ;
      RECT  126150.0 43500.0 124950.0 44700.0 ;
      RECT  117150.0 7800.0 115950.0 9000.0 ;
      RECT  120150.0 5100.0 118950.0 6300.0 ;
      RECT  123150.0 19800.0 121950.0 21000.0 ;
      RECT  120150.0 22500.0 118950.0 23700.0 ;
      RECT  117150.0 35400.0 115950.0 36600.0 ;
      RECT  126150.0 32700.0 124950.0 33900.0 ;
      RECT  123150.0 47400.0 121950.0 48600.0 ;
      RECT  126150.0 50100.0 124950.0 51300.0 ;
      RECT  97500.0 600.0 98400.0 54000.0 ;
      RECT  100500.0 600.0 101400.0 54000.0 ;
      RECT  221400.0 289650.0 231600.0 338550.0 ;
      RECT  262200.0 289650.0 272400.0 338550.0 ;
      RECT  303000.0 289650.0 313200.0 338550.0 ;
      RECT  343800.0 289650.0 354000.0 338550.0 ;
      RECT  384600.0 289650.0 394800.0 338550.0 ;
      RECT  425400.0 289650.0 435600.0 338550.0 ;
      RECT  466200.0 289650.0 476400.0 338550.0 ;
      RECT  507000.0 289650.0 517200.0 338550.0 ;
      RECT  547800.0 289650.0 558000.0 338550.0 ;
      RECT  588600.0 289650.0 598800.0 338550.0 ;
      RECT  629400.0 289650.0 639600.0 338550.0 ;
      RECT  670200.0 289650.0 680400.0 338550.0 ;
      RECT  711000.0 289650.0 721200.0 338550.0 ;
      RECT  751800.0 289650.0 762000.0 338550.0 ;
      RECT  792600.0 289650.0 802800.0 338550.0 ;
      RECT  833400.0 289650.0 843600.0 338550.0 ;
      RECT  874200.0 289650.0 884400.0 338550.0 ;
      RECT  915000.0 289650.0 925200.0 338550.0 ;
      RECT  955800.0 289650.0 966000.0 338550.0 ;
      RECT  996600.0 289650.0 1006800.0 338550.0 ;
      RECT  1037400.0 289650.0 1047600.0 338550.0 ;
      RECT  1078200.0 289650.0 1088400.0 338550.0 ;
      RECT  1119000.0 289650.0 1129200.0 338550.0 ;
      RECT  1159800.0 289650.0 1170000.0 338550.0 ;
      RECT  1200600.0 289650.0 1210800.0 338550.0 ;
      RECT  1241400.0 289650.0 1251600.0 338550.0 ;
      RECT  1282200.0 289650.0 1292400.0 338550.0 ;
      RECT  1323000.0 289650.0 1333200.0 338550.0 ;
      RECT  1363800.0 289650.0 1374000.0 338550.0 ;
      RECT  1404600.0 289650.0 1414800.0 338550.0 ;
      RECT  1445400.0 289650.0 1455600.0 338550.0 ;
      RECT  1486200.0 289650.0 1496400.0 338550.0 ;
      RECT  224400.0 289650.0 225600.0 302850.0 ;
      RECT  227400.0 289650.0 228600.0 302850.0 ;
      RECT  265200.0 289650.0 266400.0 302850.0 ;
      RECT  268200.0 289650.0 269400.0 302850.0 ;
      RECT  306000.0 289650.0 307200.0 302850.0 ;
      RECT  309000.0 289650.0 310200.0 302850.0 ;
      RECT  346800.0 289650.0 348000.0 302850.0 ;
      RECT  349800.0 289650.0 351000.0 302850.0 ;
      RECT  387600.0 289650.0 388800.0 302850.0 ;
      RECT  390600.0 289650.0 391800.0 302850.0 ;
      RECT  428400.0 289650.0 429600.0 302850.0 ;
      RECT  431400.0 289650.0 432600.0 302850.0 ;
      RECT  469200.0 289650.0 470400.0 302850.0 ;
      RECT  472200.0 289650.0 473400.0 302850.0 ;
      RECT  510000.0 289650.0 511200.0 302850.0 ;
      RECT  513000.0 289650.0 514200.0 302850.0 ;
      RECT  550800.0 289650.0 552000.0 302850.0 ;
      RECT  553800.0 289650.0 555000.0 302850.0 ;
      RECT  591600.0 289650.0 592800.0 302850.0 ;
      RECT  594600.0 289650.0 595800.0 302850.0 ;
      RECT  632400.0 289650.0 633600.0 302850.0 ;
      RECT  635400.0 289650.0 636600.0 302850.0 ;
      RECT  673200.0 289650.0 674400.0 302850.0 ;
      RECT  676200.0 289650.0 677400.0 302850.0 ;
      RECT  714000.0 289650.0 715200.0 302850.0 ;
      RECT  717000.0 289650.0 718200.0 302850.0 ;
      RECT  754800.0 289650.0 756000.0 302850.0 ;
      RECT  757800.0 289650.0 759000.0 302850.0 ;
      RECT  795600.0 289650.0 796800.0 302850.0 ;
      RECT  798600.0 289650.0 799800.0 302850.0 ;
      RECT  836400.0 289650.0 837600.0 302850.0 ;
      RECT  839400.0 289650.0 840600.0 302850.0 ;
      RECT  877200.0 289650.0 878400.0 302850.0 ;
      RECT  880200.0 289650.0 881400.0 302850.0 ;
      RECT  918000.0 289650.0 919200.0 302850.0 ;
      RECT  921000.0 289650.0 922200.0 302850.0 ;
      RECT  958800.0 289650.0 960000.0 302850.0 ;
      RECT  961800.0 289650.0 963000.0 302850.0 ;
      RECT  999600.0 289650.0 1000800.0 302850.0 ;
      RECT  1002600.0 289650.0 1003800.0 302850.0 ;
      RECT  1040400.0 289650.0 1041600.0 302850.0 ;
      RECT  1043400.0 289650.0 1044600.0 302850.0 ;
      RECT  1081200.0 289650.0 1082400.0 302850.0 ;
      RECT  1084200.0 289650.0 1085400.0 302850.0 ;
      RECT  1122000.0 289650.0 1123200.0 302850.0 ;
      RECT  1125000.0 289650.0 1126200.0 302850.0 ;
      RECT  1162800.0 289650.0 1164000.0 302850.0 ;
      RECT  1165800.0 289650.0 1167000.0 302850.0 ;
      RECT  1203600.0 289650.0 1204800.0 302850.0 ;
      RECT  1206600.0 289650.0 1207800.0 302850.0 ;
      RECT  1244400.0 289650.0 1245600.0 302850.0 ;
      RECT  1247400.0 289650.0 1248600.0 302850.0 ;
      RECT  1285200.0 289650.0 1286400.0 302850.0 ;
      RECT  1288200.0 289650.0 1289400.0 302850.0 ;
      RECT  1326000.0 289650.0 1327200.0 302850.0 ;
      RECT  1329000.0 289650.0 1330200.0 302850.0 ;
      RECT  1366800.0 289650.0 1368000.0 302850.0 ;
      RECT  1369800.0 289650.0 1371000.0 302850.0 ;
      RECT  1407600.0 289650.0 1408800.0 302850.0 ;
      RECT  1410600.0 289650.0 1411800.0 302850.0 ;
      RECT  1448400.0 289650.0 1449600.0 302850.0 ;
      RECT  1451400.0 289650.0 1452600.0 302850.0 ;
      RECT  1489200.0 289650.0 1490400.0 302850.0 ;
      RECT  1492200.0 289650.0 1493400.0 302850.0 ;
      RECT  221400.0 229050.0 231600.0 289650.0 ;
      RECT  262200.0 229050.0 272400.0 289650.0 ;
      RECT  303000.0 229050.0 313200.0 289650.0 ;
      RECT  343800.0 229050.0 354000.0 289650.0 ;
      RECT  384600.0 229050.0 394800.0 289650.0 ;
      RECT  425400.0 229050.0 435600.0 289650.0 ;
      RECT  466200.0 229050.0 476400.0 289650.0 ;
      RECT  507000.0 229050.0 517200.0 289650.0 ;
      RECT  547800.0 229050.0 558000.0 289650.0 ;
      RECT  588600.0 229050.0 598800.0 289650.0 ;
      RECT  629400.0 229050.0 639600.0 289650.0 ;
      RECT  670200.0 229050.0 680400.0 289650.0 ;
      RECT  711000.0 229050.0 721200.0 289650.0 ;
      RECT  751800.0 229050.0 762000.0 289650.0 ;
      RECT  792600.0 229050.0 802800.0 289650.0 ;
      RECT  833400.0 229050.0 843600.0 289650.0 ;
      RECT  874200.0 229050.0 884400.0 289650.0 ;
      RECT  915000.0 229050.0 925200.0 289650.0 ;
      RECT  955800.0 229050.0 966000.0 289650.0 ;
      RECT  996600.0 229050.0 1006800.0 289650.0 ;
      RECT  1037400.0 229050.0 1047600.0 289650.0 ;
      RECT  1078200.0 229050.0 1088400.0 289650.0 ;
      RECT  1119000.0 229050.0 1129200.0 289650.0 ;
      RECT  1159800.0 229050.0 1170000.0 289650.0 ;
      RECT  1200600.0 229050.0 1210800.0 289650.0 ;
      RECT  1241400.0 229050.0 1251600.0 289650.0 ;
      RECT  1282200.0 229050.0 1292400.0 289650.0 ;
      RECT  1323000.0 229050.0 1333200.0 289650.0 ;
      RECT  1363800.0 229050.0 1374000.0 289650.0 ;
      RECT  1404600.0 229050.0 1414800.0 289650.0 ;
      RECT  1445400.0 229050.0 1455600.0 289650.0 ;
      RECT  1486200.0 229050.0 1496400.0 289650.0 ;
      RECT  225900.0 229050.0 227100.0 232050.0 ;
      RECT  266700.0 229050.0 267900.0 232050.0 ;
      RECT  307500.0 229050.0 308700.0 232050.0 ;
      RECT  348300.0 229050.0 349500.0 232050.0 ;
      RECT  389100.0 229050.0 390300.0 232050.0 ;
      RECT  429900.0 229050.0 431100.0 232050.0 ;
      RECT  470700.0 229050.0 471900.0 232050.0 ;
      RECT  511500.0 229050.0 512700.0 232050.0 ;
      RECT  552300.0 229050.0 553500.0 232050.0 ;
      RECT  593100.0 229050.0 594300.0 232050.0 ;
      RECT  633900.0 229050.0 635100.0 232050.0 ;
      RECT  674700.0 229050.0 675900.0 232050.0 ;
      RECT  715500.0 229050.0 716700.0 232050.0 ;
      RECT  756300.0 229050.0 757500.0 232050.0 ;
      RECT  797100.0 229050.0 798300.0 232050.0 ;
      RECT  837900.0 229050.0 839100.0 232050.0 ;
      RECT  878700.0 229050.0 879900.0 232050.0 ;
      RECT  919500.0 229050.0 920700.0 232050.0 ;
      RECT  960300.0 229050.0 961500.0 232050.0 ;
      RECT  1001100.0 229050.0 1002300.0 232050.0 ;
      RECT  1041900.0 229050.0 1043100.0 232050.0 ;
      RECT  1082700.0 229050.0 1083900.0 232050.0 ;
      RECT  1123500.0 229050.0 1124700.0 232050.0 ;
      RECT  1164300.0 229050.0 1165500.0 232050.0 ;
      RECT  1205100.0 229050.0 1206300.0 232050.0 ;
      RECT  1245900.0 229050.0 1247100.0 232050.0 ;
      RECT  1286700.0 229050.0 1287900.0 232050.0 ;
      RECT  1327500.0 229050.0 1328700.0 232050.0 ;
      RECT  1368300.0 229050.0 1369500.0 232050.0 ;
      RECT  1409100.0 229050.0 1410300.0 232050.0 ;
      RECT  1449900.0 229050.0 1451100.0 232050.0 ;
      RECT  1490700.0 229050.0 1491900.0 232050.0 ;
      RECT  224400.0 287550.0 225600.0 289650.0 ;
      RECT  227400.0 282150.0 228600.0 289650.0 ;
      RECT  265200.0 287550.0 266400.0 289650.0 ;
      RECT  268200.0 282150.0 269400.0 289650.0 ;
      RECT  306000.0 287550.0 307200.0 289650.0 ;
      RECT  309000.0 282150.0 310200.0 289650.0 ;
      RECT  346800.0 287550.0 348000.0 289650.0 ;
      RECT  349800.0 282150.0 351000.0 289650.0 ;
      RECT  387600.0 287550.0 388800.0 289650.0 ;
      RECT  390600.0 282150.0 391800.0 289650.0 ;
      RECT  428400.0 287550.0 429600.0 289650.0 ;
      RECT  431400.0 282150.0 432600.0 289650.0 ;
      RECT  469200.0 287550.0 470400.0 289650.0 ;
      RECT  472200.0 282150.0 473400.0 289650.0 ;
      RECT  510000.0 287550.0 511200.0 289650.0 ;
      RECT  513000.0 282150.0 514200.0 289650.0 ;
      RECT  550800.0 287550.0 552000.0 289650.0 ;
      RECT  553800.0 282150.0 555000.0 289650.0 ;
      RECT  591600.0 287550.0 592800.0 289650.0 ;
      RECT  594600.0 282150.0 595800.0 289650.0 ;
      RECT  632400.0 287550.0 633600.0 289650.0 ;
      RECT  635400.0 282150.0 636600.0 289650.0 ;
      RECT  673200.0 287550.0 674400.0 289650.0 ;
      RECT  676200.0 282150.0 677400.0 289650.0 ;
      RECT  714000.0 287550.0 715200.0 289650.0 ;
      RECT  717000.0 282150.0 718200.0 289650.0 ;
      RECT  754800.0 287550.0 756000.0 289650.0 ;
      RECT  757800.0 282150.0 759000.0 289650.0 ;
      RECT  795600.0 287550.0 796800.0 289650.0 ;
      RECT  798600.0 282150.0 799800.0 289650.0 ;
      RECT  836400.0 287550.0 837600.0 289650.0 ;
      RECT  839400.0 282150.0 840600.0 289650.0 ;
      RECT  877200.0 287550.0 878400.0 289650.0 ;
      RECT  880200.0 282150.0 881400.0 289650.0 ;
      RECT  918000.0 287550.0 919200.0 289650.0 ;
      RECT  921000.0 282150.0 922200.0 289650.0 ;
      RECT  958800.0 287550.0 960000.0 289650.0 ;
      RECT  961800.0 282150.0 963000.0 289650.0 ;
      RECT  999600.0 287550.0 1000800.0 289650.0 ;
      RECT  1002600.0 282150.0 1003800.0 289650.0 ;
      RECT  1040400.0 287550.0 1041600.0 289650.0 ;
      RECT  1043400.0 282150.0 1044600.0 289650.0 ;
      RECT  1081200.0 287550.0 1082400.0 289650.0 ;
      RECT  1084200.0 282150.0 1085400.0 289650.0 ;
      RECT  1122000.0 287550.0 1123200.0 289650.0 ;
      RECT  1125000.0 282150.0 1126200.0 289650.0 ;
      RECT  1162800.0 287550.0 1164000.0 289650.0 ;
      RECT  1165800.0 282150.0 1167000.0 289650.0 ;
      RECT  1203600.0 287550.0 1204800.0 289650.0 ;
      RECT  1206600.0 282150.0 1207800.0 289650.0 ;
      RECT  1244400.0 287550.0 1245600.0 289650.0 ;
      RECT  1247400.0 282150.0 1248600.0 289650.0 ;
      RECT  1285200.0 287550.0 1286400.0 289650.0 ;
      RECT  1288200.0 282150.0 1289400.0 289650.0 ;
      RECT  1326000.0 287550.0 1327200.0 289650.0 ;
      RECT  1329000.0 282150.0 1330200.0 289650.0 ;
      RECT  1366800.0 287550.0 1368000.0 289650.0 ;
      RECT  1369800.0 282150.0 1371000.0 289650.0 ;
      RECT  1407600.0 287550.0 1408800.0 289650.0 ;
      RECT  1410600.0 282150.0 1411800.0 289650.0 ;
      RECT  1448400.0 287550.0 1449600.0 289650.0 ;
      RECT  1451400.0 282150.0 1452600.0 289650.0 ;
      RECT  1489200.0 287550.0 1490400.0 289650.0 ;
      RECT  1492200.0 282150.0 1493400.0 289650.0 ;
      RECT  221400.0 169050.0 231600.0 229050.0 ;
      RECT  262200.0 169050.0 272400.0 229050.0 ;
      RECT  303000.0 169050.0 313200.0 229050.0 ;
      RECT  343800.0 169050.0 354000.0 229050.0 ;
      RECT  384600.0 169050.0 394800.0 229050.0 ;
      RECT  425400.0 169050.0 435600.0 229050.0 ;
      RECT  466200.0 169050.0 476400.0 229050.0 ;
      RECT  507000.0 169050.0 517200.0 229050.0 ;
      RECT  547800.0 169050.0 558000.0 229050.0 ;
      RECT  588600.0 169050.0 598800.0 229050.0 ;
      RECT  629400.0 169050.0 639600.0 229050.0 ;
      RECT  670200.0 169050.0 680400.0 229050.0 ;
      RECT  711000.0 169050.0 721200.0 229050.0 ;
      RECT  751800.0 169050.0 762000.0 229050.0 ;
      RECT  792600.0 169050.0 802800.0 229050.0 ;
      RECT  833400.0 169050.0 843600.0 229050.0 ;
      RECT  874200.0 169050.0 884400.0 229050.0 ;
      RECT  915000.0 169050.0 925200.0 229050.0 ;
      RECT  955800.0 169050.0 966000.0 229050.0 ;
      RECT  996600.0 169050.0 1006800.0 229050.0 ;
      RECT  1037400.0 169050.0 1047600.0 229050.0 ;
      RECT  1078200.0 169050.0 1088400.0 229050.0 ;
      RECT  1119000.0 169050.0 1129200.0 229050.0 ;
      RECT  1159800.0 169050.0 1170000.0 229050.0 ;
      RECT  1200600.0 169050.0 1210800.0 229050.0 ;
      RECT  1241400.0 169050.0 1251600.0 229050.0 ;
      RECT  1282200.0 169050.0 1292400.0 229050.0 ;
      RECT  1323000.0 169050.0 1333200.0 229050.0 ;
      RECT  1363800.0 169050.0 1374000.0 229050.0 ;
      RECT  1404600.0 169050.0 1414800.0 229050.0 ;
      RECT  1445400.0 169050.0 1455600.0 229050.0 ;
      RECT  1486200.0 169050.0 1496400.0 229050.0 ;
      RECT  225900.0 226650.0 228600.0 227850.0 ;
      RECT  223200.0 224550.0 224400.0 229050.0 ;
      RECT  266700.0 226650.0 269400.0 227850.0 ;
      RECT  264000.0 224550.0 265200.0 229050.0 ;
      RECT  307500.0 226650.0 310200.0 227850.0 ;
      RECT  304800.0 224550.0 306000.0 229050.0 ;
      RECT  348300.0 226650.0 351000.0 227850.0 ;
      RECT  345600.0 224550.0 346800.0 229050.0 ;
      RECT  389100.0 226650.0 391800.0 227850.0 ;
      RECT  386400.0 224550.0 387600.0 229050.0 ;
      RECT  429900.0 226650.0 432600.0 227850.0 ;
      RECT  427200.0 224550.0 428400.0 229050.0 ;
      RECT  470700.0 226650.0 473400.0 227850.0 ;
      RECT  468000.0 224550.0 469200.0 229050.0 ;
      RECT  511500.0 226650.0 514200.0 227850.0 ;
      RECT  508800.0 224550.0 510000.0 229050.0 ;
      RECT  552300.0 226650.0 555000.0 227850.0 ;
      RECT  549600.0 224550.0 550800.0 229050.0 ;
      RECT  593100.0 226650.0 595800.0 227850.0 ;
      RECT  590400.0 224550.0 591600.0 229050.0 ;
      RECT  633900.0 226650.0 636600.0 227850.0 ;
      RECT  631200.0 224550.0 632400.0 229050.0 ;
      RECT  674700.0 226650.0 677400.0 227850.0 ;
      RECT  672000.0 224550.0 673200.0 229050.0 ;
      RECT  715500.0 226650.0 718200.0 227850.0 ;
      RECT  712800.0 224550.0 714000.0 229050.0 ;
      RECT  756300.0 226650.0 759000.0 227850.0 ;
      RECT  753600.0 224550.0 754800.0 229050.0 ;
      RECT  797100.0 226650.0 799800.0 227850.0 ;
      RECT  794400.0 224550.0 795600.0 229050.0 ;
      RECT  837900.0 226650.0 840600.0 227850.0 ;
      RECT  835200.0 224550.0 836400.0 229050.0 ;
      RECT  878700.0 226650.0 881400.0 227850.0 ;
      RECT  876000.0 224550.0 877200.0 229050.0 ;
      RECT  919500.0 226650.0 922200.0 227850.0 ;
      RECT  916800.0 224550.0 918000.0 229050.0 ;
      RECT  960300.0 226650.0 963000.0 227850.0 ;
      RECT  957600.0 224550.0 958800.0 229050.0 ;
      RECT  1001100.0 226650.0 1003800.0 227850.0 ;
      RECT  998400.0 224550.0 999600.0 229050.0 ;
      RECT  1041900.0 226650.0 1044600.0 227850.0 ;
      RECT  1039200.0 224550.0 1040400.0 229050.0 ;
      RECT  1082700.0 226650.0 1085400.0 227850.0 ;
      RECT  1080000.0 224550.0 1081200.0 229050.0 ;
      RECT  1123500.0 226650.0 1126200.0 227850.0 ;
      RECT  1120800.0 224550.0 1122000.0 229050.0 ;
      RECT  1164300.0 226650.0 1167000.0 227850.0 ;
      RECT  1161600.0 224550.0 1162800.0 229050.0 ;
      RECT  1205100.0 226650.0 1207800.0 227850.0 ;
      RECT  1202400.0 224550.0 1203600.0 229050.0 ;
      RECT  1245900.0 226650.0 1248600.0 227850.0 ;
      RECT  1243200.0 224550.0 1244400.0 229050.0 ;
      RECT  1286700.0 226650.0 1289400.0 227850.0 ;
      RECT  1284000.0 224550.0 1285200.0 229050.0 ;
      RECT  1327500.0 226650.0 1330200.0 227850.0 ;
      RECT  1324800.0 224550.0 1326000.0 229050.0 ;
      RECT  1368300.0 226650.0 1371000.0 227850.0 ;
      RECT  1365600.0 224550.0 1366800.0 229050.0 ;
      RECT  1409100.0 226650.0 1411800.0 227850.0 ;
      RECT  1406400.0 224550.0 1407600.0 229050.0 ;
      RECT  1449900.0 226650.0 1452600.0 227850.0 ;
      RECT  1447200.0 224550.0 1448400.0 229050.0 ;
      RECT  1490700.0 226650.0 1493400.0 227850.0 ;
      RECT  1488000.0 224550.0 1489200.0 229050.0 ;
      RECT  231000.0 169050.0 232200.0 229050.0 ;
      RECT  271800.0 169050.0 273000.0 229050.0 ;
      RECT  312600.0 169050.0 313800.0 229050.0 ;
      RECT  353400.0 169050.0 354600.0 229050.0 ;
      RECT  394200.0 169050.0 395400.0 229050.0 ;
      RECT  435000.0 169050.0 436200.0 229050.0 ;
      RECT  475800.0 169050.0 477000.0 229050.0 ;
      RECT  516600.0 169050.0 517800.0 229050.0 ;
      RECT  557400.0 169050.0 558600.0 229050.0 ;
      RECT  598200.0 169050.0 599400.0 229050.0 ;
      RECT  639000.0 169050.0 640200.0 229050.0 ;
      RECT  679800.0 169050.0 681000.0 229050.0 ;
      RECT  720600.0 169050.0 721800.0 229050.0 ;
      RECT  761400.0 169050.0 762600.0 229050.0 ;
      RECT  802200.0 169050.0 803400.0 229050.0 ;
      RECT  843000.0 169050.0 844200.0 229050.0 ;
      RECT  883800.0 169050.0 885000.0 229050.0 ;
      RECT  924600.0 169050.0 925800.0 229050.0 ;
      RECT  965400.0 169050.0 966600.0 229050.0 ;
      RECT  1006200.0 169050.0 1007400.0 229050.0 ;
      RECT  1047000.0 169050.0 1048200.0 229050.0 ;
      RECT  1087800.0 169050.0 1089000.0 229050.0 ;
      RECT  1128600.0 169050.0 1129800.0 229050.0 ;
      RECT  1169400.0 169050.0 1170600.0 229050.0 ;
      RECT  1210200.0 169050.0 1211400.0 229050.0 ;
      RECT  1251000.0 169050.0 1252200.0 229050.0 ;
      RECT  1291800.0 169050.0 1293000.0 229050.0 ;
      RECT  1332600.0 169050.0 1333800.0 229050.0 ;
      RECT  1373400.0 169050.0 1374600.0 229050.0 ;
      RECT  1414200.0 169050.0 1415400.0 229050.0 ;
      RECT  1455000.0 169050.0 1456200.0 229050.0 ;
      RECT  1495800.0 169050.0 1497000.0 229050.0 ;
      RECT  221400.0 169050.0 231600.0 147150.0 ;
      RECT  262200.0 169050.0 272400.0 147150.0 ;
      RECT  303000.0 169050.0 313200.0 147150.0 ;
      RECT  343800.0 169050.0 354000.0 147150.0 ;
      RECT  384600.0 169050.0 394800.0 147150.0 ;
      RECT  425400.0 169050.0 435600.0 147150.0 ;
      RECT  466200.0 169050.0 476400.0 147150.0 ;
      RECT  507000.0 169050.0 517200.0 147150.0 ;
      RECT  547800.0 169050.0 558000.0 147150.0 ;
      RECT  588600.0 169050.0 598800.0 147150.0 ;
      RECT  629400.0 169050.0 639600.0 147150.0 ;
      RECT  670200.0 169050.0 680400.0 147150.0 ;
      RECT  711000.0 169050.0 721200.0 147150.0 ;
      RECT  751800.0 169050.0 762000.0 147150.0 ;
      RECT  792600.0 169050.0 802800.0 147150.0 ;
      RECT  833400.0 169050.0 843600.0 147150.0 ;
      RECT  874200.0 169050.0 884400.0 147150.0 ;
      RECT  915000.0 169050.0 925200.0 147150.0 ;
      RECT  955800.0 169050.0 966000.0 147150.0 ;
      RECT  996600.0 169050.0 1006800.0 147150.0 ;
      RECT  1037400.0 169050.0 1047600.0 147150.0 ;
      RECT  1078200.0 169050.0 1088400.0 147150.0 ;
      RECT  1119000.0 169050.0 1129200.0 147150.0 ;
      RECT  1159800.0 169050.0 1170000.0 147150.0 ;
      RECT  1200600.0 169050.0 1210800.0 147150.0 ;
      RECT  1241400.0 169050.0 1251600.0 147150.0 ;
      RECT  1282200.0 169050.0 1292400.0 147150.0 ;
      RECT  1323000.0 169050.0 1333200.0 147150.0 ;
      RECT  1363800.0 169050.0 1374000.0 147150.0 ;
      RECT  1404600.0 169050.0 1414800.0 147150.0 ;
      RECT  1445400.0 169050.0 1455600.0 147150.0 ;
      RECT  1486200.0 169050.0 1496400.0 147150.0 ;
      RECT  225900.0 154050.0 227100.0 147150.0 ;
      RECT  266700.0 154050.0 267900.0 147150.0 ;
      RECT  307500.0 154050.0 308700.0 147150.0 ;
      RECT  348300.0 154050.0 349500.0 147150.0 ;
      RECT  389100.0 154050.0 390300.0 147150.0 ;
      RECT  429900.0 154050.0 431100.0 147150.0 ;
      RECT  470700.0 154050.0 471900.0 147150.0 ;
      RECT  511500.0 154050.0 512700.0 147150.0 ;
      RECT  552300.0 154050.0 553500.0 147150.0 ;
      RECT  593100.0 154050.0 594300.0 147150.0 ;
      RECT  633900.0 154050.0 635100.0 147150.0 ;
      RECT  674700.0 154050.0 675900.0 147150.0 ;
      RECT  715500.0 154050.0 716700.0 147150.0 ;
      RECT  756300.0 154050.0 757500.0 147150.0 ;
      RECT  797100.0 154050.0 798300.0 147150.0 ;
      RECT  837900.0 154050.0 839100.0 147150.0 ;
      RECT  878700.0 154050.0 879900.0 147150.0 ;
      RECT  919500.0 154050.0 920700.0 147150.0 ;
      RECT  960300.0 154050.0 961500.0 147150.0 ;
      RECT  1001100.0 154050.0 1002300.0 147150.0 ;
      RECT  1041900.0 154050.0 1043100.0 147150.0 ;
      RECT  1082700.0 154050.0 1083900.0 147150.0 ;
      RECT  1123500.0 154050.0 1124700.0 147150.0 ;
      RECT  1164300.0 154050.0 1165500.0 147150.0 ;
      RECT  1205100.0 154050.0 1206300.0 147150.0 ;
      RECT  1245900.0 154050.0 1247100.0 147150.0 ;
      RECT  1286700.0 154050.0 1287900.0 147150.0 ;
      RECT  1327500.0 154050.0 1328700.0 147150.0 ;
      RECT  1368300.0 154050.0 1369500.0 147150.0 ;
      RECT  1409100.0 154050.0 1410300.0 147150.0 ;
      RECT  1449900.0 154050.0 1451100.0 147150.0 ;
      RECT  1490700.0 154050.0 1491900.0 147150.0 ;
      RECT  225900.0 169050.0 227100.0 167550.0 ;
      RECT  266700.0 169050.0 267900.0 167550.0 ;
      RECT  307500.0 169050.0 308700.0 167550.0 ;
      RECT  348300.0 169050.0 349500.0 167550.0 ;
      RECT  389100.0 169050.0 390300.0 167550.0 ;
      RECT  429900.0 169050.0 431100.0 167550.0 ;
      RECT  470700.0 169050.0 471900.0 167550.0 ;
      RECT  511500.0 169050.0 512700.0 167550.0 ;
      RECT  552300.0 169050.0 553500.0 167550.0 ;
      RECT  593100.0 169050.0 594300.0 167550.0 ;
      RECT  633900.0 169050.0 635100.0 167550.0 ;
      RECT  674700.0 169050.0 675900.0 167550.0 ;
      RECT  715500.0 169050.0 716700.0 167550.0 ;
      RECT  756300.0 169050.0 757500.0 167550.0 ;
      RECT  797100.0 169050.0 798300.0 167550.0 ;
      RECT  837900.0 169050.0 839100.0 167550.0 ;
      RECT  878700.0 169050.0 879900.0 167550.0 ;
      RECT  919500.0 169050.0 920700.0 167550.0 ;
      RECT  960300.0 169050.0 961500.0 167550.0 ;
      RECT  1001100.0 169050.0 1002300.0 167550.0 ;
      RECT  1041900.0 169050.0 1043100.0 167550.0 ;
      RECT  1082700.0 169050.0 1083900.0 167550.0 ;
      RECT  1123500.0 169050.0 1124700.0 167550.0 ;
      RECT  1164300.0 169050.0 1165500.0 167550.0 ;
      RECT  1205100.0 169050.0 1206300.0 167550.0 ;
      RECT  1245900.0 169050.0 1247100.0 167550.0 ;
      RECT  1286700.0 169050.0 1287900.0 167550.0 ;
      RECT  1327500.0 169050.0 1328700.0 167550.0 ;
      RECT  1368300.0 169050.0 1369500.0 167550.0 ;
      RECT  1409100.0 169050.0 1410300.0 167550.0 ;
      RECT  1449900.0 169050.0 1451100.0 167550.0 ;
      RECT  1490700.0 169050.0 1491900.0 167550.0 ;
      RECT  59100.0 158400.0 60000.0 2145600.0 ;
      RECT  61200.0 158400.0 62100.0 2145600.0 ;
      RECT  63300.0 158400.0 64200.0 2145600.0 ;
      RECT  65400.0 158400.0 66300.0 2145600.0 ;
      RECT  67500.0 158400.0 68400.0 2145600.0 ;
      RECT  69600.0 158400.0 70500.0 2145600.0 ;
      RECT  71700.0 158400.0 72600.0 2145600.0 ;
      RECT  73800.0 158400.0 74700.0 2145600.0 ;
      RECT  75900.0 158400.0 76800.0 2145600.0 ;
      RECT  78000.0 158400.0 78900.0 2145600.0 ;
      RECT  80100.0 158400.0 81000.0 2145600.0 ;
      RECT  82200.0 158400.0 83100.0 2145600.0 ;
      RECT  84300.0 158400.0 85200.0 2145600.0 ;
      RECT  86400.0 158400.0 87300.0 2145600.0 ;
      RECT  88500.0 158400.0 89400.0 2145600.0 ;
      RECT  90600.0 158400.0 91500.0 2145600.0 ;
      RECT  122700.0 158400.0 121800.0 211800.0 ;
      RECT  119700.0 158400.0 118800.0 211800.0 ;
      RECT  128700.0 158400.0 127800.0 211800.0 ;
      RECT  125700.0 158400.0 124800.0 211800.0 ;
      RECT  112350.0 165750.0 111450.0 166650.0 ;
      RECT  109950.0 165750.0 109050.0 166650.0 ;
      RECT  112350.0 166200.0 111450.0 169050.0 ;
      RECT  111900.0 165750.0 109500.0 166650.0 ;
      RECT  109950.0 161550.0 109050.0 166200.0 ;
      RECT  112500.0 169050.0 111300.0 170250.0 ;
      RECT  110100.0 160350.0 108900.0 161550.0 ;
      RECT  108900.0 165600.0 110100.0 166800.0 ;
      RECT  112350.0 178650.0 111450.0 177750.0 ;
      RECT  109950.0 178650.0 109050.0 177750.0 ;
      RECT  112350.0 178200.0 111450.0 175350.0 ;
      RECT  111900.0 178650.0 109500.0 177750.0 ;
      RECT  109950.0 182850.0 109050.0 178200.0 ;
      RECT  112500.0 175350.0 111300.0 174150.0 ;
      RECT  110100.0 184050.0 108900.0 182850.0 ;
      RECT  108900.0 178800.0 110100.0 177600.0 ;
      RECT  112350.0 193350.0 111450.0 194250.0 ;
      RECT  109950.0 193350.0 109050.0 194250.0 ;
      RECT  112350.0 193800.0 111450.0 196650.0 ;
      RECT  111900.0 193350.0 109500.0 194250.0 ;
      RECT  109950.0 189150.0 109050.0 193800.0 ;
      RECT  112500.0 196650.0 111300.0 197850.0 ;
      RECT  110100.0 187950.0 108900.0 189150.0 ;
      RECT  108900.0 193200.0 110100.0 194400.0 ;
      RECT  112350.0 206250.0 111450.0 205350.0 ;
      RECT  109950.0 206250.0 109050.0 205350.0 ;
      RECT  112350.0 205800.0 111450.0 202950.0 ;
      RECT  111900.0 206250.0 109500.0 205350.0 ;
      RECT  109950.0 210450.0 109050.0 205800.0 ;
      RECT  112500.0 202950.0 111300.0 201750.0 ;
      RECT  110100.0 211650.0 108900.0 210450.0 ;
      RECT  108900.0 206400.0 110100.0 205200.0 ;
      RECT  127650.0 168900.0 128850.0 170100.0 ;
      RECT  146250.0 164400.0 147450.0 165600.0 ;
      RECT  124650.0 182700.0 125850.0 183900.0 ;
      RECT  143250.0 178800.0 144450.0 180000.0 ;
      RECT  146250.0 187500.0 147450.0 188700.0 ;
      RECT  121650.0 187500.0 122850.0 188700.0 ;
      RECT  143250.0 201300.0 144450.0 202500.0 ;
      RECT  118650.0 201300.0 119850.0 202500.0 ;
      RECT  127650.0 165600.0 128850.0 166800.0 ;
      RECT  124650.0 162900.0 125850.0 164100.0 ;
      RECT  121650.0 177600.0 122850.0 178800.0 ;
      RECT  124650.0 180300.0 125850.0 181500.0 ;
      RECT  127650.0 193200.0 128850.0 194400.0 ;
      RECT  118650.0 190500.0 119850.0 191700.0 ;
      RECT  121650.0 205200.0 122850.0 206400.0 ;
      RECT  118650.0 207900.0 119850.0 209100.0 ;
      RECT  147300.0 158400.0 146400.0 211800.0 ;
      RECT  144300.0 158400.0 143400.0 211800.0 ;
      RECT  122700.0 213600.0 121800.0 267000.0 ;
      RECT  119700.0 213600.0 118800.0 267000.0 ;
      RECT  128700.0 213600.0 127800.0 267000.0 ;
      RECT  125700.0 213600.0 124800.0 267000.0 ;
      RECT  112350.0 220950.0 111450.0 221850.0 ;
      RECT  109950.0 220950.0 109050.0 221850.0 ;
      RECT  112350.0 221400.0 111450.0 224250.0 ;
      RECT  111900.0 220950.0 109500.0 221850.0 ;
      RECT  109950.0 216750.0 109050.0 221400.0 ;
      RECT  112500.0 224250.0 111300.0 225450.0 ;
      RECT  110100.0 215550.0 108900.0 216750.0 ;
      RECT  108900.0 220800.0 110100.0 222000.0 ;
      RECT  112350.0 233850.0 111450.0 232950.0 ;
      RECT  109950.0 233850.0 109050.0 232950.0 ;
      RECT  112350.0 233400.0 111450.0 230550.0 ;
      RECT  111900.0 233850.0 109500.0 232950.0 ;
      RECT  109950.0 238050.0 109050.0 233400.0 ;
      RECT  112500.0 230550.0 111300.0 229350.0 ;
      RECT  110100.0 239250.0 108900.0 238050.0 ;
      RECT  108900.0 234000.0 110100.0 232800.0 ;
      RECT  112350.0 248550.0 111450.0 249450.0 ;
      RECT  109950.0 248550.0 109050.0 249450.0 ;
      RECT  112350.0 249000.0 111450.0 251850.0 ;
      RECT  111900.0 248550.0 109500.0 249450.0 ;
      RECT  109950.0 244350.0 109050.0 249000.0 ;
      RECT  112500.0 251850.0 111300.0 253050.0 ;
      RECT  110100.0 243150.0 108900.0 244350.0 ;
      RECT  108900.0 248400.0 110100.0 249600.0 ;
      RECT  112350.0 261450.0 111450.0 260550.0 ;
      RECT  109950.0 261450.0 109050.0 260550.0 ;
      RECT  112350.0 261000.0 111450.0 258150.0 ;
      RECT  111900.0 261450.0 109500.0 260550.0 ;
      RECT  109950.0 265650.0 109050.0 261000.0 ;
      RECT  112500.0 258150.0 111300.0 256950.0 ;
      RECT  110100.0 266850.0 108900.0 265650.0 ;
      RECT  108900.0 261600.0 110100.0 260400.0 ;
      RECT  127650.0 224100.0 128850.0 225300.0 ;
      RECT  146250.0 219600.0 147450.0 220800.0 ;
      RECT  124650.0 237900.0 125850.0 239100.0 ;
      RECT  143250.0 234000.0 144450.0 235200.0 ;
      RECT  146250.0 242700.0 147450.0 243900.0 ;
      RECT  121650.0 242700.0 122850.0 243900.0 ;
      RECT  143250.0 256500.0 144450.0 257700.0 ;
      RECT  118650.0 256500.0 119850.0 257700.0 ;
      RECT  127650.0 220800.0 128850.0 222000.0 ;
      RECT  124650.0 218100.0 125850.0 219300.0 ;
      RECT  121650.0 232800.0 122850.0 234000.0 ;
      RECT  124650.0 235500.0 125850.0 236700.0 ;
      RECT  127650.0 248400.0 128850.0 249600.0 ;
      RECT  118650.0 245700.0 119850.0 246900.0 ;
      RECT  121650.0 260400.0 122850.0 261600.0 ;
      RECT  118650.0 263100.0 119850.0 264300.0 ;
      RECT  147300.0 213600.0 146400.0 267000.0 ;
      RECT  144300.0 213600.0 143400.0 267000.0 ;
      RECT  129900.0 268800.0 129000.0 377400.0 ;
      RECT  126900.0 268800.0 126000.0 377400.0 ;
      RECT  123900.0 268800.0 123000.0 377400.0 ;
      RECT  135900.0 268800.0 135000.0 377400.0 ;
      RECT  132900.0 268800.0 132000.0 377400.0 ;
      RECT  120900.0 268800.0 120000.0 377400.0 ;
      RECT  108750.0 271950.0 107850.0 279450.0 ;
      RECT  113550.0 276900.0 112650.0 277800.0 ;
      RECT  108750.0 276900.0 107850.0 277800.0 ;
      RECT  113550.0 277350.0 112650.0 279450.0 ;
      RECT  113100.0 276900.0 108300.0 277800.0 ;
      RECT  108750.0 271950.0 107850.0 277350.0 ;
      RECT  113700.0 279450.0 112500.0 280650.0 ;
      RECT  108900.0 279450.0 107700.0 280650.0 ;
      RECT  108900.0 270750.0 107700.0 271950.0 ;
      RECT  108900.0 276750.0 107700.0 277950.0 ;
      RECT  108750.0 293250.0 107850.0 285750.0 ;
      RECT  113550.0 288300.0 112650.0 287400.0 ;
      RECT  108750.0 288300.0 107850.0 287400.0 ;
      RECT  113550.0 287850.0 112650.0 285750.0 ;
      RECT  113100.0 288300.0 108300.0 287400.0 ;
      RECT  108750.0 293250.0 107850.0 287850.0 ;
      RECT  113700.0 285750.0 112500.0 284550.0 ;
      RECT  108900.0 285750.0 107700.0 284550.0 ;
      RECT  108900.0 294450.0 107700.0 293250.0 ;
      RECT  108900.0 288450.0 107700.0 287250.0 ;
      RECT  108750.0 299550.0 107850.0 307050.0 ;
      RECT  113550.0 304500.0 112650.0 305400.0 ;
      RECT  108750.0 304500.0 107850.0 305400.0 ;
      RECT  113550.0 304950.0 112650.0 307050.0 ;
      RECT  113100.0 304500.0 108300.0 305400.0 ;
      RECT  108750.0 299550.0 107850.0 304950.0 ;
      RECT  113700.0 307050.0 112500.0 308250.0 ;
      RECT  108900.0 307050.0 107700.0 308250.0 ;
      RECT  108900.0 298350.0 107700.0 299550.0 ;
      RECT  108900.0 304350.0 107700.0 305550.0 ;
      RECT  108750.0 320850.0 107850.0 313350.0 ;
      RECT  113550.0 315900.0 112650.0 315000.0 ;
      RECT  108750.0 315900.0 107850.0 315000.0 ;
      RECT  113550.0 315450.0 112650.0 313350.0 ;
      RECT  113100.0 315900.0 108300.0 315000.0 ;
      RECT  108750.0 320850.0 107850.0 315450.0 ;
      RECT  113700.0 313350.0 112500.0 312150.0 ;
      RECT  108900.0 313350.0 107700.0 312150.0 ;
      RECT  108900.0 322050.0 107700.0 320850.0 ;
      RECT  108900.0 316050.0 107700.0 314850.0 ;
      RECT  108750.0 327150.0 107850.0 334650.0 ;
      RECT  113550.0 332100.0 112650.0 333000.0 ;
      RECT  108750.0 332100.0 107850.0 333000.0 ;
      RECT  113550.0 332550.0 112650.0 334650.0 ;
      RECT  113100.0 332100.0 108300.0 333000.0 ;
      RECT  108750.0 327150.0 107850.0 332550.0 ;
      RECT  113700.0 334650.0 112500.0 335850.0 ;
      RECT  108900.0 334650.0 107700.0 335850.0 ;
      RECT  108900.0 325950.0 107700.0 327150.0 ;
      RECT  108900.0 331950.0 107700.0 333150.0 ;
      RECT  108750.0 348450.0 107850.0 340950.0 ;
      RECT  113550.0 343500.0 112650.0 342600.0 ;
      RECT  108750.0 343500.0 107850.0 342600.0 ;
      RECT  113550.0 343050.0 112650.0 340950.0 ;
      RECT  113100.0 343500.0 108300.0 342600.0 ;
      RECT  108750.0 348450.0 107850.0 343050.0 ;
      RECT  113700.0 340950.0 112500.0 339750.0 ;
      RECT  108900.0 340950.0 107700.0 339750.0 ;
      RECT  108900.0 349650.0 107700.0 348450.0 ;
      RECT  108900.0 343650.0 107700.0 342450.0 ;
      RECT  108750.0 354750.0 107850.0 362250.0 ;
      RECT  113550.0 359700.0 112650.0 360600.0 ;
      RECT  108750.0 359700.0 107850.0 360600.0 ;
      RECT  113550.0 360150.0 112650.0 362250.0 ;
      RECT  113100.0 359700.0 108300.0 360600.0 ;
      RECT  108750.0 354750.0 107850.0 360150.0 ;
      RECT  113700.0 362250.0 112500.0 363450.0 ;
      RECT  108900.0 362250.0 107700.0 363450.0 ;
      RECT  108900.0 353550.0 107700.0 354750.0 ;
      RECT  108900.0 359550.0 107700.0 360750.0 ;
      RECT  108750.0 376050.0 107850.0 368550.0 ;
      RECT  113550.0 371100.0 112650.0 370200.0 ;
      RECT  108750.0 371100.0 107850.0 370200.0 ;
      RECT  113550.0 370650.0 112650.0 368550.0 ;
      RECT  113100.0 371100.0 108300.0 370200.0 ;
      RECT  108750.0 376050.0 107850.0 370650.0 ;
      RECT  113700.0 368550.0 112500.0 367350.0 ;
      RECT  108900.0 368550.0 107700.0 367350.0 ;
      RECT  108900.0 377250.0 107700.0 376050.0 ;
      RECT  108900.0 371250.0 107700.0 370050.0 ;
      RECT  134850.0 279300.0 136050.0 280500.0 ;
      RECT  156450.0 274800.0 157650.0 276000.0 ;
      RECT  131850.0 293100.0 133050.0 294300.0 ;
      RECT  153450.0 289200.0 154650.0 290400.0 ;
      RECT  128850.0 306900.0 130050.0 308100.0 ;
      RECT  150450.0 302400.0 151650.0 303600.0 ;
      RECT  156450.0 311700.0 157650.0 312900.0 ;
      RECT  125850.0 311700.0 127050.0 312900.0 ;
      RECT  153450.0 325500.0 154650.0 326700.0 ;
      RECT  122850.0 325500.0 124050.0 326700.0 ;
      RECT  150450.0 339300.0 151650.0 340500.0 ;
      RECT  119850.0 339300.0 121050.0 340500.0 ;
      RECT  134850.0 276750.0 136050.0 277950.0 ;
      RECT  131850.0 274800.0 133050.0 276000.0 ;
      RECT  128850.0 272850.0 130050.0 274050.0 ;
      RECT  125850.0 287250.0 127050.0 288450.0 ;
      RECT  131850.0 289200.0 133050.0 290400.0 ;
      RECT  128850.0 291150.0 130050.0 292350.0 ;
      RECT  134850.0 304350.0 136050.0 305550.0 ;
      RECT  122850.0 302400.0 124050.0 303600.0 ;
      RECT  128850.0 300450.0 130050.0 301650.0 ;
      RECT  125850.0 314850.0 127050.0 316050.0 ;
      RECT  122850.0 316800.0 124050.0 318000.0 ;
      RECT  128850.0 318750.0 130050.0 319950.0 ;
      RECT  134850.0 331950.0 136050.0 333150.0 ;
      RECT  131850.0 330000.0 133050.0 331200.0 ;
      RECT  119850.0 328050.0 121050.0 329250.0 ;
      RECT  125850.0 342450.0 127050.0 343650.0 ;
      RECT  131850.0 344400.0 133050.0 345600.0 ;
      RECT  119850.0 346350.0 121050.0 347550.0 ;
      RECT  134850.0 359550.0 136050.0 360750.0 ;
      RECT  122850.0 357600.0 124050.0 358800.0 ;
      RECT  119850.0 355650.0 121050.0 356850.0 ;
      RECT  125850.0 370050.0 127050.0 371250.0 ;
      RECT  122850.0 372000.0 124050.0 373200.0 ;
      RECT  119850.0 373950.0 121050.0 375150.0 ;
      RECT  157500.0 268800.0 156600.0 377400.0 ;
      RECT  154500.0 268800.0 153600.0 377400.0 ;
      RECT  151500.0 268800.0 150600.0 377400.0 ;
      RECT  101850.0 382350.0 102750.0 389850.0 ;
      RECT  97050.0 387300.0 97950.0 388200.0 ;
      RECT  101850.0 387300.0 102750.0 388200.0 ;
      RECT  97050.0 387750.0 97950.0 389850.0 ;
      RECT  97500.0 387300.0 102300.0 388200.0 ;
      RECT  101850.0 382350.0 102750.0 387750.0 ;
      RECT  96900.0 389850.0 98100.0 391050.0 ;
      RECT  101700.0 389850.0 102900.0 391050.0 ;
      RECT  101700.0 381150.0 102900.0 382350.0 ;
      RECT  101700.0 387150.0 102900.0 388350.0 ;
      RECT  101850.0 403650.0 102750.0 396150.0 ;
      RECT  97050.0 398700.0 97950.0 397800.0 ;
      RECT  101850.0 398700.0 102750.0 397800.0 ;
      RECT  97050.0 398250.0 97950.0 396150.0 ;
      RECT  97500.0 398700.0 102300.0 397800.0 ;
      RECT  101850.0 403650.0 102750.0 398250.0 ;
      RECT  96900.0 396150.0 98100.0 394950.0 ;
      RECT  101700.0 396150.0 102900.0 394950.0 ;
      RECT  101700.0 404850.0 102900.0 403650.0 ;
      RECT  101700.0 398850.0 102900.0 397650.0 ;
      RECT  101850.0 409950.0 102750.0 417450.0 ;
      RECT  97050.0 414900.0 97950.0 415800.0 ;
      RECT  101850.0 414900.0 102750.0 415800.0 ;
      RECT  97050.0 415350.0 97950.0 417450.0 ;
      RECT  97500.0 414900.0 102300.0 415800.0 ;
      RECT  101850.0 409950.0 102750.0 415350.0 ;
      RECT  96900.0 417450.0 98100.0 418650.0 ;
      RECT  101700.0 417450.0 102900.0 418650.0 ;
      RECT  101700.0 408750.0 102900.0 409950.0 ;
      RECT  101700.0 414750.0 102900.0 415950.0 ;
      RECT  101850.0 431250.0 102750.0 423750.0 ;
      RECT  97050.0 426300.0 97950.0 425400.0 ;
      RECT  101850.0 426300.0 102750.0 425400.0 ;
      RECT  97050.0 425850.0 97950.0 423750.0 ;
      RECT  97500.0 426300.0 102300.0 425400.0 ;
      RECT  101850.0 431250.0 102750.0 425850.0 ;
      RECT  96900.0 423750.0 98100.0 422550.0 ;
      RECT  101700.0 423750.0 102900.0 422550.0 ;
      RECT  101700.0 432450.0 102900.0 431250.0 ;
      RECT  101700.0 426450.0 102900.0 425250.0 ;
      RECT  101850.0 437550.0 102750.0 445050.0 ;
      RECT  97050.0 442500.0 97950.0 443400.0 ;
      RECT  101850.0 442500.0 102750.0 443400.0 ;
      RECT  97050.0 442950.0 97950.0 445050.0 ;
      RECT  97500.0 442500.0 102300.0 443400.0 ;
      RECT  101850.0 437550.0 102750.0 442950.0 ;
      RECT  96900.0 445050.0 98100.0 446250.0 ;
      RECT  101700.0 445050.0 102900.0 446250.0 ;
      RECT  101700.0 436350.0 102900.0 437550.0 ;
      RECT  101700.0 442350.0 102900.0 443550.0 ;
      RECT  101850.0 458850.0 102750.0 451350.0 ;
      RECT  97050.0 453900.0 97950.0 453000.0 ;
      RECT  101850.0 453900.0 102750.0 453000.0 ;
      RECT  97050.0 453450.0 97950.0 451350.0 ;
      RECT  97500.0 453900.0 102300.0 453000.0 ;
      RECT  101850.0 458850.0 102750.0 453450.0 ;
      RECT  96900.0 451350.0 98100.0 450150.0 ;
      RECT  101700.0 451350.0 102900.0 450150.0 ;
      RECT  101700.0 460050.0 102900.0 458850.0 ;
      RECT  101700.0 454050.0 102900.0 452850.0 ;
      RECT  101850.0 465150.0 102750.0 472650.0 ;
      RECT  97050.0 470100.0 97950.0 471000.0 ;
      RECT  101850.0 470100.0 102750.0 471000.0 ;
      RECT  97050.0 470550.0 97950.0 472650.0 ;
      RECT  97500.0 470100.0 102300.0 471000.0 ;
      RECT  101850.0 465150.0 102750.0 470550.0 ;
      RECT  96900.0 472650.0 98100.0 473850.0 ;
      RECT  101700.0 472650.0 102900.0 473850.0 ;
      RECT  101700.0 463950.0 102900.0 465150.0 ;
      RECT  101700.0 469950.0 102900.0 471150.0 ;
      RECT  101850.0 486450.0 102750.0 478950.0 ;
      RECT  97050.0 481500.0 97950.0 480600.0 ;
      RECT  101850.0 481500.0 102750.0 480600.0 ;
      RECT  97050.0 481050.0 97950.0 478950.0 ;
      RECT  97500.0 481500.0 102300.0 480600.0 ;
      RECT  101850.0 486450.0 102750.0 481050.0 ;
      RECT  96900.0 478950.0 98100.0 477750.0 ;
      RECT  101700.0 478950.0 102900.0 477750.0 ;
      RECT  101700.0 487650.0 102900.0 486450.0 ;
      RECT  101700.0 481650.0 102900.0 480450.0 ;
      RECT  101850.0 492750.0 102750.0 500250.0 ;
      RECT  97050.0 497700.0 97950.0 498600.0 ;
      RECT  101850.0 497700.0 102750.0 498600.0 ;
      RECT  97050.0 498150.0 97950.0 500250.0 ;
      RECT  97500.0 497700.0 102300.0 498600.0 ;
      RECT  101850.0 492750.0 102750.0 498150.0 ;
      RECT  96900.0 500250.0 98100.0 501450.0 ;
      RECT  101700.0 500250.0 102900.0 501450.0 ;
      RECT  101700.0 491550.0 102900.0 492750.0 ;
      RECT  101700.0 497550.0 102900.0 498750.0 ;
      RECT  101850.0 514050.0 102750.0 506550.0 ;
      RECT  97050.0 509100.0 97950.0 508200.0 ;
      RECT  101850.0 509100.0 102750.0 508200.0 ;
      RECT  97050.0 508650.0 97950.0 506550.0 ;
      RECT  97500.0 509100.0 102300.0 508200.0 ;
      RECT  101850.0 514050.0 102750.0 508650.0 ;
      RECT  96900.0 506550.0 98100.0 505350.0 ;
      RECT  101700.0 506550.0 102900.0 505350.0 ;
      RECT  101700.0 515250.0 102900.0 514050.0 ;
      RECT  101700.0 509250.0 102900.0 508050.0 ;
      RECT  101850.0 520350.0 102750.0 527850.0 ;
      RECT  97050.0 525300.0 97950.0 526200.0 ;
      RECT  101850.0 525300.0 102750.0 526200.0 ;
      RECT  97050.0 525750.0 97950.0 527850.0 ;
      RECT  97500.0 525300.0 102300.0 526200.0 ;
      RECT  101850.0 520350.0 102750.0 525750.0 ;
      RECT  96900.0 527850.0 98100.0 529050.0 ;
      RECT  101700.0 527850.0 102900.0 529050.0 ;
      RECT  101700.0 519150.0 102900.0 520350.0 ;
      RECT  101700.0 525150.0 102900.0 526350.0 ;
      RECT  101850.0 541650.0 102750.0 534150.0 ;
      RECT  97050.0 536700.0 97950.0 535800.0 ;
      RECT  101850.0 536700.0 102750.0 535800.0 ;
      RECT  97050.0 536250.0 97950.0 534150.0 ;
      RECT  97500.0 536700.0 102300.0 535800.0 ;
      RECT  101850.0 541650.0 102750.0 536250.0 ;
      RECT  96900.0 534150.0 98100.0 532950.0 ;
      RECT  101700.0 534150.0 102900.0 532950.0 ;
      RECT  101700.0 542850.0 102900.0 541650.0 ;
      RECT  101700.0 536850.0 102900.0 535650.0 ;
      RECT  101850.0 547950.0 102750.0 555450.0 ;
      RECT  97050.0 552900.0 97950.0 553800.0 ;
      RECT  101850.0 552900.0 102750.0 553800.0 ;
      RECT  97050.0 553350.0 97950.0 555450.0 ;
      RECT  97500.0 552900.0 102300.0 553800.0 ;
      RECT  101850.0 547950.0 102750.0 553350.0 ;
      RECT  96900.0 555450.0 98100.0 556650.0 ;
      RECT  101700.0 555450.0 102900.0 556650.0 ;
      RECT  101700.0 546750.0 102900.0 547950.0 ;
      RECT  101700.0 552750.0 102900.0 553950.0 ;
      RECT  101850.0 569250.0 102750.0 561750.0 ;
      RECT  97050.0 564300.0 97950.0 563400.0 ;
      RECT  101850.0 564300.0 102750.0 563400.0 ;
      RECT  97050.0 563850.0 97950.0 561750.0 ;
      RECT  97500.0 564300.0 102300.0 563400.0 ;
      RECT  101850.0 569250.0 102750.0 563850.0 ;
      RECT  96900.0 561750.0 98100.0 560550.0 ;
      RECT  101700.0 561750.0 102900.0 560550.0 ;
      RECT  101700.0 570450.0 102900.0 569250.0 ;
      RECT  101700.0 564450.0 102900.0 563250.0 ;
      RECT  101850.0 575550.0 102750.0 583050.0 ;
      RECT  97050.0 580500.0 97950.0 581400.0 ;
      RECT  101850.0 580500.0 102750.0 581400.0 ;
      RECT  97050.0 580950.0 97950.0 583050.0 ;
      RECT  97500.0 580500.0 102300.0 581400.0 ;
      RECT  101850.0 575550.0 102750.0 580950.0 ;
      RECT  96900.0 583050.0 98100.0 584250.0 ;
      RECT  101700.0 583050.0 102900.0 584250.0 ;
      RECT  101700.0 574350.0 102900.0 575550.0 ;
      RECT  101700.0 580350.0 102900.0 581550.0 ;
      RECT  101850.0 596850.0 102750.0 589350.0 ;
      RECT  97050.0 591900.0 97950.0 591000.0 ;
      RECT  101850.0 591900.0 102750.0 591000.0 ;
      RECT  97050.0 591450.0 97950.0 589350.0 ;
      RECT  97500.0 591900.0 102300.0 591000.0 ;
      RECT  101850.0 596850.0 102750.0 591450.0 ;
      RECT  96900.0 589350.0 98100.0 588150.0 ;
      RECT  101700.0 589350.0 102900.0 588150.0 ;
      RECT  101700.0 598050.0 102900.0 596850.0 ;
      RECT  101700.0 592050.0 102900.0 590850.0 ;
      RECT  101850.0 603150.0 102750.0 610650.0 ;
      RECT  97050.0 608100.0 97950.0 609000.0 ;
      RECT  101850.0 608100.0 102750.0 609000.0 ;
      RECT  97050.0 608550.0 97950.0 610650.0 ;
      RECT  97500.0 608100.0 102300.0 609000.0 ;
      RECT  101850.0 603150.0 102750.0 608550.0 ;
      RECT  96900.0 610650.0 98100.0 611850.0 ;
      RECT  101700.0 610650.0 102900.0 611850.0 ;
      RECT  101700.0 601950.0 102900.0 603150.0 ;
      RECT  101700.0 607950.0 102900.0 609150.0 ;
      RECT  101850.0 624450.0 102750.0 616950.0 ;
      RECT  97050.0 619500.0 97950.0 618600.0 ;
      RECT  101850.0 619500.0 102750.0 618600.0 ;
      RECT  97050.0 619050.0 97950.0 616950.0 ;
      RECT  97500.0 619500.0 102300.0 618600.0 ;
      RECT  101850.0 624450.0 102750.0 619050.0 ;
      RECT  96900.0 616950.0 98100.0 615750.0 ;
      RECT  101700.0 616950.0 102900.0 615750.0 ;
      RECT  101700.0 625650.0 102900.0 624450.0 ;
      RECT  101700.0 619650.0 102900.0 618450.0 ;
      RECT  101850.0 630750.0 102750.0 638250.0 ;
      RECT  97050.0 635700.0 97950.0 636600.0 ;
      RECT  101850.0 635700.0 102750.0 636600.0 ;
      RECT  97050.0 636150.0 97950.0 638250.0 ;
      RECT  97500.0 635700.0 102300.0 636600.0 ;
      RECT  101850.0 630750.0 102750.0 636150.0 ;
      RECT  96900.0 638250.0 98100.0 639450.0 ;
      RECT  101700.0 638250.0 102900.0 639450.0 ;
      RECT  101700.0 629550.0 102900.0 630750.0 ;
      RECT  101700.0 635550.0 102900.0 636750.0 ;
      RECT  101850.0 652050.0 102750.0 644550.0 ;
      RECT  97050.0 647100.0 97950.0 646200.0 ;
      RECT  101850.0 647100.0 102750.0 646200.0 ;
      RECT  97050.0 646650.0 97950.0 644550.0 ;
      RECT  97500.0 647100.0 102300.0 646200.0 ;
      RECT  101850.0 652050.0 102750.0 646650.0 ;
      RECT  96900.0 644550.0 98100.0 643350.0 ;
      RECT  101700.0 644550.0 102900.0 643350.0 ;
      RECT  101700.0 653250.0 102900.0 652050.0 ;
      RECT  101700.0 647250.0 102900.0 646050.0 ;
      RECT  101850.0 658350.0 102750.0 665850.0 ;
      RECT  97050.0 663300.0 97950.0 664200.0 ;
      RECT  101850.0 663300.0 102750.0 664200.0 ;
      RECT  97050.0 663750.0 97950.0 665850.0 ;
      RECT  97500.0 663300.0 102300.0 664200.0 ;
      RECT  101850.0 658350.0 102750.0 663750.0 ;
      RECT  96900.0 665850.0 98100.0 667050.0 ;
      RECT  101700.0 665850.0 102900.0 667050.0 ;
      RECT  101700.0 657150.0 102900.0 658350.0 ;
      RECT  101700.0 663150.0 102900.0 664350.0 ;
      RECT  101850.0 679650.0 102750.0 672150.0 ;
      RECT  97050.0 674700.0 97950.0 673800.0 ;
      RECT  101850.0 674700.0 102750.0 673800.0 ;
      RECT  97050.0 674250.0 97950.0 672150.0 ;
      RECT  97500.0 674700.0 102300.0 673800.0 ;
      RECT  101850.0 679650.0 102750.0 674250.0 ;
      RECT  96900.0 672150.0 98100.0 670950.0 ;
      RECT  101700.0 672150.0 102900.0 670950.0 ;
      RECT  101700.0 680850.0 102900.0 679650.0 ;
      RECT  101700.0 674850.0 102900.0 673650.0 ;
      RECT  101850.0 685950.0 102750.0 693450.0 ;
      RECT  97050.0 690900.0 97950.0 691800.0 ;
      RECT  101850.0 690900.0 102750.0 691800.0 ;
      RECT  97050.0 691350.0 97950.0 693450.0 ;
      RECT  97500.0 690900.0 102300.0 691800.0 ;
      RECT  101850.0 685950.0 102750.0 691350.0 ;
      RECT  96900.0 693450.0 98100.0 694650.0 ;
      RECT  101700.0 693450.0 102900.0 694650.0 ;
      RECT  101700.0 684750.0 102900.0 685950.0 ;
      RECT  101700.0 690750.0 102900.0 691950.0 ;
      RECT  101850.0 707250.0 102750.0 699750.0 ;
      RECT  97050.0 702300.0 97950.0 701400.0 ;
      RECT  101850.0 702300.0 102750.0 701400.0 ;
      RECT  97050.0 701850.0 97950.0 699750.0 ;
      RECT  97500.0 702300.0 102300.0 701400.0 ;
      RECT  101850.0 707250.0 102750.0 701850.0 ;
      RECT  96900.0 699750.0 98100.0 698550.0 ;
      RECT  101700.0 699750.0 102900.0 698550.0 ;
      RECT  101700.0 708450.0 102900.0 707250.0 ;
      RECT  101700.0 702450.0 102900.0 701250.0 ;
      RECT  101850.0 713550.0 102750.0 721050.0 ;
      RECT  97050.0 718500.0 97950.0 719400.0 ;
      RECT  101850.0 718500.0 102750.0 719400.0 ;
      RECT  97050.0 718950.0 97950.0 721050.0 ;
      RECT  97500.0 718500.0 102300.0 719400.0 ;
      RECT  101850.0 713550.0 102750.0 718950.0 ;
      RECT  96900.0 721050.0 98100.0 722250.0 ;
      RECT  101700.0 721050.0 102900.0 722250.0 ;
      RECT  101700.0 712350.0 102900.0 713550.0 ;
      RECT  101700.0 718350.0 102900.0 719550.0 ;
      RECT  101850.0 734850.0 102750.0 727350.0 ;
      RECT  97050.0 729900.0 97950.0 729000.0 ;
      RECT  101850.0 729900.0 102750.0 729000.0 ;
      RECT  97050.0 729450.0 97950.0 727350.0 ;
      RECT  97500.0 729900.0 102300.0 729000.0 ;
      RECT  101850.0 734850.0 102750.0 729450.0 ;
      RECT  96900.0 727350.0 98100.0 726150.0 ;
      RECT  101700.0 727350.0 102900.0 726150.0 ;
      RECT  101700.0 736050.0 102900.0 734850.0 ;
      RECT  101700.0 730050.0 102900.0 728850.0 ;
      RECT  101850.0 741150.0 102750.0 748650.0 ;
      RECT  97050.0 746100.0 97950.0 747000.0 ;
      RECT  101850.0 746100.0 102750.0 747000.0 ;
      RECT  97050.0 746550.0 97950.0 748650.0 ;
      RECT  97500.0 746100.0 102300.0 747000.0 ;
      RECT  101850.0 741150.0 102750.0 746550.0 ;
      RECT  96900.0 748650.0 98100.0 749850.0 ;
      RECT  101700.0 748650.0 102900.0 749850.0 ;
      RECT  101700.0 739950.0 102900.0 741150.0 ;
      RECT  101700.0 745950.0 102900.0 747150.0 ;
      RECT  101850.0 762450.0 102750.0 754950.0 ;
      RECT  97050.0 757500.0 97950.0 756600.0 ;
      RECT  101850.0 757500.0 102750.0 756600.0 ;
      RECT  97050.0 757050.0 97950.0 754950.0 ;
      RECT  97500.0 757500.0 102300.0 756600.0 ;
      RECT  101850.0 762450.0 102750.0 757050.0 ;
      RECT  96900.0 754950.0 98100.0 753750.0 ;
      RECT  101700.0 754950.0 102900.0 753750.0 ;
      RECT  101700.0 763650.0 102900.0 762450.0 ;
      RECT  101700.0 757650.0 102900.0 756450.0 ;
      RECT  101850.0 768750.0 102750.0 776250.0 ;
      RECT  97050.0 773700.0 97950.0 774600.0 ;
      RECT  101850.0 773700.0 102750.0 774600.0 ;
      RECT  97050.0 774150.0 97950.0 776250.0 ;
      RECT  97500.0 773700.0 102300.0 774600.0 ;
      RECT  101850.0 768750.0 102750.0 774150.0 ;
      RECT  96900.0 776250.0 98100.0 777450.0 ;
      RECT  101700.0 776250.0 102900.0 777450.0 ;
      RECT  101700.0 767550.0 102900.0 768750.0 ;
      RECT  101700.0 773550.0 102900.0 774750.0 ;
      RECT  101850.0 790050.0 102750.0 782550.0 ;
      RECT  97050.0 785100.0 97950.0 784200.0 ;
      RECT  101850.0 785100.0 102750.0 784200.0 ;
      RECT  97050.0 784650.0 97950.0 782550.0 ;
      RECT  97500.0 785100.0 102300.0 784200.0 ;
      RECT  101850.0 790050.0 102750.0 784650.0 ;
      RECT  96900.0 782550.0 98100.0 781350.0 ;
      RECT  101700.0 782550.0 102900.0 781350.0 ;
      RECT  101700.0 791250.0 102900.0 790050.0 ;
      RECT  101700.0 785250.0 102900.0 784050.0 ;
      RECT  101850.0 796350.0 102750.0 803850.0 ;
      RECT  97050.0 801300.0 97950.0 802200.0 ;
      RECT  101850.0 801300.0 102750.0 802200.0 ;
      RECT  97050.0 801750.0 97950.0 803850.0 ;
      RECT  97500.0 801300.0 102300.0 802200.0 ;
      RECT  101850.0 796350.0 102750.0 801750.0 ;
      RECT  96900.0 803850.0 98100.0 805050.0 ;
      RECT  101700.0 803850.0 102900.0 805050.0 ;
      RECT  101700.0 795150.0 102900.0 796350.0 ;
      RECT  101700.0 801150.0 102900.0 802350.0 ;
      RECT  101850.0 817650.0 102750.0 810150.0 ;
      RECT  97050.0 812700.0 97950.0 811800.0 ;
      RECT  101850.0 812700.0 102750.0 811800.0 ;
      RECT  97050.0 812250.0 97950.0 810150.0 ;
      RECT  97500.0 812700.0 102300.0 811800.0 ;
      RECT  101850.0 817650.0 102750.0 812250.0 ;
      RECT  96900.0 810150.0 98100.0 808950.0 ;
      RECT  101700.0 810150.0 102900.0 808950.0 ;
      RECT  101700.0 818850.0 102900.0 817650.0 ;
      RECT  101700.0 812850.0 102900.0 811650.0 ;
      RECT  101850.0 823950.0 102750.0 831450.0 ;
      RECT  97050.0 828900.0 97950.0 829800.0 ;
      RECT  101850.0 828900.0 102750.0 829800.0 ;
      RECT  97050.0 829350.0 97950.0 831450.0 ;
      RECT  97500.0 828900.0 102300.0 829800.0 ;
      RECT  101850.0 823950.0 102750.0 829350.0 ;
      RECT  96900.0 831450.0 98100.0 832650.0 ;
      RECT  101700.0 831450.0 102900.0 832650.0 ;
      RECT  101700.0 822750.0 102900.0 823950.0 ;
      RECT  101700.0 828750.0 102900.0 829950.0 ;
      RECT  101850.0 845250.0 102750.0 837750.0 ;
      RECT  97050.0 840300.0 97950.0 839400.0 ;
      RECT  101850.0 840300.0 102750.0 839400.0 ;
      RECT  97050.0 839850.0 97950.0 837750.0 ;
      RECT  97500.0 840300.0 102300.0 839400.0 ;
      RECT  101850.0 845250.0 102750.0 839850.0 ;
      RECT  96900.0 837750.0 98100.0 836550.0 ;
      RECT  101700.0 837750.0 102900.0 836550.0 ;
      RECT  101700.0 846450.0 102900.0 845250.0 ;
      RECT  101700.0 840450.0 102900.0 839250.0 ;
      RECT  101850.0 851550.0 102750.0 859050.0 ;
      RECT  97050.0 856500.0 97950.0 857400.0 ;
      RECT  101850.0 856500.0 102750.0 857400.0 ;
      RECT  97050.0 856950.0 97950.0 859050.0 ;
      RECT  97500.0 856500.0 102300.0 857400.0 ;
      RECT  101850.0 851550.0 102750.0 856950.0 ;
      RECT  96900.0 859050.0 98100.0 860250.0 ;
      RECT  101700.0 859050.0 102900.0 860250.0 ;
      RECT  101700.0 850350.0 102900.0 851550.0 ;
      RECT  101700.0 856350.0 102900.0 857550.0 ;
      RECT  101850.0 872850.0 102750.0 865350.0 ;
      RECT  97050.0 867900.0 97950.0 867000.0 ;
      RECT  101850.0 867900.0 102750.0 867000.0 ;
      RECT  97050.0 867450.0 97950.0 865350.0 ;
      RECT  97500.0 867900.0 102300.0 867000.0 ;
      RECT  101850.0 872850.0 102750.0 867450.0 ;
      RECT  96900.0 865350.0 98100.0 864150.0 ;
      RECT  101700.0 865350.0 102900.0 864150.0 ;
      RECT  101700.0 874050.0 102900.0 872850.0 ;
      RECT  101700.0 868050.0 102900.0 866850.0 ;
      RECT  101850.0 879150.0 102750.0 886650.0 ;
      RECT  97050.0 884100.0 97950.0 885000.0 ;
      RECT  101850.0 884100.0 102750.0 885000.0 ;
      RECT  97050.0 884550.0 97950.0 886650.0 ;
      RECT  97500.0 884100.0 102300.0 885000.0 ;
      RECT  101850.0 879150.0 102750.0 884550.0 ;
      RECT  96900.0 886650.0 98100.0 887850.0 ;
      RECT  101700.0 886650.0 102900.0 887850.0 ;
      RECT  101700.0 877950.0 102900.0 879150.0 ;
      RECT  101700.0 883950.0 102900.0 885150.0 ;
      RECT  101850.0 900450.0 102750.0 892950.0 ;
      RECT  97050.0 895500.0 97950.0 894600.0 ;
      RECT  101850.0 895500.0 102750.0 894600.0 ;
      RECT  97050.0 895050.0 97950.0 892950.0 ;
      RECT  97500.0 895500.0 102300.0 894600.0 ;
      RECT  101850.0 900450.0 102750.0 895050.0 ;
      RECT  96900.0 892950.0 98100.0 891750.0 ;
      RECT  101700.0 892950.0 102900.0 891750.0 ;
      RECT  101700.0 901650.0 102900.0 900450.0 ;
      RECT  101700.0 895650.0 102900.0 894450.0 ;
      RECT  101850.0 906750.0 102750.0 914250.0 ;
      RECT  97050.0 911700.0 97950.0 912600.0 ;
      RECT  101850.0 911700.0 102750.0 912600.0 ;
      RECT  97050.0 912150.0 97950.0 914250.0 ;
      RECT  97500.0 911700.0 102300.0 912600.0 ;
      RECT  101850.0 906750.0 102750.0 912150.0 ;
      RECT  96900.0 914250.0 98100.0 915450.0 ;
      RECT  101700.0 914250.0 102900.0 915450.0 ;
      RECT  101700.0 905550.0 102900.0 906750.0 ;
      RECT  101700.0 911550.0 102900.0 912750.0 ;
      RECT  101850.0 928050.0 102750.0 920550.0 ;
      RECT  97050.0 923100.0 97950.0 922200.0 ;
      RECT  101850.0 923100.0 102750.0 922200.0 ;
      RECT  97050.0 922650.0 97950.0 920550.0 ;
      RECT  97500.0 923100.0 102300.0 922200.0 ;
      RECT  101850.0 928050.0 102750.0 922650.0 ;
      RECT  96900.0 920550.0 98100.0 919350.0 ;
      RECT  101700.0 920550.0 102900.0 919350.0 ;
      RECT  101700.0 929250.0 102900.0 928050.0 ;
      RECT  101700.0 923250.0 102900.0 922050.0 ;
      RECT  101850.0 934350.0 102750.0 941850.0 ;
      RECT  97050.0 939300.0 97950.0 940200.0 ;
      RECT  101850.0 939300.0 102750.0 940200.0 ;
      RECT  97050.0 939750.0 97950.0 941850.0 ;
      RECT  97500.0 939300.0 102300.0 940200.0 ;
      RECT  101850.0 934350.0 102750.0 939750.0 ;
      RECT  96900.0 941850.0 98100.0 943050.0 ;
      RECT  101700.0 941850.0 102900.0 943050.0 ;
      RECT  101700.0 933150.0 102900.0 934350.0 ;
      RECT  101700.0 939150.0 102900.0 940350.0 ;
      RECT  101850.0 955650.0 102750.0 948150.0 ;
      RECT  97050.0 950700.0 97950.0 949800.0 ;
      RECT  101850.0 950700.0 102750.0 949800.0 ;
      RECT  97050.0 950250.0 97950.0 948150.0 ;
      RECT  97500.0 950700.0 102300.0 949800.0 ;
      RECT  101850.0 955650.0 102750.0 950250.0 ;
      RECT  96900.0 948150.0 98100.0 946950.0 ;
      RECT  101700.0 948150.0 102900.0 946950.0 ;
      RECT  101700.0 956850.0 102900.0 955650.0 ;
      RECT  101700.0 950850.0 102900.0 949650.0 ;
      RECT  101850.0 961950.0 102750.0 969450.0 ;
      RECT  97050.0 966900.0 97950.0 967800.0 ;
      RECT  101850.0 966900.0 102750.0 967800.0 ;
      RECT  97050.0 967350.0 97950.0 969450.0 ;
      RECT  97500.0 966900.0 102300.0 967800.0 ;
      RECT  101850.0 961950.0 102750.0 967350.0 ;
      RECT  96900.0 969450.0 98100.0 970650.0 ;
      RECT  101700.0 969450.0 102900.0 970650.0 ;
      RECT  101700.0 960750.0 102900.0 961950.0 ;
      RECT  101700.0 966750.0 102900.0 967950.0 ;
      RECT  101850.0 983250.0 102750.0 975750.0 ;
      RECT  97050.0 978300.0 97950.0 977400.0 ;
      RECT  101850.0 978300.0 102750.0 977400.0 ;
      RECT  97050.0 977850.0 97950.0 975750.0 ;
      RECT  97500.0 978300.0 102300.0 977400.0 ;
      RECT  101850.0 983250.0 102750.0 977850.0 ;
      RECT  96900.0 975750.0 98100.0 974550.0 ;
      RECT  101700.0 975750.0 102900.0 974550.0 ;
      RECT  101700.0 984450.0 102900.0 983250.0 ;
      RECT  101700.0 978450.0 102900.0 977250.0 ;
      RECT  101850.0 989550.0 102750.0 997050.0 ;
      RECT  97050.0 994500.0 97950.0 995400.0 ;
      RECT  101850.0 994500.0 102750.0 995400.0 ;
      RECT  97050.0 994950.0 97950.0 997050.0 ;
      RECT  97500.0 994500.0 102300.0 995400.0 ;
      RECT  101850.0 989550.0 102750.0 994950.0 ;
      RECT  96900.0 997050.0 98100.0 998250.0 ;
      RECT  101700.0 997050.0 102900.0 998250.0 ;
      RECT  101700.0 988350.0 102900.0 989550.0 ;
      RECT  101700.0 994350.0 102900.0 995550.0 ;
      RECT  101850.0 1010850.0 102750.0 1003350.0 ;
      RECT  97050.0 1005900.0 97950.0 1005000.0 ;
      RECT  101850.0 1005900.0 102750.0 1005000.0 ;
      RECT  97050.0 1005450.0 97950.0 1003350.0 ;
      RECT  97500.0 1005900.0 102300.0 1005000.0 ;
      RECT  101850.0 1010850.0 102750.0 1005450.0 ;
      RECT  96900.0 1003350.0 98100.0 1002150.0 ;
      RECT  101700.0 1003350.0 102900.0 1002150.0 ;
      RECT  101700.0 1012050.0 102900.0 1010850.0 ;
      RECT  101700.0 1006050.0 102900.0 1004850.0 ;
      RECT  101850.0 1017150.0 102750.0 1024650.0 ;
      RECT  97050.0 1022100.0 97950.0 1023000.0 ;
      RECT  101850.0 1022100.0 102750.0 1023000.0 ;
      RECT  97050.0 1022550.0 97950.0 1024650.0 ;
      RECT  97500.0 1022100.0 102300.0 1023000.0 ;
      RECT  101850.0 1017150.0 102750.0 1022550.0 ;
      RECT  96900.0 1024650.0 98100.0 1025850.0 ;
      RECT  101700.0 1024650.0 102900.0 1025850.0 ;
      RECT  101700.0 1015950.0 102900.0 1017150.0 ;
      RECT  101700.0 1021950.0 102900.0 1023150.0 ;
      RECT  101850.0 1038450.0 102750.0 1030950.0 ;
      RECT  97050.0 1033500.0 97950.0 1032600.0 ;
      RECT  101850.0 1033500.0 102750.0 1032600.0 ;
      RECT  97050.0 1033050.0 97950.0 1030950.0 ;
      RECT  97500.0 1033500.0 102300.0 1032600.0 ;
      RECT  101850.0 1038450.0 102750.0 1033050.0 ;
      RECT  96900.0 1030950.0 98100.0 1029750.0 ;
      RECT  101700.0 1030950.0 102900.0 1029750.0 ;
      RECT  101700.0 1039650.0 102900.0 1038450.0 ;
      RECT  101700.0 1033650.0 102900.0 1032450.0 ;
      RECT  101850.0 1044750.0 102750.0 1052250.0 ;
      RECT  97050.0 1049700.0 97950.0 1050600.0 ;
      RECT  101850.0 1049700.0 102750.0 1050600.0 ;
      RECT  97050.0 1050150.0 97950.0 1052250.0 ;
      RECT  97500.0 1049700.0 102300.0 1050600.0 ;
      RECT  101850.0 1044750.0 102750.0 1050150.0 ;
      RECT  96900.0 1052250.0 98100.0 1053450.0 ;
      RECT  101700.0 1052250.0 102900.0 1053450.0 ;
      RECT  101700.0 1043550.0 102900.0 1044750.0 ;
      RECT  101700.0 1049550.0 102900.0 1050750.0 ;
      RECT  101850.0 1066050.0 102750.0 1058550.0 ;
      RECT  97050.0 1061100.0 97950.0 1060200.0 ;
      RECT  101850.0 1061100.0 102750.0 1060200.0 ;
      RECT  97050.0 1060650.0 97950.0 1058550.0 ;
      RECT  97500.0 1061100.0 102300.0 1060200.0 ;
      RECT  101850.0 1066050.0 102750.0 1060650.0 ;
      RECT  96900.0 1058550.0 98100.0 1057350.0 ;
      RECT  101700.0 1058550.0 102900.0 1057350.0 ;
      RECT  101700.0 1067250.0 102900.0 1066050.0 ;
      RECT  101700.0 1061250.0 102900.0 1060050.0 ;
      RECT  101850.0 1072350.0 102750.0 1079850.0 ;
      RECT  97050.0 1077300.0 97950.0 1078200.0 ;
      RECT  101850.0 1077300.0 102750.0 1078200.0 ;
      RECT  97050.0 1077750.0 97950.0 1079850.0 ;
      RECT  97500.0 1077300.0 102300.0 1078200.0 ;
      RECT  101850.0 1072350.0 102750.0 1077750.0 ;
      RECT  96900.0 1079850.0 98100.0 1081050.0 ;
      RECT  101700.0 1079850.0 102900.0 1081050.0 ;
      RECT  101700.0 1071150.0 102900.0 1072350.0 ;
      RECT  101700.0 1077150.0 102900.0 1078350.0 ;
      RECT  101850.0 1093650.0 102750.0 1086150.0 ;
      RECT  97050.0 1088700.0 97950.0 1087800.0 ;
      RECT  101850.0 1088700.0 102750.0 1087800.0 ;
      RECT  97050.0 1088250.0 97950.0 1086150.0 ;
      RECT  97500.0 1088700.0 102300.0 1087800.0 ;
      RECT  101850.0 1093650.0 102750.0 1088250.0 ;
      RECT  96900.0 1086150.0 98100.0 1084950.0 ;
      RECT  101700.0 1086150.0 102900.0 1084950.0 ;
      RECT  101700.0 1094850.0 102900.0 1093650.0 ;
      RECT  101700.0 1088850.0 102900.0 1087650.0 ;
      RECT  101850.0 1099950.0 102750.0 1107450.0 ;
      RECT  97050.0 1104900.0 97950.0 1105800.0 ;
      RECT  101850.0 1104900.0 102750.0 1105800.0 ;
      RECT  97050.0 1105350.0 97950.0 1107450.0 ;
      RECT  97500.0 1104900.0 102300.0 1105800.0 ;
      RECT  101850.0 1099950.0 102750.0 1105350.0 ;
      RECT  96900.0 1107450.0 98100.0 1108650.0 ;
      RECT  101700.0 1107450.0 102900.0 1108650.0 ;
      RECT  101700.0 1098750.0 102900.0 1099950.0 ;
      RECT  101700.0 1104750.0 102900.0 1105950.0 ;
      RECT  101850.0 1121250.0 102750.0 1113750.0 ;
      RECT  97050.0 1116300.0 97950.0 1115400.0 ;
      RECT  101850.0 1116300.0 102750.0 1115400.0 ;
      RECT  97050.0 1115850.0 97950.0 1113750.0 ;
      RECT  97500.0 1116300.0 102300.0 1115400.0 ;
      RECT  101850.0 1121250.0 102750.0 1115850.0 ;
      RECT  96900.0 1113750.0 98100.0 1112550.0 ;
      RECT  101700.0 1113750.0 102900.0 1112550.0 ;
      RECT  101700.0 1122450.0 102900.0 1121250.0 ;
      RECT  101700.0 1116450.0 102900.0 1115250.0 ;
      RECT  101850.0 1127550.0 102750.0 1135050.0 ;
      RECT  97050.0 1132500.0 97950.0 1133400.0 ;
      RECT  101850.0 1132500.0 102750.0 1133400.0 ;
      RECT  97050.0 1132950.0 97950.0 1135050.0 ;
      RECT  97500.0 1132500.0 102300.0 1133400.0 ;
      RECT  101850.0 1127550.0 102750.0 1132950.0 ;
      RECT  96900.0 1135050.0 98100.0 1136250.0 ;
      RECT  101700.0 1135050.0 102900.0 1136250.0 ;
      RECT  101700.0 1126350.0 102900.0 1127550.0 ;
      RECT  101700.0 1132350.0 102900.0 1133550.0 ;
      RECT  101850.0 1148850.0 102750.0 1141350.0 ;
      RECT  97050.0 1143900.0 97950.0 1143000.0 ;
      RECT  101850.0 1143900.0 102750.0 1143000.0 ;
      RECT  97050.0 1143450.0 97950.0 1141350.0 ;
      RECT  97500.0 1143900.0 102300.0 1143000.0 ;
      RECT  101850.0 1148850.0 102750.0 1143450.0 ;
      RECT  96900.0 1141350.0 98100.0 1140150.0 ;
      RECT  101700.0 1141350.0 102900.0 1140150.0 ;
      RECT  101700.0 1150050.0 102900.0 1148850.0 ;
      RECT  101700.0 1144050.0 102900.0 1142850.0 ;
      RECT  101850.0 1155150.0 102750.0 1162650.0 ;
      RECT  97050.0 1160100.0 97950.0 1161000.0 ;
      RECT  101850.0 1160100.0 102750.0 1161000.0 ;
      RECT  97050.0 1160550.0 97950.0 1162650.0 ;
      RECT  97500.0 1160100.0 102300.0 1161000.0 ;
      RECT  101850.0 1155150.0 102750.0 1160550.0 ;
      RECT  96900.0 1162650.0 98100.0 1163850.0 ;
      RECT  101700.0 1162650.0 102900.0 1163850.0 ;
      RECT  101700.0 1153950.0 102900.0 1155150.0 ;
      RECT  101700.0 1159950.0 102900.0 1161150.0 ;
      RECT  101850.0 1176450.0 102750.0 1168950.0 ;
      RECT  97050.0 1171500.0 97950.0 1170600.0 ;
      RECT  101850.0 1171500.0 102750.0 1170600.0 ;
      RECT  97050.0 1171050.0 97950.0 1168950.0 ;
      RECT  97500.0 1171500.0 102300.0 1170600.0 ;
      RECT  101850.0 1176450.0 102750.0 1171050.0 ;
      RECT  96900.0 1168950.0 98100.0 1167750.0 ;
      RECT  101700.0 1168950.0 102900.0 1167750.0 ;
      RECT  101700.0 1177650.0 102900.0 1176450.0 ;
      RECT  101700.0 1171650.0 102900.0 1170450.0 ;
      RECT  101850.0 1182750.0 102750.0 1190250.0 ;
      RECT  97050.0 1187700.0 97950.0 1188600.0 ;
      RECT  101850.0 1187700.0 102750.0 1188600.0 ;
      RECT  97050.0 1188150.0 97950.0 1190250.0 ;
      RECT  97500.0 1187700.0 102300.0 1188600.0 ;
      RECT  101850.0 1182750.0 102750.0 1188150.0 ;
      RECT  96900.0 1190250.0 98100.0 1191450.0 ;
      RECT  101700.0 1190250.0 102900.0 1191450.0 ;
      RECT  101700.0 1181550.0 102900.0 1182750.0 ;
      RECT  101700.0 1187550.0 102900.0 1188750.0 ;
      RECT  101850.0 1204050.0 102750.0 1196550.0 ;
      RECT  97050.0 1199100.0 97950.0 1198200.0 ;
      RECT  101850.0 1199100.0 102750.0 1198200.0 ;
      RECT  97050.0 1198650.0 97950.0 1196550.0 ;
      RECT  97500.0 1199100.0 102300.0 1198200.0 ;
      RECT  101850.0 1204050.0 102750.0 1198650.0 ;
      RECT  96900.0 1196550.0 98100.0 1195350.0 ;
      RECT  101700.0 1196550.0 102900.0 1195350.0 ;
      RECT  101700.0 1205250.0 102900.0 1204050.0 ;
      RECT  101700.0 1199250.0 102900.0 1198050.0 ;
      RECT  101850.0 1210350.0 102750.0 1217850.0 ;
      RECT  97050.0 1215300.0 97950.0 1216200.0 ;
      RECT  101850.0 1215300.0 102750.0 1216200.0 ;
      RECT  97050.0 1215750.0 97950.0 1217850.0 ;
      RECT  97500.0 1215300.0 102300.0 1216200.0 ;
      RECT  101850.0 1210350.0 102750.0 1215750.0 ;
      RECT  96900.0 1217850.0 98100.0 1219050.0 ;
      RECT  101700.0 1217850.0 102900.0 1219050.0 ;
      RECT  101700.0 1209150.0 102900.0 1210350.0 ;
      RECT  101700.0 1215150.0 102900.0 1216350.0 ;
      RECT  101850.0 1231650.0 102750.0 1224150.0 ;
      RECT  97050.0 1226700.0 97950.0 1225800.0 ;
      RECT  101850.0 1226700.0 102750.0 1225800.0 ;
      RECT  97050.0 1226250.0 97950.0 1224150.0 ;
      RECT  97500.0 1226700.0 102300.0 1225800.0 ;
      RECT  101850.0 1231650.0 102750.0 1226250.0 ;
      RECT  96900.0 1224150.0 98100.0 1222950.0 ;
      RECT  101700.0 1224150.0 102900.0 1222950.0 ;
      RECT  101700.0 1232850.0 102900.0 1231650.0 ;
      RECT  101700.0 1226850.0 102900.0 1225650.0 ;
      RECT  101850.0 1237950.0 102750.0 1245450.0 ;
      RECT  97050.0 1242900.0 97950.0 1243800.0 ;
      RECT  101850.0 1242900.0 102750.0 1243800.0 ;
      RECT  97050.0 1243350.0 97950.0 1245450.0 ;
      RECT  97500.0 1242900.0 102300.0 1243800.0 ;
      RECT  101850.0 1237950.0 102750.0 1243350.0 ;
      RECT  96900.0 1245450.0 98100.0 1246650.0 ;
      RECT  101700.0 1245450.0 102900.0 1246650.0 ;
      RECT  101700.0 1236750.0 102900.0 1237950.0 ;
      RECT  101700.0 1242750.0 102900.0 1243950.0 ;
      RECT  101850.0 1259250.0 102750.0 1251750.0 ;
      RECT  97050.0 1254300.0 97950.0 1253400.0 ;
      RECT  101850.0 1254300.0 102750.0 1253400.0 ;
      RECT  97050.0 1253850.0 97950.0 1251750.0 ;
      RECT  97500.0 1254300.0 102300.0 1253400.0 ;
      RECT  101850.0 1259250.0 102750.0 1253850.0 ;
      RECT  96900.0 1251750.0 98100.0 1250550.0 ;
      RECT  101700.0 1251750.0 102900.0 1250550.0 ;
      RECT  101700.0 1260450.0 102900.0 1259250.0 ;
      RECT  101700.0 1254450.0 102900.0 1253250.0 ;
      RECT  101850.0 1265550.0 102750.0 1273050.0 ;
      RECT  97050.0 1270500.0 97950.0 1271400.0 ;
      RECT  101850.0 1270500.0 102750.0 1271400.0 ;
      RECT  97050.0 1270950.0 97950.0 1273050.0 ;
      RECT  97500.0 1270500.0 102300.0 1271400.0 ;
      RECT  101850.0 1265550.0 102750.0 1270950.0 ;
      RECT  96900.0 1273050.0 98100.0 1274250.0 ;
      RECT  101700.0 1273050.0 102900.0 1274250.0 ;
      RECT  101700.0 1264350.0 102900.0 1265550.0 ;
      RECT  101700.0 1270350.0 102900.0 1271550.0 ;
      RECT  101850.0 1286850.0 102750.0 1279350.0 ;
      RECT  97050.0 1281900.0 97950.0 1281000.0 ;
      RECT  101850.0 1281900.0 102750.0 1281000.0 ;
      RECT  97050.0 1281450.0 97950.0 1279350.0 ;
      RECT  97500.0 1281900.0 102300.0 1281000.0 ;
      RECT  101850.0 1286850.0 102750.0 1281450.0 ;
      RECT  96900.0 1279350.0 98100.0 1278150.0 ;
      RECT  101700.0 1279350.0 102900.0 1278150.0 ;
      RECT  101700.0 1288050.0 102900.0 1286850.0 ;
      RECT  101700.0 1282050.0 102900.0 1280850.0 ;
      RECT  101850.0 1293150.0 102750.0 1300650.0 ;
      RECT  97050.0 1298100.0 97950.0 1299000.0 ;
      RECT  101850.0 1298100.0 102750.0 1299000.0 ;
      RECT  97050.0 1298550.0 97950.0 1300650.0 ;
      RECT  97500.0 1298100.0 102300.0 1299000.0 ;
      RECT  101850.0 1293150.0 102750.0 1298550.0 ;
      RECT  96900.0 1300650.0 98100.0 1301850.0 ;
      RECT  101700.0 1300650.0 102900.0 1301850.0 ;
      RECT  101700.0 1291950.0 102900.0 1293150.0 ;
      RECT  101700.0 1297950.0 102900.0 1299150.0 ;
      RECT  101850.0 1314450.0 102750.0 1306950.0 ;
      RECT  97050.0 1309500.0 97950.0 1308600.0 ;
      RECT  101850.0 1309500.0 102750.0 1308600.0 ;
      RECT  97050.0 1309050.0 97950.0 1306950.0 ;
      RECT  97500.0 1309500.0 102300.0 1308600.0 ;
      RECT  101850.0 1314450.0 102750.0 1309050.0 ;
      RECT  96900.0 1306950.0 98100.0 1305750.0 ;
      RECT  101700.0 1306950.0 102900.0 1305750.0 ;
      RECT  101700.0 1315650.0 102900.0 1314450.0 ;
      RECT  101700.0 1309650.0 102900.0 1308450.0 ;
      RECT  101850.0 1320750.0 102750.0 1328250.0 ;
      RECT  97050.0 1325700.0 97950.0 1326600.0 ;
      RECT  101850.0 1325700.0 102750.0 1326600.0 ;
      RECT  97050.0 1326150.0 97950.0 1328250.0 ;
      RECT  97500.0 1325700.0 102300.0 1326600.0 ;
      RECT  101850.0 1320750.0 102750.0 1326150.0 ;
      RECT  96900.0 1328250.0 98100.0 1329450.0 ;
      RECT  101700.0 1328250.0 102900.0 1329450.0 ;
      RECT  101700.0 1319550.0 102900.0 1320750.0 ;
      RECT  101700.0 1325550.0 102900.0 1326750.0 ;
      RECT  101850.0 1342050.0 102750.0 1334550.0 ;
      RECT  97050.0 1337100.0 97950.0 1336200.0 ;
      RECT  101850.0 1337100.0 102750.0 1336200.0 ;
      RECT  97050.0 1336650.0 97950.0 1334550.0 ;
      RECT  97500.0 1337100.0 102300.0 1336200.0 ;
      RECT  101850.0 1342050.0 102750.0 1336650.0 ;
      RECT  96900.0 1334550.0 98100.0 1333350.0 ;
      RECT  101700.0 1334550.0 102900.0 1333350.0 ;
      RECT  101700.0 1343250.0 102900.0 1342050.0 ;
      RECT  101700.0 1337250.0 102900.0 1336050.0 ;
      RECT  101850.0 1348350.0 102750.0 1355850.0 ;
      RECT  97050.0 1353300.0 97950.0 1354200.0 ;
      RECT  101850.0 1353300.0 102750.0 1354200.0 ;
      RECT  97050.0 1353750.0 97950.0 1355850.0 ;
      RECT  97500.0 1353300.0 102300.0 1354200.0 ;
      RECT  101850.0 1348350.0 102750.0 1353750.0 ;
      RECT  96900.0 1355850.0 98100.0 1357050.0 ;
      RECT  101700.0 1355850.0 102900.0 1357050.0 ;
      RECT  101700.0 1347150.0 102900.0 1348350.0 ;
      RECT  101700.0 1353150.0 102900.0 1354350.0 ;
      RECT  101850.0 1369650.0 102750.0 1362150.0 ;
      RECT  97050.0 1364700.0 97950.0 1363800.0 ;
      RECT  101850.0 1364700.0 102750.0 1363800.0 ;
      RECT  97050.0 1364250.0 97950.0 1362150.0 ;
      RECT  97500.0 1364700.0 102300.0 1363800.0 ;
      RECT  101850.0 1369650.0 102750.0 1364250.0 ;
      RECT  96900.0 1362150.0 98100.0 1360950.0 ;
      RECT  101700.0 1362150.0 102900.0 1360950.0 ;
      RECT  101700.0 1370850.0 102900.0 1369650.0 ;
      RECT  101700.0 1364850.0 102900.0 1363650.0 ;
      RECT  101850.0 1375950.0 102750.0 1383450.0 ;
      RECT  97050.0 1380900.0 97950.0 1381800.0 ;
      RECT  101850.0 1380900.0 102750.0 1381800.0 ;
      RECT  97050.0 1381350.0 97950.0 1383450.0 ;
      RECT  97500.0 1380900.0 102300.0 1381800.0 ;
      RECT  101850.0 1375950.0 102750.0 1381350.0 ;
      RECT  96900.0 1383450.0 98100.0 1384650.0 ;
      RECT  101700.0 1383450.0 102900.0 1384650.0 ;
      RECT  101700.0 1374750.0 102900.0 1375950.0 ;
      RECT  101700.0 1380750.0 102900.0 1381950.0 ;
      RECT  101850.0 1397250.0 102750.0 1389750.0 ;
      RECT  97050.0 1392300.0 97950.0 1391400.0 ;
      RECT  101850.0 1392300.0 102750.0 1391400.0 ;
      RECT  97050.0 1391850.0 97950.0 1389750.0 ;
      RECT  97500.0 1392300.0 102300.0 1391400.0 ;
      RECT  101850.0 1397250.0 102750.0 1391850.0 ;
      RECT  96900.0 1389750.0 98100.0 1388550.0 ;
      RECT  101700.0 1389750.0 102900.0 1388550.0 ;
      RECT  101700.0 1398450.0 102900.0 1397250.0 ;
      RECT  101700.0 1392450.0 102900.0 1391250.0 ;
      RECT  101850.0 1403550.0 102750.0 1411050.0 ;
      RECT  97050.0 1408500.0 97950.0 1409400.0 ;
      RECT  101850.0 1408500.0 102750.0 1409400.0 ;
      RECT  97050.0 1408950.0 97950.0 1411050.0 ;
      RECT  97500.0 1408500.0 102300.0 1409400.0 ;
      RECT  101850.0 1403550.0 102750.0 1408950.0 ;
      RECT  96900.0 1411050.0 98100.0 1412250.0 ;
      RECT  101700.0 1411050.0 102900.0 1412250.0 ;
      RECT  101700.0 1402350.0 102900.0 1403550.0 ;
      RECT  101700.0 1408350.0 102900.0 1409550.0 ;
      RECT  101850.0 1424850.0 102750.0 1417350.0 ;
      RECT  97050.0 1419900.0 97950.0 1419000.0 ;
      RECT  101850.0 1419900.0 102750.0 1419000.0 ;
      RECT  97050.0 1419450.0 97950.0 1417350.0 ;
      RECT  97500.0 1419900.0 102300.0 1419000.0 ;
      RECT  101850.0 1424850.0 102750.0 1419450.0 ;
      RECT  96900.0 1417350.0 98100.0 1416150.0 ;
      RECT  101700.0 1417350.0 102900.0 1416150.0 ;
      RECT  101700.0 1426050.0 102900.0 1424850.0 ;
      RECT  101700.0 1420050.0 102900.0 1418850.0 ;
      RECT  101850.0 1431150.0 102750.0 1438650.0 ;
      RECT  97050.0 1436100.0 97950.0 1437000.0 ;
      RECT  101850.0 1436100.0 102750.0 1437000.0 ;
      RECT  97050.0 1436550.0 97950.0 1438650.0 ;
      RECT  97500.0 1436100.0 102300.0 1437000.0 ;
      RECT  101850.0 1431150.0 102750.0 1436550.0 ;
      RECT  96900.0 1438650.0 98100.0 1439850.0 ;
      RECT  101700.0 1438650.0 102900.0 1439850.0 ;
      RECT  101700.0 1429950.0 102900.0 1431150.0 ;
      RECT  101700.0 1435950.0 102900.0 1437150.0 ;
      RECT  101850.0 1452450.0 102750.0 1444950.0 ;
      RECT  97050.0 1447500.0 97950.0 1446600.0 ;
      RECT  101850.0 1447500.0 102750.0 1446600.0 ;
      RECT  97050.0 1447050.0 97950.0 1444950.0 ;
      RECT  97500.0 1447500.0 102300.0 1446600.0 ;
      RECT  101850.0 1452450.0 102750.0 1447050.0 ;
      RECT  96900.0 1444950.0 98100.0 1443750.0 ;
      RECT  101700.0 1444950.0 102900.0 1443750.0 ;
      RECT  101700.0 1453650.0 102900.0 1452450.0 ;
      RECT  101700.0 1447650.0 102900.0 1446450.0 ;
      RECT  101850.0 1458750.0 102750.0 1466250.0 ;
      RECT  97050.0 1463700.0 97950.0 1464600.0 ;
      RECT  101850.0 1463700.0 102750.0 1464600.0 ;
      RECT  97050.0 1464150.0 97950.0 1466250.0 ;
      RECT  97500.0 1463700.0 102300.0 1464600.0 ;
      RECT  101850.0 1458750.0 102750.0 1464150.0 ;
      RECT  96900.0 1466250.0 98100.0 1467450.0 ;
      RECT  101700.0 1466250.0 102900.0 1467450.0 ;
      RECT  101700.0 1457550.0 102900.0 1458750.0 ;
      RECT  101700.0 1463550.0 102900.0 1464750.0 ;
      RECT  101850.0 1480050.0 102750.0 1472550.0 ;
      RECT  97050.0 1475100.0 97950.0 1474200.0 ;
      RECT  101850.0 1475100.0 102750.0 1474200.0 ;
      RECT  97050.0 1474650.0 97950.0 1472550.0 ;
      RECT  97500.0 1475100.0 102300.0 1474200.0 ;
      RECT  101850.0 1480050.0 102750.0 1474650.0 ;
      RECT  96900.0 1472550.0 98100.0 1471350.0 ;
      RECT  101700.0 1472550.0 102900.0 1471350.0 ;
      RECT  101700.0 1481250.0 102900.0 1480050.0 ;
      RECT  101700.0 1475250.0 102900.0 1474050.0 ;
      RECT  101850.0 1486350.0 102750.0 1493850.0 ;
      RECT  97050.0 1491300.0 97950.0 1492200.0 ;
      RECT  101850.0 1491300.0 102750.0 1492200.0 ;
      RECT  97050.0 1491750.0 97950.0 1493850.0 ;
      RECT  97500.0 1491300.0 102300.0 1492200.0 ;
      RECT  101850.0 1486350.0 102750.0 1491750.0 ;
      RECT  96900.0 1493850.0 98100.0 1495050.0 ;
      RECT  101700.0 1493850.0 102900.0 1495050.0 ;
      RECT  101700.0 1485150.0 102900.0 1486350.0 ;
      RECT  101700.0 1491150.0 102900.0 1492350.0 ;
      RECT  101850.0 1507650.0 102750.0 1500150.0 ;
      RECT  97050.0 1502700.0 97950.0 1501800.0 ;
      RECT  101850.0 1502700.0 102750.0 1501800.0 ;
      RECT  97050.0 1502250.0 97950.0 1500150.0 ;
      RECT  97500.0 1502700.0 102300.0 1501800.0 ;
      RECT  101850.0 1507650.0 102750.0 1502250.0 ;
      RECT  96900.0 1500150.0 98100.0 1498950.0 ;
      RECT  101700.0 1500150.0 102900.0 1498950.0 ;
      RECT  101700.0 1508850.0 102900.0 1507650.0 ;
      RECT  101700.0 1502850.0 102900.0 1501650.0 ;
      RECT  101850.0 1513950.0 102750.0 1521450.0 ;
      RECT  97050.0 1518900.0 97950.0 1519800.0 ;
      RECT  101850.0 1518900.0 102750.0 1519800.0 ;
      RECT  97050.0 1519350.0 97950.0 1521450.0 ;
      RECT  97500.0 1518900.0 102300.0 1519800.0 ;
      RECT  101850.0 1513950.0 102750.0 1519350.0 ;
      RECT  96900.0 1521450.0 98100.0 1522650.0 ;
      RECT  101700.0 1521450.0 102900.0 1522650.0 ;
      RECT  101700.0 1512750.0 102900.0 1513950.0 ;
      RECT  101700.0 1518750.0 102900.0 1519950.0 ;
      RECT  101850.0 1535250.0 102750.0 1527750.0 ;
      RECT  97050.0 1530300.0 97950.0 1529400.0 ;
      RECT  101850.0 1530300.0 102750.0 1529400.0 ;
      RECT  97050.0 1529850.0 97950.0 1527750.0 ;
      RECT  97500.0 1530300.0 102300.0 1529400.0 ;
      RECT  101850.0 1535250.0 102750.0 1529850.0 ;
      RECT  96900.0 1527750.0 98100.0 1526550.0 ;
      RECT  101700.0 1527750.0 102900.0 1526550.0 ;
      RECT  101700.0 1536450.0 102900.0 1535250.0 ;
      RECT  101700.0 1530450.0 102900.0 1529250.0 ;
      RECT  101850.0 1541550.0 102750.0 1549050.0 ;
      RECT  97050.0 1546500.0 97950.0 1547400.0 ;
      RECT  101850.0 1546500.0 102750.0 1547400.0 ;
      RECT  97050.0 1546950.0 97950.0 1549050.0 ;
      RECT  97500.0 1546500.0 102300.0 1547400.0 ;
      RECT  101850.0 1541550.0 102750.0 1546950.0 ;
      RECT  96900.0 1549050.0 98100.0 1550250.0 ;
      RECT  101700.0 1549050.0 102900.0 1550250.0 ;
      RECT  101700.0 1540350.0 102900.0 1541550.0 ;
      RECT  101700.0 1546350.0 102900.0 1547550.0 ;
      RECT  101850.0 1562850.0 102750.0 1555350.0 ;
      RECT  97050.0 1557900.0 97950.0 1557000.0 ;
      RECT  101850.0 1557900.0 102750.0 1557000.0 ;
      RECT  97050.0 1557450.0 97950.0 1555350.0 ;
      RECT  97500.0 1557900.0 102300.0 1557000.0 ;
      RECT  101850.0 1562850.0 102750.0 1557450.0 ;
      RECT  96900.0 1555350.0 98100.0 1554150.0 ;
      RECT  101700.0 1555350.0 102900.0 1554150.0 ;
      RECT  101700.0 1564050.0 102900.0 1562850.0 ;
      RECT  101700.0 1558050.0 102900.0 1556850.0 ;
      RECT  101850.0 1569150.0 102750.0 1576650.0 ;
      RECT  97050.0 1574100.0 97950.0 1575000.0 ;
      RECT  101850.0 1574100.0 102750.0 1575000.0 ;
      RECT  97050.0 1574550.0 97950.0 1576650.0 ;
      RECT  97500.0 1574100.0 102300.0 1575000.0 ;
      RECT  101850.0 1569150.0 102750.0 1574550.0 ;
      RECT  96900.0 1576650.0 98100.0 1577850.0 ;
      RECT  101700.0 1576650.0 102900.0 1577850.0 ;
      RECT  101700.0 1567950.0 102900.0 1569150.0 ;
      RECT  101700.0 1573950.0 102900.0 1575150.0 ;
      RECT  101850.0 1590450.0 102750.0 1582950.0 ;
      RECT  97050.0 1585500.0 97950.0 1584600.0 ;
      RECT  101850.0 1585500.0 102750.0 1584600.0 ;
      RECT  97050.0 1585050.0 97950.0 1582950.0 ;
      RECT  97500.0 1585500.0 102300.0 1584600.0 ;
      RECT  101850.0 1590450.0 102750.0 1585050.0 ;
      RECT  96900.0 1582950.0 98100.0 1581750.0 ;
      RECT  101700.0 1582950.0 102900.0 1581750.0 ;
      RECT  101700.0 1591650.0 102900.0 1590450.0 ;
      RECT  101700.0 1585650.0 102900.0 1584450.0 ;
      RECT  101850.0 1596750.0 102750.0 1604250.0 ;
      RECT  97050.0 1601700.0 97950.0 1602600.0 ;
      RECT  101850.0 1601700.0 102750.0 1602600.0 ;
      RECT  97050.0 1602150.0 97950.0 1604250.0 ;
      RECT  97500.0 1601700.0 102300.0 1602600.0 ;
      RECT  101850.0 1596750.0 102750.0 1602150.0 ;
      RECT  96900.0 1604250.0 98100.0 1605450.0 ;
      RECT  101700.0 1604250.0 102900.0 1605450.0 ;
      RECT  101700.0 1595550.0 102900.0 1596750.0 ;
      RECT  101700.0 1601550.0 102900.0 1602750.0 ;
      RECT  101850.0 1618050.0 102750.0 1610550.0 ;
      RECT  97050.0 1613100.0 97950.0 1612200.0 ;
      RECT  101850.0 1613100.0 102750.0 1612200.0 ;
      RECT  97050.0 1612650.0 97950.0 1610550.0 ;
      RECT  97500.0 1613100.0 102300.0 1612200.0 ;
      RECT  101850.0 1618050.0 102750.0 1612650.0 ;
      RECT  96900.0 1610550.0 98100.0 1609350.0 ;
      RECT  101700.0 1610550.0 102900.0 1609350.0 ;
      RECT  101700.0 1619250.0 102900.0 1618050.0 ;
      RECT  101700.0 1613250.0 102900.0 1612050.0 ;
      RECT  101850.0 1624350.0 102750.0 1631850.0 ;
      RECT  97050.0 1629300.0 97950.0 1630200.0 ;
      RECT  101850.0 1629300.0 102750.0 1630200.0 ;
      RECT  97050.0 1629750.0 97950.0 1631850.0 ;
      RECT  97500.0 1629300.0 102300.0 1630200.0 ;
      RECT  101850.0 1624350.0 102750.0 1629750.0 ;
      RECT  96900.0 1631850.0 98100.0 1633050.0 ;
      RECT  101700.0 1631850.0 102900.0 1633050.0 ;
      RECT  101700.0 1623150.0 102900.0 1624350.0 ;
      RECT  101700.0 1629150.0 102900.0 1630350.0 ;
      RECT  101850.0 1645650.0 102750.0 1638150.0 ;
      RECT  97050.0 1640700.0 97950.0 1639800.0 ;
      RECT  101850.0 1640700.0 102750.0 1639800.0 ;
      RECT  97050.0 1640250.0 97950.0 1638150.0 ;
      RECT  97500.0 1640700.0 102300.0 1639800.0 ;
      RECT  101850.0 1645650.0 102750.0 1640250.0 ;
      RECT  96900.0 1638150.0 98100.0 1636950.0 ;
      RECT  101700.0 1638150.0 102900.0 1636950.0 ;
      RECT  101700.0 1646850.0 102900.0 1645650.0 ;
      RECT  101700.0 1640850.0 102900.0 1639650.0 ;
      RECT  101850.0 1651950.0 102750.0 1659450.0 ;
      RECT  97050.0 1656900.0 97950.0 1657800.0 ;
      RECT  101850.0 1656900.0 102750.0 1657800.0 ;
      RECT  97050.0 1657350.0 97950.0 1659450.0 ;
      RECT  97500.0 1656900.0 102300.0 1657800.0 ;
      RECT  101850.0 1651950.0 102750.0 1657350.0 ;
      RECT  96900.0 1659450.0 98100.0 1660650.0 ;
      RECT  101700.0 1659450.0 102900.0 1660650.0 ;
      RECT  101700.0 1650750.0 102900.0 1651950.0 ;
      RECT  101700.0 1656750.0 102900.0 1657950.0 ;
      RECT  101850.0 1673250.0 102750.0 1665750.0 ;
      RECT  97050.0 1668300.0 97950.0 1667400.0 ;
      RECT  101850.0 1668300.0 102750.0 1667400.0 ;
      RECT  97050.0 1667850.0 97950.0 1665750.0 ;
      RECT  97500.0 1668300.0 102300.0 1667400.0 ;
      RECT  101850.0 1673250.0 102750.0 1667850.0 ;
      RECT  96900.0 1665750.0 98100.0 1664550.0 ;
      RECT  101700.0 1665750.0 102900.0 1664550.0 ;
      RECT  101700.0 1674450.0 102900.0 1673250.0 ;
      RECT  101700.0 1668450.0 102900.0 1667250.0 ;
      RECT  101850.0 1679550.0 102750.0 1687050.0 ;
      RECT  97050.0 1684500.0 97950.0 1685400.0 ;
      RECT  101850.0 1684500.0 102750.0 1685400.0 ;
      RECT  97050.0 1684950.0 97950.0 1687050.0 ;
      RECT  97500.0 1684500.0 102300.0 1685400.0 ;
      RECT  101850.0 1679550.0 102750.0 1684950.0 ;
      RECT  96900.0 1687050.0 98100.0 1688250.0 ;
      RECT  101700.0 1687050.0 102900.0 1688250.0 ;
      RECT  101700.0 1678350.0 102900.0 1679550.0 ;
      RECT  101700.0 1684350.0 102900.0 1685550.0 ;
      RECT  101850.0 1700850.0 102750.0 1693350.0 ;
      RECT  97050.0 1695900.0 97950.0 1695000.0 ;
      RECT  101850.0 1695900.0 102750.0 1695000.0 ;
      RECT  97050.0 1695450.0 97950.0 1693350.0 ;
      RECT  97500.0 1695900.0 102300.0 1695000.0 ;
      RECT  101850.0 1700850.0 102750.0 1695450.0 ;
      RECT  96900.0 1693350.0 98100.0 1692150.0 ;
      RECT  101700.0 1693350.0 102900.0 1692150.0 ;
      RECT  101700.0 1702050.0 102900.0 1700850.0 ;
      RECT  101700.0 1696050.0 102900.0 1694850.0 ;
      RECT  101850.0 1707150.0 102750.0 1714650.0 ;
      RECT  97050.0 1712100.0 97950.0 1713000.0 ;
      RECT  101850.0 1712100.0 102750.0 1713000.0 ;
      RECT  97050.0 1712550.0 97950.0 1714650.0 ;
      RECT  97500.0 1712100.0 102300.0 1713000.0 ;
      RECT  101850.0 1707150.0 102750.0 1712550.0 ;
      RECT  96900.0 1714650.0 98100.0 1715850.0 ;
      RECT  101700.0 1714650.0 102900.0 1715850.0 ;
      RECT  101700.0 1705950.0 102900.0 1707150.0 ;
      RECT  101700.0 1711950.0 102900.0 1713150.0 ;
      RECT  101850.0 1728450.0 102750.0 1720950.0 ;
      RECT  97050.0 1723500.0 97950.0 1722600.0 ;
      RECT  101850.0 1723500.0 102750.0 1722600.0 ;
      RECT  97050.0 1723050.0 97950.0 1720950.0 ;
      RECT  97500.0 1723500.0 102300.0 1722600.0 ;
      RECT  101850.0 1728450.0 102750.0 1723050.0 ;
      RECT  96900.0 1720950.0 98100.0 1719750.0 ;
      RECT  101700.0 1720950.0 102900.0 1719750.0 ;
      RECT  101700.0 1729650.0 102900.0 1728450.0 ;
      RECT  101700.0 1723650.0 102900.0 1722450.0 ;
      RECT  101850.0 1734750.0 102750.0 1742250.0 ;
      RECT  97050.0 1739700.0 97950.0 1740600.0 ;
      RECT  101850.0 1739700.0 102750.0 1740600.0 ;
      RECT  97050.0 1740150.0 97950.0 1742250.0 ;
      RECT  97500.0 1739700.0 102300.0 1740600.0 ;
      RECT  101850.0 1734750.0 102750.0 1740150.0 ;
      RECT  96900.0 1742250.0 98100.0 1743450.0 ;
      RECT  101700.0 1742250.0 102900.0 1743450.0 ;
      RECT  101700.0 1733550.0 102900.0 1734750.0 ;
      RECT  101700.0 1739550.0 102900.0 1740750.0 ;
      RECT  101850.0 1756050.0 102750.0 1748550.0 ;
      RECT  97050.0 1751100.0 97950.0 1750200.0 ;
      RECT  101850.0 1751100.0 102750.0 1750200.0 ;
      RECT  97050.0 1750650.0 97950.0 1748550.0 ;
      RECT  97500.0 1751100.0 102300.0 1750200.0 ;
      RECT  101850.0 1756050.0 102750.0 1750650.0 ;
      RECT  96900.0 1748550.0 98100.0 1747350.0 ;
      RECT  101700.0 1748550.0 102900.0 1747350.0 ;
      RECT  101700.0 1757250.0 102900.0 1756050.0 ;
      RECT  101700.0 1751250.0 102900.0 1750050.0 ;
      RECT  101850.0 1762350.0 102750.0 1769850.0 ;
      RECT  97050.0 1767300.0 97950.0 1768200.0 ;
      RECT  101850.0 1767300.0 102750.0 1768200.0 ;
      RECT  97050.0 1767750.0 97950.0 1769850.0 ;
      RECT  97500.0 1767300.0 102300.0 1768200.0 ;
      RECT  101850.0 1762350.0 102750.0 1767750.0 ;
      RECT  96900.0 1769850.0 98100.0 1771050.0 ;
      RECT  101700.0 1769850.0 102900.0 1771050.0 ;
      RECT  101700.0 1761150.0 102900.0 1762350.0 ;
      RECT  101700.0 1767150.0 102900.0 1768350.0 ;
      RECT  101850.0 1783650.0 102750.0 1776150.0 ;
      RECT  97050.0 1778700.0 97950.0 1777800.0 ;
      RECT  101850.0 1778700.0 102750.0 1777800.0 ;
      RECT  97050.0 1778250.0 97950.0 1776150.0 ;
      RECT  97500.0 1778700.0 102300.0 1777800.0 ;
      RECT  101850.0 1783650.0 102750.0 1778250.0 ;
      RECT  96900.0 1776150.0 98100.0 1774950.0 ;
      RECT  101700.0 1776150.0 102900.0 1774950.0 ;
      RECT  101700.0 1784850.0 102900.0 1783650.0 ;
      RECT  101700.0 1778850.0 102900.0 1777650.0 ;
      RECT  101850.0 1789950.0 102750.0 1797450.0 ;
      RECT  97050.0 1794900.0 97950.0 1795800.0 ;
      RECT  101850.0 1794900.0 102750.0 1795800.0 ;
      RECT  97050.0 1795350.0 97950.0 1797450.0 ;
      RECT  97500.0 1794900.0 102300.0 1795800.0 ;
      RECT  101850.0 1789950.0 102750.0 1795350.0 ;
      RECT  96900.0 1797450.0 98100.0 1798650.0 ;
      RECT  101700.0 1797450.0 102900.0 1798650.0 ;
      RECT  101700.0 1788750.0 102900.0 1789950.0 ;
      RECT  101700.0 1794750.0 102900.0 1795950.0 ;
      RECT  101850.0 1811250.0 102750.0 1803750.0 ;
      RECT  97050.0 1806300.0 97950.0 1805400.0 ;
      RECT  101850.0 1806300.0 102750.0 1805400.0 ;
      RECT  97050.0 1805850.0 97950.0 1803750.0 ;
      RECT  97500.0 1806300.0 102300.0 1805400.0 ;
      RECT  101850.0 1811250.0 102750.0 1805850.0 ;
      RECT  96900.0 1803750.0 98100.0 1802550.0 ;
      RECT  101700.0 1803750.0 102900.0 1802550.0 ;
      RECT  101700.0 1812450.0 102900.0 1811250.0 ;
      RECT  101700.0 1806450.0 102900.0 1805250.0 ;
      RECT  101850.0 1817550.0 102750.0 1825050.0 ;
      RECT  97050.0 1822500.0 97950.0 1823400.0 ;
      RECT  101850.0 1822500.0 102750.0 1823400.0 ;
      RECT  97050.0 1822950.0 97950.0 1825050.0 ;
      RECT  97500.0 1822500.0 102300.0 1823400.0 ;
      RECT  101850.0 1817550.0 102750.0 1822950.0 ;
      RECT  96900.0 1825050.0 98100.0 1826250.0 ;
      RECT  101700.0 1825050.0 102900.0 1826250.0 ;
      RECT  101700.0 1816350.0 102900.0 1817550.0 ;
      RECT  101700.0 1822350.0 102900.0 1823550.0 ;
      RECT  101850.0 1838850.0 102750.0 1831350.0 ;
      RECT  97050.0 1833900.0 97950.0 1833000.0 ;
      RECT  101850.0 1833900.0 102750.0 1833000.0 ;
      RECT  97050.0 1833450.0 97950.0 1831350.0 ;
      RECT  97500.0 1833900.0 102300.0 1833000.0 ;
      RECT  101850.0 1838850.0 102750.0 1833450.0 ;
      RECT  96900.0 1831350.0 98100.0 1830150.0 ;
      RECT  101700.0 1831350.0 102900.0 1830150.0 ;
      RECT  101700.0 1840050.0 102900.0 1838850.0 ;
      RECT  101700.0 1834050.0 102900.0 1832850.0 ;
      RECT  101850.0 1845150.0 102750.0 1852650.0 ;
      RECT  97050.0 1850100.0 97950.0 1851000.0 ;
      RECT  101850.0 1850100.0 102750.0 1851000.0 ;
      RECT  97050.0 1850550.0 97950.0 1852650.0 ;
      RECT  97500.0 1850100.0 102300.0 1851000.0 ;
      RECT  101850.0 1845150.0 102750.0 1850550.0 ;
      RECT  96900.0 1852650.0 98100.0 1853850.0 ;
      RECT  101700.0 1852650.0 102900.0 1853850.0 ;
      RECT  101700.0 1843950.0 102900.0 1845150.0 ;
      RECT  101700.0 1849950.0 102900.0 1851150.0 ;
      RECT  101850.0 1866450.0 102750.0 1858950.0 ;
      RECT  97050.0 1861500.0 97950.0 1860600.0 ;
      RECT  101850.0 1861500.0 102750.0 1860600.0 ;
      RECT  97050.0 1861050.0 97950.0 1858950.0 ;
      RECT  97500.0 1861500.0 102300.0 1860600.0 ;
      RECT  101850.0 1866450.0 102750.0 1861050.0 ;
      RECT  96900.0 1858950.0 98100.0 1857750.0 ;
      RECT  101700.0 1858950.0 102900.0 1857750.0 ;
      RECT  101700.0 1867650.0 102900.0 1866450.0 ;
      RECT  101700.0 1861650.0 102900.0 1860450.0 ;
      RECT  101850.0 1872750.0 102750.0 1880250.0 ;
      RECT  97050.0 1877700.0 97950.0 1878600.0 ;
      RECT  101850.0 1877700.0 102750.0 1878600.0 ;
      RECT  97050.0 1878150.0 97950.0 1880250.0 ;
      RECT  97500.0 1877700.0 102300.0 1878600.0 ;
      RECT  101850.0 1872750.0 102750.0 1878150.0 ;
      RECT  96900.0 1880250.0 98100.0 1881450.0 ;
      RECT  101700.0 1880250.0 102900.0 1881450.0 ;
      RECT  101700.0 1871550.0 102900.0 1872750.0 ;
      RECT  101700.0 1877550.0 102900.0 1878750.0 ;
      RECT  101850.0 1894050.0 102750.0 1886550.0 ;
      RECT  97050.0 1889100.0 97950.0 1888200.0 ;
      RECT  101850.0 1889100.0 102750.0 1888200.0 ;
      RECT  97050.0 1888650.0 97950.0 1886550.0 ;
      RECT  97500.0 1889100.0 102300.0 1888200.0 ;
      RECT  101850.0 1894050.0 102750.0 1888650.0 ;
      RECT  96900.0 1886550.0 98100.0 1885350.0 ;
      RECT  101700.0 1886550.0 102900.0 1885350.0 ;
      RECT  101700.0 1895250.0 102900.0 1894050.0 ;
      RECT  101700.0 1889250.0 102900.0 1888050.0 ;
      RECT  101850.0 1900350.0 102750.0 1907850.0 ;
      RECT  97050.0 1905300.0 97950.0 1906200.0 ;
      RECT  101850.0 1905300.0 102750.0 1906200.0 ;
      RECT  97050.0 1905750.0 97950.0 1907850.0 ;
      RECT  97500.0 1905300.0 102300.0 1906200.0 ;
      RECT  101850.0 1900350.0 102750.0 1905750.0 ;
      RECT  96900.0 1907850.0 98100.0 1909050.0 ;
      RECT  101700.0 1907850.0 102900.0 1909050.0 ;
      RECT  101700.0 1899150.0 102900.0 1900350.0 ;
      RECT  101700.0 1905150.0 102900.0 1906350.0 ;
      RECT  101850.0 1921650.0 102750.0 1914150.0 ;
      RECT  97050.0 1916700.0 97950.0 1915800.0 ;
      RECT  101850.0 1916700.0 102750.0 1915800.0 ;
      RECT  97050.0 1916250.0 97950.0 1914150.0 ;
      RECT  97500.0 1916700.0 102300.0 1915800.0 ;
      RECT  101850.0 1921650.0 102750.0 1916250.0 ;
      RECT  96900.0 1914150.0 98100.0 1912950.0 ;
      RECT  101700.0 1914150.0 102900.0 1912950.0 ;
      RECT  101700.0 1922850.0 102900.0 1921650.0 ;
      RECT  101700.0 1916850.0 102900.0 1915650.0 ;
      RECT  101850.0 1927950.0 102750.0 1935450.0 ;
      RECT  97050.0 1932900.0 97950.0 1933800.0 ;
      RECT  101850.0 1932900.0 102750.0 1933800.0 ;
      RECT  97050.0 1933350.0 97950.0 1935450.0 ;
      RECT  97500.0 1932900.0 102300.0 1933800.0 ;
      RECT  101850.0 1927950.0 102750.0 1933350.0 ;
      RECT  96900.0 1935450.0 98100.0 1936650.0 ;
      RECT  101700.0 1935450.0 102900.0 1936650.0 ;
      RECT  101700.0 1926750.0 102900.0 1927950.0 ;
      RECT  101700.0 1932750.0 102900.0 1933950.0 ;
      RECT  101850.0 1949250.0 102750.0 1941750.0 ;
      RECT  97050.0 1944300.0 97950.0 1943400.0 ;
      RECT  101850.0 1944300.0 102750.0 1943400.0 ;
      RECT  97050.0 1943850.0 97950.0 1941750.0 ;
      RECT  97500.0 1944300.0 102300.0 1943400.0 ;
      RECT  101850.0 1949250.0 102750.0 1943850.0 ;
      RECT  96900.0 1941750.0 98100.0 1940550.0 ;
      RECT  101700.0 1941750.0 102900.0 1940550.0 ;
      RECT  101700.0 1950450.0 102900.0 1949250.0 ;
      RECT  101700.0 1944450.0 102900.0 1943250.0 ;
      RECT  101850.0 1955550.0 102750.0 1963050.0 ;
      RECT  97050.0 1960500.0 97950.0 1961400.0 ;
      RECT  101850.0 1960500.0 102750.0 1961400.0 ;
      RECT  97050.0 1960950.0 97950.0 1963050.0 ;
      RECT  97500.0 1960500.0 102300.0 1961400.0 ;
      RECT  101850.0 1955550.0 102750.0 1960950.0 ;
      RECT  96900.0 1963050.0 98100.0 1964250.0 ;
      RECT  101700.0 1963050.0 102900.0 1964250.0 ;
      RECT  101700.0 1954350.0 102900.0 1955550.0 ;
      RECT  101700.0 1960350.0 102900.0 1961550.0 ;
      RECT  101850.0 1976850.0 102750.0 1969350.0 ;
      RECT  97050.0 1971900.0 97950.0 1971000.0 ;
      RECT  101850.0 1971900.0 102750.0 1971000.0 ;
      RECT  97050.0 1971450.0 97950.0 1969350.0 ;
      RECT  97500.0 1971900.0 102300.0 1971000.0 ;
      RECT  101850.0 1976850.0 102750.0 1971450.0 ;
      RECT  96900.0 1969350.0 98100.0 1968150.0 ;
      RECT  101700.0 1969350.0 102900.0 1968150.0 ;
      RECT  101700.0 1978050.0 102900.0 1976850.0 ;
      RECT  101700.0 1972050.0 102900.0 1970850.0 ;
      RECT  101850.0 1983150.0 102750.0 1990650.0 ;
      RECT  97050.0 1988100.0 97950.0 1989000.0 ;
      RECT  101850.0 1988100.0 102750.0 1989000.0 ;
      RECT  97050.0 1988550.0 97950.0 1990650.0 ;
      RECT  97500.0 1988100.0 102300.0 1989000.0 ;
      RECT  101850.0 1983150.0 102750.0 1988550.0 ;
      RECT  96900.0 1990650.0 98100.0 1991850.0 ;
      RECT  101700.0 1990650.0 102900.0 1991850.0 ;
      RECT  101700.0 1981950.0 102900.0 1983150.0 ;
      RECT  101700.0 1987950.0 102900.0 1989150.0 ;
      RECT  101850.0 2004450.0 102750.0 1996950.0 ;
      RECT  97050.0 1999500.0 97950.0 1998600.0 ;
      RECT  101850.0 1999500.0 102750.0 1998600.0 ;
      RECT  97050.0 1999050.0 97950.0 1996950.0 ;
      RECT  97500.0 1999500.0 102300.0 1998600.0 ;
      RECT  101850.0 2004450.0 102750.0 1999050.0 ;
      RECT  96900.0 1996950.0 98100.0 1995750.0 ;
      RECT  101700.0 1996950.0 102900.0 1995750.0 ;
      RECT  101700.0 2005650.0 102900.0 2004450.0 ;
      RECT  101700.0 1999650.0 102900.0 1998450.0 ;
      RECT  101850.0 2010750.0 102750.0 2018250.0 ;
      RECT  97050.0 2015700.0 97950.0 2016600.0 ;
      RECT  101850.0 2015700.0 102750.0 2016600.0 ;
      RECT  97050.0 2016150.0 97950.0 2018250.0 ;
      RECT  97500.0 2015700.0 102300.0 2016600.0 ;
      RECT  101850.0 2010750.0 102750.0 2016150.0 ;
      RECT  96900.0 2018250.0 98100.0 2019450.0 ;
      RECT  101700.0 2018250.0 102900.0 2019450.0 ;
      RECT  101700.0 2009550.0 102900.0 2010750.0 ;
      RECT  101700.0 2015550.0 102900.0 2016750.0 ;
      RECT  101850.0 2032050.0 102750.0 2024550.0 ;
      RECT  97050.0 2027100.0 97950.0 2026200.0 ;
      RECT  101850.0 2027100.0 102750.0 2026200.0 ;
      RECT  97050.0 2026650.0 97950.0 2024550.0 ;
      RECT  97500.0 2027100.0 102300.0 2026200.0 ;
      RECT  101850.0 2032050.0 102750.0 2026650.0 ;
      RECT  96900.0 2024550.0 98100.0 2023350.0 ;
      RECT  101700.0 2024550.0 102900.0 2023350.0 ;
      RECT  101700.0 2033250.0 102900.0 2032050.0 ;
      RECT  101700.0 2027250.0 102900.0 2026050.0 ;
      RECT  101850.0 2038350.0 102750.0 2045850.0 ;
      RECT  97050.0 2043300.0 97950.0 2044200.0 ;
      RECT  101850.0 2043300.0 102750.0 2044200.0 ;
      RECT  97050.0 2043750.0 97950.0 2045850.0 ;
      RECT  97500.0 2043300.0 102300.0 2044200.0 ;
      RECT  101850.0 2038350.0 102750.0 2043750.0 ;
      RECT  96900.0 2045850.0 98100.0 2047050.0 ;
      RECT  101700.0 2045850.0 102900.0 2047050.0 ;
      RECT  101700.0 2037150.0 102900.0 2038350.0 ;
      RECT  101700.0 2043150.0 102900.0 2044350.0 ;
      RECT  101850.0 2059650.0 102750.0 2052150.0 ;
      RECT  97050.0 2054700.0 97950.0 2053800.0 ;
      RECT  101850.0 2054700.0 102750.0 2053800.0 ;
      RECT  97050.0 2054250.0 97950.0 2052150.0 ;
      RECT  97500.0 2054700.0 102300.0 2053800.0 ;
      RECT  101850.0 2059650.0 102750.0 2054250.0 ;
      RECT  96900.0 2052150.0 98100.0 2050950.0 ;
      RECT  101700.0 2052150.0 102900.0 2050950.0 ;
      RECT  101700.0 2060850.0 102900.0 2059650.0 ;
      RECT  101700.0 2054850.0 102900.0 2053650.0 ;
      RECT  101850.0 2065950.0 102750.0 2073450.0 ;
      RECT  97050.0 2070900.0 97950.0 2071800.0 ;
      RECT  101850.0 2070900.0 102750.0 2071800.0 ;
      RECT  97050.0 2071350.0 97950.0 2073450.0 ;
      RECT  97500.0 2070900.0 102300.0 2071800.0 ;
      RECT  101850.0 2065950.0 102750.0 2071350.0 ;
      RECT  96900.0 2073450.0 98100.0 2074650.0 ;
      RECT  101700.0 2073450.0 102900.0 2074650.0 ;
      RECT  101700.0 2064750.0 102900.0 2065950.0 ;
      RECT  101700.0 2070750.0 102900.0 2071950.0 ;
      RECT  101850.0 2087250.0 102750.0 2079750.0 ;
      RECT  97050.0 2082300.0 97950.0 2081400.0 ;
      RECT  101850.0 2082300.0 102750.0 2081400.0 ;
      RECT  97050.0 2081850.0 97950.0 2079750.0 ;
      RECT  97500.0 2082300.0 102300.0 2081400.0 ;
      RECT  101850.0 2087250.0 102750.0 2081850.0 ;
      RECT  96900.0 2079750.0 98100.0 2078550.0 ;
      RECT  101700.0 2079750.0 102900.0 2078550.0 ;
      RECT  101700.0 2088450.0 102900.0 2087250.0 ;
      RECT  101700.0 2082450.0 102900.0 2081250.0 ;
      RECT  101850.0 2093550.0 102750.0 2101050.0 ;
      RECT  97050.0 2098500.0 97950.0 2099400.0 ;
      RECT  101850.0 2098500.0 102750.0 2099400.0 ;
      RECT  97050.0 2098950.0 97950.0 2101050.0 ;
      RECT  97500.0 2098500.0 102300.0 2099400.0 ;
      RECT  101850.0 2093550.0 102750.0 2098950.0 ;
      RECT  96900.0 2101050.0 98100.0 2102250.0 ;
      RECT  101700.0 2101050.0 102900.0 2102250.0 ;
      RECT  101700.0 2092350.0 102900.0 2093550.0 ;
      RECT  101700.0 2098350.0 102900.0 2099550.0 ;
      RECT  101850.0 2114850.0 102750.0 2107350.0 ;
      RECT  97050.0 2109900.0 97950.0 2109000.0 ;
      RECT  101850.0 2109900.0 102750.0 2109000.0 ;
      RECT  97050.0 2109450.0 97950.0 2107350.0 ;
      RECT  97500.0 2109900.0 102300.0 2109000.0 ;
      RECT  101850.0 2114850.0 102750.0 2109450.0 ;
      RECT  96900.0 2107350.0 98100.0 2106150.0 ;
      RECT  101700.0 2107350.0 102900.0 2106150.0 ;
      RECT  101700.0 2116050.0 102900.0 2114850.0 ;
      RECT  101700.0 2110050.0 102900.0 2108850.0 ;
      RECT  101850.0 2121150.0 102750.0 2128650.0 ;
      RECT  97050.0 2126100.0 97950.0 2127000.0 ;
      RECT  101850.0 2126100.0 102750.0 2127000.0 ;
      RECT  97050.0 2126550.0 97950.0 2128650.0 ;
      RECT  97500.0 2126100.0 102300.0 2127000.0 ;
      RECT  101850.0 2121150.0 102750.0 2126550.0 ;
      RECT  96900.0 2128650.0 98100.0 2129850.0 ;
      RECT  101700.0 2128650.0 102900.0 2129850.0 ;
      RECT  101700.0 2119950.0 102900.0 2121150.0 ;
      RECT  101700.0 2125950.0 102900.0 2127150.0 ;
      RECT  101850.0 2142450.0 102750.0 2134950.0 ;
      RECT  97050.0 2137500.0 97950.0 2136600.0 ;
      RECT  101850.0 2137500.0 102750.0 2136600.0 ;
      RECT  97050.0 2137050.0 97950.0 2134950.0 ;
      RECT  97500.0 2137500.0 102300.0 2136600.0 ;
      RECT  101850.0 2142450.0 102750.0 2137050.0 ;
      RECT  96900.0 2134950.0 98100.0 2133750.0 ;
      RECT  101700.0 2134950.0 102900.0 2133750.0 ;
      RECT  101700.0 2143650.0 102900.0 2142450.0 ;
      RECT  101700.0 2137650.0 102900.0 2136450.0 ;
      RECT  60150.0 164400.0 58950.0 165600.0 ;
      RECT  62250.0 178800.0 61050.0 180000.0 ;
      RECT  64350.0 192000.0 63150.0 193200.0 ;
      RECT  66450.0 206400.0 65250.0 207600.0 ;
      RECT  68550.0 219600.0 67350.0 220800.0 ;
      RECT  70650.0 234000.0 69450.0 235200.0 ;
      RECT  72750.0 247200.0 71550.0 248400.0 ;
      RECT  74850.0 261600.0 73650.0 262800.0 ;
      RECT  76950.0 274800.0 75750.0 276000.0 ;
      RECT  79050.0 289200.0 77850.0 290400.0 ;
      RECT  81150.0 302400.0 79950.0 303600.0 ;
      RECT  83250.0 316800.0 82050.0 318000.0 ;
      RECT  85350.0 330000.0 84150.0 331200.0 ;
      RECT  87450.0 344400.0 86250.0 345600.0 ;
      RECT  89550.0 357600.0 88350.0 358800.0 ;
      RECT  91650.0 372000.0 90450.0 373200.0 ;
      RECT  60150.0 387150.0 58950.0 388350.0 ;
      RECT  68550.0 385200.0 67350.0 386400.0 ;
      RECT  76950.0 383250.0 75750.0 384450.0 ;
      RECT  60150.0 397650.0 58950.0 398850.0 ;
      RECT  68550.0 399600.0 67350.0 400800.0 ;
      RECT  79050.0 401550.0 77850.0 402750.0 ;
      RECT  60150.0 414750.0 58950.0 415950.0 ;
      RECT  68550.0 412800.0 67350.0 414000.0 ;
      RECT  81150.0 410850.0 79950.0 412050.0 ;
      RECT  60150.0 425250.0 58950.0 426450.0 ;
      RECT  68550.0 427200.0 67350.0 428400.0 ;
      RECT  83250.0 429150.0 82050.0 430350.0 ;
      RECT  60150.0 442350.0 58950.0 443550.0 ;
      RECT  68550.0 440400.0 67350.0 441600.0 ;
      RECT  85350.0 438450.0 84150.0 439650.0 ;
      RECT  60150.0 452850.0 58950.0 454050.0 ;
      RECT  68550.0 454800.0 67350.0 456000.0 ;
      RECT  87450.0 456750.0 86250.0 457950.0 ;
      RECT  60150.0 469950.0 58950.0 471150.0 ;
      RECT  68550.0 468000.0 67350.0 469200.0 ;
      RECT  89550.0 466050.0 88350.0 467250.0 ;
      RECT  60150.0 480450.0 58950.0 481650.0 ;
      RECT  68550.0 482400.0 67350.0 483600.0 ;
      RECT  91650.0 484350.0 90450.0 485550.0 ;
      RECT  60150.0 497550.0 58950.0 498750.0 ;
      RECT  70650.0 495600.0 69450.0 496800.0 ;
      RECT  76950.0 493650.0 75750.0 494850.0 ;
      RECT  60150.0 508050.0 58950.0 509250.0 ;
      RECT  70650.0 510000.0 69450.0 511200.0 ;
      RECT  79050.0 511950.0 77850.0 513150.0 ;
      RECT  60150.0 525150.0 58950.0 526350.0 ;
      RECT  70650.0 523200.0 69450.0 524400.0 ;
      RECT  81150.0 521250.0 79950.0 522450.0 ;
      RECT  60150.0 535650.0 58950.0 536850.0 ;
      RECT  70650.0 537600.0 69450.0 538800.0 ;
      RECT  83250.0 539550.0 82050.0 540750.0 ;
      RECT  60150.0 552750.0 58950.0 553950.0 ;
      RECT  70650.0 550800.0 69450.0 552000.0 ;
      RECT  85350.0 548850.0 84150.0 550050.0 ;
      RECT  60150.0 563250.0 58950.0 564450.0 ;
      RECT  70650.0 565200.0 69450.0 566400.0 ;
      RECT  87450.0 567150.0 86250.0 568350.0 ;
      RECT  60150.0 580350.0 58950.0 581550.0 ;
      RECT  70650.0 578400.0 69450.0 579600.0 ;
      RECT  89550.0 576450.0 88350.0 577650.0 ;
      RECT  60150.0 590850.0 58950.0 592050.0 ;
      RECT  70650.0 592800.0 69450.0 594000.0 ;
      RECT  91650.0 594750.0 90450.0 595950.0 ;
      RECT  60150.0 607950.0 58950.0 609150.0 ;
      RECT  72750.0 606000.0 71550.0 607200.0 ;
      RECT  76950.0 604050.0 75750.0 605250.0 ;
      RECT  60150.0 618450.0 58950.0 619650.0 ;
      RECT  72750.0 620400.0 71550.0 621600.0 ;
      RECT  79050.0 622350.0 77850.0 623550.0 ;
      RECT  60150.0 635550.0 58950.0 636750.0 ;
      RECT  72750.0 633600.0 71550.0 634800.0 ;
      RECT  81150.0 631650.0 79950.0 632850.0 ;
      RECT  60150.0 646050.0 58950.0 647250.0 ;
      RECT  72750.0 648000.0 71550.0 649200.0 ;
      RECT  83250.0 649950.0 82050.0 651150.0 ;
      RECT  60150.0 663150.0 58950.0 664350.0 ;
      RECT  72750.0 661200.0 71550.0 662400.0 ;
      RECT  85350.0 659250.0 84150.0 660450.0 ;
      RECT  60150.0 673650.0 58950.0 674850.0 ;
      RECT  72750.0 675600.0 71550.0 676800.0 ;
      RECT  87450.0 677550.0 86250.0 678750.0 ;
      RECT  60150.0 690750.0 58950.0 691950.0 ;
      RECT  72750.0 688800.0 71550.0 690000.0 ;
      RECT  89550.0 686850.0 88350.0 688050.0 ;
      RECT  60150.0 701250.0 58950.0 702450.0 ;
      RECT  72750.0 703200.0 71550.0 704400.0 ;
      RECT  91650.0 705150.0 90450.0 706350.0 ;
      RECT  60150.0 718350.0 58950.0 719550.0 ;
      RECT  74850.0 716400.0 73650.0 717600.0 ;
      RECT  76950.0 714450.0 75750.0 715650.0 ;
      RECT  60150.0 728850.0 58950.0 730050.0 ;
      RECT  74850.0 730800.0 73650.0 732000.0 ;
      RECT  79050.0 732750.0 77850.0 733950.0 ;
      RECT  60150.0 745950.0 58950.0 747150.0 ;
      RECT  74850.0 744000.0 73650.0 745200.0 ;
      RECT  81150.0 742050.0 79950.0 743250.0 ;
      RECT  60150.0 756450.0 58950.0 757650.0 ;
      RECT  74850.0 758400.0 73650.0 759600.0 ;
      RECT  83250.0 760350.0 82050.0 761550.0 ;
      RECT  60150.0 773550.0 58950.0 774750.0 ;
      RECT  74850.0 771600.0 73650.0 772800.0 ;
      RECT  85350.0 769650.0 84150.0 770850.0 ;
      RECT  60150.0 784050.0 58950.0 785250.0 ;
      RECT  74850.0 786000.0 73650.0 787200.0 ;
      RECT  87450.0 787950.0 86250.0 789150.0 ;
      RECT  60150.0 801150.0 58950.0 802350.0 ;
      RECT  74850.0 799200.0 73650.0 800400.0 ;
      RECT  89550.0 797250.0 88350.0 798450.0 ;
      RECT  60150.0 811650.0 58950.0 812850.0 ;
      RECT  74850.0 813600.0 73650.0 814800.0 ;
      RECT  91650.0 815550.0 90450.0 816750.0 ;
      RECT  62250.0 828750.0 61050.0 829950.0 ;
      RECT  68550.0 826800.0 67350.0 828000.0 ;
      RECT  76950.0 824850.0 75750.0 826050.0 ;
      RECT  62250.0 839250.0 61050.0 840450.0 ;
      RECT  68550.0 841200.0 67350.0 842400.0 ;
      RECT  79050.0 843150.0 77850.0 844350.0 ;
      RECT  62250.0 856350.0 61050.0 857550.0 ;
      RECT  68550.0 854400.0 67350.0 855600.0 ;
      RECT  81150.0 852450.0 79950.0 853650.0 ;
      RECT  62250.0 866850.0 61050.0 868050.0 ;
      RECT  68550.0 868800.0 67350.0 870000.0 ;
      RECT  83250.0 870750.0 82050.0 871950.0 ;
      RECT  62250.0 883950.0 61050.0 885150.0 ;
      RECT  68550.0 882000.0 67350.0 883200.0 ;
      RECT  85350.0 880050.0 84150.0 881250.0 ;
      RECT  62250.0 894450.0 61050.0 895650.0 ;
      RECT  68550.0 896400.0 67350.0 897600.0 ;
      RECT  87450.0 898350.0 86250.0 899550.0 ;
      RECT  62250.0 911550.0 61050.0 912750.0 ;
      RECT  68550.0 909600.0 67350.0 910800.0 ;
      RECT  89550.0 907650.0 88350.0 908850.0 ;
      RECT  62250.0 922050.0 61050.0 923250.0 ;
      RECT  68550.0 924000.0 67350.0 925200.0 ;
      RECT  91650.0 925950.0 90450.0 927150.0 ;
      RECT  62250.0 939150.0 61050.0 940350.0 ;
      RECT  70650.0 937200.0 69450.0 938400.0 ;
      RECT  76950.0 935250.0 75750.0 936450.0 ;
      RECT  62250.0 949650.0 61050.0 950850.0 ;
      RECT  70650.0 951600.0 69450.0 952800.0 ;
      RECT  79050.0 953550.0 77850.0 954750.0 ;
      RECT  62250.0 966750.0 61050.0 967950.0 ;
      RECT  70650.0 964800.0 69450.0 966000.0 ;
      RECT  81150.0 962850.0 79950.0 964050.0 ;
      RECT  62250.0 977250.0 61050.0 978450.0 ;
      RECT  70650.0 979200.0 69450.0 980400.0 ;
      RECT  83250.0 981150.0 82050.0 982350.0 ;
      RECT  62250.0 994350.0 61050.0 995550.0 ;
      RECT  70650.0 992400.0 69450.0 993600.0 ;
      RECT  85350.0 990450.0 84150.0 991650.0 ;
      RECT  62250.0 1004850.0 61050.0 1006050.0 ;
      RECT  70650.0 1006800.0 69450.0 1008000.0 ;
      RECT  87450.0 1008750.0 86250.0 1009950.0 ;
      RECT  62250.0 1021950.0 61050.0 1023150.0 ;
      RECT  70650.0 1020000.0 69450.0 1021200.0 ;
      RECT  89550.0 1018050.0 88350.0 1019250.0 ;
      RECT  62250.0 1032450.0 61050.0 1033650.0 ;
      RECT  70650.0 1034400.0 69450.0 1035600.0 ;
      RECT  91650.0 1036350.0 90450.0 1037550.0 ;
      RECT  62250.0 1049550.0 61050.0 1050750.0 ;
      RECT  72750.0 1047600.0 71550.0 1048800.0 ;
      RECT  76950.0 1045650.0 75750.0 1046850.0 ;
      RECT  62250.0 1060050.0 61050.0 1061250.0 ;
      RECT  72750.0 1062000.0 71550.0 1063200.0 ;
      RECT  79050.0 1063950.0 77850.0 1065150.0 ;
      RECT  62250.0 1077150.0 61050.0 1078350.0 ;
      RECT  72750.0 1075200.0 71550.0 1076400.0 ;
      RECT  81150.0 1073250.0 79950.0 1074450.0 ;
      RECT  62250.0 1087650.0 61050.0 1088850.0 ;
      RECT  72750.0 1089600.0 71550.0 1090800.0 ;
      RECT  83250.0 1091550.0 82050.0 1092750.0 ;
      RECT  62250.0 1104750.0 61050.0 1105950.0 ;
      RECT  72750.0 1102800.0 71550.0 1104000.0 ;
      RECT  85350.0 1100850.0 84150.0 1102050.0 ;
      RECT  62250.0 1115250.0 61050.0 1116450.0 ;
      RECT  72750.0 1117200.0 71550.0 1118400.0 ;
      RECT  87450.0 1119150.0 86250.0 1120350.0 ;
      RECT  62250.0 1132350.0 61050.0 1133550.0 ;
      RECT  72750.0 1130400.0 71550.0 1131600.0 ;
      RECT  89550.0 1128450.0 88350.0 1129650.0 ;
      RECT  62250.0 1142850.0 61050.0 1144050.0 ;
      RECT  72750.0 1144800.0 71550.0 1146000.0 ;
      RECT  91650.0 1146750.0 90450.0 1147950.0 ;
      RECT  62250.0 1159950.0 61050.0 1161150.0 ;
      RECT  74850.0 1158000.0 73650.0 1159200.0 ;
      RECT  76950.0 1156050.0 75750.0 1157250.0 ;
      RECT  62250.0 1170450.0 61050.0 1171650.0 ;
      RECT  74850.0 1172400.0 73650.0 1173600.0 ;
      RECT  79050.0 1174350.0 77850.0 1175550.0 ;
      RECT  62250.0 1187550.0 61050.0 1188750.0 ;
      RECT  74850.0 1185600.0 73650.0 1186800.0 ;
      RECT  81150.0 1183650.0 79950.0 1184850.0 ;
      RECT  62250.0 1198050.0 61050.0 1199250.0 ;
      RECT  74850.0 1200000.0 73650.0 1201200.0 ;
      RECT  83250.0 1201950.0 82050.0 1203150.0 ;
      RECT  62250.0 1215150.0 61050.0 1216350.0 ;
      RECT  74850.0 1213200.0 73650.0 1214400.0 ;
      RECT  85350.0 1211250.0 84150.0 1212450.0 ;
      RECT  62250.0 1225650.0 61050.0 1226850.0 ;
      RECT  74850.0 1227600.0 73650.0 1228800.0 ;
      RECT  87450.0 1229550.0 86250.0 1230750.0 ;
      RECT  62250.0 1242750.0 61050.0 1243950.0 ;
      RECT  74850.0 1240800.0 73650.0 1242000.0 ;
      RECT  89550.0 1238850.0 88350.0 1240050.0 ;
      RECT  62250.0 1253250.0 61050.0 1254450.0 ;
      RECT  74850.0 1255200.0 73650.0 1256400.0 ;
      RECT  91650.0 1257150.0 90450.0 1258350.0 ;
      RECT  64350.0 1270350.0 63150.0 1271550.0 ;
      RECT  68550.0 1268400.0 67350.0 1269600.0 ;
      RECT  76950.0 1266450.0 75750.0 1267650.0 ;
      RECT  64350.0 1280850.0 63150.0 1282050.0 ;
      RECT  68550.0 1282800.0 67350.0 1284000.0 ;
      RECT  79050.0 1284750.0 77850.0 1285950.0 ;
      RECT  64350.0 1297950.0 63150.0 1299150.0 ;
      RECT  68550.0 1296000.0 67350.0 1297200.0 ;
      RECT  81150.0 1294050.0 79950.0 1295250.0 ;
      RECT  64350.0 1308450.0 63150.0 1309650.0 ;
      RECT  68550.0 1310400.0 67350.0 1311600.0 ;
      RECT  83250.0 1312350.0 82050.0 1313550.0 ;
      RECT  64350.0 1325550.0 63150.0 1326750.0 ;
      RECT  68550.0 1323600.0 67350.0 1324800.0 ;
      RECT  85350.0 1321650.0 84150.0 1322850.0 ;
      RECT  64350.0 1336050.0 63150.0 1337250.0 ;
      RECT  68550.0 1338000.0 67350.0 1339200.0 ;
      RECT  87450.0 1339950.0 86250.0 1341150.0 ;
      RECT  64350.0 1353150.0 63150.0 1354350.0 ;
      RECT  68550.0 1351200.0 67350.0 1352400.0 ;
      RECT  89550.0 1349250.0 88350.0 1350450.0 ;
      RECT  64350.0 1363650.0 63150.0 1364850.0 ;
      RECT  68550.0 1365600.0 67350.0 1366800.0 ;
      RECT  91650.0 1367550.0 90450.0 1368750.0 ;
      RECT  64350.0 1380750.0 63150.0 1381950.0 ;
      RECT  70650.0 1378800.0 69450.0 1380000.0 ;
      RECT  76950.0 1376850.0 75750.0 1378050.0 ;
      RECT  64350.0 1391250.0 63150.0 1392450.0 ;
      RECT  70650.0 1393200.0 69450.0 1394400.0 ;
      RECT  79050.0 1395150.0 77850.0 1396350.0 ;
      RECT  64350.0 1408350.0 63150.0 1409550.0 ;
      RECT  70650.0 1406400.0 69450.0 1407600.0 ;
      RECT  81150.0 1404450.0 79950.0 1405650.0 ;
      RECT  64350.0 1418850.0 63150.0 1420050.0 ;
      RECT  70650.0 1420800.0 69450.0 1422000.0 ;
      RECT  83250.0 1422750.0 82050.0 1423950.0 ;
      RECT  64350.0 1435950.0 63150.0 1437150.0 ;
      RECT  70650.0 1434000.0 69450.0 1435200.0 ;
      RECT  85350.0 1432050.0 84150.0 1433250.0 ;
      RECT  64350.0 1446450.0 63150.0 1447650.0 ;
      RECT  70650.0 1448400.0 69450.0 1449600.0 ;
      RECT  87450.0 1450350.0 86250.0 1451550.0 ;
      RECT  64350.0 1463550.0 63150.0 1464750.0 ;
      RECT  70650.0 1461600.0 69450.0 1462800.0 ;
      RECT  89550.0 1459650.0 88350.0 1460850.0 ;
      RECT  64350.0 1474050.0 63150.0 1475250.0 ;
      RECT  70650.0 1476000.0 69450.0 1477200.0 ;
      RECT  91650.0 1477950.0 90450.0 1479150.0 ;
      RECT  64350.0 1491150.0 63150.0 1492350.0 ;
      RECT  72750.0 1489200.0 71550.0 1490400.0 ;
      RECT  76950.0 1487250.0 75750.0 1488450.0 ;
      RECT  64350.0 1501650.0 63150.0 1502850.0 ;
      RECT  72750.0 1503600.0 71550.0 1504800.0 ;
      RECT  79050.0 1505550.0 77850.0 1506750.0 ;
      RECT  64350.0 1518750.0 63150.0 1519950.0 ;
      RECT  72750.0 1516800.0 71550.0 1518000.0 ;
      RECT  81150.0 1514850.0 79950.0 1516050.0 ;
      RECT  64350.0 1529250.0 63150.0 1530450.0 ;
      RECT  72750.0 1531200.0 71550.0 1532400.0 ;
      RECT  83250.0 1533150.0 82050.0 1534350.0 ;
      RECT  64350.0 1546350.0 63150.0 1547550.0 ;
      RECT  72750.0 1544400.0 71550.0 1545600.0 ;
      RECT  85350.0 1542450.0 84150.0 1543650.0 ;
      RECT  64350.0 1556850.0 63150.0 1558050.0 ;
      RECT  72750.0 1558800.0 71550.0 1560000.0 ;
      RECT  87450.0 1560750.0 86250.0 1561950.0 ;
      RECT  64350.0 1573950.0 63150.0 1575150.0 ;
      RECT  72750.0 1572000.0 71550.0 1573200.0 ;
      RECT  89550.0 1570050.0 88350.0 1571250.0 ;
      RECT  64350.0 1584450.0 63150.0 1585650.0 ;
      RECT  72750.0 1586400.0 71550.0 1587600.0 ;
      RECT  91650.0 1588350.0 90450.0 1589550.0 ;
      RECT  64350.0 1601550.0 63150.0 1602750.0 ;
      RECT  74850.0 1599600.0 73650.0 1600800.0 ;
      RECT  76950.0 1597650.0 75750.0 1598850.0 ;
      RECT  64350.0 1612050.0 63150.0 1613250.0 ;
      RECT  74850.0 1614000.0 73650.0 1615200.0 ;
      RECT  79050.0 1615950.0 77850.0 1617150.0 ;
      RECT  64350.0 1629150.0 63150.0 1630350.0 ;
      RECT  74850.0 1627200.0 73650.0 1628400.0 ;
      RECT  81150.0 1625250.0 79950.0 1626450.0 ;
      RECT  64350.0 1639650.0 63150.0 1640850.0 ;
      RECT  74850.0 1641600.0 73650.0 1642800.0 ;
      RECT  83250.0 1643550.0 82050.0 1644750.0 ;
      RECT  64350.0 1656750.0 63150.0 1657950.0 ;
      RECT  74850.0 1654800.0 73650.0 1656000.0 ;
      RECT  85350.0 1652850.0 84150.0 1654050.0 ;
      RECT  64350.0 1667250.0 63150.0 1668450.0 ;
      RECT  74850.0 1669200.0 73650.0 1670400.0 ;
      RECT  87450.0 1671150.0 86250.0 1672350.0 ;
      RECT  64350.0 1684350.0 63150.0 1685550.0 ;
      RECT  74850.0 1682400.0 73650.0 1683600.0 ;
      RECT  89550.0 1680450.0 88350.0 1681650.0 ;
      RECT  64350.0 1694850.0 63150.0 1696050.0 ;
      RECT  74850.0 1696800.0 73650.0 1698000.0 ;
      RECT  91650.0 1698750.0 90450.0 1699950.0 ;
      RECT  66450.0 1711950.0 65250.0 1713150.0 ;
      RECT  68550.0 1710000.0 67350.0 1711200.0 ;
      RECT  76950.0 1708050.0 75750.0 1709250.0 ;
      RECT  66450.0 1722450.0 65250.0 1723650.0 ;
      RECT  68550.0 1724400.0 67350.0 1725600.0 ;
      RECT  79050.0 1726350.0 77850.0 1727550.0 ;
      RECT  66450.0 1739550.0 65250.0 1740750.0 ;
      RECT  68550.0 1737600.0 67350.0 1738800.0 ;
      RECT  81150.0 1735650.0 79950.0 1736850.0 ;
      RECT  66450.0 1750050.0 65250.0 1751250.0 ;
      RECT  68550.0 1752000.0 67350.0 1753200.0 ;
      RECT  83250.0 1753950.0 82050.0 1755150.0 ;
      RECT  66450.0 1767150.0 65250.0 1768350.0 ;
      RECT  68550.0 1765200.0 67350.0 1766400.0 ;
      RECT  85350.0 1763250.0 84150.0 1764450.0 ;
      RECT  66450.0 1777650.0 65250.0 1778850.0 ;
      RECT  68550.0 1779600.0 67350.0 1780800.0 ;
      RECT  87450.0 1781550.0 86250.0 1782750.0 ;
      RECT  66450.0 1794750.0 65250.0 1795950.0 ;
      RECT  68550.0 1792800.0 67350.0 1794000.0 ;
      RECT  89550.0 1790850.0 88350.0 1792050.0 ;
      RECT  66450.0 1805250.0 65250.0 1806450.0 ;
      RECT  68550.0 1807200.0 67350.0 1808400.0 ;
      RECT  91650.0 1809150.0 90450.0 1810350.0 ;
      RECT  66450.0 1822350.0 65250.0 1823550.0 ;
      RECT  70650.0 1820400.0 69450.0 1821600.0 ;
      RECT  76950.0 1818450.0 75750.0 1819650.0 ;
      RECT  66450.0 1832850.0 65250.0 1834050.0 ;
      RECT  70650.0 1834800.0 69450.0 1836000.0 ;
      RECT  79050.0 1836750.0 77850.0 1837950.0 ;
      RECT  66450.0 1849950.0 65250.0 1851150.0 ;
      RECT  70650.0 1848000.0 69450.0 1849200.0 ;
      RECT  81150.0 1846050.0 79950.0 1847250.0 ;
      RECT  66450.0 1860450.0 65250.0 1861650.0 ;
      RECT  70650.0 1862400.0 69450.0 1863600.0 ;
      RECT  83250.0 1864350.0 82050.0 1865550.0 ;
      RECT  66450.0 1877550.0 65250.0 1878750.0 ;
      RECT  70650.0 1875600.0 69450.0 1876800.0 ;
      RECT  85350.0 1873650.0 84150.0 1874850.0 ;
      RECT  66450.0 1888050.0 65250.0 1889250.0 ;
      RECT  70650.0 1890000.0 69450.0 1891200.0 ;
      RECT  87450.0 1891950.0 86250.0 1893150.0 ;
      RECT  66450.0 1905150.0 65250.0 1906350.0 ;
      RECT  70650.0 1903200.0 69450.0 1904400.0 ;
      RECT  89550.0 1901250.0 88350.0 1902450.0 ;
      RECT  66450.0 1915650.0 65250.0 1916850.0 ;
      RECT  70650.0 1917600.0 69450.0 1918800.0 ;
      RECT  91650.0 1919550.0 90450.0 1920750.0 ;
      RECT  66450.0 1932750.0 65250.0 1933950.0 ;
      RECT  72750.0 1930800.0 71550.0 1932000.0 ;
      RECT  76950.0 1928850.0 75750.0 1930050.0 ;
      RECT  66450.0 1943250.0 65250.0 1944450.0 ;
      RECT  72750.0 1945200.0 71550.0 1946400.0 ;
      RECT  79050.0 1947150.0 77850.0 1948350.0 ;
      RECT  66450.0 1960350.0 65250.0 1961550.0 ;
      RECT  72750.0 1958400.0 71550.0 1959600.0 ;
      RECT  81150.0 1956450.0 79950.0 1957650.0 ;
      RECT  66450.0 1970850.0 65250.0 1972050.0 ;
      RECT  72750.0 1972800.0 71550.0 1974000.0 ;
      RECT  83250.0 1974750.0 82050.0 1975950.0 ;
      RECT  66450.0 1987950.0 65250.0 1989150.0 ;
      RECT  72750.0 1986000.0 71550.0 1987200.0 ;
      RECT  85350.0 1984050.0 84150.0 1985250.0 ;
      RECT  66450.0 1998450.0 65250.0 1999650.0 ;
      RECT  72750.0 2000400.0 71550.0 2001600.0 ;
      RECT  87450.0 2002350.0 86250.0 2003550.0 ;
      RECT  66450.0 2015550.0 65250.0 2016750.0 ;
      RECT  72750.0 2013600.0 71550.0 2014800.0 ;
      RECT  89550.0 2011650.0 88350.0 2012850.0 ;
      RECT  66450.0 2026050.0 65250.0 2027250.0 ;
      RECT  72750.0 2028000.0 71550.0 2029200.0 ;
      RECT  91650.0 2029950.0 90450.0 2031150.0 ;
      RECT  66450.0 2043150.0 65250.0 2044350.0 ;
      RECT  74850.0 2041200.0 73650.0 2042400.0 ;
      RECT  76950.0 2039250.0 75750.0 2040450.0 ;
      RECT  66450.0 2053650.0 65250.0 2054850.0 ;
      RECT  74850.0 2055600.0 73650.0 2056800.0 ;
      RECT  79050.0 2057550.0 77850.0 2058750.0 ;
      RECT  66450.0 2070750.0 65250.0 2071950.0 ;
      RECT  74850.0 2068800.0 73650.0 2070000.0 ;
      RECT  81150.0 2066850.0 79950.0 2068050.0 ;
      RECT  66450.0 2081250.0 65250.0 2082450.0 ;
      RECT  74850.0 2083200.0 73650.0 2084400.0 ;
      RECT  83250.0 2085150.0 82050.0 2086350.0 ;
      RECT  66450.0 2098350.0 65250.0 2099550.0 ;
      RECT  74850.0 2096400.0 73650.0 2097600.0 ;
      RECT  85350.0 2094450.0 84150.0 2095650.0 ;
      RECT  66450.0 2108850.0 65250.0 2110050.0 ;
      RECT  74850.0 2110800.0 73650.0 2112000.0 ;
      RECT  87450.0 2112750.0 86250.0 2113950.0 ;
      RECT  66450.0 2125950.0 65250.0 2127150.0 ;
      RECT  74850.0 2124000.0 73650.0 2125200.0 ;
      RECT  89550.0 2122050.0 88350.0 2123250.0 ;
      RECT  66450.0 2136450.0 65250.0 2137650.0 ;
      RECT  74850.0 2138400.0 73650.0 2139600.0 ;
      RECT  91650.0 2140350.0 90450.0 2141550.0 ;
      RECT  146400.0 158400.0 147300.0 211800.0 ;
      RECT  143400.0 158400.0 144300.0 211800.0 ;
      RECT  146400.0 213600.0 147300.0 267000.0 ;
      RECT  143400.0 213600.0 144300.0 267000.0 ;
      RECT  156600.0 268800.0 157500.0 377400.0 ;
      RECT  153600.0 268800.0 154500.0 377400.0 ;
      RECT  150600.0 268800.0 151500.0 377400.0 ;
      RECT  122550.0 383850.0 123450.0 384750.0 ;
      RECT  122550.0 383400.0 123450.0 384300.0 ;
      RECT  123000.0 383850.0 139200.0 384750.0 ;
      RECT  122550.0 401250.0 123450.0 402150.0 ;
      RECT  122550.0 401700.0 123450.0 402600.0 ;
      RECT  123000.0 401250.0 139200.0 402150.0 ;
      RECT  122550.0 411450.0 123450.0 412350.0 ;
      RECT  122550.0 411000.0 123450.0 411900.0 ;
      RECT  123000.0 411450.0 139200.0 412350.0 ;
      RECT  122550.0 428850.0 123450.0 429750.0 ;
      RECT  122550.0 429300.0 123450.0 430200.0 ;
      RECT  123000.0 428850.0 139200.0 429750.0 ;
      RECT  122550.0 439050.0 123450.0 439950.0 ;
      RECT  122550.0 438600.0 123450.0 439500.0 ;
      RECT  123000.0 439050.0 139200.0 439950.0 ;
      RECT  122550.0 456450.0 123450.0 457350.0 ;
      RECT  122550.0 456900.0 123450.0 457800.0 ;
      RECT  123000.0 456450.0 139200.0 457350.0 ;
      RECT  122550.0 466650.0 123450.0 467550.0 ;
      RECT  122550.0 466200.0 123450.0 467100.0 ;
      RECT  123000.0 466650.0 139200.0 467550.0 ;
      RECT  122550.0 484050.0 123450.0 484950.0 ;
      RECT  122550.0 484500.0 123450.0 485400.0 ;
      RECT  123000.0 484050.0 139200.0 484950.0 ;
      RECT  122550.0 494250.0 123450.0 495150.0 ;
      RECT  122550.0 493800.0 123450.0 494700.0 ;
      RECT  123000.0 494250.0 139200.0 495150.0 ;
      RECT  122550.0 511650.0 123450.0 512550.0 ;
      RECT  122550.0 512100.0 123450.0 513000.0 ;
      RECT  123000.0 511650.0 139200.0 512550.0 ;
      RECT  122550.0 521850.0 123450.0 522750.0 ;
      RECT  122550.0 521400.0 123450.0 522300.0 ;
      RECT  123000.0 521850.0 139200.0 522750.0 ;
      RECT  122550.0 539250.0 123450.0 540150.0 ;
      RECT  122550.0 539700.0 123450.0 540600.0 ;
      RECT  123000.0 539250.0 139200.0 540150.0 ;
      RECT  122550.0 549450.0 123450.0 550350.0 ;
      RECT  122550.0 549000.0 123450.0 549900.0 ;
      RECT  123000.0 549450.0 139200.0 550350.0 ;
      RECT  122550.0 566850.0 123450.0 567750.0 ;
      RECT  122550.0 567300.0 123450.0 568200.0 ;
      RECT  123000.0 566850.0 139200.0 567750.0 ;
      RECT  122550.0 577050.0 123450.0 577950.0 ;
      RECT  122550.0 576600.0 123450.0 577500.0 ;
      RECT  123000.0 577050.0 139200.0 577950.0 ;
      RECT  122550.0 594450.0 123450.0 595350.0 ;
      RECT  122550.0 594900.0 123450.0 595800.0 ;
      RECT  123000.0 594450.0 139200.0 595350.0 ;
      RECT  122550.0 604650.0 123450.0 605550.0 ;
      RECT  122550.0 604200.0 123450.0 605100.0 ;
      RECT  123000.0 604650.0 139200.0 605550.0 ;
      RECT  122550.0 622050.0 123450.0 622950.0 ;
      RECT  122550.0 622500.0 123450.0 623400.0 ;
      RECT  123000.0 622050.0 139200.0 622950.0 ;
      RECT  122550.0 632250.0 123450.0 633150.0 ;
      RECT  122550.0 631800.0 123450.0 632700.0 ;
      RECT  123000.0 632250.0 139200.0 633150.0 ;
      RECT  122550.0 649650.0 123450.0 650550.0 ;
      RECT  122550.0 650100.0 123450.0 651000.0 ;
      RECT  123000.0 649650.0 139200.0 650550.0 ;
      RECT  122550.0 659850.0 123450.0 660750.0 ;
      RECT  122550.0 659400.0 123450.0 660300.0 ;
      RECT  123000.0 659850.0 139200.0 660750.0 ;
      RECT  122550.0 677250.0 123450.0 678150.0 ;
      RECT  122550.0 677700.0 123450.0 678600.0 ;
      RECT  123000.0 677250.0 139200.0 678150.0 ;
      RECT  122550.0 687450.0 123450.0 688350.0 ;
      RECT  122550.0 687000.0 123450.0 687900.0 ;
      RECT  123000.0 687450.0 139200.0 688350.0 ;
      RECT  122550.0 704850.0 123450.0 705750.0 ;
      RECT  122550.0 705300.0 123450.0 706200.0 ;
      RECT  123000.0 704850.0 139200.0 705750.0 ;
      RECT  122550.0 715050.0 123450.0 715950.0 ;
      RECT  122550.0 714600.0 123450.0 715500.0 ;
      RECT  123000.0 715050.0 139200.0 715950.0 ;
      RECT  122550.0 732450.0 123450.0 733350.0 ;
      RECT  122550.0 732900.0 123450.0 733800.0 ;
      RECT  123000.0 732450.0 139200.0 733350.0 ;
      RECT  122550.0 742650.0 123450.0 743550.0 ;
      RECT  122550.0 742200.0 123450.0 743100.0 ;
      RECT  123000.0 742650.0 139200.0 743550.0 ;
      RECT  122550.0 760050.0 123450.0 760950.0 ;
      RECT  122550.0 760500.0 123450.0 761400.0 ;
      RECT  123000.0 760050.0 139200.0 760950.0 ;
      RECT  122550.0 770250.0 123450.0 771150.0 ;
      RECT  122550.0 769800.0 123450.0 770700.0 ;
      RECT  123000.0 770250.0 139200.0 771150.0 ;
      RECT  122550.0 787650.0 123450.0 788550.0 ;
      RECT  122550.0 788100.0 123450.0 789000.0 ;
      RECT  123000.0 787650.0 139200.0 788550.0 ;
      RECT  122550.0 797850.0 123450.0 798750.0 ;
      RECT  122550.0 797400.0 123450.0 798300.0 ;
      RECT  123000.0 797850.0 139200.0 798750.0 ;
      RECT  122550.0 815250.0 123450.0 816150.0 ;
      RECT  122550.0 815700.0 123450.0 816600.0 ;
      RECT  123000.0 815250.0 139200.0 816150.0 ;
      RECT  122550.0 825450.0 123450.0 826350.0 ;
      RECT  122550.0 825000.0 123450.0 825900.0 ;
      RECT  123000.0 825450.0 139200.0 826350.0 ;
      RECT  122550.0 842850.0 123450.0 843750.0 ;
      RECT  122550.0 843300.0 123450.0 844200.0 ;
      RECT  123000.0 842850.0 139200.0 843750.0 ;
      RECT  122550.0 853050.0 123450.0 853950.0 ;
      RECT  122550.0 852600.0 123450.0 853500.0 ;
      RECT  123000.0 853050.0 139200.0 853950.0 ;
      RECT  122550.0 870450.0 123450.0 871350.0 ;
      RECT  122550.0 870900.0 123450.0 871800.0 ;
      RECT  123000.0 870450.0 139200.0 871350.0 ;
      RECT  122550.0 880650.0 123450.0 881550.0 ;
      RECT  122550.0 880200.0 123450.0 881100.0 ;
      RECT  123000.0 880650.0 139200.0 881550.0 ;
      RECT  122550.0 898050.0 123450.0 898950.0 ;
      RECT  122550.0 898500.0 123450.0 899400.0 ;
      RECT  123000.0 898050.0 139200.0 898950.0 ;
      RECT  122550.0 908250.0 123450.0 909150.0 ;
      RECT  122550.0 907800.0 123450.0 908700.0 ;
      RECT  123000.0 908250.0 139200.0 909150.0 ;
      RECT  122550.0 925650.0 123450.0 926550.0 ;
      RECT  122550.0 926100.0 123450.0 927000.0 ;
      RECT  123000.0 925650.0 139200.0 926550.0 ;
      RECT  122550.0 935850.0 123450.0 936750.0 ;
      RECT  122550.0 935400.0 123450.0 936300.0 ;
      RECT  123000.0 935850.0 139200.0 936750.0 ;
      RECT  122550.0 953250.0 123450.0 954150.0 ;
      RECT  122550.0 953700.0 123450.0 954600.0 ;
      RECT  123000.0 953250.0 139200.0 954150.0 ;
      RECT  122550.0 963450.0 123450.0 964350.0 ;
      RECT  122550.0 963000.0 123450.0 963900.0 ;
      RECT  123000.0 963450.0 139200.0 964350.0 ;
      RECT  122550.0 980850.0 123450.0 981750.0 ;
      RECT  122550.0 981300.0 123450.0 982200.0 ;
      RECT  123000.0 980850.0 139200.0 981750.0 ;
      RECT  122550.0 991050.0 123450.0 991950.0 ;
      RECT  122550.0 990600.0 123450.0 991500.0 ;
      RECT  123000.0 991050.0 139200.0 991950.0 ;
      RECT  122550.0 1008450.0 123450.0 1009350.0 ;
      RECT  122550.0 1008900.0 123450.0 1009800.0 ;
      RECT  123000.0 1008450.0 139200.0 1009350.0 ;
      RECT  122550.0 1018650.0 123450.0 1019550.0 ;
      RECT  122550.0 1018200.0 123450.0 1019100.0 ;
      RECT  123000.0 1018650.0 139200.0 1019550.0 ;
      RECT  122550.0 1036050.0 123450.0 1036950.0 ;
      RECT  122550.0 1036500.0 123450.0 1037400.0 ;
      RECT  123000.0 1036050.0 139200.0 1036950.0 ;
      RECT  122550.0 1046250.0 123450.0 1047150.0 ;
      RECT  122550.0 1045800.0 123450.0 1046700.0 ;
      RECT  123000.0 1046250.0 139200.0 1047150.0 ;
      RECT  122550.0 1063650.0 123450.0 1064550.0 ;
      RECT  122550.0 1064100.0 123450.0 1065000.0 ;
      RECT  123000.0 1063650.0 139200.0 1064550.0 ;
      RECT  122550.0 1073850.0 123450.0 1074750.0 ;
      RECT  122550.0 1073400.0 123450.0 1074300.0 ;
      RECT  123000.0 1073850.0 139200.0 1074750.0 ;
      RECT  122550.0 1091250.0 123450.0 1092150.0 ;
      RECT  122550.0 1091700.0 123450.0 1092600.0 ;
      RECT  123000.0 1091250.0 139200.0 1092150.0 ;
      RECT  122550.0 1101450.0 123450.0 1102350.0 ;
      RECT  122550.0 1101000.0 123450.0 1101900.0 ;
      RECT  123000.0 1101450.0 139200.0 1102350.0 ;
      RECT  122550.0 1118850.0 123450.0 1119750.0 ;
      RECT  122550.0 1119300.0 123450.0 1120200.0 ;
      RECT  123000.0 1118850.0 139200.0 1119750.0 ;
      RECT  122550.0 1129050.0 123450.0 1129950.0 ;
      RECT  122550.0 1128600.0 123450.0 1129500.0 ;
      RECT  123000.0 1129050.0 139200.0 1129950.0 ;
      RECT  122550.0 1146450.0 123450.0 1147350.0 ;
      RECT  122550.0 1146900.0 123450.0 1147800.0 ;
      RECT  123000.0 1146450.0 139200.0 1147350.0 ;
      RECT  122550.0 1156650.0 123450.0 1157550.0 ;
      RECT  122550.0 1156200.0 123450.0 1157100.0 ;
      RECT  123000.0 1156650.0 139200.0 1157550.0 ;
      RECT  122550.0 1174050.0 123450.0 1174950.0 ;
      RECT  122550.0 1174500.0 123450.0 1175400.0 ;
      RECT  123000.0 1174050.0 139200.0 1174950.0 ;
      RECT  122550.0 1184250.0 123450.0 1185150.0 ;
      RECT  122550.0 1183800.0 123450.0 1184700.0 ;
      RECT  123000.0 1184250.0 139200.0 1185150.0 ;
      RECT  122550.0 1201650.0 123450.0 1202550.0 ;
      RECT  122550.0 1202100.0 123450.0 1203000.0 ;
      RECT  123000.0 1201650.0 139200.0 1202550.0 ;
      RECT  122550.0 1211850.0 123450.0 1212750.0 ;
      RECT  122550.0 1211400.0 123450.0 1212300.0 ;
      RECT  123000.0 1211850.0 139200.0 1212750.0 ;
      RECT  122550.0 1229250.0 123450.0 1230150.0 ;
      RECT  122550.0 1229700.0 123450.0 1230600.0 ;
      RECT  123000.0 1229250.0 139200.0 1230150.0 ;
      RECT  122550.0 1239450.0 123450.0 1240350.0 ;
      RECT  122550.0 1239000.0 123450.0 1239900.0 ;
      RECT  123000.0 1239450.0 139200.0 1240350.0 ;
      RECT  122550.0 1256850.0 123450.0 1257750.0 ;
      RECT  122550.0 1257300.0 123450.0 1258200.0 ;
      RECT  123000.0 1256850.0 139200.0 1257750.0 ;
      RECT  122550.0 1267050.0 123450.0 1267950.0 ;
      RECT  122550.0 1266600.0 123450.0 1267500.0 ;
      RECT  123000.0 1267050.0 139200.0 1267950.0 ;
      RECT  122550.0 1284450.0 123450.0 1285350.0 ;
      RECT  122550.0 1284900.0 123450.0 1285800.0 ;
      RECT  123000.0 1284450.0 139200.0 1285350.0 ;
      RECT  122550.0 1294650.0 123450.0 1295550.0 ;
      RECT  122550.0 1294200.0 123450.0 1295100.0 ;
      RECT  123000.0 1294650.0 139200.0 1295550.0 ;
      RECT  122550.0 1312050.0 123450.0 1312950.0 ;
      RECT  122550.0 1312500.0 123450.0 1313400.0 ;
      RECT  123000.0 1312050.0 139200.0 1312950.0 ;
      RECT  122550.0 1322250.0 123450.0 1323150.0 ;
      RECT  122550.0 1321800.0 123450.0 1322700.0 ;
      RECT  123000.0 1322250.0 139200.0 1323150.0 ;
      RECT  122550.0 1339650.0 123450.0 1340550.0 ;
      RECT  122550.0 1340100.0 123450.0 1341000.0 ;
      RECT  123000.0 1339650.0 139200.0 1340550.0 ;
      RECT  122550.0 1349850.0 123450.0 1350750.0 ;
      RECT  122550.0 1349400.0 123450.0 1350300.0 ;
      RECT  123000.0 1349850.0 139200.0 1350750.0 ;
      RECT  122550.0 1367250.0 123450.0 1368150.0 ;
      RECT  122550.0 1367700.0 123450.0 1368600.0 ;
      RECT  123000.0 1367250.0 139200.0 1368150.0 ;
      RECT  122550.0 1377450.0 123450.0 1378350.0 ;
      RECT  122550.0 1377000.0 123450.0 1377900.0 ;
      RECT  123000.0 1377450.0 139200.0 1378350.0 ;
      RECT  122550.0 1394850.0 123450.0 1395750.0 ;
      RECT  122550.0 1395300.0 123450.0 1396200.0 ;
      RECT  123000.0 1394850.0 139200.0 1395750.0 ;
      RECT  122550.0 1405050.0 123450.0 1405950.0 ;
      RECT  122550.0 1404600.0 123450.0 1405500.0 ;
      RECT  123000.0 1405050.0 139200.0 1405950.0 ;
      RECT  122550.0 1422450.0 123450.0 1423350.0 ;
      RECT  122550.0 1422900.0 123450.0 1423800.0 ;
      RECT  123000.0 1422450.0 139200.0 1423350.0 ;
      RECT  122550.0 1432650.0 123450.0 1433550.0 ;
      RECT  122550.0 1432200.0 123450.0 1433100.0 ;
      RECT  123000.0 1432650.0 139200.0 1433550.0 ;
      RECT  122550.0 1450050.0 123450.0 1450950.0 ;
      RECT  122550.0 1450500.0 123450.0 1451400.0 ;
      RECT  123000.0 1450050.0 139200.0 1450950.0 ;
      RECT  122550.0 1460250.0 123450.0 1461150.0 ;
      RECT  122550.0 1459800.0 123450.0 1460700.0 ;
      RECT  123000.0 1460250.0 139200.0 1461150.0 ;
      RECT  122550.0 1477650.0 123450.0 1478550.0 ;
      RECT  122550.0 1478100.0 123450.0 1479000.0 ;
      RECT  123000.0 1477650.0 139200.0 1478550.0 ;
      RECT  122550.0 1487850.0 123450.0 1488750.0 ;
      RECT  122550.0 1487400.0 123450.0 1488300.0 ;
      RECT  123000.0 1487850.0 139200.0 1488750.0 ;
      RECT  122550.0 1505250.0 123450.0 1506150.0 ;
      RECT  122550.0 1505700.0 123450.0 1506600.0 ;
      RECT  123000.0 1505250.0 139200.0 1506150.0 ;
      RECT  122550.0 1515450.0 123450.0 1516350.0 ;
      RECT  122550.0 1515000.0 123450.0 1515900.0 ;
      RECT  123000.0 1515450.0 139200.0 1516350.0 ;
      RECT  122550.0 1532850.0 123450.0 1533750.0 ;
      RECT  122550.0 1533300.0 123450.0 1534200.0 ;
      RECT  123000.0 1532850.0 139200.0 1533750.0 ;
      RECT  122550.0 1543050.0 123450.0 1543950.0 ;
      RECT  122550.0 1542600.0 123450.0 1543500.0 ;
      RECT  123000.0 1543050.0 139200.0 1543950.0 ;
      RECT  122550.0 1560450.0 123450.0 1561350.0 ;
      RECT  122550.0 1560900.0 123450.0 1561800.0 ;
      RECT  123000.0 1560450.0 139200.0 1561350.0 ;
      RECT  122550.0 1570650.0 123450.0 1571550.0 ;
      RECT  122550.0 1570200.0 123450.0 1571100.0 ;
      RECT  123000.0 1570650.0 139200.0 1571550.0 ;
      RECT  122550.0 1588050.0 123450.0 1588950.0 ;
      RECT  122550.0 1588500.0 123450.0 1589400.0 ;
      RECT  123000.0 1588050.0 139200.0 1588950.0 ;
      RECT  122550.0 1598250.0 123450.0 1599150.0 ;
      RECT  122550.0 1597800.0 123450.0 1598700.0 ;
      RECT  123000.0 1598250.0 139200.0 1599150.0 ;
      RECT  122550.0 1615650.0 123450.0 1616550.0 ;
      RECT  122550.0 1616100.0 123450.0 1617000.0 ;
      RECT  123000.0 1615650.0 139200.0 1616550.0 ;
      RECT  122550.0 1625850.0 123450.0 1626750.0 ;
      RECT  122550.0 1625400.0 123450.0 1626300.0 ;
      RECT  123000.0 1625850.0 139200.0 1626750.0 ;
      RECT  122550.0 1643250.0 123450.0 1644150.0 ;
      RECT  122550.0 1643700.0 123450.0 1644600.0 ;
      RECT  123000.0 1643250.0 139200.0 1644150.0 ;
      RECT  122550.0 1653450.0 123450.0 1654350.0 ;
      RECT  122550.0 1653000.0 123450.0 1653900.0 ;
      RECT  123000.0 1653450.0 139200.0 1654350.0 ;
      RECT  122550.0 1670850.0 123450.0 1671750.0 ;
      RECT  122550.0 1671300.0 123450.0 1672200.0 ;
      RECT  123000.0 1670850.0 139200.0 1671750.0 ;
      RECT  122550.0 1681050.0 123450.0 1681950.0 ;
      RECT  122550.0 1680600.0 123450.0 1681500.0 ;
      RECT  123000.0 1681050.0 139200.0 1681950.0 ;
      RECT  122550.0 1698450.0 123450.0 1699350.0 ;
      RECT  122550.0 1698900.0 123450.0 1699800.0 ;
      RECT  123000.0 1698450.0 139200.0 1699350.0 ;
      RECT  122550.0 1708650.0 123450.0 1709550.0 ;
      RECT  122550.0 1708200.0 123450.0 1709100.0 ;
      RECT  123000.0 1708650.0 139200.0 1709550.0 ;
      RECT  122550.0 1726050.0 123450.0 1726950.0 ;
      RECT  122550.0 1726500.0 123450.0 1727400.0 ;
      RECT  123000.0 1726050.0 139200.0 1726950.0 ;
      RECT  122550.0 1736250.0 123450.0 1737150.0 ;
      RECT  122550.0 1735800.0 123450.0 1736700.0 ;
      RECT  123000.0 1736250.0 139200.0 1737150.0 ;
      RECT  122550.0 1753650.0 123450.0 1754550.0 ;
      RECT  122550.0 1754100.0 123450.0 1755000.0 ;
      RECT  123000.0 1753650.0 139200.0 1754550.0 ;
      RECT  122550.0 1763850.0 123450.0 1764750.0 ;
      RECT  122550.0 1763400.0 123450.0 1764300.0 ;
      RECT  123000.0 1763850.0 139200.0 1764750.0 ;
      RECT  122550.0 1781250.0 123450.0 1782150.0 ;
      RECT  122550.0 1781700.0 123450.0 1782600.0 ;
      RECT  123000.0 1781250.0 139200.0 1782150.0 ;
      RECT  122550.0 1791450.0 123450.0 1792350.0 ;
      RECT  122550.0 1791000.0 123450.0 1791900.0 ;
      RECT  123000.0 1791450.0 139200.0 1792350.0 ;
      RECT  122550.0 1808850.0 123450.0 1809750.0 ;
      RECT  122550.0 1809300.0 123450.0 1810200.0 ;
      RECT  123000.0 1808850.0 139200.0 1809750.0 ;
      RECT  122550.0 1819050.0 123450.0 1819950.0 ;
      RECT  122550.0 1818600.0 123450.0 1819500.0 ;
      RECT  123000.0 1819050.0 139200.0 1819950.0 ;
      RECT  122550.0 1836450.0 123450.0 1837350.0 ;
      RECT  122550.0 1836900.0 123450.0 1837800.0 ;
      RECT  123000.0 1836450.0 139200.0 1837350.0 ;
      RECT  122550.0 1846650.0 123450.0 1847550.0 ;
      RECT  122550.0 1846200.0 123450.0 1847100.0 ;
      RECT  123000.0 1846650.0 139200.0 1847550.0 ;
      RECT  122550.0 1864050.0 123450.0 1864950.0 ;
      RECT  122550.0 1864500.0 123450.0 1865400.0 ;
      RECT  123000.0 1864050.0 139200.0 1864950.0 ;
      RECT  122550.0 1874250.0 123450.0 1875150.0 ;
      RECT  122550.0 1873800.0 123450.0 1874700.0 ;
      RECT  123000.0 1874250.0 139200.0 1875150.0 ;
      RECT  122550.0 1891650.0 123450.0 1892550.0 ;
      RECT  122550.0 1892100.0 123450.0 1893000.0 ;
      RECT  123000.0 1891650.0 139200.0 1892550.0 ;
      RECT  122550.0 1901850.0 123450.0 1902750.0 ;
      RECT  122550.0 1901400.0 123450.0 1902300.0 ;
      RECT  123000.0 1901850.0 139200.0 1902750.0 ;
      RECT  122550.0 1919250.0 123450.0 1920150.0 ;
      RECT  122550.0 1919700.0 123450.0 1920600.0 ;
      RECT  123000.0 1919250.0 139200.0 1920150.0 ;
      RECT  122550.0 1929450.0 123450.0 1930350.0 ;
      RECT  122550.0 1929000.0 123450.0 1929900.0 ;
      RECT  123000.0 1929450.0 139200.0 1930350.0 ;
      RECT  122550.0 1946850.0 123450.0 1947750.0 ;
      RECT  122550.0 1947300.0 123450.0 1948200.0 ;
      RECT  123000.0 1946850.0 139200.0 1947750.0 ;
      RECT  122550.0 1957050.0 123450.0 1957950.0 ;
      RECT  122550.0 1956600.0 123450.0 1957500.0 ;
      RECT  123000.0 1957050.0 139200.0 1957950.0 ;
      RECT  122550.0 1974450.0 123450.0 1975350.0 ;
      RECT  122550.0 1974900.0 123450.0 1975800.0 ;
      RECT  123000.0 1974450.0 139200.0 1975350.0 ;
      RECT  122550.0 1984650.0 123450.0 1985550.0 ;
      RECT  122550.0 1984200.0 123450.0 1985100.0 ;
      RECT  123000.0 1984650.0 139200.0 1985550.0 ;
      RECT  122550.0 2002050.0 123450.0 2002950.0 ;
      RECT  122550.0 2002500.0 123450.0 2003400.0 ;
      RECT  123000.0 2002050.0 139200.0 2002950.0 ;
      RECT  122550.0 2012250.0 123450.0 2013150.0 ;
      RECT  122550.0 2011800.0 123450.0 2012700.0 ;
      RECT  123000.0 2012250.0 139200.0 2013150.0 ;
      RECT  122550.0 2029650.0 123450.0 2030550.0 ;
      RECT  122550.0 2030100.0 123450.0 2031000.0 ;
      RECT  123000.0 2029650.0 139200.0 2030550.0 ;
      RECT  122550.0 2039850.0 123450.0 2040750.0 ;
      RECT  122550.0 2039400.0 123450.0 2040300.0 ;
      RECT  123000.0 2039850.0 139200.0 2040750.0 ;
      RECT  122550.0 2057250.0 123450.0 2058150.0 ;
      RECT  122550.0 2057700.0 123450.0 2058600.0 ;
      RECT  123000.0 2057250.0 139200.0 2058150.0 ;
      RECT  122550.0 2067450.0 123450.0 2068350.0 ;
      RECT  122550.0 2067000.0 123450.0 2067900.0 ;
      RECT  123000.0 2067450.0 139200.0 2068350.0 ;
      RECT  122550.0 2084850.0 123450.0 2085750.0 ;
      RECT  122550.0 2085300.0 123450.0 2086200.0 ;
      RECT  123000.0 2084850.0 139200.0 2085750.0 ;
      RECT  122550.0 2095050.0 123450.0 2095950.0 ;
      RECT  122550.0 2094600.0 123450.0 2095500.0 ;
      RECT  123000.0 2095050.0 139200.0 2095950.0 ;
      RECT  122550.0 2112450.0 123450.0 2113350.0 ;
      RECT  122550.0 2112900.0 123450.0 2113800.0 ;
      RECT  123000.0 2112450.0 139200.0 2113350.0 ;
      RECT  122550.0 2122650.0 123450.0 2123550.0 ;
      RECT  122550.0 2122200.0 123450.0 2123100.0 ;
      RECT  123000.0 2122650.0 139200.0 2123550.0 ;
      RECT  122550.0 2140050.0 123450.0 2140950.0 ;
      RECT  122550.0 2140500.0 123450.0 2141400.0 ;
      RECT  123000.0 2140050.0 139200.0 2140950.0 ;
      RECT  138150.0 386550.0 139050.0 387450.0 ;
      RECT  140550.0 386550.0 141450.0 387450.0 ;
      RECT  138150.0 387000.0 139050.0 389850.0 ;
      RECT  138600.0 386550.0 141000.0 387450.0 ;
      RECT  140550.0 382350.0 141450.0 387000.0 ;
      RECT  138000.0 389850.0 139200.0 391050.0 ;
      RECT  140400.0 381150.0 141600.0 382350.0 ;
      RECT  141600.0 386400.0 140400.0 387600.0 ;
      RECT  120450.0 385200.0 121650.0 386400.0 ;
      RECT  122400.0 382800.0 123600.0 384000.0 ;
      RECT  139200.0 383700.0 138000.0 384900.0 ;
      RECT  138150.0 399450.0 139050.0 398550.0 ;
      RECT  140550.0 399450.0 141450.0 398550.0 ;
      RECT  138150.0 399000.0 139050.0 396150.0 ;
      RECT  138600.0 399450.0 141000.0 398550.0 ;
      RECT  140550.0 403650.0 141450.0 399000.0 ;
      RECT  138000.0 396150.0 139200.0 394950.0 ;
      RECT  140400.0 404850.0 141600.0 403650.0 ;
      RECT  141600.0 399600.0 140400.0 398400.0 ;
      RECT  120450.0 399600.0 121650.0 400800.0 ;
      RECT  122400.0 402000.0 123600.0 403200.0 ;
      RECT  139200.0 401100.0 138000.0 402300.0 ;
      RECT  138150.0 414150.0 139050.0 415050.0 ;
      RECT  140550.0 414150.0 141450.0 415050.0 ;
      RECT  138150.0 414600.0 139050.0 417450.0 ;
      RECT  138600.0 414150.0 141000.0 415050.0 ;
      RECT  140550.0 409950.0 141450.0 414600.0 ;
      RECT  138000.0 417450.0 139200.0 418650.0 ;
      RECT  140400.0 408750.0 141600.0 409950.0 ;
      RECT  141600.0 414000.0 140400.0 415200.0 ;
      RECT  120450.0 412800.0 121650.0 414000.0 ;
      RECT  122400.0 410400.0 123600.0 411600.0 ;
      RECT  139200.0 411300.0 138000.0 412500.0 ;
      RECT  138150.0 427050.0 139050.0 426150.0 ;
      RECT  140550.0 427050.0 141450.0 426150.0 ;
      RECT  138150.0 426600.0 139050.0 423750.0 ;
      RECT  138600.0 427050.0 141000.0 426150.0 ;
      RECT  140550.0 431250.0 141450.0 426600.0 ;
      RECT  138000.0 423750.0 139200.0 422550.0 ;
      RECT  140400.0 432450.0 141600.0 431250.0 ;
      RECT  141600.0 427200.0 140400.0 426000.0 ;
      RECT  120450.0 427200.0 121650.0 428400.0 ;
      RECT  122400.0 429600.0 123600.0 430800.0 ;
      RECT  139200.0 428700.0 138000.0 429900.0 ;
      RECT  138150.0 441750.0 139050.0 442650.0 ;
      RECT  140550.0 441750.0 141450.0 442650.0 ;
      RECT  138150.0 442200.0 139050.0 445050.0 ;
      RECT  138600.0 441750.0 141000.0 442650.0 ;
      RECT  140550.0 437550.0 141450.0 442200.0 ;
      RECT  138000.0 445050.0 139200.0 446250.0 ;
      RECT  140400.0 436350.0 141600.0 437550.0 ;
      RECT  141600.0 441600.0 140400.0 442800.0 ;
      RECT  120450.0 440400.0 121650.0 441600.0 ;
      RECT  122400.0 438000.0 123600.0 439200.0 ;
      RECT  139200.0 438900.0 138000.0 440100.0 ;
      RECT  138150.0 454650.0 139050.0 453750.0 ;
      RECT  140550.0 454650.0 141450.0 453750.0 ;
      RECT  138150.0 454200.0 139050.0 451350.0 ;
      RECT  138600.0 454650.0 141000.0 453750.0 ;
      RECT  140550.0 458850.0 141450.0 454200.0 ;
      RECT  138000.0 451350.0 139200.0 450150.0 ;
      RECT  140400.0 460050.0 141600.0 458850.0 ;
      RECT  141600.0 454800.0 140400.0 453600.0 ;
      RECT  120450.0 454800.0 121650.0 456000.0 ;
      RECT  122400.0 457200.0 123600.0 458400.0 ;
      RECT  139200.0 456300.0 138000.0 457500.0 ;
      RECT  138150.0 469350.0 139050.0 470250.0 ;
      RECT  140550.0 469350.0 141450.0 470250.0 ;
      RECT  138150.0 469800.0 139050.0 472650.0 ;
      RECT  138600.0 469350.0 141000.0 470250.0 ;
      RECT  140550.0 465150.0 141450.0 469800.0 ;
      RECT  138000.0 472650.0 139200.0 473850.0 ;
      RECT  140400.0 463950.0 141600.0 465150.0 ;
      RECT  141600.0 469200.0 140400.0 470400.0 ;
      RECT  120450.0 468000.0 121650.0 469200.0 ;
      RECT  122400.0 465600.0 123600.0 466800.0 ;
      RECT  139200.0 466500.0 138000.0 467700.0 ;
      RECT  138150.0 482250.0 139050.0 481350.0 ;
      RECT  140550.0 482250.0 141450.0 481350.0 ;
      RECT  138150.0 481800.0 139050.0 478950.0 ;
      RECT  138600.0 482250.0 141000.0 481350.0 ;
      RECT  140550.0 486450.0 141450.0 481800.0 ;
      RECT  138000.0 478950.0 139200.0 477750.0 ;
      RECT  140400.0 487650.0 141600.0 486450.0 ;
      RECT  141600.0 482400.0 140400.0 481200.0 ;
      RECT  120450.0 482400.0 121650.0 483600.0 ;
      RECT  122400.0 484800.0 123600.0 486000.0 ;
      RECT  139200.0 483900.0 138000.0 485100.0 ;
      RECT  138150.0 496950.0 139050.0 497850.0 ;
      RECT  140550.0 496950.0 141450.0 497850.0 ;
      RECT  138150.0 497400.0 139050.0 500250.0 ;
      RECT  138600.0 496950.0 141000.0 497850.0 ;
      RECT  140550.0 492750.0 141450.0 497400.0 ;
      RECT  138000.0 500250.0 139200.0 501450.0 ;
      RECT  140400.0 491550.0 141600.0 492750.0 ;
      RECT  141600.0 496800.0 140400.0 498000.0 ;
      RECT  120450.0 495600.0 121650.0 496800.0 ;
      RECT  122400.0 493200.0 123600.0 494400.0 ;
      RECT  139200.0 494100.0 138000.0 495300.0 ;
      RECT  138150.0 509850.0 139050.0 508950.0 ;
      RECT  140550.0 509850.0 141450.0 508950.0 ;
      RECT  138150.0 509400.0 139050.0 506550.0 ;
      RECT  138600.0 509850.0 141000.0 508950.0 ;
      RECT  140550.0 514050.0 141450.0 509400.0 ;
      RECT  138000.0 506550.0 139200.0 505350.0 ;
      RECT  140400.0 515250.0 141600.0 514050.0 ;
      RECT  141600.0 510000.0 140400.0 508800.0 ;
      RECT  120450.0 510000.0 121650.0 511200.0 ;
      RECT  122400.0 512400.0 123600.0 513600.0 ;
      RECT  139200.0 511500.0 138000.0 512700.0 ;
      RECT  138150.0 524550.0 139050.0 525450.0 ;
      RECT  140550.0 524550.0 141450.0 525450.0 ;
      RECT  138150.0 525000.0 139050.0 527850.0 ;
      RECT  138600.0 524550.0 141000.0 525450.0 ;
      RECT  140550.0 520350.0 141450.0 525000.0 ;
      RECT  138000.0 527850.0 139200.0 529050.0 ;
      RECT  140400.0 519150.0 141600.0 520350.0 ;
      RECT  141600.0 524400.0 140400.0 525600.0 ;
      RECT  120450.0 523200.0 121650.0 524400.0 ;
      RECT  122400.0 520800.0 123600.0 522000.0 ;
      RECT  139200.0 521700.0 138000.0 522900.0 ;
      RECT  138150.0 537450.0 139050.0 536550.0 ;
      RECT  140550.0 537450.0 141450.0 536550.0 ;
      RECT  138150.0 537000.0 139050.0 534150.0 ;
      RECT  138600.0 537450.0 141000.0 536550.0 ;
      RECT  140550.0 541650.0 141450.0 537000.0 ;
      RECT  138000.0 534150.0 139200.0 532950.0 ;
      RECT  140400.0 542850.0 141600.0 541650.0 ;
      RECT  141600.0 537600.0 140400.0 536400.0 ;
      RECT  120450.0 537600.0 121650.0 538800.0 ;
      RECT  122400.0 540000.0 123600.0 541200.0 ;
      RECT  139200.0 539100.0 138000.0 540300.0 ;
      RECT  138150.0 552150.0 139050.0 553050.0 ;
      RECT  140550.0 552150.0 141450.0 553050.0 ;
      RECT  138150.0 552600.0 139050.0 555450.0 ;
      RECT  138600.0 552150.0 141000.0 553050.0 ;
      RECT  140550.0 547950.0 141450.0 552600.0 ;
      RECT  138000.0 555450.0 139200.0 556650.0 ;
      RECT  140400.0 546750.0 141600.0 547950.0 ;
      RECT  141600.0 552000.0 140400.0 553200.0 ;
      RECT  120450.0 550800.0 121650.0 552000.0 ;
      RECT  122400.0 548400.0 123600.0 549600.0 ;
      RECT  139200.0 549300.0 138000.0 550500.0 ;
      RECT  138150.0 565050.0 139050.0 564150.0 ;
      RECT  140550.0 565050.0 141450.0 564150.0 ;
      RECT  138150.0 564600.0 139050.0 561750.0 ;
      RECT  138600.0 565050.0 141000.0 564150.0 ;
      RECT  140550.0 569250.0 141450.0 564600.0 ;
      RECT  138000.0 561750.0 139200.0 560550.0 ;
      RECT  140400.0 570450.0 141600.0 569250.0 ;
      RECT  141600.0 565200.0 140400.0 564000.0 ;
      RECT  120450.0 565200.0 121650.0 566400.0 ;
      RECT  122400.0 567600.0 123600.0 568800.0 ;
      RECT  139200.0 566700.0 138000.0 567900.0 ;
      RECT  138150.0 579750.0 139050.0 580650.0 ;
      RECT  140550.0 579750.0 141450.0 580650.0 ;
      RECT  138150.0 580200.0 139050.0 583050.0 ;
      RECT  138600.0 579750.0 141000.0 580650.0 ;
      RECT  140550.0 575550.0 141450.0 580200.0 ;
      RECT  138000.0 583050.0 139200.0 584250.0 ;
      RECT  140400.0 574350.0 141600.0 575550.0 ;
      RECT  141600.0 579600.0 140400.0 580800.0 ;
      RECT  120450.0 578400.0 121650.0 579600.0 ;
      RECT  122400.0 576000.0 123600.0 577200.0 ;
      RECT  139200.0 576900.0 138000.0 578100.0 ;
      RECT  138150.0 592650.0 139050.0 591750.0 ;
      RECT  140550.0 592650.0 141450.0 591750.0 ;
      RECT  138150.0 592200.0 139050.0 589350.0 ;
      RECT  138600.0 592650.0 141000.0 591750.0 ;
      RECT  140550.0 596850.0 141450.0 592200.0 ;
      RECT  138000.0 589350.0 139200.0 588150.0 ;
      RECT  140400.0 598050.0 141600.0 596850.0 ;
      RECT  141600.0 592800.0 140400.0 591600.0 ;
      RECT  120450.0 592800.0 121650.0 594000.0 ;
      RECT  122400.0 595200.0 123600.0 596400.0 ;
      RECT  139200.0 594300.0 138000.0 595500.0 ;
      RECT  138150.0 607350.0 139050.0 608250.0 ;
      RECT  140550.0 607350.0 141450.0 608250.0 ;
      RECT  138150.0 607800.0 139050.0 610650.0 ;
      RECT  138600.0 607350.0 141000.0 608250.0 ;
      RECT  140550.0 603150.0 141450.0 607800.0 ;
      RECT  138000.0 610650.0 139200.0 611850.0 ;
      RECT  140400.0 601950.0 141600.0 603150.0 ;
      RECT  141600.0 607200.0 140400.0 608400.0 ;
      RECT  120450.0 606000.0 121650.0 607200.0 ;
      RECT  122400.0 603600.0 123600.0 604800.0 ;
      RECT  139200.0 604500.0 138000.0 605700.0 ;
      RECT  138150.0 620250.0 139050.0 619350.0 ;
      RECT  140550.0 620250.0 141450.0 619350.0 ;
      RECT  138150.0 619800.0 139050.0 616950.0 ;
      RECT  138600.0 620250.0 141000.0 619350.0 ;
      RECT  140550.0 624450.0 141450.0 619800.0 ;
      RECT  138000.0 616950.0 139200.0 615750.0 ;
      RECT  140400.0 625650.0 141600.0 624450.0 ;
      RECT  141600.0 620400.0 140400.0 619200.0 ;
      RECT  120450.0 620400.0 121650.0 621600.0 ;
      RECT  122400.0 622800.0 123600.0 624000.0 ;
      RECT  139200.0 621900.0 138000.0 623100.0 ;
      RECT  138150.0 634950.0 139050.0 635850.0 ;
      RECT  140550.0 634950.0 141450.0 635850.0 ;
      RECT  138150.0 635400.0 139050.0 638250.0 ;
      RECT  138600.0 634950.0 141000.0 635850.0 ;
      RECT  140550.0 630750.0 141450.0 635400.0 ;
      RECT  138000.0 638250.0 139200.0 639450.0 ;
      RECT  140400.0 629550.0 141600.0 630750.0 ;
      RECT  141600.0 634800.0 140400.0 636000.0 ;
      RECT  120450.0 633600.0 121650.0 634800.0 ;
      RECT  122400.0 631200.0 123600.0 632400.0 ;
      RECT  139200.0 632100.0 138000.0 633300.0 ;
      RECT  138150.0 647850.0 139050.0 646950.0 ;
      RECT  140550.0 647850.0 141450.0 646950.0 ;
      RECT  138150.0 647400.0 139050.0 644550.0 ;
      RECT  138600.0 647850.0 141000.0 646950.0 ;
      RECT  140550.0 652050.0 141450.0 647400.0 ;
      RECT  138000.0 644550.0 139200.0 643350.0 ;
      RECT  140400.0 653250.0 141600.0 652050.0 ;
      RECT  141600.0 648000.0 140400.0 646800.0 ;
      RECT  120450.0 648000.0 121650.0 649200.0 ;
      RECT  122400.0 650400.0 123600.0 651600.0 ;
      RECT  139200.0 649500.0 138000.0 650700.0 ;
      RECT  138150.0 662550.0 139050.0 663450.0 ;
      RECT  140550.0 662550.0 141450.0 663450.0 ;
      RECT  138150.0 663000.0 139050.0 665850.0 ;
      RECT  138600.0 662550.0 141000.0 663450.0 ;
      RECT  140550.0 658350.0 141450.0 663000.0 ;
      RECT  138000.0 665850.0 139200.0 667050.0 ;
      RECT  140400.0 657150.0 141600.0 658350.0 ;
      RECT  141600.0 662400.0 140400.0 663600.0 ;
      RECT  120450.0 661200.0 121650.0 662400.0 ;
      RECT  122400.0 658800.0 123600.0 660000.0 ;
      RECT  139200.0 659700.0 138000.0 660900.0 ;
      RECT  138150.0 675450.0 139050.0 674550.0 ;
      RECT  140550.0 675450.0 141450.0 674550.0 ;
      RECT  138150.0 675000.0 139050.0 672150.0 ;
      RECT  138600.0 675450.0 141000.0 674550.0 ;
      RECT  140550.0 679650.0 141450.0 675000.0 ;
      RECT  138000.0 672150.0 139200.0 670950.0 ;
      RECT  140400.0 680850.0 141600.0 679650.0 ;
      RECT  141600.0 675600.0 140400.0 674400.0 ;
      RECT  120450.0 675600.0 121650.0 676800.0 ;
      RECT  122400.0 678000.0 123600.0 679200.0 ;
      RECT  139200.0 677100.0 138000.0 678300.0 ;
      RECT  138150.0 690150.0 139050.0 691050.0 ;
      RECT  140550.0 690150.0 141450.0 691050.0 ;
      RECT  138150.0 690600.0 139050.0 693450.0 ;
      RECT  138600.0 690150.0 141000.0 691050.0 ;
      RECT  140550.0 685950.0 141450.0 690600.0 ;
      RECT  138000.0 693450.0 139200.0 694650.0 ;
      RECT  140400.0 684750.0 141600.0 685950.0 ;
      RECT  141600.0 690000.0 140400.0 691200.0 ;
      RECT  120450.0 688800.0 121650.0 690000.0 ;
      RECT  122400.0 686400.0 123600.0 687600.0 ;
      RECT  139200.0 687300.0 138000.0 688500.0 ;
      RECT  138150.0 703050.0 139050.0 702150.0 ;
      RECT  140550.0 703050.0 141450.0 702150.0 ;
      RECT  138150.0 702600.0 139050.0 699750.0 ;
      RECT  138600.0 703050.0 141000.0 702150.0 ;
      RECT  140550.0 707250.0 141450.0 702600.0 ;
      RECT  138000.0 699750.0 139200.0 698550.0 ;
      RECT  140400.0 708450.0 141600.0 707250.0 ;
      RECT  141600.0 703200.0 140400.0 702000.0 ;
      RECT  120450.0 703200.0 121650.0 704400.0 ;
      RECT  122400.0 705600.0 123600.0 706800.0 ;
      RECT  139200.0 704700.0 138000.0 705900.0 ;
      RECT  138150.0 717750.0 139050.0 718650.0 ;
      RECT  140550.0 717750.0 141450.0 718650.0 ;
      RECT  138150.0 718200.0 139050.0 721050.0 ;
      RECT  138600.0 717750.0 141000.0 718650.0 ;
      RECT  140550.0 713550.0 141450.0 718200.0 ;
      RECT  138000.0 721050.0 139200.0 722250.0 ;
      RECT  140400.0 712350.0 141600.0 713550.0 ;
      RECT  141600.0 717600.0 140400.0 718800.0 ;
      RECT  120450.0 716400.0 121650.0 717600.0 ;
      RECT  122400.0 714000.0 123600.0 715200.0 ;
      RECT  139200.0 714900.0 138000.0 716100.0 ;
      RECT  138150.0 730650.0 139050.0 729750.0 ;
      RECT  140550.0 730650.0 141450.0 729750.0 ;
      RECT  138150.0 730200.0 139050.0 727350.0 ;
      RECT  138600.0 730650.0 141000.0 729750.0 ;
      RECT  140550.0 734850.0 141450.0 730200.0 ;
      RECT  138000.0 727350.0 139200.0 726150.0 ;
      RECT  140400.0 736050.0 141600.0 734850.0 ;
      RECT  141600.0 730800.0 140400.0 729600.0 ;
      RECT  120450.0 730800.0 121650.0 732000.0 ;
      RECT  122400.0 733200.0 123600.0 734400.0 ;
      RECT  139200.0 732300.0 138000.0 733500.0 ;
      RECT  138150.0 745350.0 139050.0 746250.0 ;
      RECT  140550.0 745350.0 141450.0 746250.0 ;
      RECT  138150.0 745800.0 139050.0 748650.0 ;
      RECT  138600.0 745350.0 141000.0 746250.0 ;
      RECT  140550.0 741150.0 141450.0 745800.0 ;
      RECT  138000.0 748650.0 139200.0 749850.0 ;
      RECT  140400.0 739950.0 141600.0 741150.0 ;
      RECT  141600.0 745200.0 140400.0 746400.0 ;
      RECT  120450.0 744000.0 121650.0 745200.0 ;
      RECT  122400.0 741600.0 123600.0 742800.0 ;
      RECT  139200.0 742500.0 138000.0 743700.0 ;
      RECT  138150.0 758250.0 139050.0 757350.0 ;
      RECT  140550.0 758250.0 141450.0 757350.0 ;
      RECT  138150.0 757800.0 139050.0 754950.0 ;
      RECT  138600.0 758250.0 141000.0 757350.0 ;
      RECT  140550.0 762450.0 141450.0 757800.0 ;
      RECT  138000.0 754950.0 139200.0 753750.0 ;
      RECT  140400.0 763650.0 141600.0 762450.0 ;
      RECT  141600.0 758400.0 140400.0 757200.0 ;
      RECT  120450.0 758400.0 121650.0 759600.0 ;
      RECT  122400.0 760800.0 123600.0 762000.0 ;
      RECT  139200.0 759900.0 138000.0 761100.0 ;
      RECT  138150.0 772950.0 139050.0 773850.0 ;
      RECT  140550.0 772950.0 141450.0 773850.0 ;
      RECT  138150.0 773400.0 139050.0 776250.0 ;
      RECT  138600.0 772950.0 141000.0 773850.0 ;
      RECT  140550.0 768750.0 141450.0 773400.0 ;
      RECT  138000.0 776250.0 139200.0 777450.0 ;
      RECT  140400.0 767550.0 141600.0 768750.0 ;
      RECT  141600.0 772800.0 140400.0 774000.0 ;
      RECT  120450.0 771600.0 121650.0 772800.0 ;
      RECT  122400.0 769200.0 123600.0 770400.0 ;
      RECT  139200.0 770100.0 138000.0 771300.0 ;
      RECT  138150.0 785850.0 139050.0 784950.0 ;
      RECT  140550.0 785850.0 141450.0 784950.0 ;
      RECT  138150.0 785400.0 139050.0 782550.0 ;
      RECT  138600.0 785850.0 141000.0 784950.0 ;
      RECT  140550.0 790050.0 141450.0 785400.0 ;
      RECT  138000.0 782550.0 139200.0 781350.0 ;
      RECT  140400.0 791250.0 141600.0 790050.0 ;
      RECT  141600.0 786000.0 140400.0 784800.0 ;
      RECT  120450.0 786000.0 121650.0 787200.0 ;
      RECT  122400.0 788400.0 123600.0 789600.0 ;
      RECT  139200.0 787500.0 138000.0 788700.0 ;
      RECT  138150.0 800550.0 139050.0 801450.0 ;
      RECT  140550.0 800550.0 141450.0 801450.0 ;
      RECT  138150.0 801000.0 139050.0 803850.0 ;
      RECT  138600.0 800550.0 141000.0 801450.0 ;
      RECT  140550.0 796350.0 141450.0 801000.0 ;
      RECT  138000.0 803850.0 139200.0 805050.0 ;
      RECT  140400.0 795150.0 141600.0 796350.0 ;
      RECT  141600.0 800400.0 140400.0 801600.0 ;
      RECT  120450.0 799200.0 121650.0 800400.0 ;
      RECT  122400.0 796800.0 123600.0 798000.0 ;
      RECT  139200.0 797700.0 138000.0 798900.0 ;
      RECT  138150.0 813450.0 139050.0 812550.0 ;
      RECT  140550.0 813450.0 141450.0 812550.0 ;
      RECT  138150.0 813000.0 139050.0 810150.0 ;
      RECT  138600.0 813450.0 141000.0 812550.0 ;
      RECT  140550.0 817650.0 141450.0 813000.0 ;
      RECT  138000.0 810150.0 139200.0 808950.0 ;
      RECT  140400.0 818850.0 141600.0 817650.0 ;
      RECT  141600.0 813600.0 140400.0 812400.0 ;
      RECT  120450.0 813600.0 121650.0 814800.0 ;
      RECT  122400.0 816000.0 123600.0 817200.0 ;
      RECT  139200.0 815100.0 138000.0 816300.0 ;
      RECT  138150.0 828150.0 139050.0 829050.0 ;
      RECT  140550.0 828150.0 141450.0 829050.0 ;
      RECT  138150.0 828600.0 139050.0 831450.0 ;
      RECT  138600.0 828150.0 141000.0 829050.0 ;
      RECT  140550.0 823950.0 141450.0 828600.0 ;
      RECT  138000.0 831450.0 139200.0 832650.0 ;
      RECT  140400.0 822750.0 141600.0 823950.0 ;
      RECT  141600.0 828000.0 140400.0 829200.0 ;
      RECT  120450.0 826800.0 121650.0 828000.0 ;
      RECT  122400.0 824400.0 123600.0 825600.0 ;
      RECT  139200.0 825300.0 138000.0 826500.0 ;
      RECT  138150.0 841050.0 139050.0 840150.0 ;
      RECT  140550.0 841050.0 141450.0 840150.0 ;
      RECT  138150.0 840600.0 139050.0 837750.0 ;
      RECT  138600.0 841050.0 141000.0 840150.0 ;
      RECT  140550.0 845250.0 141450.0 840600.0 ;
      RECT  138000.0 837750.0 139200.0 836550.0 ;
      RECT  140400.0 846450.0 141600.0 845250.0 ;
      RECT  141600.0 841200.0 140400.0 840000.0 ;
      RECT  120450.0 841200.0 121650.0 842400.0 ;
      RECT  122400.0 843600.0 123600.0 844800.0 ;
      RECT  139200.0 842700.0 138000.0 843900.0 ;
      RECT  138150.0 855750.0 139050.0 856650.0 ;
      RECT  140550.0 855750.0 141450.0 856650.0 ;
      RECT  138150.0 856200.0 139050.0 859050.0 ;
      RECT  138600.0 855750.0 141000.0 856650.0 ;
      RECT  140550.0 851550.0 141450.0 856200.0 ;
      RECT  138000.0 859050.0 139200.0 860250.0 ;
      RECT  140400.0 850350.0 141600.0 851550.0 ;
      RECT  141600.0 855600.0 140400.0 856800.0 ;
      RECT  120450.0 854400.0 121650.0 855600.0 ;
      RECT  122400.0 852000.0 123600.0 853200.0 ;
      RECT  139200.0 852900.0 138000.0 854100.0 ;
      RECT  138150.0 868650.0 139050.0 867750.0 ;
      RECT  140550.0 868650.0 141450.0 867750.0 ;
      RECT  138150.0 868200.0 139050.0 865350.0 ;
      RECT  138600.0 868650.0 141000.0 867750.0 ;
      RECT  140550.0 872850.0 141450.0 868200.0 ;
      RECT  138000.0 865350.0 139200.0 864150.0 ;
      RECT  140400.0 874050.0 141600.0 872850.0 ;
      RECT  141600.0 868800.0 140400.0 867600.0 ;
      RECT  120450.0 868800.0 121650.0 870000.0 ;
      RECT  122400.0 871200.0 123600.0 872400.0 ;
      RECT  139200.0 870300.0 138000.0 871500.0 ;
      RECT  138150.0 883350.0 139050.0 884250.0 ;
      RECT  140550.0 883350.0 141450.0 884250.0 ;
      RECT  138150.0 883800.0 139050.0 886650.0 ;
      RECT  138600.0 883350.0 141000.0 884250.0 ;
      RECT  140550.0 879150.0 141450.0 883800.0 ;
      RECT  138000.0 886650.0 139200.0 887850.0 ;
      RECT  140400.0 877950.0 141600.0 879150.0 ;
      RECT  141600.0 883200.0 140400.0 884400.0 ;
      RECT  120450.0 882000.0 121650.0 883200.0 ;
      RECT  122400.0 879600.0 123600.0 880800.0 ;
      RECT  139200.0 880500.0 138000.0 881700.0 ;
      RECT  138150.0 896250.0 139050.0 895350.0 ;
      RECT  140550.0 896250.0 141450.0 895350.0 ;
      RECT  138150.0 895800.0 139050.0 892950.0 ;
      RECT  138600.0 896250.0 141000.0 895350.0 ;
      RECT  140550.0 900450.0 141450.0 895800.0 ;
      RECT  138000.0 892950.0 139200.0 891750.0 ;
      RECT  140400.0 901650.0 141600.0 900450.0 ;
      RECT  141600.0 896400.0 140400.0 895200.0 ;
      RECT  120450.0 896400.0 121650.0 897600.0 ;
      RECT  122400.0 898800.0 123600.0 900000.0 ;
      RECT  139200.0 897900.0 138000.0 899100.0 ;
      RECT  138150.0 910950.0 139050.0 911850.0 ;
      RECT  140550.0 910950.0 141450.0 911850.0 ;
      RECT  138150.0 911400.0 139050.0 914250.0 ;
      RECT  138600.0 910950.0 141000.0 911850.0 ;
      RECT  140550.0 906750.0 141450.0 911400.0 ;
      RECT  138000.0 914250.0 139200.0 915450.0 ;
      RECT  140400.0 905550.0 141600.0 906750.0 ;
      RECT  141600.0 910800.0 140400.0 912000.0 ;
      RECT  120450.0 909600.0 121650.0 910800.0 ;
      RECT  122400.0 907200.0 123600.0 908400.0 ;
      RECT  139200.0 908100.0 138000.0 909300.0 ;
      RECT  138150.0 923850.0 139050.0 922950.0 ;
      RECT  140550.0 923850.0 141450.0 922950.0 ;
      RECT  138150.0 923400.0 139050.0 920550.0 ;
      RECT  138600.0 923850.0 141000.0 922950.0 ;
      RECT  140550.0 928050.0 141450.0 923400.0 ;
      RECT  138000.0 920550.0 139200.0 919350.0 ;
      RECT  140400.0 929250.0 141600.0 928050.0 ;
      RECT  141600.0 924000.0 140400.0 922800.0 ;
      RECT  120450.0 924000.0 121650.0 925200.0 ;
      RECT  122400.0 926400.0 123600.0 927600.0 ;
      RECT  139200.0 925500.0 138000.0 926700.0 ;
      RECT  138150.0 938550.0 139050.0 939450.0 ;
      RECT  140550.0 938550.0 141450.0 939450.0 ;
      RECT  138150.0 939000.0 139050.0 941850.0 ;
      RECT  138600.0 938550.0 141000.0 939450.0 ;
      RECT  140550.0 934350.0 141450.0 939000.0 ;
      RECT  138000.0 941850.0 139200.0 943050.0 ;
      RECT  140400.0 933150.0 141600.0 934350.0 ;
      RECT  141600.0 938400.0 140400.0 939600.0 ;
      RECT  120450.0 937200.0 121650.0 938400.0 ;
      RECT  122400.0 934800.0 123600.0 936000.0 ;
      RECT  139200.0 935700.0 138000.0 936900.0 ;
      RECT  138150.0 951450.0 139050.0 950550.0 ;
      RECT  140550.0 951450.0 141450.0 950550.0 ;
      RECT  138150.0 951000.0 139050.0 948150.0 ;
      RECT  138600.0 951450.0 141000.0 950550.0 ;
      RECT  140550.0 955650.0 141450.0 951000.0 ;
      RECT  138000.0 948150.0 139200.0 946950.0 ;
      RECT  140400.0 956850.0 141600.0 955650.0 ;
      RECT  141600.0 951600.0 140400.0 950400.0 ;
      RECT  120450.0 951600.0 121650.0 952800.0 ;
      RECT  122400.0 954000.0 123600.0 955200.0 ;
      RECT  139200.0 953100.0 138000.0 954300.0 ;
      RECT  138150.0 966150.0 139050.0 967050.0 ;
      RECT  140550.0 966150.0 141450.0 967050.0 ;
      RECT  138150.0 966600.0 139050.0 969450.0 ;
      RECT  138600.0 966150.0 141000.0 967050.0 ;
      RECT  140550.0 961950.0 141450.0 966600.0 ;
      RECT  138000.0 969450.0 139200.0 970650.0 ;
      RECT  140400.0 960750.0 141600.0 961950.0 ;
      RECT  141600.0 966000.0 140400.0 967200.0 ;
      RECT  120450.0 964800.0 121650.0 966000.0 ;
      RECT  122400.0 962400.0 123600.0 963600.0 ;
      RECT  139200.0 963300.0 138000.0 964500.0 ;
      RECT  138150.0 979050.0 139050.0 978150.0 ;
      RECT  140550.0 979050.0 141450.0 978150.0 ;
      RECT  138150.0 978600.0 139050.0 975750.0 ;
      RECT  138600.0 979050.0 141000.0 978150.0 ;
      RECT  140550.0 983250.0 141450.0 978600.0 ;
      RECT  138000.0 975750.0 139200.0 974550.0 ;
      RECT  140400.0 984450.0 141600.0 983250.0 ;
      RECT  141600.0 979200.0 140400.0 978000.0 ;
      RECT  120450.0 979200.0 121650.0 980400.0 ;
      RECT  122400.0 981600.0 123600.0 982800.0 ;
      RECT  139200.0 980700.0 138000.0 981900.0 ;
      RECT  138150.0 993750.0 139050.0 994650.0 ;
      RECT  140550.0 993750.0 141450.0 994650.0 ;
      RECT  138150.0 994200.0 139050.0 997050.0 ;
      RECT  138600.0 993750.0 141000.0 994650.0 ;
      RECT  140550.0 989550.0 141450.0 994200.0 ;
      RECT  138000.0 997050.0 139200.0 998250.0 ;
      RECT  140400.0 988350.0 141600.0 989550.0 ;
      RECT  141600.0 993600.0 140400.0 994800.0 ;
      RECT  120450.0 992400.0 121650.0 993600.0 ;
      RECT  122400.0 990000.0 123600.0 991200.0 ;
      RECT  139200.0 990900.0 138000.0 992100.0 ;
      RECT  138150.0 1006650.0 139050.0 1005750.0 ;
      RECT  140550.0 1006650.0 141450.0 1005750.0 ;
      RECT  138150.0 1006200.0 139050.0 1003350.0 ;
      RECT  138600.0 1006650.0 141000.0 1005750.0 ;
      RECT  140550.0 1010850.0 141450.0 1006200.0 ;
      RECT  138000.0 1003350.0 139200.0 1002150.0 ;
      RECT  140400.0 1012050.0 141600.0 1010850.0 ;
      RECT  141600.0 1006800.0 140400.0 1005600.0 ;
      RECT  120450.0 1006800.0 121650.0 1008000.0 ;
      RECT  122400.0 1009200.0 123600.0 1010400.0 ;
      RECT  139200.0 1008300.0 138000.0 1009500.0 ;
      RECT  138150.0 1021350.0 139050.0 1022250.0 ;
      RECT  140550.0 1021350.0 141450.0 1022250.0 ;
      RECT  138150.0 1021800.0 139050.0 1024650.0 ;
      RECT  138600.0 1021350.0 141000.0 1022250.0 ;
      RECT  140550.0 1017150.0 141450.0 1021800.0 ;
      RECT  138000.0 1024650.0 139200.0 1025850.0 ;
      RECT  140400.0 1015950.0 141600.0 1017150.0 ;
      RECT  141600.0 1021200.0 140400.0 1022400.0 ;
      RECT  120450.0 1020000.0 121650.0 1021200.0 ;
      RECT  122400.0 1017600.0 123600.0 1018800.0 ;
      RECT  139200.0 1018500.0 138000.0 1019700.0 ;
      RECT  138150.0 1034250.0 139050.0 1033350.0 ;
      RECT  140550.0 1034250.0 141450.0 1033350.0 ;
      RECT  138150.0 1033800.0 139050.0 1030950.0 ;
      RECT  138600.0 1034250.0 141000.0 1033350.0 ;
      RECT  140550.0 1038450.0 141450.0 1033800.0 ;
      RECT  138000.0 1030950.0 139200.0 1029750.0 ;
      RECT  140400.0 1039650.0 141600.0 1038450.0 ;
      RECT  141600.0 1034400.0 140400.0 1033200.0 ;
      RECT  120450.0 1034400.0 121650.0 1035600.0 ;
      RECT  122400.0 1036800.0 123600.0 1038000.0 ;
      RECT  139200.0 1035900.0 138000.0 1037100.0 ;
      RECT  138150.0 1048950.0 139050.0 1049850.0 ;
      RECT  140550.0 1048950.0 141450.0 1049850.0 ;
      RECT  138150.0 1049400.0 139050.0 1052250.0 ;
      RECT  138600.0 1048950.0 141000.0 1049850.0 ;
      RECT  140550.0 1044750.0 141450.0 1049400.0 ;
      RECT  138000.0 1052250.0 139200.0 1053450.0 ;
      RECT  140400.0 1043550.0 141600.0 1044750.0 ;
      RECT  141600.0 1048800.0 140400.0 1050000.0 ;
      RECT  120450.0 1047600.0 121650.0 1048800.0 ;
      RECT  122400.0 1045200.0 123600.0 1046400.0 ;
      RECT  139200.0 1046100.0 138000.0 1047300.0 ;
      RECT  138150.0 1061850.0 139050.0 1060950.0 ;
      RECT  140550.0 1061850.0 141450.0 1060950.0 ;
      RECT  138150.0 1061400.0 139050.0 1058550.0 ;
      RECT  138600.0 1061850.0 141000.0 1060950.0 ;
      RECT  140550.0 1066050.0 141450.0 1061400.0 ;
      RECT  138000.0 1058550.0 139200.0 1057350.0 ;
      RECT  140400.0 1067250.0 141600.0 1066050.0 ;
      RECT  141600.0 1062000.0 140400.0 1060800.0 ;
      RECT  120450.0 1062000.0 121650.0 1063200.0 ;
      RECT  122400.0 1064400.0 123600.0 1065600.0 ;
      RECT  139200.0 1063500.0 138000.0 1064700.0 ;
      RECT  138150.0 1076550.0 139050.0 1077450.0 ;
      RECT  140550.0 1076550.0 141450.0 1077450.0 ;
      RECT  138150.0 1077000.0 139050.0 1079850.0 ;
      RECT  138600.0 1076550.0 141000.0 1077450.0 ;
      RECT  140550.0 1072350.0 141450.0 1077000.0 ;
      RECT  138000.0 1079850.0 139200.0 1081050.0 ;
      RECT  140400.0 1071150.0 141600.0 1072350.0 ;
      RECT  141600.0 1076400.0 140400.0 1077600.0 ;
      RECT  120450.0 1075200.0 121650.0 1076400.0 ;
      RECT  122400.0 1072800.0 123600.0 1074000.0 ;
      RECT  139200.0 1073700.0 138000.0 1074900.0 ;
      RECT  138150.0 1089450.0 139050.0 1088550.0 ;
      RECT  140550.0 1089450.0 141450.0 1088550.0 ;
      RECT  138150.0 1089000.0 139050.0 1086150.0 ;
      RECT  138600.0 1089450.0 141000.0 1088550.0 ;
      RECT  140550.0 1093650.0 141450.0 1089000.0 ;
      RECT  138000.0 1086150.0 139200.0 1084950.0 ;
      RECT  140400.0 1094850.0 141600.0 1093650.0 ;
      RECT  141600.0 1089600.0 140400.0 1088400.0 ;
      RECT  120450.0 1089600.0 121650.0 1090800.0 ;
      RECT  122400.0 1092000.0 123600.0 1093200.0 ;
      RECT  139200.0 1091100.0 138000.0 1092300.0 ;
      RECT  138150.0 1104150.0 139050.0 1105050.0 ;
      RECT  140550.0 1104150.0 141450.0 1105050.0 ;
      RECT  138150.0 1104600.0 139050.0 1107450.0 ;
      RECT  138600.0 1104150.0 141000.0 1105050.0 ;
      RECT  140550.0 1099950.0 141450.0 1104600.0 ;
      RECT  138000.0 1107450.0 139200.0 1108650.0 ;
      RECT  140400.0 1098750.0 141600.0 1099950.0 ;
      RECT  141600.0 1104000.0 140400.0 1105200.0 ;
      RECT  120450.0 1102800.0 121650.0 1104000.0 ;
      RECT  122400.0 1100400.0 123600.0 1101600.0 ;
      RECT  139200.0 1101300.0 138000.0 1102500.0 ;
      RECT  138150.0 1117050.0 139050.0 1116150.0 ;
      RECT  140550.0 1117050.0 141450.0 1116150.0 ;
      RECT  138150.0 1116600.0 139050.0 1113750.0 ;
      RECT  138600.0 1117050.0 141000.0 1116150.0 ;
      RECT  140550.0 1121250.0 141450.0 1116600.0 ;
      RECT  138000.0 1113750.0 139200.0 1112550.0 ;
      RECT  140400.0 1122450.0 141600.0 1121250.0 ;
      RECT  141600.0 1117200.0 140400.0 1116000.0 ;
      RECT  120450.0 1117200.0 121650.0 1118400.0 ;
      RECT  122400.0 1119600.0 123600.0 1120800.0 ;
      RECT  139200.0 1118700.0 138000.0 1119900.0 ;
      RECT  138150.0 1131750.0 139050.0 1132650.0 ;
      RECT  140550.0 1131750.0 141450.0 1132650.0 ;
      RECT  138150.0 1132200.0 139050.0 1135050.0 ;
      RECT  138600.0 1131750.0 141000.0 1132650.0 ;
      RECT  140550.0 1127550.0 141450.0 1132200.0 ;
      RECT  138000.0 1135050.0 139200.0 1136250.0 ;
      RECT  140400.0 1126350.0 141600.0 1127550.0 ;
      RECT  141600.0 1131600.0 140400.0 1132800.0 ;
      RECT  120450.0 1130400.0 121650.0 1131600.0 ;
      RECT  122400.0 1128000.0 123600.0 1129200.0 ;
      RECT  139200.0 1128900.0 138000.0 1130100.0 ;
      RECT  138150.0 1144650.0 139050.0 1143750.0 ;
      RECT  140550.0 1144650.0 141450.0 1143750.0 ;
      RECT  138150.0 1144200.0 139050.0 1141350.0 ;
      RECT  138600.0 1144650.0 141000.0 1143750.0 ;
      RECT  140550.0 1148850.0 141450.0 1144200.0 ;
      RECT  138000.0 1141350.0 139200.0 1140150.0 ;
      RECT  140400.0 1150050.0 141600.0 1148850.0 ;
      RECT  141600.0 1144800.0 140400.0 1143600.0 ;
      RECT  120450.0 1144800.0 121650.0 1146000.0 ;
      RECT  122400.0 1147200.0 123600.0 1148400.0 ;
      RECT  139200.0 1146300.0 138000.0 1147500.0 ;
      RECT  138150.0 1159350.0 139050.0 1160250.0 ;
      RECT  140550.0 1159350.0 141450.0 1160250.0 ;
      RECT  138150.0 1159800.0 139050.0 1162650.0 ;
      RECT  138600.0 1159350.0 141000.0 1160250.0 ;
      RECT  140550.0 1155150.0 141450.0 1159800.0 ;
      RECT  138000.0 1162650.0 139200.0 1163850.0 ;
      RECT  140400.0 1153950.0 141600.0 1155150.0 ;
      RECT  141600.0 1159200.0 140400.0 1160400.0 ;
      RECT  120450.0 1158000.0 121650.0 1159200.0 ;
      RECT  122400.0 1155600.0 123600.0 1156800.0 ;
      RECT  139200.0 1156500.0 138000.0 1157700.0 ;
      RECT  138150.0 1172250.0 139050.0 1171350.0 ;
      RECT  140550.0 1172250.0 141450.0 1171350.0 ;
      RECT  138150.0 1171800.0 139050.0 1168950.0 ;
      RECT  138600.0 1172250.0 141000.0 1171350.0 ;
      RECT  140550.0 1176450.0 141450.0 1171800.0 ;
      RECT  138000.0 1168950.0 139200.0 1167750.0 ;
      RECT  140400.0 1177650.0 141600.0 1176450.0 ;
      RECT  141600.0 1172400.0 140400.0 1171200.0 ;
      RECT  120450.0 1172400.0 121650.0 1173600.0 ;
      RECT  122400.0 1174800.0 123600.0 1176000.0 ;
      RECT  139200.0 1173900.0 138000.0 1175100.0 ;
      RECT  138150.0 1186950.0 139050.0 1187850.0 ;
      RECT  140550.0 1186950.0 141450.0 1187850.0 ;
      RECT  138150.0 1187400.0 139050.0 1190250.0 ;
      RECT  138600.0 1186950.0 141000.0 1187850.0 ;
      RECT  140550.0 1182750.0 141450.0 1187400.0 ;
      RECT  138000.0 1190250.0 139200.0 1191450.0 ;
      RECT  140400.0 1181550.0 141600.0 1182750.0 ;
      RECT  141600.0 1186800.0 140400.0 1188000.0 ;
      RECT  120450.0 1185600.0 121650.0 1186800.0 ;
      RECT  122400.0 1183200.0 123600.0 1184400.0 ;
      RECT  139200.0 1184100.0 138000.0 1185300.0 ;
      RECT  138150.0 1199850.0 139050.0 1198950.0 ;
      RECT  140550.0 1199850.0 141450.0 1198950.0 ;
      RECT  138150.0 1199400.0 139050.0 1196550.0 ;
      RECT  138600.0 1199850.0 141000.0 1198950.0 ;
      RECT  140550.0 1204050.0 141450.0 1199400.0 ;
      RECT  138000.0 1196550.0 139200.0 1195350.0 ;
      RECT  140400.0 1205250.0 141600.0 1204050.0 ;
      RECT  141600.0 1200000.0 140400.0 1198800.0 ;
      RECT  120450.0 1200000.0 121650.0 1201200.0 ;
      RECT  122400.0 1202400.0 123600.0 1203600.0 ;
      RECT  139200.0 1201500.0 138000.0 1202700.0 ;
      RECT  138150.0 1214550.0 139050.0 1215450.0 ;
      RECT  140550.0 1214550.0 141450.0 1215450.0 ;
      RECT  138150.0 1215000.0 139050.0 1217850.0 ;
      RECT  138600.0 1214550.0 141000.0 1215450.0 ;
      RECT  140550.0 1210350.0 141450.0 1215000.0 ;
      RECT  138000.0 1217850.0 139200.0 1219050.0 ;
      RECT  140400.0 1209150.0 141600.0 1210350.0 ;
      RECT  141600.0 1214400.0 140400.0 1215600.0 ;
      RECT  120450.0 1213200.0 121650.0 1214400.0 ;
      RECT  122400.0 1210800.0 123600.0 1212000.0 ;
      RECT  139200.0 1211700.0 138000.0 1212900.0 ;
      RECT  138150.0 1227450.0 139050.0 1226550.0 ;
      RECT  140550.0 1227450.0 141450.0 1226550.0 ;
      RECT  138150.0 1227000.0 139050.0 1224150.0 ;
      RECT  138600.0 1227450.0 141000.0 1226550.0 ;
      RECT  140550.0 1231650.0 141450.0 1227000.0 ;
      RECT  138000.0 1224150.0 139200.0 1222950.0 ;
      RECT  140400.0 1232850.0 141600.0 1231650.0 ;
      RECT  141600.0 1227600.0 140400.0 1226400.0 ;
      RECT  120450.0 1227600.0 121650.0 1228800.0 ;
      RECT  122400.0 1230000.0 123600.0 1231200.0 ;
      RECT  139200.0 1229100.0 138000.0 1230300.0 ;
      RECT  138150.0 1242150.0 139050.0 1243050.0 ;
      RECT  140550.0 1242150.0 141450.0 1243050.0 ;
      RECT  138150.0 1242600.0 139050.0 1245450.0 ;
      RECT  138600.0 1242150.0 141000.0 1243050.0 ;
      RECT  140550.0 1237950.0 141450.0 1242600.0 ;
      RECT  138000.0 1245450.0 139200.0 1246650.0 ;
      RECT  140400.0 1236750.0 141600.0 1237950.0 ;
      RECT  141600.0 1242000.0 140400.0 1243200.0 ;
      RECT  120450.0 1240800.0 121650.0 1242000.0 ;
      RECT  122400.0 1238400.0 123600.0 1239600.0 ;
      RECT  139200.0 1239300.0 138000.0 1240500.0 ;
      RECT  138150.0 1255050.0 139050.0 1254150.0 ;
      RECT  140550.0 1255050.0 141450.0 1254150.0 ;
      RECT  138150.0 1254600.0 139050.0 1251750.0 ;
      RECT  138600.0 1255050.0 141000.0 1254150.0 ;
      RECT  140550.0 1259250.0 141450.0 1254600.0 ;
      RECT  138000.0 1251750.0 139200.0 1250550.0 ;
      RECT  140400.0 1260450.0 141600.0 1259250.0 ;
      RECT  141600.0 1255200.0 140400.0 1254000.0 ;
      RECT  120450.0 1255200.0 121650.0 1256400.0 ;
      RECT  122400.0 1257600.0 123600.0 1258800.0 ;
      RECT  139200.0 1256700.0 138000.0 1257900.0 ;
      RECT  138150.0 1269750.0 139050.0 1270650.0 ;
      RECT  140550.0 1269750.0 141450.0 1270650.0 ;
      RECT  138150.0 1270200.0 139050.0 1273050.0 ;
      RECT  138600.0 1269750.0 141000.0 1270650.0 ;
      RECT  140550.0 1265550.0 141450.0 1270200.0 ;
      RECT  138000.0 1273050.0 139200.0 1274250.0 ;
      RECT  140400.0 1264350.0 141600.0 1265550.0 ;
      RECT  141600.0 1269600.0 140400.0 1270800.0 ;
      RECT  120450.0 1268400.0 121650.0 1269600.0 ;
      RECT  122400.0 1266000.0 123600.0 1267200.0 ;
      RECT  139200.0 1266900.0 138000.0 1268100.0 ;
      RECT  138150.0 1282650.0 139050.0 1281750.0 ;
      RECT  140550.0 1282650.0 141450.0 1281750.0 ;
      RECT  138150.0 1282200.0 139050.0 1279350.0 ;
      RECT  138600.0 1282650.0 141000.0 1281750.0 ;
      RECT  140550.0 1286850.0 141450.0 1282200.0 ;
      RECT  138000.0 1279350.0 139200.0 1278150.0 ;
      RECT  140400.0 1288050.0 141600.0 1286850.0 ;
      RECT  141600.0 1282800.0 140400.0 1281600.0 ;
      RECT  120450.0 1282800.0 121650.0 1284000.0 ;
      RECT  122400.0 1285200.0 123600.0 1286400.0 ;
      RECT  139200.0 1284300.0 138000.0 1285500.0 ;
      RECT  138150.0 1297350.0 139050.0 1298250.0 ;
      RECT  140550.0 1297350.0 141450.0 1298250.0 ;
      RECT  138150.0 1297800.0 139050.0 1300650.0 ;
      RECT  138600.0 1297350.0 141000.0 1298250.0 ;
      RECT  140550.0 1293150.0 141450.0 1297800.0 ;
      RECT  138000.0 1300650.0 139200.0 1301850.0 ;
      RECT  140400.0 1291950.0 141600.0 1293150.0 ;
      RECT  141600.0 1297200.0 140400.0 1298400.0 ;
      RECT  120450.0 1296000.0 121650.0 1297200.0 ;
      RECT  122400.0 1293600.0 123600.0 1294800.0 ;
      RECT  139200.0 1294500.0 138000.0 1295700.0 ;
      RECT  138150.0 1310250.0 139050.0 1309350.0 ;
      RECT  140550.0 1310250.0 141450.0 1309350.0 ;
      RECT  138150.0 1309800.0 139050.0 1306950.0 ;
      RECT  138600.0 1310250.0 141000.0 1309350.0 ;
      RECT  140550.0 1314450.0 141450.0 1309800.0 ;
      RECT  138000.0 1306950.0 139200.0 1305750.0 ;
      RECT  140400.0 1315650.0 141600.0 1314450.0 ;
      RECT  141600.0 1310400.0 140400.0 1309200.0 ;
      RECT  120450.0 1310400.0 121650.0 1311600.0 ;
      RECT  122400.0 1312800.0 123600.0 1314000.0 ;
      RECT  139200.0 1311900.0 138000.0 1313100.0 ;
      RECT  138150.0 1324950.0 139050.0 1325850.0 ;
      RECT  140550.0 1324950.0 141450.0 1325850.0 ;
      RECT  138150.0 1325400.0 139050.0 1328250.0 ;
      RECT  138600.0 1324950.0 141000.0 1325850.0 ;
      RECT  140550.0 1320750.0 141450.0 1325400.0 ;
      RECT  138000.0 1328250.0 139200.0 1329450.0 ;
      RECT  140400.0 1319550.0 141600.0 1320750.0 ;
      RECT  141600.0 1324800.0 140400.0 1326000.0 ;
      RECT  120450.0 1323600.0 121650.0 1324800.0 ;
      RECT  122400.0 1321200.0 123600.0 1322400.0 ;
      RECT  139200.0 1322100.0 138000.0 1323300.0 ;
      RECT  138150.0 1337850.0 139050.0 1336950.0 ;
      RECT  140550.0 1337850.0 141450.0 1336950.0 ;
      RECT  138150.0 1337400.0 139050.0 1334550.0 ;
      RECT  138600.0 1337850.0 141000.0 1336950.0 ;
      RECT  140550.0 1342050.0 141450.0 1337400.0 ;
      RECT  138000.0 1334550.0 139200.0 1333350.0 ;
      RECT  140400.0 1343250.0 141600.0 1342050.0 ;
      RECT  141600.0 1338000.0 140400.0 1336800.0 ;
      RECT  120450.0 1338000.0 121650.0 1339200.0 ;
      RECT  122400.0 1340400.0 123600.0 1341600.0 ;
      RECT  139200.0 1339500.0 138000.0 1340700.0 ;
      RECT  138150.0 1352550.0 139050.0 1353450.0 ;
      RECT  140550.0 1352550.0 141450.0 1353450.0 ;
      RECT  138150.0 1353000.0 139050.0 1355850.0 ;
      RECT  138600.0 1352550.0 141000.0 1353450.0 ;
      RECT  140550.0 1348350.0 141450.0 1353000.0 ;
      RECT  138000.0 1355850.0 139200.0 1357050.0 ;
      RECT  140400.0 1347150.0 141600.0 1348350.0 ;
      RECT  141600.0 1352400.0 140400.0 1353600.0 ;
      RECT  120450.0 1351200.0 121650.0 1352400.0 ;
      RECT  122400.0 1348800.0 123600.0 1350000.0 ;
      RECT  139200.0 1349700.0 138000.0 1350900.0 ;
      RECT  138150.0 1365450.0 139050.0 1364550.0 ;
      RECT  140550.0 1365450.0 141450.0 1364550.0 ;
      RECT  138150.0 1365000.0 139050.0 1362150.0 ;
      RECT  138600.0 1365450.0 141000.0 1364550.0 ;
      RECT  140550.0 1369650.0 141450.0 1365000.0 ;
      RECT  138000.0 1362150.0 139200.0 1360950.0 ;
      RECT  140400.0 1370850.0 141600.0 1369650.0 ;
      RECT  141600.0 1365600.0 140400.0 1364400.0 ;
      RECT  120450.0 1365600.0 121650.0 1366800.0 ;
      RECT  122400.0 1368000.0 123600.0 1369200.0 ;
      RECT  139200.0 1367100.0 138000.0 1368300.0 ;
      RECT  138150.0 1380150.0 139050.0 1381050.0 ;
      RECT  140550.0 1380150.0 141450.0 1381050.0 ;
      RECT  138150.0 1380600.0 139050.0 1383450.0 ;
      RECT  138600.0 1380150.0 141000.0 1381050.0 ;
      RECT  140550.0 1375950.0 141450.0 1380600.0 ;
      RECT  138000.0 1383450.0 139200.0 1384650.0 ;
      RECT  140400.0 1374750.0 141600.0 1375950.0 ;
      RECT  141600.0 1380000.0 140400.0 1381200.0 ;
      RECT  120450.0 1378800.0 121650.0 1380000.0 ;
      RECT  122400.0 1376400.0 123600.0 1377600.0 ;
      RECT  139200.0 1377300.0 138000.0 1378500.0 ;
      RECT  138150.0 1393050.0 139050.0 1392150.0 ;
      RECT  140550.0 1393050.0 141450.0 1392150.0 ;
      RECT  138150.0 1392600.0 139050.0 1389750.0 ;
      RECT  138600.0 1393050.0 141000.0 1392150.0 ;
      RECT  140550.0 1397250.0 141450.0 1392600.0 ;
      RECT  138000.0 1389750.0 139200.0 1388550.0 ;
      RECT  140400.0 1398450.0 141600.0 1397250.0 ;
      RECT  141600.0 1393200.0 140400.0 1392000.0 ;
      RECT  120450.0 1393200.0 121650.0 1394400.0 ;
      RECT  122400.0 1395600.0 123600.0 1396800.0 ;
      RECT  139200.0 1394700.0 138000.0 1395900.0 ;
      RECT  138150.0 1407750.0 139050.0 1408650.0 ;
      RECT  140550.0 1407750.0 141450.0 1408650.0 ;
      RECT  138150.0 1408200.0 139050.0 1411050.0 ;
      RECT  138600.0 1407750.0 141000.0 1408650.0 ;
      RECT  140550.0 1403550.0 141450.0 1408200.0 ;
      RECT  138000.0 1411050.0 139200.0 1412250.0 ;
      RECT  140400.0 1402350.0 141600.0 1403550.0 ;
      RECT  141600.0 1407600.0 140400.0 1408800.0 ;
      RECT  120450.0 1406400.0 121650.0 1407600.0 ;
      RECT  122400.0 1404000.0 123600.0 1405200.0 ;
      RECT  139200.0 1404900.0 138000.0 1406100.0 ;
      RECT  138150.0 1420650.0 139050.0 1419750.0 ;
      RECT  140550.0 1420650.0 141450.0 1419750.0 ;
      RECT  138150.0 1420200.0 139050.0 1417350.0 ;
      RECT  138600.0 1420650.0 141000.0 1419750.0 ;
      RECT  140550.0 1424850.0 141450.0 1420200.0 ;
      RECT  138000.0 1417350.0 139200.0 1416150.0 ;
      RECT  140400.0 1426050.0 141600.0 1424850.0 ;
      RECT  141600.0 1420800.0 140400.0 1419600.0 ;
      RECT  120450.0 1420800.0 121650.0 1422000.0 ;
      RECT  122400.0 1423200.0 123600.0 1424400.0 ;
      RECT  139200.0 1422300.0 138000.0 1423500.0 ;
      RECT  138150.0 1435350.0 139050.0 1436250.0 ;
      RECT  140550.0 1435350.0 141450.0 1436250.0 ;
      RECT  138150.0 1435800.0 139050.0 1438650.0 ;
      RECT  138600.0 1435350.0 141000.0 1436250.0 ;
      RECT  140550.0 1431150.0 141450.0 1435800.0 ;
      RECT  138000.0 1438650.0 139200.0 1439850.0 ;
      RECT  140400.0 1429950.0 141600.0 1431150.0 ;
      RECT  141600.0 1435200.0 140400.0 1436400.0 ;
      RECT  120450.0 1434000.0 121650.0 1435200.0 ;
      RECT  122400.0 1431600.0 123600.0 1432800.0 ;
      RECT  139200.0 1432500.0 138000.0 1433700.0 ;
      RECT  138150.0 1448250.0 139050.0 1447350.0 ;
      RECT  140550.0 1448250.0 141450.0 1447350.0 ;
      RECT  138150.0 1447800.0 139050.0 1444950.0 ;
      RECT  138600.0 1448250.0 141000.0 1447350.0 ;
      RECT  140550.0 1452450.0 141450.0 1447800.0 ;
      RECT  138000.0 1444950.0 139200.0 1443750.0 ;
      RECT  140400.0 1453650.0 141600.0 1452450.0 ;
      RECT  141600.0 1448400.0 140400.0 1447200.0 ;
      RECT  120450.0 1448400.0 121650.0 1449600.0 ;
      RECT  122400.0 1450800.0 123600.0 1452000.0 ;
      RECT  139200.0 1449900.0 138000.0 1451100.0 ;
      RECT  138150.0 1462950.0 139050.0 1463850.0 ;
      RECT  140550.0 1462950.0 141450.0 1463850.0 ;
      RECT  138150.0 1463400.0 139050.0 1466250.0 ;
      RECT  138600.0 1462950.0 141000.0 1463850.0 ;
      RECT  140550.0 1458750.0 141450.0 1463400.0 ;
      RECT  138000.0 1466250.0 139200.0 1467450.0 ;
      RECT  140400.0 1457550.0 141600.0 1458750.0 ;
      RECT  141600.0 1462800.0 140400.0 1464000.0 ;
      RECT  120450.0 1461600.0 121650.0 1462800.0 ;
      RECT  122400.0 1459200.0 123600.0 1460400.0 ;
      RECT  139200.0 1460100.0 138000.0 1461300.0 ;
      RECT  138150.0 1475850.0 139050.0 1474950.0 ;
      RECT  140550.0 1475850.0 141450.0 1474950.0 ;
      RECT  138150.0 1475400.0 139050.0 1472550.0 ;
      RECT  138600.0 1475850.0 141000.0 1474950.0 ;
      RECT  140550.0 1480050.0 141450.0 1475400.0 ;
      RECT  138000.0 1472550.0 139200.0 1471350.0 ;
      RECT  140400.0 1481250.0 141600.0 1480050.0 ;
      RECT  141600.0 1476000.0 140400.0 1474800.0 ;
      RECT  120450.0 1476000.0 121650.0 1477200.0 ;
      RECT  122400.0 1478400.0 123600.0 1479600.0 ;
      RECT  139200.0 1477500.0 138000.0 1478700.0 ;
      RECT  138150.0 1490550.0 139050.0 1491450.0 ;
      RECT  140550.0 1490550.0 141450.0 1491450.0 ;
      RECT  138150.0 1491000.0 139050.0 1493850.0 ;
      RECT  138600.0 1490550.0 141000.0 1491450.0 ;
      RECT  140550.0 1486350.0 141450.0 1491000.0 ;
      RECT  138000.0 1493850.0 139200.0 1495050.0 ;
      RECT  140400.0 1485150.0 141600.0 1486350.0 ;
      RECT  141600.0 1490400.0 140400.0 1491600.0 ;
      RECT  120450.0 1489200.0 121650.0 1490400.0 ;
      RECT  122400.0 1486800.0 123600.0 1488000.0 ;
      RECT  139200.0 1487700.0 138000.0 1488900.0 ;
      RECT  138150.0 1503450.0 139050.0 1502550.0 ;
      RECT  140550.0 1503450.0 141450.0 1502550.0 ;
      RECT  138150.0 1503000.0 139050.0 1500150.0 ;
      RECT  138600.0 1503450.0 141000.0 1502550.0 ;
      RECT  140550.0 1507650.0 141450.0 1503000.0 ;
      RECT  138000.0 1500150.0 139200.0 1498950.0 ;
      RECT  140400.0 1508850.0 141600.0 1507650.0 ;
      RECT  141600.0 1503600.0 140400.0 1502400.0 ;
      RECT  120450.0 1503600.0 121650.0 1504800.0 ;
      RECT  122400.0 1506000.0 123600.0 1507200.0 ;
      RECT  139200.0 1505100.0 138000.0 1506300.0 ;
      RECT  138150.0 1518150.0 139050.0 1519050.0 ;
      RECT  140550.0 1518150.0 141450.0 1519050.0 ;
      RECT  138150.0 1518600.0 139050.0 1521450.0 ;
      RECT  138600.0 1518150.0 141000.0 1519050.0 ;
      RECT  140550.0 1513950.0 141450.0 1518600.0 ;
      RECT  138000.0 1521450.0 139200.0 1522650.0 ;
      RECT  140400.0 1512750.0 141600.0 1513950.0 ;
      RECT  141600.0 1518000.0 140400.0 1519200.0 ;
      RECT  120450.0 1516800.0 121650.0 1518000.0 ;
      RECT  122400.0 1514400.0 123600.0 1515600.0 ;
      RECT  139200.0 1515300.0 138000.0 1516500.0 ;
      RECT  138150.0 1531050.0 139050.0 1530150.0 ;
      RECT  140550.0 1531050.0 141450.0 1530150.0 ;
      RECT  138150.0 1530600.0 139050.0 1527750.0 ;
      RECT  138600.0 1531050.0 141000.0 1530150.0 ;
      RECT  140550.0 1535250.0 141450.0 1530600.0 ;
      RECT  138000.0 1527750.0 139200.0 1526550.0 ;
      RECT  140400.0 1536450.0 141600.0 1535250.0 ;
      RECT  141600.0 1531200.0 140400.0 1530000.0 ;
      RECT  120450.0 1531200.0 121650.0 1532400.0 ;
      RECT  122400.0 1533600.0 123600.0 1534800.0 ;
      RECT  139200.0 1532700.0 138000.0 1533900.0 ;
      RECT  138150.0 1545750.0 139050.0 1546650.0 ;
      RECT  140550.0 1545750.0 141450.0 1546650.0 ;
      RECT  138150.0 1546200.0 139050.0 1549050.0 ;
      RECT  138600.0 1545750.0 141000.0 1546650.0 ;
      RECT  140550.0 1541550.0 141450.0 1546200.0 ;
      RECT  138000.0 1549050.0 139200.0 1550250.0 ;
      RECT  140400.0 1540350.0 141600.0 1541550.0 ;
      RECT  141600.0 1545600.0 140400.0 1546800.0 ;
      RECT  120450.0 1544400.0 121650.0 1545600.0 ;
      RECT  122400.0 1542000.0 123600.0 1543200.0 ;
      RECT  139200.0 1542900.0 138000.0 1544100.0 ;
      RECT  138150.0 1558650.0 139050.0 1557750.0 ;
      RECT  140550.0 1558650.0 141450.0 1557750.0 ;
      RECT  138150.0 1558200.0 139050.0 1555350.0 ;
      RECT  138600.0 1558650.0 141000.0 1557750.0 ;
      RECT  140550.0 1562850.0 141450.0 1558200.0 ;
      RECT  138000.0 1555350.0 139200.0 1554150.0 ;
      RECT  140400.0 1564050.0 141600.0 1562850.0 ;
      RECT  141600.0 1558800.0 140400.0 1557600.0 ;
      RECT  120450.0 1558800.0 121650.0 1560000.0 ;
      RECT  122400.0 1561200.0 123600.0 1562400.0 ;
      RECT  139200.0 1560300.0 138000.0 1561500.0 ;
      RECT  138150.0 1573350.0 139050.0 1574250.0 ;
      RECT  140550.0 1573350.0 141450.0 1574250.0 ;
      RECT  138150.0 1573800.0 139050.0 1576650.0 ;
      RECT  138600.0 1573350.0 141000.0 1574250.0 ;
      RECT  140550.0 1569150.0 141450.0 1573800.0 ;
      RECT  138000.0 1576650.0 139200.0 1577850.0 ;
      RECT  140400.0 1567950.0 141600.0 1569150.0 ;
      RECT  141600.0 1573200.0 140400.0 1574400.0 ;
      RECT  120450.0 1572000.0 121650.0 1573200.0 ;
      RECT  122400.0 1569600.0 123600.0 1570800.0 ;
      RECT  139200.0 1570500.0 138000.0 1571700.0 ;
      RECT  138150.0 1586250.0 139050.0 1585350.0 ;
      RECT  140550.0 1586250.0 141450.0 1585350.0 ;
      RECT  138150.0 1585800.0 139050.0 1582950.0 ;
      RECT  138600.0 1586250.0 141000.0 1585350.0 ;
      RECT  140550.0 1590450.0 141450.0 1585800.0 ;
      RECT  138000.0 1582950.0 139200.0 1581750.0 ;
      RECT  140400.0 1591650.0 141600.0 1590450.0 ;
      RECT  141600.0 1586400.0 140400.0 1585200.0 ;
      RECT  120450.0 1586400.0 121650.0 1587600.0 ;
      RECT  122400.0 1588800.0 123600.0 1590000.0 ;
      RECT  139200.0 1587900.0 138000.0 1589100.0 ;
      RECT  138150.0 1600950.0 139050.0 1601850.0 ;
      RECT  140550.0 1600950.0 141450.0 1601850.0 ;
      RECT  138150.0 1601400.0 139050.0 1604250.0 ;
      RECT  138600.0 1600950.0 141000.0 1601850.0 ;
      RECT  140550.0 1596750.0 141450.0 1601400.0 ;
      RECT  138000.0 1604250.0 139200.0 1605450.0 ;
      RECT  140400.0 1595550.0 141600.0 1596750.0 ;
      RECT  141600.0 1600800.0 140400.0 1602000.0 ;
      RECT  120450.0 1599600.0 121650.0 1600800.0 ;
      RECT  122400.0 1597200.0 123600.0 1598400.0 ;
      RECT  139200.0 1598100.0 138000.0 1599300.0 ;
      RECT  138150.0 1613850.0 139050.0 1612950.0 ;
      RECT  140550.0 1613850.0 141450.0 1612950.0 ;
      RECT  138150.0 1613400.0 139050.0 1610550.0 ;
      RECT  138600.0 1613850.0 141000.0 1612950.0 ;
      RECT  140550.0 1618050.0 141450.0 1613400.0 ;
      RECT  138000.0 1610550.0 139200.0 1609350.0 ;
      RECT  140400.0 1619250.0 141600.0 1618050.0 ;
      RECT  141600.0 1614000.0 140400.0 1612800.0 ;
      RECT  120450.0 1614000.0 121650.0 1615200.0 ;
      RECT  122400.0 1616400.0 123600.0 1617600.0 ;
      RECT  139200.0 1615500.0 138000.0 1616700.0 ;
      RECT  138150.0 1628550.0 139050.0 1629450.0 ;
      RECT  140550.0 1628550.0 141450.0 1629450.0 ;
      RECT  138150.0 1629000.0 139050.0 1631850.0 ;
      RECT  138600.0 1628550.0 141000.0 1629450.0 ;
      RECT  140550.0 1624350.0 141450.0 1629000.0 ;
      RECT  138000.0 1631850.0 139200.0 1633050.0 ;
      RECT  140400.0 1623150.0 141600.0 1624350.0 ;
      RECT  141600.0 1628400.0 140400.0 1629600.0 ;
      RECT  120450.0 1627200.0 121650.0 1628400.0 ;
      RECT  122400.0 1624800.0 123600.0 1626000.0 ;
      RECT  139200.0 1625700.0 138000.0 1626900.0 ;
      RECT  138150.0 1641450.0 139050.0 1640550.0 ;
      RECT  140550.0 1641450.0 141450.0 1640550.0 ;
      RECT  138150.0 1641000.0 139050.0 1638150.0 ;
      RECT  138600.0 1641450.0 141000.0 1640550.0 ;
      RECT  140550.0 1645650.0 141450.0 1641000.0 ;
      RECT  138000.0 1638150.0 139200.0 1636950.0 ;
      RECT  140400.0 1646850.0 141600.0 1645650.0 ;
      RECT  141600.0 1641600.0 140400.0 1640400.0 ;
      RECT  120450.0 1641600.0 121650.0 1642800.0 ;
      RECT  122400.0 1644000.0 123600.0 1645200.0 ;
      RECT  139200.0 1643100.0 138000.0 1644300.0 ;
      RECT  138150.0 1656150.0 139050.0 1657050.0 ;
      RECT  140550.0 1656150.0 141450.0 1657050.0 ;
      RECT  138150.0 1656600.0 139050.0 1659450.0 ;
      RECT  138600.0 1656150.0 141000.0 1657050.0 ;
      RECT  140550.0 1651950.0 141450.0 1656600.0 ;
      RECT  138000.0 1659450.0 139200.0 1660650.0 ;
      RECT  140400.0 1650750.0 141600.0 1651950.0 ;
      RECT  141600.0 1656000.0 140400.0 1657200.0 ;
      RECT  120450.0 1654800.0 121650.0 1656000.0 ;
      RECT  122400.0 1652400.0 123600.0 1653600.0 ;
      RECT  139200.0 1653300.0 138000.0 1654500.0 ;
      RECT  138150.0 1669050.0 139050.0 1668150.0 ;
      RECT  140550.0 1669050.0 141450.0 1668150.0 ;
      RECT  138150.0 1668600.0 139050.0 1665750.0 ;
      RECT  138600.0 1669050.0 141000.0 1668150.0 ;
      RECT  140550.0 1673250.0 141450.0 1668600.0 ;
      RECT  138000.0 1665750.0 139200.0 1664550.0 ;
      RECT  140400.0 1674450.0 141600.0 1673250.0 ;
      RECT  141600.0 1669200.0 140400.0 1668000.0 ;
      RECT  120450.0 1669200.0 121650.0 1670400.0 ;
      RECT  122400.0 1671600.0 123600.0 1672800.0 ;
      RECT  139200.0 1670700.0 138000.0 1671900.0 ;
      RECT  138150.0 1683750.0 139050.0 1684650.0 ;
      RECT  140550.0 1683750.0 141450.0 1684650.0 ;
      RECT  138150.0 1684200.0 139050.0 1687050.0 ;
      RECT  138600.0 1683750.0 141000.0 1684650.0 ;
      RECT  140550.0 1679550.0 141450.0 1684200.0 ;
      RECT  138000.0 1687050.0 139200.0 1688250.0 ;
      RECT  140400.0 1678350.0 141600.0 1679550.0 ;
      RECT  141600.0 1683600.0 140400.0 1684800.0 ;
      RECT  120450.0 1682400.0 121650.0 1683600.0 ;
      RECT  122400.0 1680000.0 123600.0 1681200.0 ;
      RECT  139200.0 1680900.0 138000.0 1682100.0 ;
      RECT  138150.0 1696650.0 139050.0 1695750.0 ;
      RECT  140550.0 1696650.0 141450.0 1695750.0 ;
      RECT  138150.0 1696200.0 139050.0 1693350.0 ;
      RECT  138600.0 1696650.0 141000.0 1695750.0 ;
      RECT  140550.0 1700850.0 141450.0 1696200.0 ;
      RECT  138000.0 1693350.0 139200.0 1692150.0 ;
      RECT  140400.0 1702050.0 141600.0 1700850.0 ;
      RECT  141600.0 1696800.0 140400.0 1695600.0 ;
      RECT  120450.0 1696800.0 121650.0 1698000.0 ;
      RECT  122400.0 1699200.0 123600.0 1700400.0 ;
      RECT  139200.0 1698300.0 138000.0 1699500.0 ;
      RECT  138150.0 1711350.0 139050.0 1712250.0 ;
      RECT  140550.0 1711350.0 141450.0 1712250.0 ;
      RECT  138150.0 1711800.0 139050.0 1714650.0 ;
      RECT  138600.0 1711350.0 141000.0 1712250.0 ;
      RECT  140550.0 1707150.0 141450.0 1711800.0 ;
      RECT  138000.0 1714650.0 139200.0 1715850.0 ;
      RECT  140400.0 1705950.0 141600.0 1707150.0 ;
      RECT  141600.0 1711200.0 140400.0 1712400.0 ;
      RECT  120450.0 1710000.0 121650.0 1711200.0 ;
      RECT  122400.0 1707600.0 123600.0 1708800.0 ;
      RECT  139200.0 1708500.0 138000.0 1709700.0 ;
      RECT  138150.0 1724250.0 139050.0 1723350.0 ;
      RECT  140550.0 1724250.0 141450.0 1723350.0 ;
      RECT  138150.0 1723800.0 139050.0 1720950.0 ;
      RECT  138600.0 1724250.0 141000.0 1723350.0 ;
      RECT  140550.0 1728450.0 141450.0 1723800.0 ;
      RECT  138000.0 1720950.0 139200.0 1719750.0 ;
      RECT  140400.0 1729650.0 141600.0 1728450.0 ;
      RECT  141600.0 1724400.0 140400.0 1723200.0 ;
      RECT  120450.0 1724400.0 121650.0 1725600.0 ;
      RECT  122400.0 1726800.0 123600.0 1728000.0 ;
      RECT  139200.0 1725900.0 138000.0 1727100.0 ;
      RECT  138150.0 1738950.0 139050.0 1739850.0 ;
      RECT  140550.0 1738950.0 141450.0 1739850.0 ;
      RECT  138150.0 1739400.0 139050.0 1742250.0 ;
      RECT  138600.0 1738950.0 141000.0 1739850.0 ;
      RECT  140550.0 1734750.0 141450.0 1739400.0 ;
      RECT  138000.0 1742250.0 139200.0 1743450.0 ;
      RECT  140400.0 1733550.0 141600.0 1734750.0 ;
      RECT  141600.0 1738800.0 140400.0 1740000.0 ;
      RECT  120450.0 1737600.0 121650.0 1738800.0 ;
      RECT  122400.0 1735200.0 123600.0 1736400.0 ;
      RECT  139200.0 1736100.0 138000.0 1737300.0 ;
      RECT  138150.0 1751850.0 139050.0 1750950.0 ;
      RECT  140550.0 1751850.0 141450.0 1750950.0 ;
      RECT  138150.0 1751400.0 139050.0 1748550.0 ;
      RECT  138600.0 1751850.0 141000.0 1750950.0 ;
      RECT  140550.0 1756050.0 141450.0 1751400.0 ;
      RECT  138000.0 1748550.0 139200.0 1747350.0 ;
      RECT  140400.0 1757250.0 141600.0 1756050.0 ;
      RECT  141600.0 1752000.0 140400.0 1750800.0 ;
      RECT  120450.0 1752000.0 121650.0 1753200.0 ;
      RECT  122400.0 1754400.0 123600.0 1755600.0 ;
      RECT  139200.0 1753500.0 138000.0 1754700.0 ;
      RECT  138150.0 1766550.0 139050.0 1767450.0 ;
      RECT  140550.0 1766550.0 141450.0 1767450.0 ;
      RECT  138150.0 1767000.0 139050.0 1769850.0 ;
      RECT  138600.0 1766550.0 141000.0 1767450.0 ;
      RECT  140550.0 1762350.0 141450.0 1767000.0 ;
      RECT  138000.0 1769850.0 139200.0 1771050.0 ;
      RECT  140400.0 1761150.0 141600.0 1762350.0 ;
      RECT  141600.0 1766400.0 140400.0 1767600.0 ;
      RECT  120450.0 1765200.0 121650.0 1766400.0 ;
      RECT  122400.0 1762800.0 123600.0 1764000.0 ;
      RECT  139200.0 1763700.0 138000.0 1764900.0 ;
      RECT  138150.0 1779450.0 139050.0 1778550.0 ;
      RECT  140550.0 1779450.0 141450.0 1778550.0 ;
      RECT  138150.0 1779000.0 139050.0 1776150.0 ;
      RECT  138600.0 1779450.0 141000.0 1778550.0 ;
      RECT  140550.0 1783650.0 141450.0 1779000.0 ;
      RECT  138000.0 1776150.0 139200.0 1774950.0 ;
      RECT  140400.0 1784850.0 141600.0 1783650.0 ;
      RECT  141600.0 1779600.0 140400.0 1778400.0 ;
      RECT  120450.0 1779600.0 121650.0 1780800.0 ;
      RECT  122400.0 1782000.0 123600.0 1783200.0 ;
      RECT  139200.0 1781100.0 138000.0 1782300.0 ;
      RECT  138150.0 1794150.0 139050.0 1795050.0 ;
      RECT  140550.0 1794150.0 141450.0 1795050.0 ;
      RECT  138150.0 1794600.0 139050.0 1797450.0 ;
      RECT  138600.0 1794150.0 141000.0 1795050.0 ;
      RECT  140550.0 1789950.0 141450.0 1794600.0 ;
      RECT  138000.0 1797450.0 139200.0 1798650.0 ;
      RECT  140400.0 1788750.0 141600.0 1789950.0 ;
      RECT  141600.0 1794000.0 140400.0 1795200.0 ;
      RECT  120450.0 1792800.0 121650.0 1794000.0 ;
      RECT  122400.0 1790400.0 123600.0 1791600.0 ;
      RECT  139200.0 1791300.0 138000.0 1792500.0 ;
      RECT  138150.0 1807050.0 139050.0 1806150.0 ;
      RECT  140550.0 1807050.0 141450.0 1806150.0 ;
      RECT  138150.0 1806600.0 139050.0 1803750.0 ;
      RECT  138600.0 1807050.0 141000.0 1806150.0 ;
      RECT  140550.0 1811250.0 141450.0 1806600.0 ;
      RECT  138000.0 1803750.0 139200.0 1802550.0 ;
      RECT  140400.0 1812450.0 141600.0 1811250.0 ;
      RECT  141600.0 1807200.0 140400.0 1806000.0 ;
      RECT  120450.0 1807200.0 121650.0 1808400.0 ;
      RECT  122400.0 1809600.0 123600.0 1810800.0 ;
      RECT  139200.0 1808700.0 138000.0 1809900.0 ;
      RECT  138150.0 1821750.0 139050.0 1822650.0 ;
      RECT  140550.0 1821750.0 141450.0 1822650.0 ;
      RECT  138150.0 1822200.0 139050.0 1825050.0 ;
      RECT  138600.0 1821750.0 141000.0 1822650.0 ;
      RECT  140550.0 1817550.0 141450.0 1822200.0 ;
      RECT  138000.0 1825050.0 139200.0 1826250.0 ;
      RECT  140400.0 1816350.0 141600.0 1817550.0 ;
      RECT  141600.0 1821600.0 140400.0 1822800.0 ;
      RECT  120450.0 1820400.0 121650.0 1821600.0 ;
      RECT  122400.0 1818000.0 123600.0 1819200.0 ;
      RECT  139200.0 1818900.0 138000.0 1820100.0 ;
      RECT  138150.0 1834650.0 139050.0 1833750.0 ;
      RECT  140550.0 1834650.0 141450.0 1833750.0 ;
      RECT  138150.0 1834200.0 139050.0 1831350.0 ;
      RECT  138600.0 1834650.0 141000.0 1833750.0 ;
      RECT  140550.0 1838850.0 141450.0 1834200.0 ;
      RECT  138000.0 1831350.0 139200.0 1830150.0 ;
      RECT  140400.0 1840050.0 141600.0 1838850.0 ;
      RECT  141600.0 1834800.0 140400.0 1833600.0 ;
      RECT  120450.0 1834800.0 121650.0 1836000.0 ;
      RECT  122400.0 1837200.0 123600.0 1838400.0 ;
      RECT  139200.0 1836300.0 138000.0 1837500.0 ;
      RECT  138150.0 1849350.0 139050.0 1850250.0 ;
      RECT  140550.0 1849350.0 141450.0 1850250.0 ;
      RECT  138150.0 1849800.0 139050.0 1852650.0 ;
      RECT  138600.0 1849350.0 141000.0 1850250.0 ;
      RECT  140550.0 1845150.0 141450.0 1849800.0 ;
      RECT  138000.0 1852650.0 139200.0 1853850.0 ;
      RECT  140400.0 1843950.0 141600.0 1845150.0 ;
      RECT  141600.0 1849200.0 140400.0 1850400.0 ;
      RECT  120450.0 1848000.0 121650.0 1849200.0 ;
      RECT  122400.0 1845600.0 123600.0 1846800.0 ;
      RECT  139200.0 1846500.0 138000.0 1847700.0 ;
      RECT  138150.0 1862250.0 139050.0 1861350.0 ;
      RECT  140550.0 1862250.0 141450.0 1861350.0 ;
      RECT  138150.0 1861800.0 139050.0 1858950.0 ;
      RECT  138600.0 1862250.0 141000.0 1861350.0 ;
      RECT  140550.0 1866450.0 141450.0 1861800.0 ;
      RECT  138000.0 1858950.0 139200.0 1857750.0 ;
      RECT  140400.0 1867650.0 141600.0 1866450.0 ;
      RECT  141600.0 1862400.0 140400.0 1861200.0 ;
      RECT  120450.0 1862400.0 121650.0 1863600.0 ;
      RECT  122400.0 1864800.0 123600.0 1866000.0 ;
      RECT  139200.0 1863900.0 138000.0 1865100.0 ;
      RECT  138150.0 1876950.0 139050.0 1877850.0 ;
      RECT  140550.0 1876950.0 141450.0 1877850.0 ;
      RECT  138150.0 1877400.0 139050.0 1880250.0 ;
      RECT  138600.0 1876950.0 141000.0 1877850.0 ;
      RECT  140550.0 1872750.0 141450.0 1877400.0 ;
      RECT  138000.0 1880250.0 139200.0 1881450.0 ;
      RECT  140400.0 1871550.0 141600.0 1872750.0 ;
      RECT  141600.0 1876800.0 140400.0 1878000.0 ;
      RECT  120450.0 1875600.0 121650.0 1876800.0 ;
      RECT  122400.0 1873200.0 123600.0 1874400.0 ;
      RECT  139200.0 1874100.0 138000.0 1875300.0 ;
      RECT  138150.0 1889850.0 139050.0 1888950.0 ;
      RECT  140550.0 1889850.0 141450.0 1888950.0 ;
      RECT  138150.0 1889400.0 139050.0 1886550.0 ;
      RECT  138600.0 1889850.0 141000.0 1888950.0 ;
      RECT  140550.0 1894050.0 141450.0 1889400.0 ;
      RECT  138000.0 1886550.0 139200.0 1885350.0 ;
      RECT  140400.0 1895250.0 141600.0 1894050.0 ;
      RECT  141600.0 1890000.0 140400.0 1888800.0 ;
      RECT  120450.0 1890000.0 121650.0 1891200.0 ;
      RECT  122400.0 1892400.0 123600.0 1893600.0 ;
      RECT  139200.0 1891500.0 138000.0 1892700.0 ;
      RECT  138150.0 1904550.0 139050.0 1905450.0 ;
      RECT  140550.0 1904550.0 141450.0 1905450.0 ;
      RECT  138150.0 1905000.0 139050.0 1907850.0 ;
      RECT  138600.0 1904550.0 141000.0 1905450.0 ;
      RECT  140550.0 1900350.0 141450.0 1905000.0 ;
      RECT  138000.0 1907850.0 139200.0 1909050.0 ;
      RECT  140400.0 1899150.0 141600.0 1900350.0 ;
      RECT  141600.0 1904400.0 140400.0 1905600.0 ;
      RECT  120450.0 1903200.0 121650.0 1904400.0 ;
      RECT  122400.0 1900800.0 123600.0 1902000.0 ;
      RECT  139200.0 1901700.0 138000.0 1902900.0 ;
      RECT  138150.0 1917450.0 139050.0 1916550.0 ;
      RECT  140550.0 1917450.0 141450.0 1916550.0 ;
      RECT  138150.0 1917000.0 139050.0 1914150.0 ;
      RECT  138600.0 1917450.0 141000.0 1916550.0 ;
      RECT  140550.0 1921650.0 141450.0 1917000.0 ;
      RECT  138000.0 1914150.0 139200.0 1912950.0 ;
      RECT  140400.0 1922850.0 141600.0 1921650.0 ;
      RECT  141600.0 1917600.0 140400.0 1916400.0 ;
      RECT  120450.0 1917600.0 121650.0 1918800.0 ;
      RECT  122400.0 1920000.0 123600.0 1921200.0 ;
      RECT  139200.0 1919100.0 138000.0 1920300.0 ;
      RECT  138150.0 1932150.0 139050.0 1933050.0 ;
      RECT  140550.0 1932150.0 141450.0 1933050.0 ;
      RECT  138150.0 1932600.0 139050.0 1935450.0 ;
      RECT  138600.0 1932150.0 141000.0 1933050.0 ;
      RECT  140550.0 1927950.0 141450.0 1932600.0 ;
      RECT  138000.0 1935450.0 139200.0 1936650.0 ;
      RECT  140400.0 1926750.0 141600.0 1927950.0 ;
      RECT  141600.0 1932000.0 140400.0 1933200.0 ;
      RECT  120450.0 1930800.0 121650.0 1932000.0 ;
      RECT  122400.0 1928400.0 123600.0 1929600.0 ;
      RECT  139200.0 1929300.0 138000.0 1930500.0 ;
      RECT  138150.0 1945050.0 139050.0 1944150.0 ;
      RECT  140550.0 1945050.0 141450.0 1944150.0 ;
      RECT  138150.0 1944600.0 139050.0 1941750.0 ;
      RECT  138600.0 1945050.0 141000.0 1944150.0 ;
      RECT  140550.0 1949250.0 141450.0 1944600.0 ;
      RECT  138000.0 1941750.0 139200.0 1940550.0 ;
      RECT  140400.0 1950450.0 141600.0 1949250.0 ;
      RECT  141600.0 1945200.0 140400.0 1944000.0 ;
      RECT  120450.0 1945200.0 121650.0 1946400.0 ;
      RECT  122400.0 1947600.0 123600.0 1948800.0 ;
      RECT  139200.0 1946700.0 138000.0 1947900.0 ;
      RECT  138150.0 1959750.0 139050.0 1960650.0 ;
      RECT  140550.0 1959750.0 141450.0 1960650.0 ;
      RECT  138150.0 1960200.0 139050.0 1963050.0 ;
      RECT  138600.0 1959750.0 141000.0 1960650.0 ;
      RECT  140550.0 1955550.0 141450.0 1960200.0 ;
      RECT  138000.0 1963050.0 139200.0 1964250.0 ;
      RECT  140400.0 1954350.0 141600.0 1955550.0 ;
      RECT  141600.0 1959600.0 140400.0 1960800.0 ;
      RECT  120450.0 1958400.0 121650.0 1959600.0 ;
      RECT  122400.0 1956000.0 123600.0 1957200.0 ;
      RECT  139200.0 1956900.0 138000.0 1958100.0 ;
      RECT  138150.0 1972650.0 139050.0 1971750.0 ;
      RECT  140550.0 1972650.0 141450.0 1971750.0 ;
      RECT  138150.0 1972200.0 139050.0 1969350.0 ;
      RECT  138600.0 1972650.0 141000.0 1971750.0 ;
      RECT  140550.0 1976850.0 141450.0 1972200.0 ;
      RECT  138000.0 1969350.0 139200.0 1968150.0 ;
      RECT  140400.0 1978050.0 141600.0 1976850.0 ;
      RECT  141600.0 1972800.0 140400.0 1971600.0 ;
      RECT  120450.0 1972800.0 121650.0 1974000.0 ;
      RECT  122400.0 1975200.0 123600.0 1976400.0 ;
      RECT  139200.0 1974300.0 138000.0 1975500.0 ;
      RECT  138150.0 1987350.0 139050.0 1988250.0 ;
      RECT  140550.0 1987350.0 141450.0 1988250.0 ;
      RECT  138150.0 1987800.0 139050.0 1990650.0 ;
      RECT  138600.0 1987350.0 141000.0 1988250.0 ;
      RECT  140550.0 1983150.0 141450.0 1987800.0 ;
      RECT  138000.0 1990650.0 139200.0 1991850.0 ;
      RECT  140400.0 1981950.0 141600.0 1983150.0 ;
      RECT  141600.0 1987200.0 140400.0 1988400.0 ;
      RECT  120450.0 1986000.0 121650.0 1987200.0 ;
      RECT  122400.0 1983600.0 123600.0 1984800.0 ;
      RECT  139200.0 1984500.0 138000.0 1985700.0 ;
      RECT  138150.0 2000250.0 139050.0 1999350.0 ;
      RECT  140550.0 2000250.0 141450.0 1999350.0 ;
      RECT  138150.0 1999800.0 139050.0 1996950.0 ;
      RECT  138600.0 2000250.0 141000.0 1999350.0 ;
      RECT  140550.0 2004450.0 141450.0 1999800.0 ;
      RECT  138000.0 1996950.0 139200.0 1995750.0 ;
      RECT  140400.0 2005650.0 141600.0 2004450.0 ;
      RECT  141600.0 2000400.0 140400.0 1999200.0 ;
      RECT  120450.0 2000400.0 121650.0 2001600.0 ;
      RECT  122400.0 2002800.0 123600.0 2004000.0 ;
      RECT  139200.0 2001900.0 138000.0 2003100.0 ;
      RECT  138150.0 2014950.0 139050.0 2015850.0 ;
      RECT  140550.0 2014950.0 141450.0 2015850.0 ;
      RECT  138150.0 2015400.0 139050.0 2018250.0 ;
      RECT  138600.0 2014950.0 141000.0 2015850.0 ;
      RECT  140550.0 2010750.0 141450.0 2015400.0 ;
      RECT  138000.0 2018250.0 139200.0 2019450.0 ;
      RECT  140400.0 2009550.0 141600.0 2010750.0 ;
      RECT  141600.0 2014800.0 140400.0 2016000.0 ;
      RECT  120450.0 2013600.0 121650.0 2014800.0 ;
      RECT  122400.0 2011200.0 123600.0 2012400.0 ;
      RECT  139200.0 2012100.0 138000.0 2013300.0 ;
      RECT  138150.0 2027850.0 139050.0 2026950.0 ;
      RECT  140550.0 2027850.0 141450.0 2026950.0 ;
      RECT  138150.0 2027400.0 139050.0 2024550.0 ;
      RECT  138600.0 2027850.0 141000.0 2026950.0 ;
      RECT  140550.0 2032050.0 141450.0 2027400.0 ;
      RECT  138000.0 2024550.0 139200.0 2023350.0 ;
      RECT  140400.0 2033250.0 141600.0 2032050.0 ;
      RECT  141600.0 2028000.0 140400.0 2026800.0 ;
      RECT  120450.0 2028000.0 121650.0 2029200.0 ;
      RECT  122400.0 2030400.0 123600.0 2031600.0 ;
      RECT  139200.0 2029500.0 138000.0 2030700.0 ;
      RECT  138150.0 2042550.0 139050.0 2043450.0 ;
      RECT  140550.0 2042550.0 141450.0 2043450.0 ;
      RECT  138150.0 2043000.0 139050.0 2045850.0 ;
      RECT  138600.0 2042550.0 141000.0 2043450.0 ;
      RECT  140550.0 2038350.0 141450.0 2043000.0 ;
      RECT  138000.0 2045850.0 139200.0 2047050.0 ;
      RECT  140400.0 2037150.0 141600.0 2038350.0 ;
      RECT  141600.0 2042400.0 140400.0 2043600.0 ;
      RECT  120450.0 2041200.0 121650.0 2042400.0 ;
      RECT  122400.0 2038800.0 123600.0 2040000.0 ;
      RECT  139200.0 2039700.0 138000.0 2040900.0 ;
      RECT  138150.0 2055450.0 139050.0 2054550.0 ;
      RECT  140550.0 2055450.0 141450.0 2054550.0 ;
      RECT  138150.0 2055000.0 139050.0 2052150.0 ;
      RECT  138600.0 2055450.0 141000.0 2054550.0 ;
      RECT  140550.0 2059650.0 141450.0 2055000.0 ;
      RECT  138000.0 2052150.0 139200.0 2050950.0 ;
      RECT  140400.0 2060850.0 141600.0 2059650.0 ;
      RECT  141600.0 2055600.0 140400.0 2054400.0 ;
      RECT  120450.0 2055600.0 121650.0 2056800.0 ;
      RECT  122400.0 2058000.0 123600.0 2059200.0 ;
      RECT  139200.0 2057100.0 138000.0 2058300.0 ;
      RECT  138150.0 2070150.0 139050.0 2071050.0 ;
      RECT  140550.0 2070150.0 141450.0 2071050.0 ;
      RECT  138150.0 2070600.0 139050.0 2073450.0 ;
      RECT  138600.0 2070150.0 141000.0 2071050.0 ;
      RECT  140550.0 2065950.0 141450.0 2070600.0 ;
      RECT  138000.0 2073450.0 139200.0 2074650.0 ;
      RECT  140400.0 2064750.0 141600.0 2065950.0 ;
      RECT  141600.0 2070000.0 140400.0 2071200.0 ;
      RECT  120450.0 2068800.0 121650.0 2070000.0 ;
      RECT  122400.0 2066400.0 123600.0 2067600.0 ;
      RECT  139200.0 2067300.0 138000.0 2068500.0 ;
      RECT  138150.0 2083050.0 139050.0 2082150.0 ;
      RECT  140550.0 2083050.0 141450.0 2082150.0 ;
      RECT  138150.0 2082600.0 139050.0 2079750.0 ;
      RECT  138600.0 2083050.0 141000.0 2082150.0 ;
      RECT  140550.0 2087250.0 141450.0 2082600.0 ;
      RECT  138000.0 2079750.0 139200.0 2078550.0 ;
      RECT  140400.0 2088450.0 141600.0 2087250.0 ;
      RECT  141600.0 2083200.0 140400.0 2082000.0 ;
      RECT  120450.0 2083200.0 121650.0 2084400.0 ;
      RECT  122400.0 2085600.0 123600.0 2086800.0 ;
      RECT  139200.0 2084700.0 138000.0 2085900.0 ;
      RECT  138150.0 2097750.0 139050.0 2098650.0 ;
      RECT  140550.0 2097750.0 141450.0 2098650.0 ;
      RECT  138150.0 2098200.0 139050.0 2101050.0 ;
      RECT  138600.0 2097750.0 141000.0 2098650.0 ;
      RECT  140550.0 2093550.0 141450.0 2098200.0 ;
      RECT  138000.0 2101050.0 139200.0 2102250.0 ;
      RECT  140400.0 2092350.0 141600.0 2093550.0 ;
      RECT  141600.0 2097600.0 140400.0 2098800.0 ;
      RECT  120450.0 2096400.0 121650.0 2097600.0 ;
      RECT  122400.0 2094000.0 123600.0 2095200.0 ;
      RECT  139200.0 2094900.0 138000.0 2096100.0 ;
      RECT  138150.0 2110650.0 139050.0 2109750.0 ;
      RECT  140550.0 2110650.0 141450.0 2109750.0 ;
      RECT  138150.0 2110200.0 139050.0 2107350.0 ;
      RECT  138600.0 2110650.0 141000.0 2109750.0 ;
      RECT  140550.0 2114850.0 141450.0 2110200.0 ;
      RECT  138000.0 2107350.0 139200.0 2106150.0 ;
      RECT  140400.0 2116050.0 141600.0 2114850.0 ;
      RECT  141600.0 2110800.0 140400.0 2109600.0 ;
      RECT  120450.0 2110800.0 121650.0 2112000.0 ;
      RECT  122400.0 2113200.0 123600.0 2114400.0 ;
      RECT  139200.0 2112300.0 138000.0 2113500.0 ;
      RECT  138150.0 2125350.0 139050.0 2126250.0 ;
      RECT  140550.0 2125350.0 141450.0 2126250.0 ;
      RECT  138150.0 2125800.0 139050.0 2128650.0 ;
      RECT  138600.0 2125350.0 141000.0 2126250.0 ;
      RECT  140550.0 2121150.0 141450.0 2125800.0 ;
      RECT  138000.0 2128650.0 139200.0 2129850.0 ;
      RECT  140400.0 2119950.0 141600.0 2121150.0 ;
      RECT  141600.0 2125200.0 140400.0 2126400.0 ;
      RECT  120450.0 2124000.0 121650.0 2125200.0 ;
      RECT  122400.0 2121600.0 123600.0 2122800.0 ;
      RECT  139200.0 2122500.0 138000.0 2123700.0 ;
      RECT  138150.0 2138250.0 139050.0 2137350.0 ;
      RECT  140550.0 2138250.0 141450.0 2137350.0 ;
      RECT  138150.0 2137800.0 139050.0 2134950.0 ;
      RECT  138600.0 2138250.0 141000.0 2137350.0 ;
      RECT  140550.0 2142450.0 141450.0 2137800.0 ;
      RECT  138000.0 2134950.0 139200.0 2133750.0 ;
      RECT  140400.0 2143650.0 141600.0 2142450.0 ;
      RECT  141600.0 2138400.0 140400.0 2137200.0 ;
      RECT  120450.0 2138400.0 121650.0 2139600.0 ;
      RECT  122400.0 2140800.0 123600.0 2142000.0 ;
      RECT  139200.0 2139900.0 138000.0 2141100.0 ;
      RECT  120600.0 379200.0 121500.0 2145600.0 ;
      RECT  59100.0 153000.0 119100.0 142800.0 ;
      RECT  59100.0 132600.0 119100.0 142800.0 ;
      RECT  59100.0 132600.0 119100.0 122400.0 ;
      RECT  59100.0 112200.0 119100.0 122400.0 ;
      RECT  59100.0 112200.0 119100.0 102000.0 ;
      RECT  59100.0 91800.0 119100.0 102000.0 ;
      RECT  59100.0 91800.0 119100.0 81600.0 ;
      RECT  59100.0 71400.0 119100.0 81600.0 ;
      RECT  59100.0 71400.0 119100.0 61200.0 ;
      RECT  116700.0 148500.0 117900.0 145800.0 ;
      RECT  114600.0 151200.0 119100.0 150000.0 ;
      RECT  116700.0 139800.0 117900.0 137100.0 ;
      RECT  114600.0 135600.0 119100.0 134400.0 ;
      RECT  116700.0 128100.0 117900.0 125400.0 ;
      RECT  114600.0 130800.0 119100.0 129600.0 ;
      RECT  116700.0 119400.0 117900.0 116700.0 ;
      RECT  114600.0 115200.0 119100.0 114000.0 ;
      RECT  116700.0 107700.0 117900.0 105000.0 ;
      RECT  114600.0 110400.0 119100.0 109200.0 ;
      RECT  116700.0 99000.0 117900.0 96300.0 ;
      RECT  114600.0 94800.0 119100.0 93600.0 ;
      RECT  116700.0 87300.0 117900.0 84600.0 ;
      RECT  114600.0 90000.0 119100.0 88800.0 ;
      RECT  116700.0 78600.0 117900.0 75900.0 ;
      RECT  114600.0 74400.0 119100.0 73200.0 ;
      RECT  116700.0 66900.0 117900.0 64200.0 ;
      RECT  114600.0 69600.0 119100.0 68400.0 ;
      RECT  59100.0 143400.0 119100.0 142200.0 ;
      RECT  59100.0 123000.0 119100.0 121800.0 ;
      RECT  59100.0 102600.0 119100.0 101400.0 ;
      RECT  59100.0 82200.0 119100.0 81000.0 ;
      RECT  59100.0 61800.0 119100.0 60600.0 ;
      RECT  222450.0 144900.0 223650.0 146100.0 ;
      RECT  263250.0 144900.0 264450.0 146100.0 ;
      RECT  304050.0 144900.0 305250.0 146100.0 ;
      RECT  344850.0 144900.0 346050.0 146100.0 ;
      RECT  385650.0 144900.0 386850.0 146100.0 ;
      RECT  426450.0 144900.0 427650.0 146100.0 ;
      RECT  467250.0 144900.0 468450.0 146100.0 ;
      RECT  508050.0 144900.0 509250.0 146100.0 ;
      RECT  548850.0 144900.0 550050.0 146100.0 ;
      RECT  589650.0 144900.0 590850.0 146100.0 ;
      RECT  630450.0 144900.0 631650.0 146100.0 ;
      RECT  671250.0 144900.0 672450.0 146100.0 ;
      RECT  712050.0 144900.0 713250.0 146100.0 ;
      RECT  752850.0 144900.0 754050.0 146100.0 ;
      RECT  793650.0 144900.0 794850.0 146100.0 ;
      RECT  834450.0 144900.0 835650.0 146100.0 ;
      RECT  875250.0 144900.0 876450.0 146100.0 ;
      RECT  916050.0 144900.0 917250.0 146100.0 ;
      RECT  956850.0 144900.0 958050.0 146100.0 ;
      RECT  997650.0 144900.0 998850.0 146100.0 ;
      RECT  1038450.0 144900.0 1039650.0 146100.0 ;
      RECT  1079250.0 144900.0 1080450.0 146100.0 ;
      RECT  1120050.0 144900.0 1121250.0 146100.0 ;
      RECT  1160850.0 144900.0 1162050.0 146100.0 ;
      RECT  1201650.0 144900.0 1202850.0 146100.0 ;
      RECT  1242450.0 144900.0 1243650.0 146100.0 ;
      RECT  1283250.0 144900.0 1284450.0 146100.0 ;
      RECT  1324050.0 144900.0 1325250.0 146100.0 ;
      RECT  1364850.0 144900.0 1366050.0 146100.0 ;
      RECT  1405650.0 144900.0 1406850.0 146100.0 ;
      RECT  1446450.0 144900.0 1447650.0 146100.0 ;
      RECT  1487250.0 144900.0 1488450.0 146100.0 ;
      RECT  226200.0 900.0 227400.0 2100.0 ;
      RECT  267000.0 900.0 268200.0 2100.0 ;
      RECT  307800.0 900.0 309000.0 2100.0 ;
      RECT  348600.0 900.0 349800.0 2100.0 ;
      RECT  389400.0 900.0 390600.0 2100.0 ;
      RECT  430200.0 900.0 431400.0 2100.0 ;
      RECT  471000.0 900.0 472200.0 2100.0 ;
      RECT  511800.0 900.0 513000.0 2100.0 ;
      RECT  552600.0 900.0 553800.0 2100.0 ;
      RECT  593400.0 900.0 594600.0 2100.0 ;
      RECT  634200.0 900.0 635400.0 2100.0 ;
      RECT  675000.0 900.0 676200.0 2100.0 ;
      RECT  715800.0 900.0 717000.0 2100.0 ;
      RECT  756600.0 900.0 757800.0 2100.0 ;
      RECT  797400.0 900.0 798600.0 2100.0 ;
      RECT  838200.0 900.0 839400.0 2100.0 ;
      RECT  879000.0 900.0 880200.0 2100.0 ;
      RECT  919800.0 900.0 921000.0 2100.0 ;
      RECT  960600.0 900.0 961800.0 2100.0 ;
      RECT  1001400.0 900.0 1002600.0 2100.0 ;
      RECT  1042200.0 900.0 1043400.0 2100.0 ;
      RECT  1083000.0 900.0 1084200.0 2100.0 ;
      RECT  1123800.0 900.0 1125000.0 2100.0 ;
      RECT  1164600.0 900.0 1165800.0 2100.0 ;
      RECT  1205400.0 900.0 1206600.0 2100.0 ;
      RECT  1246200.0 900.0 1247400.0 2100.0 ;
      RECT  1287000.0 900.0 1288200.0 2100.0 ;
      RECT  1327800.0 900.0 1329000.0 2100.0 ;
      RECT  1368600.0 900.0 1369800.0 2100.0 ;
      RECT  1409400.0 900.0 1410600.0 2100.0 ;
      RECT  1450200.0 900.0 1451400.0 2100.0 ;
      RECT  1491000.0 900.0 1492200.0 2100.0 ;
      RECT  193950.0 379800.0 195150.0 378600.0 ;
      RECT  193950.0 407400.0 195150.0 406200.0 ;
      RECT  193950.0 435000.0 195150.0 433800.0 ;
      RECT  193950.0 462600.0 195150.0 461400.0 ;
      RECT  193950.0 490200.0 195150.0 489000.0 ;
      RECT  193950.0 517800.0 195150.0 516600.0 ;
      RECT  193950.0 545400.0 195150.0 544200.0 ;
      RECT  193950.0 573000.0 195150.0 571800.0 ;
      RECT  193950.0 600600.0 195150.0 599400.0 ;
      RECT  193950.0 628200.0 195150.0 627000.0 ;
      RECT  193950.0 655800.0 195150.0 654600.0 ;
      RECT  193950.0 683400.0 195150.0 682200.0 ;
      RECT  193950.0 711000.0 195150.0 709800.0 ;
      RECT  193950.0 738600.0 195150.0 737400.0 ;
      RECT  193950.0 766200.0 195150.0 765000.0 ;
      RECT  193950.0 793800.0 195150.0 792600.0 ;
      RECT  193950.0 821400.0 195150.0 820200.0 ;
      RECT  193950.0 849000.0 195150.0 847800.0 ;
      RECT  193950.0 876600.0 195150.0 875400.0 ;
      RECT  193950.0 904200.0 195150.0 903000.0 ;
      RECT  193950.0 931800.0 195150.0 930600.0 ;
      RECT  193950.0 959400.0 195150.0 958200.0 ;
      RECT  193950.0 987000.0 195150.0 985800.0 ;
      RECT  193950.0 1014600.0 195150.0 1013400.0 ;
      RECT  193950.0 1042200.0 195150.0 1041000.0 ;
      RECT  193950.0 1069800.0 195150.0 1068600.0 ;
      RECT  193950.0 1097400.0 195150.0 1096200.0 ;
      RECT  193950.0 1125000.0 195150.0 1123800.0 ;
      RECT  193950.0 1152600.0 195150.0 1151400.0 ;
      RECT  193950.0 1180200.0 195150.0 1179000.0 ;
      RECT  193950.0 1207800.0 195150.0 1206600.0 ;
      RECT  193950.0 1235400.0 195150.0 1234200.0 ;
      RECT  193950.0 1263000.0 195150.0 1261800.0 ;
      RECT  193950.0 1290600.0 195150.0 1289400.0 ;
      RECT  193950.0 1318200.0 195150.0 1317000.0 ;
      RECT  193950.0 1345800.0 195150.0 1344600.0 ;
      RECT  193950.0 1373400.0 195150.0 1372200.0 ;
      RECT  193950.0 1401000.0 195150.0 1399800.0 ;
      RECT  193950.0 1428600.0 195150.0 1427400.0 ;
      RECT  193950.0 1456200.0 195150.0 1455000.0 ;
      RECT  193950.0 1483800.0 195150.0 1482600.0 ;
      RECT  193950.0 1511400.0 195150.0 1510200.0 ;
      RECT  193950.0 1539000.0 195150.0 1537800.0 ;
      RECT  193950.0 1566600.0 195150.0 1565400.0 ;
      RECT  193950.0 1594200.0 195150.0 1593000.0 ;
      RECT  193950.0 1621800.0 195150.0 1620600.0 ;
      RECT  193950.0 1649400.0 195150.0 1648200.0 ;
      RECT  193950.0 1677000.0 195150.0 1675800.0 ;
      RECT  193950.0 1704600.0 195150.0 1703400.0 ;
      RECT  193950.0 1732200.0 195150.0 1731000.0 ;
      RECT  193950.0 1759800.0 195150.0 1758600.0 ;
      RECT  193950.0 1787400.0 195150.0 1786200.0 ;
      RECT  193950.0 1815000.0 195150.0 1813800.0 ;
      RECT  193950.0 1842600.0 195150.0 1841400.0 ;
      RECT  193950.0 1870200.0 195150.0 1869000.0 ;
      RECT  193950.0 1897800.0 195150.0 1896600.0 ;
      RECT  193950.0 1925400.0 195150.0 1924200.0 ;
      RECT  193950.0 1953000.0 195150.0 1951800.0 ;
      RECT  193950.0 1980600.0 195150.0 1979400.0 ;
      RECT  193950.0 2008200.0 195150.0 2007000.0 ;
      RECT  193950.0 2035800.0 195150.0 2034600.0 ;
      RECT  193950.0 2063400.0 195150.0 2062200.0 ;
      RECT  193950.0 2091000.0 195150.0 2089800.0 ;
      RECT  193950.0 2118600.0 195150.0 2117400.0 ;
      RECT  193950.0 2146200.0 195150.0 2145000.0 ;
      RECT  147300.0 160650.0 146100.0 161850.0 ;
      RECT  162600.0 160500.0 161400.0 161700.0 ;
      RECT  144300.0 174450.0 143100.0 175650.0 ;
      RECT  165300.0 174300.0 164100.0 175500.0 ;
      RECT  147300.0 215850.0 146100.0 217050.0 ;
      RECT  168000.0 215700.0 166800.0 216900.0 ;
      RECT  144300.0 229650.0 143100.0 230850.0 ;
      RECT  170700.0 229500.0 169500.0 230700.0 ;
      RECT  157500.0 271050.0 156300.0 272250.0 ;
      RECT  173400.0 270900.0 172200.0 272100.0 ;
      RECT  154500.0 284850.0 153300.0 286050.0 ;
      RECT  176100.0 284700.0 174900.0 285900.0 ;
      RECT  151500.0 298650.0 150300.0 299850.0 ;
      RECT  178800.0 298500.0 177600.0 299700.0 ;
      RECT  159600.0 157800.0 158400.0 159000.0 ;
      RECT  159600.0 157800.0 158400.0 159000.0 ;
      RECT  193350.0 159000.0 194550.0 157800.0 ;
      RECT  159600.0 185400.0 158400.0 186600.0 ;
      RECT  159600.0 185400.0 158400.0 186600.0 ;
      RECT  193350.0 186600.0 194550.0 185400.0 ;
      RECT  159600.0 213000.0 158400.0 214200.0 ;
      RECT  159600.0 213000.0 158400.0 214200.0 ;
      RECT  193350.0 214200.0 194550.0 213000.0 ;
      RECT  159600.0 240600.0 158400.0 241800.0 ;
      RECT  159600.0 240600.0 158400.0 241800.0 ;
      RECT  193350.0 241800.0 194550.0 240600.0 ;
      RECT  159600.0 268200.0 158400.0 269400.0 ;
      RECT  159600.0 268200.0 158400.0 269400.0 ;
      RECT  193350.0 269400.0 194550.0 268200.0 ;
      RECT  159600.0 295800.0 158400.0 297000.0 ;
      RECT  159600.0 295800.0 158400.0 297000.0 ;
      RECT  193350.0 297000.0 194550.0 295800.0 ;
      RECT  159600.0 323400.0 158400.0 324600.0 ;
      RECT  159600.0 323400.0 158400.0 324600.0 ;
      RECT  193350.0 324600.0 194550.0 323400.0 ;
      RECT  159600.0 351000.0 158400.0 352200.0 ;
      RECT  159600.0 351000.0 158400.0 352200.0 ;
      RECT  193350.0 352200.0 194550.0 351000.0 ;
      RECT  181500.0 351150.0 180300.0 352350.0 ;
      RECT  184200.0 349050.0 183000.0 350250.0 ;
      RECT  186900.0 346950.0 185700.0 348150.0 ;
      RECT  189600.0 344850.0 188400.0 346050.0 ;
      RECT  181500.0 6600.0 180300.0 7800.0 ;
      RECT  184200.0 21000.0 183000.0 22200.0 ;
      RECT  186900.0 34200.0 185700.0 35400.0 ;
      RECT  189600.0 48600.0 188400.0 49800.0 ;
      RECT  193950.0 1200.0 195150.0 -6.83897383169e-11 ;
      RECT  193950.0 28800.0 195150.0 27600.0 ;
      RECT  193950.0 56400.0 195150.0 55200.0 ;
      RECT  118500.0 76650.0 117300.0 77850.0 ;
      RECT  97350.0 53400.0 98550.0 54600.0 ;
      RECT  118500.0 64950.0 117300.0 66150.0 ;
      RECT  100350.0 53400.0 101550.0 54600.0 ;
      RECT  118500.0 146550.0 117300.0 147750.0 ;
      RECT  162600.0 146550.0 161400.0 147750.0 ;
      RECT  118500.0 137850.0 117300.0 139050.0 ;
      RECT  165300.0 137850.0 164100.0 139050.0 ;
      RECT  118500.0 126150.0 117300.0 127350.0 ;
      RECT  168000.0 126150.0 166800.0 127350.0 ;
      RECT  118500.0 117450.0 117300.0 118650.0 ;
      RECT  170700.0 117450.0 169500.0 118650.0 ;
      RECT  118500.0 105750.0 117300.0 106950.0 ;
      RECT  173400.0 105750.0 172200.0 106950.0 ;
      RECT  118500.0 97050.0 117300.0 98250.0 ;
      RECT  176100.0 97050.0 174900.0 98250.0 ;
      RECT  118500.0 85350.0 117300.0 86550.0 ;
      RECT  178800.0 85350.0 177600.0 86550.0 ;
      RECT  120300.0 142200.0 119100.0 143400.0 ;
      RECT  195150.0 142350.0 193950.0 143550.0 ;
      RECT  120300.0 121800.0 119100.0 123000.0 ;
      RECT  195150.0 121950.0 193950.0 123150.0 ;
      RECT  120300.0 101400.0 119100.0 102600.0 ;
      RECT  195150.0 101550.0 193950.0 102750.0 ;
      RECT  120300.0 81000.0 119100.0 82200.0 ;
      RECT  195150.0 81150.0 193950.0 82350.0 ;
      RECT  120300.0 60600.0 119100.0 61800.0 ;
      RECT  195150.0 60750.0 193950.0 61950.0 ;
      RECT  210300.0 171300.0 209100.0 172500.0 ;
      RECT  204900.0 166800.0 203700.0 168000.0 ;
      RECT  207600.0 164400.0 206400.0 165600.0 ;
      RECT  210300.0 2153850.0 209100.0 2155050.0 ;
      RECT  213000.0 236100.0 211800.0 237300.0 ;
      RECT  215700.0 334200.0 214500.0 335400.0 ;
      RECT  202200.0 154500.0 201000.0 155700.0 ;
      RECT  121650.0 2147100.0 120450.0 2148300.0 ;
      RECT  202200.0 2147100.0 201000.0 2148300.0 ;
      RECT  198450.0 162450.0 197250.0 163650.0 ;
      RECT  198450.0 332250.0 197250.0 333450.0 ;
      RECT  198450.0 234150.0 197250.0 235350.0 ;
      RECT  225900.0 600.0 226800.0 2400.0 ;
      RECT  266700.0 600.0 267600.0 2400.0 ;
      RECT  307500.0 600.0 308400.0 2400.0 ;
      RECT  348300.0 600.0 349200.0 2400.0 ;
      RECT  389100.0 600.0 390000.0 2400.0 ;
      RECT  429900.0 600.0 430800.0 2400.0 ;
      RECT  470700.0 600.0 471600.0 2400.0 ;
      RECT  511500.0 600.0 512400.0 2400.0 ;
      RECT  552300.0 600.0 553200.0 2400.0 ;
      RECT  593100.0 600.0 594000.0 2400.0 ;
      RECT  633900.0 600.0 634800.0 2400.0 ;
      RECT  674700.0 600.0 675600.0 2400.0 ;
      RECT  715500.0 600.0 716400.0 2400.0 ;
      RECT  756300.0 600.0 757200.0 2400.0 ;
      RECT  797100.0 600.0 798000.0 2400.0 ;
      RECT  837900.0 600.0 838800.0 2400.0 ;
      RECT  878700.0 600.0 879600.0 2400.0 ;
      RECT  919500.0 600.0 920400.0 2400.0 ;
      RECT  960300.0 600.0 961200.0 2400.0 ;
      RECT  1001100.0 600.0 1002000.0 2400.0 ;
      RECT  1041900.0 600.0 1042800.0 2400.0 ;
      RECT  1082700.0 600.0 1083600.0 2400.0 ;
      RECT  1123500.0 600.0 1124400.0 2400.0 ;
      RECT  1164300.0 600.0 1165200.0 2400.0 ;
      RECT  1205100.0 600.0 1206000.0 2400.0 ;
      RECT  1245900.0 600.0 1246800.0 2400.0 ;
      RECT  1286700.0 600.0 1287600.0 2400.0 ;
      RECT  1327500.0 600.0 1328400.0 2400.0 ;
      RECT  1368300.0 600.0 1369200.0 2400.0 ;
      RECT  1409100.0 600.0 1410000.0 2400.0 ;
      RECT  1449900.0 600.0 1450800.0 2400.0 ;
      RECT  1490700.0 600.0 1491600.0 2400.0 ;
      RECT  214650.0 600.0 215550.0 2166000.0 ;
      RECT  211950.0 600.0 212850.0 2166000.0 ;
      RECT  203850.0 600.0 204750.0 2166000.0 ;
      RECT  206550.0 600.0 207450.0 2166000.0 ;
      RECT  209250.0 600.0 210150.0 2166000.0 ;
      RECT  201150.0 600.0 202050.0 2166000.0 ;
      RECT  193950.0 600.0 198450.0 2166000.0 ;
      RECT  49800.0 469800.0 1.42108547152e-11 470700.0 ;
      RECT  49800.0 472500.0 1.42108547152e-11 473400.0 ;
      RECT  49800.0 475200.0 1.42108547152e-11 476100.0 ;
      RECT  49800.0 480600.0 1.42108547152e-11 481500.0 ;
      RECT  43350.0 423450.0 36000.0 424350.0 ;
      RECT  33750.0 385050.0 32850.0 464850.0 ;
      RECT  49800.0 467100.0 47100.0 468000.0 ;
      RECT  38700.0 477900.0 36000.0 478800.0 ;
      RECT  24900.0 467100.0 22200.0 468000.0 ;
      RECT  11100.0 477900.0 8400.0 478800.0 ;
      RECT  7.1054273576e-12 382200.0 10200.0 442200.0 ;
      RECT  20400.0 382200.0 10200.0 442200.0 ;
      RECT  20400.0 382200.0 30600.0 442200.0 ;
      RECT  4500.0 439800.0 7200.0 441000.0 ;
      RECT  1800.0 437700.0 3000.0 442200.0 ;
      RECT  13200.0 439800.0 15900.0 441000.0 ;
      RECT  17400.0 437700.0 18600.0 442200.0 ;
      RECT  24900.0 439800.0 27600.0 441000.0 ;
      RECT  22200.0 437700.0 23400.0 442200.0 ;
      RECT  9600.0 382200.0 10800.0 442200.0 ;
      RECT  30000.0 382200.0 31200.0 442200.0 ;
      RECT  46650.0 497850.0 39150.0 498750.0 ;
      RECT  41700.0 493050.0 40800.0 493950.0 ;
      RECT  41700.0 497850.0 40800.0 498750.0 ;
      RECT  41250.0 493050.0 39150.0 493950.0 ;
      RECT  41700.0 493500.0 40800.0 498300.0 ;
      RECT  46650.0 497850.0 41250.0 498750.0 ;
      RECT  39150.0 492900.0 37950.0 494100.0 ;
      RECT  39150.0 497700.0 37950.0 498900.0 ;
      RECT  47850.0 497700.0 46650.0 498900.0 ;
      RECT  41850.0 497700.0 40650.0 498900.0 ;
      RECT  28800.0 495450.0 29700.0 496350.0 ;
      RECT  29250.0 495450.0 32250.0 496350.0 ;
      RECT  28800.0 495900.0 29700.0 496800.0 ;
      RECT  23700.0 495450.0 24600.0 496350.0 ;
      RECT  23700.0 494100.0 24600.0 495900.0 ;
      RECT  24150.0 495450.0 29250.0 496350.0 ;
      RECT  32250.0 495300.0 33450.0 496500.0 ;
      RECT  23550.0 494100.0 24750.0 492900.0 ;
      RECT  28650.0 497400.0 29850.0 496200.0 ;
      RECT  29550.0 510150.0 30450.0 511050.0 ;
      RECT  29550.0 512550.0 30450.0 513450.0 ;
      RECT  30000.0 510150.0 32850.0 511050.0 ;
      RECT  29550.0 510600.0 30450.0 513000.0 ;
      RECT  25350.0 512550.0 30000.0 513450.0 ;
      RECT  32850.0 510000.0 34050.0 511200.0 ;
      RECT  24150.0 512400.0 25350.0 513600.0 ;
      RECT  29400.0 513600.0 30600.0 512400.0 ;
      RECT  19050.0 507450.0 11550.0 508350.0 ;
      RECT  14100.0 502650.0 13200.0 503550.0 ;
      RECT  14100.0 507450.0 13200.0 508350.0 ;
      RECT  13650.0 502650.0 11550.0 503550.0 ;
      RECT  14100.0 503100.0 13200.0 507900.0 ;
      RECT  19050.0 507450.0 13650.0 508350.0 ;
      RECT  11550.0 502500.0 10350.0 503700.0 ;
      RECT  11550.0 507300.0 10350.0 508500.0 ;
      RECT  20250.0 507300.0 19050.0 508500.0 ;
      RECT  14250.0 507300.0 13050.0 508500.0 ;
      RECT  3000.0 442800.0 1800.0 441600.0 ;
      RECT  3000.0 481650.0 1800.0 480450.0 ;
      RECT  6450.0 441600.0 5250.0 440400.0 ;
      RECT  6450.0 470850.0 5250.0 469650.0 ;
      RECT  18600.0 442800.0 17400.0 441600.0 ;
      RECT  18600.0 473550.0 17400.0 472350.0 ;
      RECT  23400.0 442800.0 22200.0 441600.0 ;
      RECT  23400.0 476250.0 22200.0 475050.0 ;
      RECT  10800.0 442800.0 9600.0 441600.0 ;
      RECT  10800.0 468150.0 9600.0 466950.0 ;
      RECT  31200.0 442800.0 30000.0 441600.0 ;
      RECT  31200.0 468150.0 30000.0 466950.0 ;
      RECT  22650.0 551700.0 21750.0 941100.0 ;
      RECT  17250.0 551700.0 16350.0 936300.0 ;
      RECT  7050.0 551700.0 6150.0 936300.0 ;
      RECT  20400.0 555900.0 19500.0 564000.0 ;
      RECT  13650.0 555900.0 12750.0 560700.0 ;
      RECT  42750.0 595500.0 43650.0 602700.0 ;
      RECT  42750.0 602700.0 43650.0 612300.0 ;
      RECT  42750.0 612300.0 43650.0 621900.0 ;
      RECT  42750.0 624300.0 43650.0 631500.0 ;
      RECT  42750.0 631500.0 43650.0 641100.0 ;
      RECT  42750.0 641100.0 43650.0 650700.0 ;
      RECT  35550.0 652650.0 36450.0 653550.0 ;
      RECT  35550.0 644250.0 36450.0 645150.0 ;
      RECT  36000.0 652650.0 43200.0 653550.0 ;
      RECT  35550.0 644700.0 36450.0 653100.0 ;
      RECT  28800.0 644250.0 36000.0 645150.0 ;
      RECT  28350.0 635100.0 29250.0 644700.0 ;
      RECT  28350.0 625500.0 29250.0 635100.0 ;
      RECT  28350.0 615900.0 29250.0 623100.0 ;
      RECT  28350.0 606300.0 29250.0 615900.0 ;
      RECT  28350.0 596700.0 29250.0 606300.0 ;
      RECT  42600.0 602100.0 43800.0 603300.0 ;
      RECT  42600.0 611700.0 43800.0 612900.0 ;
      RECT  42600.0 621300.0 43800.0 622500.0 ;
      RECT  42600.0 630900.0 43800.0 632100.0 ;
      RECT  42600.0 640500.0 43800.0 641700.0 ;
      RECT  42600.0 650100.0 43800.0 651300.0 ;
      RECT  28200.0 644100.0 29400.0 645300.0 ;
      RECT  28200.0 634500.0 29400.0 635700.0 ;
      RECT  28200.0 624900.0 29400.0 626100.0 ;
      RECT  28200.0 615300.0 29400.0 616500.0 ;
      RECT  28200.0 605700.0 29400.0 606900.0 ;
      RECT  28200.0 596100.0 29400.0 597300.0 ;
      RECT  42600.0 594900.0 43800.0 596100.0 ;
      RECT  42600.0 623700.0 43800.0 624900.0 ;
      RECT  42600.0 652500.0 43800.0 653700.0 ;
      RECT  28200.0 622500.0 29400.0 623700.0 ;
      RECT  16800.0 575100.0 6600.0 561300.0 ;
      RECT  16800.0 575100.0 6600.0 588900.0 ;
      RECT  16800.0 602700.0 6600.0 588900.0 ;
      RECT  16800.0 602700.0 6600.0 616500.0 ;
      RECT  16800.0 630300.0 6600.0 616500.0 ;
      RECT  16800.0 630300.0 6600.0 644100.0 ;
      RECT  16800.0 657900.0 6600.0 644100.0 ;
      RECT  16800.0 657900.0 6600.0 671700.0 ;
      RECT  16800.0 685500.0 6600.0 671700.0 ;
      RECT  16800.0 685500.0 6600.0 699300.0 ;
      RECT  16800.0 713100.0 6600.0 699300.0 ;
      RECT  16800.0 713100.0 6600.0 726900.0 ;
      RECT  16800.0 740700.0 6600.0 726900.0 ;
      RECT  16800.0 740700.0 6600.0 754500.0 ;
      RECT  16800.0 768300.0 6600.0 754500.0 ;
      RECT  16800.0 768300.0 6600.0 782100.0 ;
      RECT  16800.0 795900.0 6600.0 782100.0 ;
      RECT  16800.0 795900.0 6600.0 809700.0 ;
      RECT  16800.0 823500.0 6600.0 809700.0 ;
      RECT  16800.0 823500.0 6600.0 837300.0 ;
      RECT  16800.0 851100.0 6600.0 837300.0 ;
      RECT  16800.0 851100.0 6600.0 864900.0 ;
      RECT  16800.0 878700.0 6600.0 864900.0 ;
      RECT  16800.0 878700.0 6600.0 892500.0 ;
      RECT  16800.0 906300.0 6600.0 892500.0 ;
      RECT  16800.0 906300.0 6600.0 920100.0 ;
      RECT  16800.0 933900.0 6600.0 920100.0 ;
      RECT  13800.0 575700.0 12600.0 937500.0 ;
      RECT  10800.0 574500.0 9600.0 936300.0 ;
      RECT  17400.0 574500.0 16200.0 936300.0 ;
      RECT  7200.0 574500.0 6000.0 936300.0 ;
      RECT  22350.0 576600.0 21150.0 577800.0 ;
      RECT  22350.0 600000.0 21150.0 601200.0 ;
      RECT  22350.0 604200.0 21150.0 605400.0 ;
      RECT  22350.0 627600.0 21150.0 628800.0 ;
      RECT  22350.0 631800.0 21150.0 633000.0 ;
      RECT  22350.0 655200.0 21150.0 656400.0 ;
      RECT  22350.0 659400.0 21150.0 660600.0 ;
      RECT  22350.0 682800.0 21150.0 684000.0 ;
      RECT  22350.0 687000.0 21150.0 688200.0 ;
      RECT  22350.0 710400.0 21150.0 711600.0 ;
      RECT  22350.0 714600.0 21150.0 715800.0 ;
      RECT  22350.0 738000.0 21150.0 739200.0 ;
      RECT  22350.0 742200.0 21150.0 743400.0 ;
      RECT  22350.0 765600.0 21150.0 766800.0 ;
      RECT  22350.0 769800.0 21150.0 771000.0 ;
      RECT  22350.0 793200.0 21150.0 794400.0 ;
      RECT  22350.0 797400.0 21150.0 798600.0 ;
      RECT  22350.0 820800.0 21150.0 822000.0 ;
      RECT  22350.0 825000.0 21150.0 826200.0 ;
      RECT  22350.0 848400.0 21150.0 849600.0 ;
      RECT  22350.0 852600.0 21150.0 853800.0 ;
      RECT  22350.0 876000.0 21150.0 877200.0 ;
      RECT  22350.0 880200.0 21150.0 881400.0 ;
      RECT  22350.0 903600.0 21150.0 904800.0 ;
      RECT  22350.0 907800.0 21150.0 909000.0 ;
      RECT  22350.0 931200.0 21150.0 932400.0 ;
      RECT  22200.0 590100.0 21000.0 591300.0 ;
      RECT  22800.0 550500.0 21600.0 551700.0 ;
      RECT  16200.0 551100.0 17400.0 552300.0 ;
      RECT  6000.0 551100.0 7200.0 552300.0 ;
      RECT  19350.0 563400.0 20550.0 564600.0 ;
      RECT  19350.0 555300.0 20550.0 556500.0 ;
      RECT  12600.0 555300.0 13800.0 556500.0 ;
      RECT  43950.0 465450.0 42750.0 464250.0 ;
      RECT  43950.0 424500.0 42750.0 423300.0 ;
      RECT  36600.0 424500.0 35400.0 423300.0 ;
      RECT  36600.0 484350.0 35400.0 483150.0 ;
      RECT  33900.0 385650.0 32700.0 384450.0 ;
      RECT  29850.0 465450.0 28650.0 464250.0 ;
      RECT  27150.0 470850.0 25950.0 469650.0 ;
      RECT  30600.0 508200.0 29400.0 507000.0 ;
      RECT  30600.0 508200.0 29400.0 507000.0 ;
      RECT  30600.0 484350.0 29400.0 483150.0 ;
      RECT  27900.0 511200.0 26700.0 510000.0 ;
      RECT  27900.0 511200.0 26700.0 510000.0 ;
      RECT  27900.0 481650.0 26700.0 480450.0 ;
      RECT  41850.0 484350.0 40650.0 483150.0 ;
      RECT  43800.0 481650.0 42600.0 480450.0 ;
      RECT  45750.0 473550.0 44550.0 472350.0 ;
      RECT  14250.0 484350.0 13050.0 483150.0 ;
      RECT  16200.0 473550.0 15000.0 472350.0 ;
      RECT  18150.0 476250.0 16950.0 475050.0 ;
      RECT  29850.0 502500.0 28650.0 503700.0 ;
      RECT  30600.0 519600.0 29400.0 520800.0 ;
      RECT  16200.0 542100.0 15000.0 543300.0 ;
      RECT  29400.0 522300.0 28200.0 523500.0 ;
      RECT  50400.0 468150.0 49200.0 466950.0 ;
      RECT  36600.0 478950.0 35400.0 477750.0 ;
      RECT  22800.0 468150.0 21600.0 466950.0 ;
      RECT  9000.0 478950.0 7800.0 477750.0 ;
      RECT  49800.0 522450.0 28800.0 523350.0 ;
      RECT  49800.0 542250.0 15600.0 543150.0 ;
      RECT  49800.0 502650.0 29250.0 503550.0 ;
      RECT  49800.0 519750.0 30000.0 520650.0 ;
      RECT  49800.0 483300.0 1.42108547152e-11 484200.0 ;
      RECT  49800.0 464400.0 1.42108547152e-11 465300.0 ;
      RECT  49800.0 477900.0 1.42108547152e-11 478800.0 ;
      RECT  49800.0 467100.0 1.42108547152e-11 468000.0 ;
      RECT  215700.0 522300.0 214500.0 523500.0 ;
      RECT  49500.0 522450.0 48300.0 523650.0 ;
      RECT  213000.0 542100.0 211800.0 543300.0 ;
      RECT  49500.0 542250.0 48300.0 543450.0 ;
      RECT  207600.0 502500.0 206400.0 503700.0 ;
      RECT  49500.0 502650.0 48300.0 503850.0 ;
      RECT  204900.0 519600.0 203700.0 520800.0 ;
      RECT  49500.0 519750.0 48300.0 520950.0 ;
      RECT  210300.0 483150.0 209100.0 484350.0 ;
      RECT  49500.0 483300.0 48300.0 484500.0 ;
      RECT  202200.0 464250.0 201000.0 465450.0 ;
      RECT  49500.0 464400.0 48300.0 465600.0 ;
      RECT  55650.0 477750.0 54450.0 478950.0 ;
      RECT  196800.0 466950.0 195600.0 468150.0 ;
      RECT  49500.0 467100.0 48300.0 468300.0 ;
   LAYER  metal3 ;
      RECT  49800.0 522150.0 215100.0 523650.0 ;
      RECT  49800.0 541950.0 212400.0 543450.0 ;
      RECT  49800.0 502350.0 207000.0 503850.0 ;
      RECT  49800.0 519450.0 204300.0 520950.0 ;
      RECT  49800.0 483000.0 209700.0 484500.0 ;
      RECT  49800.0 464100.0 201600.0 465600.0 ;
      RECT  49800.0 466800.0 196200.0 468300.0 ;
      RECT  222150.0 145350.0 223650.0 290550.0 ;
      RECT  262950.0 145350.0 264450.0 290550.0 ;
      RECT  303750.0 145350.0 305250.0 290550.0 ;
      RECT  344550.0 145350.0 346050.0 290550.0 ;
      RECT  385350.0 145350.0 386850.0 290550.0 ;
      RECT  426150.0 145350.0 427650.0 290550.0 ;
      RECT  466950.0 145350.0 468450.0 290550.0 ;
      RECT  507750.0 145350.0 509250.0 290550.0 ;
      RECT  548550.0 145350.0 550050.0 290550.0 ;
      RECT  589350.0 145350.0 590850.0 290550.0 ;
      RECT  630150.0 145350.0 631650.0 290550.0 ;
      RECT  670950.0 145350.0 672450.0 290550.0 ;
      RECT  711750.0 145350.0 713250.0 290550.0 ;
      RECT  752550.0 145350.0 754050.0 290550.0 ;
      RECT  793350.0 145350.0 794850.0 290550.0 ;
      RECT  834150.0 145350.0 835650.0 290550.0 ;
      RECT  874950.0 145350.0 876450.0 290550.0 ;
      RECT  915750.0 145350.0 917250.0 290550.0 ;
      RECT  956550.0 145350.0 958050.0 290550.0 ;
      RECT  997350.0 145350.0 998850.0 290550.0 ;
      RECT  1038150.0 145350.0 1039650.0 290550.0 ;
      RECT  1078950.0 145350.0 1080450.0 290550.0 ;
      RECT  1119750.0 145350.0 1121250.0 290550.0 ;
      RECT  1160550.0 145350.0 1162050.0 290550.0 ;
      RECT  1201350.0 145350.0 1202850.0 290550.0 ;
      RECT  1242150.0 145350.0 1243650.0 290550.0 ;
      RECT  1282950.0 145350.0 1284450.0 290550.0 ;
      RECT  1323750.0 145350.0 1325250.0 290550.0 ;
      RECT  1364550.0 145350.0 1366050.0 290550.0 ;
      RECT  1405350.0 145350.0 1406850.0 290550.0 ;
      RECT  1446150.0 145350.0 1447650.0 290550.0 ;
      RECT  1486950.0 145350.0 1488450.0 290550.0 ;
      RECT  225900.0 600.0 227400.0 169050.0 ;
      RECT  266700.0 600.0 268200.0 169050.0 ;
      RECT  307500.0 600.0 309000.0 169050.0 ;
      RECT  348300.0 600.0 349800.0 169050.0 ;
      RECT  389100.0 600.0 390600.0 169050.0 ;
      RECT  429900.0 600.0 431400.0 169050.0 ;
      RECT  470700.0 600.0 472200.0 169050.0 ;
      RECT  511500.0 600.0 513000.0 169050.0 ;
      RECT  552300.0 600.0 553800.0 169050.0 ;
      RECT  593100.0 600.0 594600.0 169050.0 ;
      RECT  633900.0 600.0 635400.0 169050.0 ;
      RECT  674700.0 600.0 676200.0 169050.0 ;
      RECT  715500.0 600.0 717000.0 169050.0 ;
      RECT  756300.0 600.0 757800.0 169050.0 ;
      RECT  797100.0 600.0 798600.0 169050.0 ;
      RECT  837900.0 600.0 839400.0 169050.0 ;
      RECT  878700.0 600.0 880200.0 169050.0 ;
      RECT  919500.0 600.0 921000.0 169050.0 ;
      RECT  960300.0 600.0 961800.0 169050.0 ;
      RECT  1001100.0 600.0 1002600.0 169050.0 ;
      RECT  1041900.0 600.0 1043400.0 169050.0 ;
      RECT  1082700.0 600.0 1084200.0 169050.0 ;
      RECT  1123500.0 600.0 1125000.0 169050.0 ;
      RECT  1164300.0 600.0 1165800.0 169050.0 ;
      RECT  1205100.0 600.0 1206600.0 169050.0 ;
      RECT  1245900.0 600.0 1247400.0 169050.0 ;
      RECT  1286700.0 600.0 1288200.0 169050.0 ;
      RECT  1327500.0 600.0 1329000.0 169050.0 ;
      RECT  1368300.0 600.0 1369800.0 169050.0 ;
      RECT  1409100.0 600.0 1410600.0 169050.0 ;
      RECT  1449900.0 600.0 1451400.0 169050.0 ;
      RECT  1490700.0 600.0 1492200.0 169050.0 ;
      RECT  159000.0 157650.0 193950.0 159150.0 ;
      RECT  159000.0 185250.0 193950.0 186750.0 ;
      RECT  159000.0 212850.0 193950.0 214350.0 ;
      RECT  159000.0 240450.0 193950.0 241950.0 ;
      RECT  159000.0 268050.0 193950.0 269550.0 ;
      RECT  159000.0 295650.0 193950.0 297150.0 ;
      RECT  159000.0 323250.0 193950.0 324750.0 ;
      RECT  159000.0 350850.0 193950.0 352350.0 ;
      RECT  97200.0 76500.0 98700.0 78000.0 ;
      RECT  97950.0 76500.0 117900.0 78000.0 ;
      RECT  97200.0 54000.0 98700.0 77250.0 ;
      RECT  100200.0 64800.0 101700.0 66300.0 ;
      RECT  100950.0 64800.0 117900.0 66300.0 ;
      RECT  100200.0 54000.0 101700.0 65550.0 ;
      RECT  222000.0 290550.0 223800.0 292350.0 ;
      RECT  262800.0 290550.0 264600.0 292350.0 ;
      RECT  303600.0 290550.0 305400.0 292350.0 ;
      RECT  344400.0 290550.0 346200.0 292350.0 ;
      RECT  385200.0 290550.0 387000.0 292350.0 ;
      RECT  426000.0 290550.0 427800.0 292350.0 ;
      RECT  466800.0 290550.0 468600.0 292350.0 ;
      RECT  507600.0 290550.0 509400.0 292350.0 ;
      RECT  548400.0 290550.0 550200.0 292350.0 ;
      RECT  589200.0 290550.0 591000.0 292350.0 ;
      RECT  630000.0 290550.0 631800.0 292350.0 ;
      RECT  670800.0 290550.0 672600.0 292350.0 ;
      RECT  711600.0 290550.0 713400.0 292350.0 ;
      RECT  752400.0 290550.0 754200.0 292350.0 ;
      RECT  793200.0 290550.0 795000.0 292350.0 ;
      RECT  834000.0 290550.0 835800.0 292350.0 ;
      RECT  874800.0 290550.0 876600.0 292350.0 ;
      RECT  915600.0 290550.0 917400.0 292350.0 ;
      RECT  956400.0 290550.0 958200.0 292350.0 ;
      RECT  997200.0 290550.0 999000.0 292350.0 ;
      RECT  1038000.0 290550.0 1039800.0 292350.0 ;
      RECT  1078800.0 290550.0 1080600.0 292350.0 ;
      RECT  1119600.0 290550.0 1121400.0 292350.0 ;
      RECT  1160400.0 290550.0 1162200.0 292350.0 ;
      RECT  1201200.0 290550.0 1203000.0 292350.0 ;
      RECT  1242000.0 290550.0 1243800.0 292350.0 ;
      RECT  1282800.0 290550.0 1284600.0 292350.0 ;
      RECT  1323600.0 290550.0 1325400.0 292350.0 ;
      RECT  1364400.0 290550.0 1366200.0 292350.0 ;
      RECT  1405200.0 290550.0 1407000.0 292350.0 ;
      RECT  1446000.0 290550.0 1447800.0 292350.0 ;
      RECT  1486800.0 290550.0 1488600.0 292350.0 ;
      RECT  225600.0 169950.0 227400.0 171750.0 ;
      RECT  266400.0 169950.0 268200.0 171750.0 ;
      RECT  307200.0 169950.0 309000.0 171750.0 ;
      RECT  348000.0 169950.0 349800.0 171750.0 ;
      RECT  388800.0 169950.0 390600.0 171750.0 ;
      RECT  429600.0 169950.0 431400.0 171750.0 ;
      RECT  470400.0 169950.0 472200.0 171750.0 ;
      RECT  511200.0 169950.0 513000.0 171750.0 ;
      RECT  552000.0 169950.0 553800.0 171750.0 ;
      RECT  592800.0 169950.0 594600.0 171750.0 ;
      RECT  633600.0 169950.0 635400.0 171750.0 ;
      RECT  674400.0 169950.0 676200.0 171750.0 ;
      RECT  715200.0 169950.0 717000.0 171750.0 ;
      RECT  756000.0 169950.0 757800.0 171750.0 ;
      RECT  796800.0 169950.0 798600.0 171750.0 ;
      RECT  837600.0 169950.0 839400.0 171750.0 ;
      RECT  878400.0 169950.0 880200.0 171750.0 ;
      RECT  919200.0 169950.0 921000.0 171750.0 ;
      RECT  960000.0 169950.0 961800.0 171750.0 ;
      RECT  1000800.0 169950.0 1002600.0 171750.0 ;
      RECT  1041600.0 169950.0 1043400.0 171750.0 ;
      RECT  1082400.0 169950.0 1084200.0 171750.0 ;
      RECT  1123200.0 169950.0 1125000.0 171750.0 ;
      RECT  1164000.0 169950.0 1165800.0 171750.0 ;
      RECT  1204800.0 169950.0 1206600.0 171750.0 ;
      RECT  1245600.0 169950.0 1247400.0 171750.0 ;
      RECT  1286400.0 169950.0 1288200.0 171750.0 ;
      RECT  1327200.0 169950.0 1329000.0 171750.0 ;
      RECT  1368000.0 169950.0 1369800.0 171750.0 ;
      RECT  1408800.0 169950.0 1410600.0 171750.0 ;
      RECT  1449600.0 169950.0 1451400.0 171750.0 ;
      RECT  1490400.0 169950.0 1492200.0 171750.0 ;
      RECT  60000.0 148800.0 61800.0 147000.0 ;
      RECT  60000.0 138600.0 61800.0 136800.0 ;
      RECT  60000.0 128400.0 61800.0 126600.0 ;
      RECT  60000.0 118200.0 61800.0 116400.0 ;
      RECT  60000.0 108000.0 61800.0 106200.0 ;
      RECT  60000.0 97800.0 61800.0 96000.0 ;
      RECT  60000.0 87600.0 61800.0 85800.0 ;
      RECT  60000.0 77400.0 61800.0 75600.0 ;
      RECT  60000.0 67200.0 61800.0 65400.0 ;
      RECT  222150.0 144600.0 223950.0 146400.0 ;
      RECT  262950.0 144600.0 264750.0 146400.0 ;
      RECT  303750.0 144600.0 305550.0 146400.0 ;
      RECT  344550.0 144600.0 346350.0 146400.0 ;
      RECT  385350.0 144600.0 387150.0 146400.0 ;
      RECT  426150.0 144600.0 427950.0 146400.0 ;
      RECT  466950.0 144600.0 468750.0 146400.0 ;
      RECT  507750.0 144600.0 509550.0 146400.0 ;
      RECT  548550.0 144600.0 550350.0 146400.0 ;
      RECT  589350.0 144600.0 591150.0 146400.0 ;
      RECT  630150.0 144600.0 631950.0 146400.0 ;
      RECT  670950.0 144600.0 672750.0 146400.0 ;
      RECT  711750.0 144600.0 713550.0 146400.0 ;
      RECT  752550.0 144600.0 754350.0 146400.0 ;
      RECT  793350.0 144600.0 795150.0 146400.0 ;
      RECT  834150.0 144600.0 835950.0 146400.0 ;
      RECT  874950.0 144600.0 876750.0 146400.0 ;
      RECT  915750.0 144600.0 917550.0 146400.0 ;
      RECT  956550.0 144600.0 958350.0 146400.0 ;
      RECT  997350.0 144600.0 999150.0 146400.0 ;
      RECT  1038150.0 144600.0 1039950.0 146400.0 ;
      RECT  1078950.0 144600.0 1080750.0 146400.0 ;
      RECT  1119750.0 144600.0 1121550.0 146400.0 ;
      RECT  1160550.0 144600.0 1162350.0 146400.0 ;
      RECT  1201350.0 144600.0 1203150.0 146400.0 ;
      RECT  1242150.0 144600.0 1243950.0 146400.0 ;
      RECT  1282950.0 144600.0 1284750.0 146400.0 ;
      RECT  1323750.0 144600.0 1325550.0 146400.0 ;
      RECT  1364550.0 144600.0 1366350.0 146400.0 ;
      RECT  1405350.0 144600.0 1407150.0 146400.0 ;
      RECT  1446150.0 144600.0 1447950.0 146400.0 ;
      RECT  1486950.0 144600.0 1488750.0 146400.0 ;
      RECT  225900.0 600.0 227700.0 2400.0 ;
      RECT  266700.0 600.0 268500.0 2400.0 ;
      RECT  307500.0 600.0 309300.0 2400.0 ;
      RECT  348300.0 600.0 350100.0 2400.0 ;
      RECT  389100.0 600.0 390900.0 2400.0 ;
      RECT  429900.0 600.0 431700.0 2400.0 ;
      RECT  470700.0 600.0 472500.0 2400.0 ;
      RECT  511500.0 600.0 513300.0 2400.0 ;
      RECT  552300.0 600.0 554100.0 2400.0 ;
      RECT  593100.0 600.0 594900.0 2400.0 ;
      RECT  633900.0 600.0 635700.0 2400.0 ;
      RECT  674700.0 600.0 676500.0 2400.0 ;
      RECT  715500.0 600.0 717300.0 2400.0 ;
      RECT  756300.0 600.0 758100.0 2400.0 ;
      RECT  797100.0 600.0 798900.0 2400.0 ;
      RECT  837900.0 600.0 839700.0 2400.0 ;
      RECT  878700.0 600.0 880500.0 2400.0 ;
      RECT  919500.0 600.0 921300.0 2400.0 ;
      RECT  960300.0 600.0 962100.0 2400.0 ;
      RECT  1001100.0 600.0 1002900.0 2400.0 ;
      RECT  1041900.0 600.0 1043700.0 2400.0 ;
      RECT  1082700.0 600.0 1084500.0 2400.0 ;
      RECT  1123500.0 600.0 1125300.0 2400.0 ;
      RECT  1164300.0 600.0 1166100.0 2400.0 ;
      RECT  1205100.0 600.0 1206900.0 2400.0 ;
      RECT  1245900.0 600.0 1247700.0 2400.0 ;
      RECT  1286700.0 600.0 1288500.0 2400.0 ;
      RECT  1327500.0 600.0 1329300.0 2400.0 ;
      RECT  1368300.0 600.0 1370100.0 2400.0 ;
      RECT  1409100.0 600.0 1410900.0 2400.0 ;
      RECT  1449900.0 600.0 1451700.0 2400.0 ;
      RECT  1490700.0 600.0 1492500.0 2400.0 ;
      RECT  159900.0 157500.0 158100.0 159300.0 ;
      RECT  193050.0 159300.0 194850.0 157500.0 ;
      RECT  159900.0 185100.0 158100.0 186900.0 ;
      RECT  193050.0 186900.0 194850.0 185100.0 ;
      RECT  159900.0 212700.0 158100.0 214500.0 ;
      RECT  193050.0 214500.0 194850.0 212700.0 ;
      RECT  159900.0 240300.0 158100.0 242100.0 ;
      RECT  193050.0 242100.0 194850.0 240300.0 ;
      RECT  159900.0 267900.0 158100.0 269700.0 ;
      RECT  193050.0 269700.0 194850.0 267900.0 ;
      RECT  159900.0 295500.0 158100.0 297300.0 ;
      RECT  193050.0 297300.0 194850.0 295500.0 ;
      RECT  159900.0 323100.0 158100.0 324900.0 ;
      RECT  193050.0 324900.0 194850.0 323100.0 ;
      RECT  159900.0 350700.0 158100.0 352500.0 ;
      RECT  193050.0 352500.0 194850.0 350700.0 ;
      RECT  118800.0 76350.0 117000.0 78150.0 ;
      RECT  97050.0 53100.0 98850.0 54900.0 ;
      RECT  118800.0 64650.0 117000.0 66450.0 ;
      RECT  100050.0 53100.0 101850.0 54900.0 ;
      RECT  52800.0 147000.0 60000.0 148500.0 ;
      RECT  52800.0 136800.0 60000.0 138300.0 ;
      RECT  52800.0 126600.0 60000.0 128100.0 ;
      RECT  52800.0 116400.0 60000.0 117900.0 ;
      RECT  52800.0 106200.0 60000.0 107700.0 ;
      RECT  52800.0 96000.0 60000.0 97500.0 ;
      RECT  52800.0 85800.0 60000.0 87300.0 ;
      RECT  52800.0 75600.0 60000.0 77100.0 ;
      RECT  52800.0 65400.0 60000.0 66900.0 ;
      RECT  3150.0 442200.0 1650.0 481050.0 ;
      RECT  6600.0 441000.0 5100.0 470250.0 ;
      RECT  18750.0 442200.0 17250.0 472950.0 ;
      RECT  23550.0 442200.0 22050.0 475650.0 ;
      RECT  10950.0 442200.0 9450.0 467550.0 ;
      RECT  31350.0 442200.0 29850.0 467550.0 ;
      RECT  36750.0 423900.0 35250.0 483750.0 ;
      RECT  30750.0 483750.0 29250.0 507600.0 ;
      RECT  28050.0 481050.0 26550.0 510600.0 ;
      RECT  4200.0 383100.0 6000.0 384900.0 ;
      RECT  14400.0 383100.0 16200.0 384900.0 ;
      RECT  24600.0 383100.0 26400.0 384900.0 ;
      RECT  3300.0 443100.0 1500.0 441300.0 ;
      RECT  3300.0 481950.0 1500.0 480150.0 ;
      RECT  6750.0 441900.0 4950.0 440100.0 ;
      RECT  6750.0 471150.0 4950.0 469350.0 ;
      RECT  18900.0 443100.0 17100.0 441300.0 ;
      RECT  18900.0 473850.0 17100.0 472050.0 ;
      RECT  23700.0 443100.0 21900.0 441300.0 ;
      RECT  23700.0 476550.0 21900.0 474750.0 ;
      RECT  11100.0 443100.0 9300.0 441300.0 ;
      RECT  11100.0 468450.0 9300.0 466650.0 ;
      RECT  31500.0 443100.0 29700.0 441300.0 ;
      RECT  31500.0 468450.0 29700.0 466650.0 ;
      RECT  36900.0 424800.0 35100.0 423000.0 ;
      RECT  36900.0 484650.0 35100.0 482850.0 ;
      RECT  30900.0 508500.0 29100.0 506700.0 ;
      RECT  30900.0 484650.0 29100.0 482850.0 ;
      RECT  28200.0 511500.0 26400.0 509700.0 ;
      RECT  28200.0 481950.0 26400.0 480150.0 ;
      RECT  16200.0 383100.0 14400.0 384900.0 ;
      RECT  26400.0 383100.0 24600.0 384900.0 ;
      RECT  6000.0 383100.0 4200.0 384900.0 ;
      RECT  216000.0 522000.0 214200.0 523800.0 ;
      RECT  49800.0 522150.0 48000.0 523950.0 ;
      RECT  213300.0 541800.0 211500.0 543600.0 ;
      RECT  49800.0 541950.0 48000.0 543750.0 ;
      RECT  207900.0 502200.0 206100.0 504000.0 ;
      RECT  49800.0 502350.0 48000.0 504150.0 ;
      RECT  205200.0 519300.0 203400.0 521100.0 ;
      RECT  49800.0 519450.0 48000.0 521250.0 ;
      RECT  210600.0 482850.0 208800.0 484650.0 ;
      RECT  49800.0 483000.0 48000.0 484800.0 ;
      RECT  202500.0 463950.0 200700.0 465750.0 ;
      RECT  49800.0 464100.0 48000.0 465900.0 ;
      RECT  197100.0 466650.0 195300.0 468450.0 ;
      RECT  49800.0 466800.0 48000.0 468600.0 ;
   END
   END    sram_1rw_32b_512w_1bank_scn3me_subm
END    LIBRARY
