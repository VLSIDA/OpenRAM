
.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dint net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dint vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dint net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dint net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dint vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n

M_8 dout_bar dint vdd vdd pmos_vtg w=180.0n l=50.0n
M_9 dout_bar dint gnd gnd nmos_vtg w=90.0n l=50.0n
M_10 dout dout_bar vdd vdd pmos_vtg w=540.0n l=50.0n
M_11 dout dout_bar gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp

