magic
tech sky130A
magscale 1 2
timestamp 1590785357
<< nwell >>
rect -152 920 656 1366
rect -152 422 654 424
rect -152 138 656 422
<< nmos >>
rect 183 1713 213 1913
rect 271 1713 301 1913
rect 183 1435 213 1507
rect 271 1435 301 1507
rect 183 736 213 846
rect 271 736 301 846
rect 115 492 145 602
rect 203 492 233 602
rect 303 530 333 602
<< pmos >>
rect 183 1219 213 1329
rect 271 1219 301 1329
rect 183 956 213 1066
rect 271 956 301 1066
rect 115 262 145 372
rect 203 262 233 372
rect 291 262 321 372
<< ndiff >>
rect 129 1901 183 1913
rect 129 1725 137 1901
rect 171 1725 183 1901
rect 129 1713 183 1725
rect 213 1901 271 1913
rect 213 1725 225 1901
rect 259 1725 271 1901
rect 213 1713 271 1725
rect 301 1901 355 1913
rect 301 1725 313 1901
rect 347 1725 355 1901
rect 301 1713 355 1725
rect 129 1495 183 1507
rect 129 1449 137 1495
rect 171 1449 183 1495
rect 129 1435 183 1449
rect 213 1495 271 1507
rect 213 1449 225 1495
rect 259 1449 271 1495
rect 213 1435 271 1449
rect 301 1495 355 1507
rect 301 1449 313 1495
rect 347 1449 355 1495
rect 301 1435 355 1449
rect 129 834 183 846
rect 129 748 137 834
rect 171 748 183 834
rect 129 736 183 748
rect 213 736 271 846
rect 301 834 359 846
rect 301 748 313 834
rect 347 748 359 834
rect 301 736 359 748
rect 61 590 115 602
rect 61 504 69 590
rect 103 504 115 590
rect 61 492 115 504
rect 145 590 203 602
rect 145 504 157 590
rect 191 504 203 590
rect 145 492 203 504
rect 233 590 303 602
rect 233 504 245 590
rect 279 530 303 590
rect 333 590 391 602
rect 333 542 345 590
rect 379 542 391 590
rect 333 530 391 542
rect 279 504 287 530
rect 233 492 287 504
<< pdiff >>
rect 129 1317 183 1329
rect 129 1232 137 1317
rect 171 1232 183 1317
rect 129 1219 183 1232
rect 213 1317 271 1329
rect 213 1232 225 1317
rect 259 1232 271 1317
rect 213 1219 271 1232
rect 301 1317 355 1329
rect 301 1232 313 1317
rect 347 1232 355 1317
rect 301 1219 355 1232
rect 129 1054 183 1066
rect 129 968 137 1054
rect 171 968 183 1054
rect 129 956 183 968
rect 213 1054 271 1066
rect 213 968 225 1054
rect 259 968 271 1054
rect 213 956 271 968
rect 301 1054 356 1066
rect 301 968 313 1054
rect 347 968 356 1054
rect 301 956 356 968
rect 61 360 115 372
rect 61 274 69 360
rect 103 274 115 360
rect 61 262 115 274
rect 145 360 203 372
rect 145 274 157 360
rect 191 274 203 360
rect 145 262 203 274
rect 233 360 291 372
rect 233 274 245 360
rect 279 274 291 360
rect 233 262 291 274
rect 321 360 376 372
rect 321 274 333 360
rect 367 274 376 360
rect 321 262 376 274
<< ndiffc >>
rect 137 1725 171 1901
rect 225 1725 259 1901
rect 313 1725 347 1901
rect 137 1449 171 1495
rect 225 1449 259 1495
rect 313 1449 347 1495
rect 137 748 171 834
rect 313 748 347 834
rect 69 504 103 590
rect 157 504 191 590
rect 245 504 279 590
rect 345 542 379 590
<< pdiffc >>
rect 137 1232 171 1317
rect 225 1232 259 1317
rect 313 1232 347 1317
rect 137 968 171 1054
rect 225 968 259 1054
rect 313 968 347 1054
rect 69 274 103 360
rect 157 274 191 360
rect 245 274 279 360
rect 333 274 367 360
<< psubdiff >>
rect 229 1561 259 1595
rect 293 1561 321 1595
rect 431 790 465 820
rect 431 728 465 756
<< nsubdiff >>
rect 225 1124 259 1158
rect 293 1124 321 1158
rect 249 174 279 208
rect 313 174 341 208
<< psubdiffcont >>
rect 259 1561 293 1595
rect 431 756 465 790
<< nsubdiffcont >>
rect 259 1124 293 1158
rect 279 174 313 208
<< poly >>
rect 183 1983 409 2011
rect 183 1981 445 1983
rect 183 1913 213 1981
rect 379 1973 445 1981
rect 379 1939 395 1973
rect 429 1939 445 1973
rect 271 1913 301 1939
rect 379 1929 445 1939
rect 183 1687 213 1713
rect 271 1641 301 1713
rect 121 1631 301 1641
rect 121 1597 137 1631
rect 171 1611 301 1631
rect 171 1597 187 1611
rect 121 1585 187 1597
rect 183 1507 213 1533
rect 271 1507 301 1533
rect 183 1329 213 1435
rect 271 1329 301 1435
rect 183 1204 213 1219
rect 78 1174 213 1204
rect 271 1204 301 1219
rect 271 1174 406 1204
rect 41 1164 108 1174
rect 41 1130 57 1164
rect 91 1130 108 1164
rect 376 1164 443 1174
rect 41 1120 108 1130
rect 376 1144 393 1164
rect 377 1130 393 1144
rect 427 1130 443 1164
rect 377 1120 443 1130
rect 183 1066 213 1092
rect 271 1066 301 1092
rect 183 846 213 956
rect 271 846 301 956
rect 183 720 213 736
rect 115 690 213 720
rect 271 720 301 736
rect 271 690 399 720
rect 115 602 145 690
rect 365 680 449 690
rect 365 660 399 680
rect 375 646 399 660
rect 433 646 449 680
rect 375 636 449 646
rect 203 602 233 628
rect 303 602 333 628
rect 115 372 145 492
rect 203 476 233 492
rect 303 476 333 530
rect 203 446 333 476
rect 203 372 233 446
rect 291 372 321 446
rect 115 150 145 262
rect 101 148 145 150
rect 101 134 155 148
rect 101 100 111 134
rect 145 100 155 134
rect 203 130 233 262
rect 291 236 321 262
rect 203 100 287 130
rect 101 84 155 100
rect 255 64 287 100
rect 255 54 317 64
rect 255 20 267 54
rect 301 20 317 54
rect 255 4 317 20
<< polycont >>
rect 395 1939 429 1973
rect 137 1597 171 1631
rect 57 1130 91 1164
rect 393 1130 427 1164
rect 399 646 433 680
rect 111 100 145 134
rect 267 20 301 54
<< locali >>
rect 381 1973 429 1989
rect 137 1901 171 1913
rect 137 1709 171 1725
rect 225 1901 259 1927
rect 117 1631 171 1647
rect 117 1597 137 1631
rect 117 1580 171 1597
rect 137 1495 171 1580
rect 137 1317 171 1449
rect 225 1595 259 1725
rect 313 1901 347 1913
rect 313 1709 347 1725
rect 381 1939 395 1973
rect 381 1923 429 1939
rect 293 1561 309 1595
rect 225 1495 259 1561
rect 225 1433 259 1449
rect 313 1495 347 1513
rect 313 1399 347 1449
rect 381 1399 415 1923
rect 313 1365 415 1399
rect 137 1216 171 1232
rect 225 1317 259 1333
rect 57 1164 103 1180
rect 91 1130 103 1164
rect 57 1114 103 1130
rect 69 590 103 1114
rect 225 1158 259 1232
rect 313 1317 347 1365
rect 313 1216 347 1232
rect 381 1164 427 1180
rect 293 1124 309 1158
rect 381 1130 393 1164
rect 137 1054 171 1070
rect 137 918 171 968
rect 225 1054 259 1124
rect 381 1114 427 1130
rect 225 952 259 968
rect 313 1054 347 1070
rect 313 918 347 968
rect 381 918 415 1114
rect 137 884 415 918
rect 137 834 171 884
rect 137 730 171 748
rect 313 834 347 850
rect 347 790 360 824
rect 394 790 471 824
rect 313 732 347 748
rect 431 740 465 756
rect 387 680 433 698
rect 387 646 399 680
rect 387 632 433 646
rect 69 444 103 504
rect 157 590 191 606
rect 157 488 191 504
rect 245 488 279 504
rect 345 622 433 632
rect 345 598 421 622
rect 345 590 391 598
rect 379 578 391 590
rect 69 410 191 444
rect 345 424 379 542
rect 69 360 103 376
rect 69 208 103 274
rect 157 360 191 410
rect 333 390 379 424
rect 157 258 191 274
rect 245 360 279 376
rect 245 208 279 274
rect 333 360 367 390
rect 333 258 367 274
rect 69 174 245 208
rect 313 174 329 208
rect 245 168 279 174
rect 94 100 111 134
rect 145 100 161 134
rect 251 20 267 54
rect 301 20 317 54
<< viali >>
rect 137 1913 171 1947
rect 313 1913 347 1947
rect 225 1561 259 1595
rect 225 1124 259 1158
rect 360 790 394 824
rect 245 590 279 624
rect 245 174 279 208
rect 111 100 145 134
rect 267 20 301 54
<< metal1 >>
rect 126 1959 156 2011
rect 328 1959 358 2011
rect 125 1947 182 1959
rect 125 1913 137 1947
rect 171 1913 182 1947
rect 125 1901 182 1913
rect 302 1947 359 1959
rect 302 1913 313 1947
rect 347 1913 359 1947
rect 302 1901 359 1913
rect 213 1595 299 1601
rect 213 1561 225 1595
rect 259 1561 321 1595
rect 213 1555 299 1561
rect 213 1158 299 1164
rect 213 1124 225 1158
rect 259 1124 299 1158
rect 213 1118 299 1124
rect 334 824 420 830
rect 334 790 360 824
rect 394 790 420 824
rect 334 789 420 790
rect 347 784 420 789
rect 219 624 305 630
rect 219 590 245 624
rect 279 590 305 624
rect 219 584 305 590
rect 233 208 319 214
rect 233 174 245 208
rect 279 174 319 208
rect 233 168 319 174
rect 99 134 157 156
rect 99 100 111 134
rect 145 128 157 134
rect 145 100 500 128
rect 99 94 500 100
rect 255 54 315 60
rect 255 20 267 54
rect 301 20 315 54
rect 255 4 315 20
<< labels >>
rlabel metal1 106 118 106 118 1 en
rlabel metal1 296 210 296 210 1 vdd
rlabel metal1 285 12 285 12 1 din
rlabel metal1 262 626 262 626 1 gnd
rlabel metal1 393 827 393 827 1 gnd
rlabel metal1 220 1140 220 1140 1 vdd
rlabel metal1 340 1973 340 1973 1 br
rlabel metal1 140 1981 140 1981 1 bl
rlabel metal1 220 1577 220 1577 1 gnd
<< properties >>
string FIXED_BBOX 0 0 500 2011
<< end >>
